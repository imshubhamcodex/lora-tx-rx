PK
     ��Z���BF BF    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0":["pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0"],"pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_1":["pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0":["pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0","pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1":["pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2":["pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3":["pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4":["pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5":["pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6":["pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7":["pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8":["pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9":["pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10":["pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11":["pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12":["pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13":["pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14":["pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15":["pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_1"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_18"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_17":[],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_18":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_19":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_27"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_20":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_26"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_21":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_25"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_22":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_24"],"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_23":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_23"],"pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_0":["pin-type-component_7e9999e8-686e-4f02-b1e7-bee04a417b43_0"],"pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_1":["pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_1"],"pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2":["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2"],"pin-type-component_7e9999e8-686e-4f02-b1e7-bee04a417b43_0":["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_0"],"pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_0":["pin-type-component_4bfdc0b0-0087-4f19-b9da-fe77fe2030bb_0"],"pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_1":["pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_1"],"pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2":["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1"],"pin-type-component_4bfdc0b0-0087-4f19-b9da-fe77fe2030bb_0":["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_0"],"pin-type-component_725c2e06-513a-456a-a054-9a1efd2410b5_0":["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_0"],"pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_0":["pin-type-component_84e67de5-59f5-4375-8901-060561a64dc9_0"],"pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_1":["pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_1"],"pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2":["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1"],"pin-type-component_84e67de5-59f5-4375-8901-060561a64dc9_0":["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_0"],"pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_0":["pin-type-component_725c2e06-513a-456a-a054-9a1efd2410b5_0"],"pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_1":["pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_1"],"pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2":["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2"],"pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_0":["pin-type-component_ad7b12e6-293b-4cf0-b5fc-2ad4811766ad_0"],"pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_1":["pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_1"],"pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2":["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0"],"pin-type-component_ad7b12e6-293b-4cf0-b5fc-2ad4811766ad_0":["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_0"],"pin-type-component_84525e3e-ef29-4e0c-a293-959707966b26_0":["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_0"],"pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_0":["pin-type-component_a4a81ac1-f999-4c5f-bf1d-d39d1364ba7e_0"],"pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_1":["pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_1"],"pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2":["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1"],"pin-type-component_a4a81ac1-f999-4c5f-bf1d-d39d1364ba7e_0":["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_0"],"pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_0":["pin-type-component_84525e3e-ef29-4e0c-a293-959707966b26_0"],"pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_1":["pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_1"],"pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2":["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2"],"pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_0":["pin-type-component_69b6c16b-f2c6-4ab0-b694-b43efd7d7efa_0"],"pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_1":["pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_1"],"pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2":["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2"],"pin-type-component_69b6c16b-f2c6-4ab0-b694-b43efd7d7efa_0":["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_0"],"pin-type-component_7fc8671b-e701-4c33-a644-f42eace24307_0":["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_0"],"pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_0":["pin-type-component_266aa6bb-5bae-4ff3-85db-bbd370178ae8_0"],"pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_1":["pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_1"],"pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2":["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1"],"pin-type-component_266aa6bb-5bae-4ff3-85db-bbd370178ae8_0":["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_0"],"pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_0":["pin-type-component_7fc8671b-e701-4c33-a644-f42eace24307_0"],"pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_1":["pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_1"],"pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2":["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2"],"pin-type-component_0af45fa8-24bc-42e4-9c24-d15187e9fbc3_0":["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_0"],"pin-type-component_5278fc75-d95d-4e4c-a86e-2e83a862e607_0":["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_0"],"pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_0":["pin-type-component_0af45fa8-24bc-42e4-9c24-d15187e9fbc3_0"],"pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1":["pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_1"],"pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2":["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2"],"pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_0":["pin-type-component_5278fc75-d95d-4e4c-a86e-2e83a862e607_0"],"pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_1":["pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_1"],"pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2":["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1"],"pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_0":["pin-type-component_e7d36833-6d1a-490c-96e9-4f178d942f47_0"],"pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_1":["pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_1"],"pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2":["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2"],"pin-type-component_e7d36833-6d1a-490c-96e9-4f178d942f47_0":["pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_0"],"pin-type-component_3d109b51-1504-4d24-a9e7-9e3fe3074724_0":["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_0"],"pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_0":["pin-type-component_34445add-d974-48d4-81af-972f5dd7934b_0"],"pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_1":["pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_1"],"pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2":["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1"],"pin-type-component_34445add-d974-48d4-81af-972f5dd7934b_0":["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_0"],"pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_0":["pin-type-component_3d109b51-1504-4d24-a9e7-9e3fe3074724_0"],"pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_1":["pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_1"],"pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2":["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2"],"pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_0":["pin-type-component_903934ae-30da-4a37-93c9-c64660e9c617_0"],"pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_1":["pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_1"],"pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2":["pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2","pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1"],"pin-type-component_903934ae-30da-4a37-93c9-c64660e9c617_0":["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_0"],"pin-type-component_5bdd54e6-172a-4994-8b34-5d8687be61e2_0":["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_0"],"pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_0":["pin-type-component_62a268f0-68fa-4016-91c7-d55a738d6b46_0"],"pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_1":["pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_1"],"pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2":["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1"],"pin-type-component_62a268f0-68fa-4016-91c7-d55a738d6b46_0":["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_0"],"pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_0":["pin-type-component_5bdd54e6-172a-4994-8b34-5d8687be61e2_0"],"pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_1":["pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_1"],"pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2":["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2"],"pin-type-component_4732636d-ea0d-4b19-877e-d2ff4ddb5e8d_0":["pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_0"],"pin-type-component_7f294ee1-7ea8-4e70-bb0a-8c8b6b15b6c9_0":["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_0"],"pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_0":["pin-type-component_4732636d-ea0d-4b19-877e-d2ff4ddb5e8d_0"],"pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_1":["pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_1"],"pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2":["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2"],"pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_0":["pin-type-component_7f294ee1-7ea8-4e70-bb0a-8c8b6b15b6c9_0"],"pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_1":["pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_1"],"pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2":["pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1"],"pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_0":["pin-type-component_b2f3a979-ce1b-444a-a7e4-6ef67b25f077_0"],"pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_1":["pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_1"],"pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2":["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1"],"pin-type-component_b2f3a979-ce1b-444a-a7e4-6ef67b25f077_0":["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_0"],"pin-type-component_0b4ba5d8-bcb4-4816-8dfe-3fa4ce9ed019_0":["pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_0"],"pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_0":["pin-type-component_29f2dcbd-c66e-4d22-9415-91c6505cd16b_0"],"pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_1":["pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_1"],"pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2":["pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1"],"pin-type-component_29f2dcbd-c66e-4d22-9415-91c6505cd16b_0":["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_0"],"pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_0":["pin-type-component_0b4ba5d8-bcb4-4816-8dfe-3fa4ce9ed019_0"],"pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_1":["pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_1"],"pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2":["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2"],"pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_0":["pin-type-component_3b6d34de-cd89-4ef4-9473-da4b3ae907df_0"],"pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_1":["pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_1"],"pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2":["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2"],"pin-type-component_3b6d34de-cd89-4ef4-9473-da4b3ae907df_0":["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_0"],"pin-type-component_dd44450f-fd4f-4059-aab9-565428093e7b_0":["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_0"],"pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_0":["pin-type-component_6d57b374-4a97-4f2c-b0da-4d4ccbef4f5a_0"],"pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_1":["pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_1"],"pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2":["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1"],"pin-type-component_6d57b374-4a97-4f2c-b0da-4d4ccbef4f5a_0":["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_0"],"pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_0":["pin-type-component_dd44450f-fd4f-4059-aab9-565428093e7b_0"],"pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_1":["pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_1"],"pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2":["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1"],"pin-type-component_0c082f01-0561-48cc-887e-4e37deace687_0":["pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_0"],"pin-type-component_d1e6942e-6a34-4356-87fa-da19b68ae6b8_0":["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_0"],"pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_0":["pin-type-component_0c082f01-0561-48cc-887e-4e37deace687_0"],"pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_1":["pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_1"],"pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2":["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1"],"pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_0":["pin-type-component_d1e6942e-6a34-4356-87fa-da19b68ae6b8_0"],"pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_1":["pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_1"],"pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2":["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1"],"pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_0":["pin-type-component_bb4a8fb4-80b5-4764-a9f6-b3d9cae671c4_0"],"pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1":["pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1"],"pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2":["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1"],"pin-type-component_bb4a8fb4-80b5-4764-a9f6-b3d9cae671c4_0":["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_0"],"pin-type-component_636bd670-72c8-425e-8740-11540fc72a9f_0":["pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_0"],"pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_0":["pin-type-component_e84ff89e-b801-43e3-905a-a7004860c743_0"],"pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1":["pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1"],"pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2":["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1"],"pin-type-component_e84ff89e-b801-43e3-905a-a7004860c743_0":["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_0"],"pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_0":["pin-type-component_636bd670-72c8-425e-8740-11540fc72a9f_0"],"pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_1":["pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_1"],"pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2":["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1"],"pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_0":["pin-type-component_edb09e16-b982-4564-8c59-d0c31b14f784_0"],"pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_1":["pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_1"],"pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2":["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1"],"pin-type-component_edb09e16-b982-4564-8c59-d0c31b14f784_0":["pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_0"],"pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0":["pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15"],"pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1":["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_0":["pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_1":["pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_2":["pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_3":["pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_4":["pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_5":["pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_6":["pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_7":["pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8":["pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9":["pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10":["pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11":["pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12":["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13":["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14":["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15":["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16":["pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_18"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_17":[],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_18":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_19":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_8"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_20":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_9"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_21":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_10"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_22":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_11"],"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_23":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_12"],"pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0":["pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14"],"pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_1":["pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_1"],"pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_0":["pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0"],"pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1":["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1"],"pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0":["pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13"],"pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_1":["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_1"],"pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_0":["pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0"],"pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_1":["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_1"],"pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_0":["pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0"],"pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_1":["pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_1"],"pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0":["pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12"],"pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_1":["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_1"],"pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_0":["pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0"],"pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_1":["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_1"],"pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0":["pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11"],"pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_1":["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_1"],"pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_0":["pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0"],"pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_1":["pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_1"],"pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0":["pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10"],"pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_1":["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_1"],"pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_0":["pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0"],"pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_1":["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_1"],"pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0":["pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9"],"pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_1":["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_1"],"pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_0":["pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0"],"pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_1":["pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_1"],"pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0":["pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8"],"pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_1":["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_1"],"pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_0":["pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0"],"pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_1":["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_1"],"pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0":["pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7"],"pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_1":["pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_1"],"pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0":["pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6"],"pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_1":["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_1"],"pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_0":["pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0"],"pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_1":["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_1"],"pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0":["pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5"],"pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_1":["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_1"],"pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_0":["pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0"],"pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_1":["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_1"],"pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_0":["pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0"],"pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_1":["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1"],"pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0":["pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4"],"pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_1":["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_1"],"pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_0":["pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0"],"pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_1":["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_1"],"pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0":["pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0"],"pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_1":["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_1"],"pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_0":["pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0"],"pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_1":["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_1"],"pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0":["pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1"],"pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_1":["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_1"],"pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_0":["pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0"],"pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_1":["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_1"],"pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0":["pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2"],"pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_1":["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_1"],"pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_0":["pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0"],"pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_1":["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_1"],"pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0":["pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3"],"pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_1":["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_1"],"pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0":["pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0"],"pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1":["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0"],"pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0":["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1"],"pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1":["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12"],"pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0":["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"],"pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1":["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0"],"pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0":["pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1"],"pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1":["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13"],"pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0":["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0"],"pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1":["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0"],"pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0":["pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1"],"pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1":["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14"],"pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0":["pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0","pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0"],"pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1":["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0"],"pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0":["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1"],"pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1":["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15"],"pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0":["pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0"],"pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_1":["pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_0"],"pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_0":["pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_1"],"pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1":["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11"],"pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0":["pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0"],"pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_1":["pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_0"],"pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_0":["pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_1"],"pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1":["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10"],"pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0":["pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0","pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0"],"pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_1":["pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_0"],"pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_0":["pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_1"],"pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1":["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9"],"pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0":["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0","pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0"],"pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_1":["pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_0"],"pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_0":["pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_1"],"pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1":["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8"],"pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0":["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0"],"pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_1":["pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_0"],"pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_0":["pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_1"],"pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1":["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_7"],"pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0":["pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0","pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0"],"pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_1":["pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_0"],"pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_0":["pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_1"],"pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1":["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_6"],"pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0":["pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0","pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_0"],"pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_1":["pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_0"],"pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_0":["pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_1"],"pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1":["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_5"],"pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_0":["pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0"],"pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_1":["pin-type-component_c107267e-960a-414d-898a-9b8f86844804_0"],"pin-type-component_c107267e-960a-414d-898a-9b8f86844804_0":["pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_1"],"pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1":["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_4"],"pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0":["pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10"],"pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1":["pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_0","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2"],"pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_0":["pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1"],"pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_1":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_0"],"pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0":["pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0"],"pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1":["pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_0","pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2"],"pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_0":["pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1"],"pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_1":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_1"],"pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0":["pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0"],"pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1":["pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_0","pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2"],"pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_0":["pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1"],"pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_1":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_2"],"pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0":["pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0"],"pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_1":["pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0"],"pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0":["pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_1","pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2"],"pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_1":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_3"],"pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0"],"pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1"],"pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2"],"pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3"],"pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4"],"pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5"],"pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6"],"pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7"],"pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8"],"pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9"],"pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10"],"pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11"],"pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12"],"pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13"],"pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14"],"pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_0":["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],"pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_1":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15"],"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0":["pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_0","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_0","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_0","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_0","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_0","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_0","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_0","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_0","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_0","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_0","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_0","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_0","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_0","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_0","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_0","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16"],"pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_6"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_0":[],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_1":[],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_2":[],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_3":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_4":[],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_5":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_9"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_6":["pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_7":["pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_4"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_8":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_19"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_9":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_20"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_10":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_21"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_11":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_22"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_12":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_23"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_13":[],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_14":[],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_15":[],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_16":[],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_17":["pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_3"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_18":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_4"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_19":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_3"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_20":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_2"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_21":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_1"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_22":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_11"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_23":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_23"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_24":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_22"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_25":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_21"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_26":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_20"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_27":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_19"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_28":[],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_29":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_12"],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_30":[],"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_31":[],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_0":[],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_1":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_21"],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_2":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_20"],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_3":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_19"],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_4":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_18"],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_5":[],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_6":[],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_7":[],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_8":[],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_9":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_5"],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_3","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0"],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_11":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_22"],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_12":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_29"],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_13":[],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_14":[],"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_15":[],"pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_0":[],"pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_1":[],"pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_2":[],"pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_3":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_17"],"pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_4":["pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_7"]},"pin_to_color":{"pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0":"#010067","pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_1":"#0076FF","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0":"#001eff","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1":"#00FFC6","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2":"#010067","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3":"#ff0066","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4":"#90FB92","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5":"#7E2DD2","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6":"#774D00","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7":"#7544B1","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8":"#FE8900","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9":"#98FF52","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10":"#683D3B","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11":"#008F9C","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12":"#6A826C","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13":"#001544","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14":"#005F39","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15":"#010067","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16":"#008F9C","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_17":"#000000","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_18":"#008F9C","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_19":"#FF029D","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_20":"#683D3B","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_21":"#FF74A3","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_22":"#968AE8","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_23":"#98FF52","pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_0":"#FF74A3","pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_1":"#0076FF","pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2":"#0E4CA1","pin-type-component_7e9999e8-686e-4f02-b1e7-bee04a417b43_0":"#FF74A3","pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_0":"#98FF52","pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_1":"#85A900","pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2":"#0E4CA1","pin-type-component_4bfdc0b0-0087-4f19-b9da-fe77fe2030bb_0":"#98FF52","pin-type-component_725c2e06-513a-456a-a054-9a1efd2410b5_0":"#01FFFE","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_0":"#BDC6FF","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_1":"#E56FFE","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2":"#9E008E","pin-type-component_84e67de5-59f5-4375-8901-060561a64dc9_0":"#BDC6FF","pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_0":"#01FFFE","pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_1":"#BDD393","pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2":"#9E008E","pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_0":"#004754","pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_1":"#0E4CA1","pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2":"#005F39","pin-type-component_ad7b12e6-293b-4cf0-b5fc-2ad4811766ad_0":"#004754","pin-type-component_84525e3e-ef29-4e0c-a293-959707966b26_0":"#774D00","pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_0":"#A5FFD2","pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_1":"#E85EBE","pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2":"#ff1100","pin-type-component_a4a81ac1-f999-4c5f-bf1d-d39d1364ba7e_0":"#A5FFD2","pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_0":"#774D00","pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_1":"#FF6E41","pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2":"#ff1100","pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_0":"#90FB92","pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_1":"#9E008E","pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2":"#005F39","pin-type-component_69b6c16b-f2c6-4ab0-b694-b43efd7d7efa_0":"#90FB92","pin-type-component_7fc8671b-e701-4c33-a644-f42eace24307_0":"#FF6E41","pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_0":"#85A900","pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_1":"#004754","pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2":"#85A900","pin-type-component_266aa6bb-5bae-4ff3-85db-bbd370178ae8_0":"#85A900","pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_0":"#FF6E41","pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_1":"#7A4782","pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2":"#85A900","pin-type-component_0af45fa8-24bc-42e4-9c24-d15187e9fbc3_0":"#00FF78","pin-type-component_5278fc75-d95d-4e4c-a86e-2e83a862e607_0":"#BDD393","pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_0":"#00FF78","pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1":"#FFB167","pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2":"#0076FF","pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_0":"#BDD393","pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_1":"#6685ff","pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2":"#0076FF","pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_0":"#005F39","pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_1":"#BB8800","pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2":"#FF6E41","pin-type-component_e7d36833-6d1a-490c-96e9-4f178d942f47_0":"#005F39","pin-type-component_3d109b51-1504-4d24-a9e7-9e3fe3074724_0":"#0E4CA1","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_0":"#010067","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_1":"#FFA6FE","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2":"#00FFC6","pin-type-component_34445add-d974-48d4-81af-972f5dd7934b_0":"#010067","pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_0":"#0E4CA1","pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_1":"#A5FFD2","pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2":"#00FFC6","pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_0":"#FF937E","pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_1":"#BDC6FF","pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2":"#FF6E41","pin-type-component_903934ae-30da-4a37-93c9-c64660e9c617_0":"#FF937E","pin-type-component_5bdd54e6-172a-4994-8b34-5d8687be61e2_0":"#5FAD4E","pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_0":"#C28C9F","pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_1":"#968AE8","pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2":"#004754","pin-type-component_62a268f0-68fa-4016-91c7-d55a738d6b46_0":"#C28C9F","pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_0":"#5FAD4E","pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_1":"#FF74A3","pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2":"#004754","pin-type-component_4732636d-ea0d-4b19-877e-d2ff4ddb5e8d_0":"#007DB5","pin-type-component_7f294ee1-7ea8-4e70-bb0a-8c8b6b15b6c9_0":"#91D0CB","pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_0":"#007DB5","pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_1":"#A75740","pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2":"#7A4782","pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_0":"#91D0CB","pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_1":"#01FFFE","pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2":"#7A4782","pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_0":"#BDD393","pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_1":"#C28C9F","pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2":"#f50a0a","pin-type-component_b2f3a979-ce1b-444a-a7e4-6ef67b25f077_0":"#BDD393","pin-type-component_0b4ba5d8-bcb4-4816-8dfe-3fa4ce9ed019_0":"#90FB92","pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_0":"#683D3B","pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_1":"#FF029D","pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2":"#B500FF","pin-type-component_29f2dcbd-c66e-4d22-9415-91c6505cd16b_0":"#683D3B","pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_0":"#90FB92","pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_1":"#5FAD4E","pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2":"#B500FF","pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_0":"#00FF78","pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_1":"#00AE7E","pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2":"#f50a0a","pin-type-component_3b6d34de-cd89-4ef4-9473-da4b3ae907df_0":"#00FF78","pin-type-component_dd44450f-fd4f-4059-aab9-565428093e7b_0":"#BB8800","pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_0":"#FE8900","pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_1":"#FF937E","pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2":"#008F9C","pin-type-component_6d57b374-4a97-4f2c-b0da-4d4ccbef4f5a_0":"#FE8900","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_0":"#BB8800","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_1":"#95003A","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2":"#008F9C","pin-type-component_0c082f01-0561-48cc-887e-4e37deace687_0":"#A75740","pin-type-component_d1e6942e-6a34-4356-87fa-da19b68ae6b8_0":"#968AE8","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_0":"#A75740","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_1":"#007DB5","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2":"#007DB5","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_0":"#968AE8","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_1":"#91D0CB","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2":"#007DB5","pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_0":"#004754","pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1":"#FF6E41","pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2":"#FE8900","pin-type-component_bb4a8fb4-80b5-4764-a9f6-b3d9cae671c4_0":"#004754","pin-type-component_636bd670-72c8-425e-8740-11540fc72a9f_0":"#774D00","pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_0":"#A5FFD2","pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1":"#00ff88","pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2":"#968AE8","pin-type-component_e84ff89e-b801-43e3-905a-a7004860c743_0":"#A5FFD2","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_0":"#774D00","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_1":"#0E4CA1","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2":"#968AE8","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_0":"#66ffa8","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_1":"#0076FF","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2":"#FE8900","pin-type-component_edb09e16-b982-4564-8c59-d0c31b14f784_0":"#66ffa8","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0":"#010067","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1":"#FF6E41","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_0":"#007DB5","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_1":"#6A826C","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_2":"#00AE7E","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_3":"#C28C9F","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_4":"#0076FF","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_5":"#85A900","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_6":"#00FFC6","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_7":"#FF6E41","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8":"#7A4782","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9":"#004754","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10":"#B500FF","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11":"#f50a0a","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12":"#007DB5","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13":"#008F9C","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14":"#968AE8","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15":"#FE8900","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16":"#5FAD4E","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_17":"#000000","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_18":"#5FAD4E","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_19":"#A75740","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_20":"#01FFFE","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_21":"#FE8900","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_22":"#BDC6FF","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_23":"#BB8800","pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0":"#005F39","pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_1":"#0E4CA1","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_0":"#005F39","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1":"#00ff88","pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0":"#001544","pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_1":"#95003A","pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_0":"#001544","pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_1":"#FF937E","pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_0":"#6A826C","pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_1":"#007DB5","pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0":"#6A826C","pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_1":"#91D0CB","pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_0":"#008F9C","pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_1":"#00AE7E","pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0":"#008F9C","pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_1":"#C28C9F","pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_0":"#683D3B","pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_1":"#5FAD4E","pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0":"#683D3B","pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_1":"#FF029D","pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_0":"#98FF52","pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_1":"#FF74A3","pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0":"#98FF52","pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_1":"#968AE8","pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_0":"#FE8900","pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_1":"#A75740","pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0":"#FE8900","pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_1":"#01FFFE","pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_0":"#7544B1","pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_1":"#BDC6FF","pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0":"#7544B1","pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_1":"#BB8800","pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0":"#774D00","pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_1":"#A5FFD2","pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_0":"#774D00","pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_1":"#FFA6FE","pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0":"#7E2DD2","pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_1":"#7A4782","pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_0":"#7E2DD2","pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_1":"#004754","pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_0":"#90FB92","pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_1":"#FFB167","pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0":"#90FB92","pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_1":"#6685ff","pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_0":"#001eff","pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_1":"#BDD393","pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0":"#001eff","pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_1":"#E56FFE","pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_0":"#00FFC6","pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_1":"#0076FF","pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0":"#00FFC6","pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_1":"#85A900","pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_0":"#010067","pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_1":"#FF6E41","pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0":"#010067","pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_1":"#E85EBE","pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_0":"#ff0066","pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_1":"#9E008E","pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0":"#ff0066","pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_1":"#0E4CA1","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0":"#7E2DD2","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1":"#91D0CB","pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0":"#91D0CB","pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1":"#007DB5","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0":"#7E2DD2","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1":"#A5FFD2","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0":"#A5FFD2","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1":"#008F9C","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0":"#7E2DD2","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1":"#FFA6FE","pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0":"#FFA6FE","pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1":"#968AE8","pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0":"#7E2DD2","pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1":"#774D00","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0":"#774D00","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1":"#FE8900","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0":"#7E2DD2","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_1":"#010067","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_0":"#010067","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1":"#f50a0a","pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0":"#7E2DD2","pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_1":"#E85EBE","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_0":"#E85EBE","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1":"#B500FF","pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0":"#7E2DD2","pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_1":"#90FB92","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_0":"#90FB92","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1":"#004754","pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0":"#7E2DD2","pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_1":"#FFDB66","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_0":"#FFDB66","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1":"#7A4782","pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0":"#7E2DD2","pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_1":"#00FF78","pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_0":"#00FF78","pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1":"#FF6E41","pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0":"#7E2DD2","pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_1":"#E56FFE","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_0":"#E56FFE","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1":"#00FFC6","pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0":"#7E2DD2","pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_1":"#BDD393","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_0":"#BDD393","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1":"#85A900","pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_0":"#7E2DD2","pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_1":"#7E2DD2","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_0":"#7E2DD2","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1":"#0076FF","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0":"#7E2DD2","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1":"#9E008E","pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_0":"#9E008E","pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_1":"#007DB5","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0":"#7E2DD2","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1":"#0E4CA1","pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_0":"#0E4CA1","pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_1":"#6A826C","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0":"#7E2DD2","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1":"#ff1100","pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_0":"#ff1100","pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_1":"#00AE7E","pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0":"#7E2DD2","pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_1":"#005F39","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0":"#005F39","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_1":"#C28C9F","pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_0":"#008F9C","pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_1":"#001eff","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_0":"#008F9C","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_1":"#00FFC6","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_0":"#008F9C","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_1":"#010067","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_0":"#008F9C","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_1":"#ff0066","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_0":"#008F9C","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_1":"#90FB92","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_0":"#008F9C","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_1":"#7E2DD2","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_0":"#008F9C","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_1":"#774D00","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_0":"#008F9C","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_1":"#7544B1","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_0":"#008F9C","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_1":"#FE8900","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_0":"#008F9C","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_1":"#98FF52","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_0":"#008F9C","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_1":"#683D3B","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_0":"#008F9C","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_1":"#008F9C","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_0":"#008F9C","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1":"#6A826C","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_0":"#008F9C","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1":"#001544","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_0":"#008F9C","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_1":"#005F39","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_0":"#008F9C","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_1":"#010067","pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0":"#008F9C","pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0":"#5FAD4E","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_0":"#000000","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_1":"#000000","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_2":"#000000","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_3":"#7E2DD2","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_4":"#000000","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_5":"#A5FFD2","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_6":"#5FAD4E","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_7":"#f73302","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_8":"#A75740","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_9":"#01FFFE","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_10":"#FE8900","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_11":"#BDC6FF","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_12":"#BB8800","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_13":"#000000","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_14":"#000000","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_15":"#000000","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_16":"#000000","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_17":"#06f40a","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_18":"#FFB167","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_19":"#B500FF","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_20":"#004754","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_21":"#e11934","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_22":"#08d46a","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_23":"#98FF52","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_24":"#968AE8","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_25":"#FF74A3","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_26":"#683D3B","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_27":"#FF029D","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_28":"#000000","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_29":"#774D00","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_30":"#000000","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_31":"#000000","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_0":"#000000","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_1":"#e11934","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_2":"#004754","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_3":"#B500FF","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_4":"#FFB167","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_5":"#000000","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_6":"#000000","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_7":"#000000","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_8":"#000000","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_9":"#A5FFD2","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10":"#7E2DD2","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_11":"#08d46a","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_12":"#774D00","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_13":"#000000","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_14":"#000000","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_15":"#000000","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_0":"#000000","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_1":"#000000","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_2":"#000000","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_3":"#06f40a","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_4":"#f73302"},"pin_to_state":{"pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0":"neutral","pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_1":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_17":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_18":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_19":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_20":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_21":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_22":"neutral","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_23":"neutral","pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_0":"neutral","pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_1":"neutral","pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2":"neutral","pin-type-component_7e9999e8-686e-4f02-b1e7-bee04a417b43_0":"neutral","pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_0":"neutral","pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_1":"neutral","pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2":"neutral","pin-type-component_4bfdc0b0-0087-4f19-b9da-fe77fe2030bb_0":"neutral","pin-type-component_725c2e06-513a-456a-a054-9a1efd2410b5_0":"neutral","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_0":"neutral","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_1":"neutral","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2":"neutral","pin-type-component_84e67de5-59f5-4375-8901-060561a64dc9_0":"neutral","pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_0":"neutral","pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_1":"neutral","pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2":"neutral","pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_0":"neutral","pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_1":"neutral","pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2":"neutral","pin-type-component_ad7b12e6-293b-4cf0-b5fc-2ad4811766ad_0":"neutral","pin-type-component_84525e3e-ef29-4e0c-a293-959707966b26_0":"neutral","pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_0":"neutral","pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_1":"neutral","pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2":"neutral","pin-type-component_a4a81ac1-f999-4c5f-bf1d-d39d1364ba7e_0":"neutral","pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_0":"neutral","pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_1":"neutral","pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2":"neutral","pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_0":"neutral","pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_1":"neutral","pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2":"neutral","pin-type-component_69b6c16b-f2c6-4ab0-b694-b43efd7d7efa_0":"neutral","pin-type-component_7fc8671b-e701-4c33-a644-f42eace24307_0":"neutral","pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_0":"neutral","pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_1":"neutral","pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2":"neutral","pin-type-component_266aa6bb-5bae-4ff3-85db-bbd370178ae8_0":"neutral","pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_0":"neutral","pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_1":"neutral","pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2":"neutral","pin-type-component_0af45fa8-24bc-42e4-9c24-d15187e9fbc3_0":"neutral","pin-type-component_5278fc75-d95d-4e4c-a86e-2e83a862e607_0":"neutral","pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_0":"neutral","pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1":"neutral","pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2":"neutral","pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_0":"neutral","pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_1":"neutral","pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2":"neutral","pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_0":"neutral","pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_1":"neutral","pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2":"neutral","pin-type-component_e7d36833-6d1a-490c-96e9-4f178d942f47_0":"neutral","pin-type-component_3d109b51-1504-4d24-a9e7-9e3fe3074724_0":"neutral","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_0":"neutral","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_1":"neutral","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2":"neutral","pin-type-component_34445add-d974-48d4-81af-972f5dd7934b_0":"neutral","pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_0":"neutral","pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_1":"neutral","pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2":"neutral","pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_0":"neutral","pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_1":"neutral","pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2":"neutral","pin-type-component_903934ae-30da-4a37-93c9-c64660e9c617_0":"neutral","pin-type-component_5bdd54e6-172a-4994-8b34-5d8687be61e2_0":"neutral","pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_0":"neutral","pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_1":"neutral","pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2":"neutral","pin-type-component_62a268f0-68fa-4016-91c7-d55a738d6b46_0":"neutral","pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_0":"neutral","pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_1":"neutral","pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2":"neutral","pin-type-component_4732636d-ea0d-4b19-877e-d2ff4ddb5e8d_0":"neutral","pin-type-component_7f294ee1-7ea8-4e70-bb0a-8c8b6b15b6c9_0":"neutral","pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_0":"neutral","pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_1":"neutral","pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2":"neutral","pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_0":"neutral","pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_1":"neutral","pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2":"neutral","pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_0":"neutral","pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_1":"neutral","pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2":"neutral","pin-type-component_b2f3a979-ce1b-444a-a7e4-6ef67b25f077_0":"neutral","pin-type-component_0b4ba5d8-bcb4-4816-8dfe-3fa4ce9ed019_0":"neutral","pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_0":"neutral","pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_1":"neutral","pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2":"neutral","pin-type-component_29f2dcbd-c66e-4d22-9415-91c6505cd16b_0":"neutral","pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_0":"neutral","pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_1":"neutral","pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2":"neutral","pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_0":"neutral","pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_1":"neutral","pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2":"neutral","pin-type-component_3b6d34de-cd89-4ef4-9473-da4b3ae907df_0":"neutral","pin-type-component_dd44450f-fd4f-4059-aab9-565428093e7b_0":"neutral","pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_0":"neutral","pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_1":"neutral","pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2":"neutral","pin-type-component_6d57b374-4a97-4f2c-b0da-4d4ccbef4f5a_0":"neutral","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_0":"neutral","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_1":"neutral","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2":"neutral","pin-type-component_0c082f01-0561-48cc-887e-4e37deace687_0":"neutral","pin-type-component_d1e6942e-6a34-4356-87fa-da19b68ae6b8_0":"neutral","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_0":"neutral","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_1":"neutral","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2":"neutral","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_0":"neutral","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_1":"neutral","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2":"neutral","pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_0":"neutral","pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1":"neutral","pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2":"neutral","pin-type-component_bb4a8fb4-80b5-4764-a9f6-b3d9cae671c4_0":"neutral","pin-type-component_636bd670-72c8-425e-8740-11540fc72a9f_0":"neutral","pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_0":"neutral","pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1":"neutral","pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2":"neutral","pin-type-component_e84ff89e-b801-43e3-905a-a7004860c743_0":"neutral","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_0":"neutral","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_1":"neutral","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2":"neutral","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_0":"neutral","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_1":"neutral","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2":"neutral","pin-type-component_edb09e16-b982-4564-8c59-d0c31b14f784_0":"neutral","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0":"neutral","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_0":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_1":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_2":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_3":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_4":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_5":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_6":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_7":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_17":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_18":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_19":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_20":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_21":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_22":"neutral","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_23":"neutral","pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0":"neutral","pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_1":"neutral","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_0":"neutral","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1":"neutral","pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0":"neutral","pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_1":"neutral","pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_0":"neutral","pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_1":"neutral","pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_0":"neutral","pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_1":"neutral","pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0":"neutral","pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_1":"neutral","pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_0":"neutral","pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_1":"neutral","pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0":"neutral","pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_1":"neutral","pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_0":"neutral","pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_1":"neutral","pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0":"neutral","pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_1":"neutral","pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_0":"neutral","pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_1":"neutral","pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0":"neutral","pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_1":"neutral","pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_0":"neutral","pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_1":"neutral","pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0":"neutral","pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_1":"neutral","pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_0":"neutral","pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_1":"neutral","pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0":"neutral","pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_1":"neutral","pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0":"neutral","pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_1":"neutral","pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_0":"neutral","pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_1":"neutral","pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0":"neutral","pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_1":"neutral","pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_0":"neutral","pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_1":"neutral","pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_0":"neutral","pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_1":"neutral","pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0":"neutral","pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_1":"neutral","pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_0":"neutral","pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_1":"neutral","pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0":"neutral","pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_1":"neutral","pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_0":"neutral","pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_1":"neutral","pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0":"neutral","pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_1":"neutral","pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_0":"neutral","pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_1":"neutral","pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0":"neutral","pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_1":"neutral","pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_0":"neutral","pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_1":"neutral","pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0":"neutral","pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_1":"neutral","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0":"neutral","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1":"neutral","pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0":"neutral","pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1":"neutral","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0":"neutral","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1":"neutral","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0":"neutral","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1":"neutral","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0":"neutral","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1":"neutral","pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0":"neutral","pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1":"neutral","pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0":"neutral","pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1":"neutral","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0":"neutral","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1":"neutral","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0":"neutral","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_1":"neutral","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_0":"neutral","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1":"neutral","pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0":"neutral","pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_1":"neutral","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_0":"neutral","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1":"neutral","pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0":"neutral","pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_1":"neutral","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_0":"neutral","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1":"neutral","pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0":"neutral","pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_1":"neutral","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_0":"neutral","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1":"neutral","pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0":"neutral","pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_1":"neutral","pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_0":"neutral","pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1":"neutral","pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0":"neutral","pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_1":"neutral","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_0":"neutral","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1":"neutral","pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0":"neutral","pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_1":"neutral","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_0":"neutral","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1":"neutral","pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_0":"neutral","pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_1":"neutral","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_0":"neutral","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1":"neutral","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0":"neutral","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1":"neutral","pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_0":"neutral","pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_1":"neutral","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0":"neutral","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1":"neutral","pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_0":"neutral","pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_1":"neutral","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0":"neutral","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1":"neutral","pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_0":"neutral","pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_1":"neutral","pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0":"neutral","pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_1":"neutral","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0":"neutral","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_1":"neutral","pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_0":"neutral","pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_1":"neutral","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_0":"neutral","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_1":"neutral","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_0":"neutral","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_1":"neutral","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_0":"neutral","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_1":"neutral","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_0":"neutral","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_1":"neutral","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_0":"neutral","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_1":"neutral","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_0":"neutral","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_1":"neutral","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_0":"neutral","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_1":"neutral","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_0":"neutral","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_1":"neutral","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_0":"neutral","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_1":"neutral","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_0":"neutral","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_1":"neutral","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_0":"neutral","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_1":"neutral","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_0":"neutral","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1":"neutral","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_0":"neutral","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1":"neutral","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_0":"neutral","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_1":"neutral","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_0":"neutral","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_1":"neutral","pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0":"neutral","pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_0":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_1":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_2":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_3":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_4":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_5":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_6":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_7":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_8":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_9":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_10":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_11":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_12":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_13":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_14":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_15":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_16":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_17":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_18":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_19":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_20":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_21":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_22":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_23":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_24":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_25":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_26":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_27":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_28":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_29":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_30":"neutral","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_31":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_0":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_1":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_2":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_3":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_4":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_5":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_6":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_7":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_8":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_9":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_11":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_12":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_13":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_14":"neutral","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_15":"neutral","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_0":"neutral","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_1":"neutral","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_2":"neutral","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_3":"neutral","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_4":"neutral"},"next_color_idx":39,"wires_placed_in_order":[["pin-type-component_3faaa76b-f816-4c9f-8694-a0742ce9c0ad_4","pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_0"],["pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_0","pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_1"],["pin-type-component_f02b596c-ca03-491a-812a-3b2807a017f7_0","pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_2"],["pin-type-component_3faaa76b-f816-4c9f-8694-a0742ce9c0ad_3","pin-type-component_b4abe5c3-7b62-43ba-bf50-bd199eacd8c2_0"],["pin-type-component_f02b596c-ca03-491a-812a-3b2807a017f7_2","pin-type-component_0a6a9ae8-6690-4443-a873-564e66f0e654_0"],["pin-type-component_b4abe5c3-7b62-43ba-bf50-bd199eacd8c2_0","pin-type-component_0a6a9ae8-6690-4443-a873-564e66f0e654_2"],["pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_3","pin-type-component_f02b596c-ca03-491a-812a-3b2807a017f7_0"],["pin-type-component_b5689c0d-8629-43ce-b194-b79107695973_2","pin-type-component_eeae5c5f-f233-4302-8f22-1b93da80a79f_2"],["pin-type-component_b5689c0d-8629-43ce-b194-b79107695973_0","pin-type-component_eeae5c5f-f233-4302-8f22-1b93da80a79f_0"],["pin-type-component_3faaa76b-f816-4c9f-8694-a0742ce9c0ad_4","pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_1"],["pin-type-component_3faaa76b-f816-4c9f-8694-a0742ce9c0ad_4","pin-type-component_f02b596c-ca03-491a-812a-3b2807a017f7_0"],["pin-type-component_49daef8d-a90d-4340-b3ab-604980de60c8_0","pin-type-component_b5689c0d-8629-43ce-b194-b79107695973_2"],["pin-type-component_49daef8d-a90d-4340-b3ab-604980de60c8_0","pin-type-component_eeae5c5f-f233-4302-8f22-1b93da80a79f_2"],["pin-type-component_b5689c0d-8629-43ce-b194-b79107695973_0","pin-type-component_3e91a306-3718-4e98-bb6f-276d56c43eeb_0"],["pin-type-component_1fbed37a-0c4e-445a-8971-de508f74e50f_0","pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_0"],["pin-type-component_7f11caa5-aeda-4da1-b237-8ef8c0d2c752_0","pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_2"],["pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_0","pin-type-component_1fbed37a-0c4e-445a-8971-de508f74e50f_0"],["pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_2","pin-type-component_7f11caa5-aeda-4da1-b237-8ef8c0d2c752_0"],["pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_1","pin-type-component_8bbfc184-10a5-446c-98f6-e71beffecd3f_0"],["pin-type-component_c86c6707-62b1-454e-8905-5c025e70ffa2_0","pin-type-component_854d4d60-1858-4ccb-99b2-38a7ca382402_0"],["pin-type-component_c86c6707-62b1-454e-8905-5c025e70ffa2_2","pin-type-component_6798c1e2-77da-48bf-b876-2e22f65ef2a4_0"],["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_0","pin-type-component_7e9999e8-686e-4f02-b1e7-bee04a417b43_0"],["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2","pin-type-component_e03f3631-cb55-4d48-bf80-427e34299dc2_0"],["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_0","pin-type-component_4bfdc0b0-0087-4f19-b9da-fe77fe2030bb_0"],["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2","pin-type-component_ada6e844-1bae-4716-870a-c40960a3bb4b_0"],["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_0","pin-type-component_725c2e06-513a-456a-a054-9a1efd2410b5_0"],["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2","pin-type-component_c9571346-472b-4672-95d7-be31dc07bc93_0"],["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_0","pin-type-component_84e67de5-59f5-4375-8901-060561a64dc9_0"],["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2","pin-type-component_5836c999-695f-47a8-8e7c-f38290544271_0"],["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2","pin-type-component_34e49cee-f08a-4772-a6d4-df82dbc6905c_0"],["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_0","pin-type-component_a4a81ac1-f999-4c5f-bf1d-d39d1364ba7e_0"],["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2","pin-type-component_e4ccca5e-2f92-4742-9f88-17c0acf9d0e5_0"],["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_0","pin-type-component_84525e3e-ef29-4e0c-a293-959707966b26_0"],["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2","pin-type-component_45b045d9-de2e-4c1e-9f03-8f59566339f3_0"],["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_0","pin-type-component_ad7b12e6-293b-4cf0-b5fc-2ad4811766ad_0"],["pin-type-component_6131d2d5-4418-42b6-aa69-5becc7f7d213_2","pin-type-component_1266203a-634e-499d-8c59-c240f96559a6_0"],["pin-type-component_6131d2d5-4418-42b6-aa69-5becc7f7d213_0","pin-type-component_222e7ad6-20c2-4c60-bcc8-d81940d5a2c1_0"],["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2","pin-type-component_1321abdf-76d2-4961-8eed-5e802ce03515_0"],["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_0","pin-type-component_69b6c16b-f2c6-4ab0-b694-b43efd7d7efa_0"],["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2","pin-type-component_80364b7e-c592-40e4-9f27-3a46aba92f9c_0"],["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_0","pin-type-component_5278fc75-d95d-4e4c-a86e-2e83a862e607_0"],["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1","pin-type-component_a3ab8da7-d370-48c7-aed7-0afc87949c1f_0"],["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_0","pin-type-component_0af45fa8-24bc-42e4-9c24-d15187e9fbc3_0"],["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2","pin-type-component_a723fcb8-a29a-44f7-91e6-b934c414e1d5_0"],["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_0","pin-type-component_266aa6bb-5bae-4ff3-85db-bbd370178ae8_0"],["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2","pin-type-component_9fb789aa-23a4-4c02-856a-7e2a62a5687c_0"],["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_0","pin-type-component_7fc8671b-e701-4c33-a644-f42eace24307_0"],["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2","pin-type-component_02c2443e-51cb-49a5-b48e-828fe43ba847_0"],["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_0","pin-type-component_34445add-d974-48d4-81af-972f5dd7934b_0"],["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2","pin-type-component_20c4afac-aed7-47a4-b18b-1cd7a3325c34_0"],["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_0","pin-type-component_3d109b51-1504-4d24-a9e7-9e3fe3074724_0"],["pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2","pin-type-component_78dc7030-f822-4db6-b90c-1a871bd2febd_0"],["pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_0","pin-type-component_e7d36833-6d1a-490c-96e9-4f178d942f47_0"],["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2","pin-type-component_d23f20e3-e8e7-4a94-b362-814ae84c95f1_0"],["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_0","pin-type-component_903934ae-30da-4a37-93c9-c64660e9c617_0"],["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2","pin-type-component_7dc8ce5e-7fe0-4560-a90a-24f57026c2ce_0"],["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_0","pin-type-component_7f294ee1-7ea8-4e70-bb0a-8c8b6b15b6c9_0"],["pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_0","pin-type-component_4732636d-ea0d-4b19-877e-d2ff4ddb5e8d_0"],["pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2","pin-type-component_f4cc5271-6fed-4fbe-b520-d7f27ca6d761_0"],["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2","pin-type-component_756a3f47-cc5c-4c12-8a88-5902936d2980_0"],["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_0","pin-type-component_62a268f0-68fa-4016-91c7-d55a738d6b46_0"],["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2","pin-type-component_5cc5144a-e27c-4a8c-a3b8-dfdff02281da_0"],["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_0","pin-type-component_5bdd54e6-172a-4994-8b34-5d8687be61e2_0"],["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2","pin-type-component_cb28eb0e-db83-4b4e-b021-b939f7a83c54_0"],["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_0","pin-type-component_29f2dcbd-c66e-4d22-9415-91c6505cd16b_0"],["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2","pin-type-component_4e5aed25-a709-4dca-a8d1-34d4dd3bbcf9_0"],["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_0","pin-type-component_d1e6942e-6a34-4356-87fa-da19b68ae6b8_0"],["pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2","pin-type-component_6544f2c2-1808-475f-8a33-efd3517c4989_0"],["pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_0","pin-type-component_0c082f01-0561-48cc-887e-4e37deace687_0"],["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2","pin-type-component_565c607a-48b0-4de4-800e-47cbf9473dce_0"],["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_0","pin-type-component_6d57b374-4a97-4f2c-b0da-4d4ccbef4f5a_0"],["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2","pin-type-component_c5d490e1-2b79-451a-b5af-757c0e65aa93_0"],["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_0","pin-type-component_dd44450f-fd4f-4059-aab9-565428093e7b_0"],["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2","pin-type-component_e808b193-47e2-4e3e-801b-fce476c62302_0"],["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_0","pin-type-component_e84ff89e-b801-43e3-905a-a7004860c743_0"],["pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2","pin-type-component_26138f80-3acc-4ecb-b94a-9f0d8ab839a6_0"],["pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_0","pin-type-component_636bd670-72c8-425e-8740-11540fc72a9f_0"],["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2","pin-type-component_7419eacb-81ea-40c7-af9f-438e4f0521b0_0"],["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_0","pin-type-component_bb4a8fb4-80b5-4764-a9f6-b3d9cae671c4_0"],["pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2","pin-type-component_a1044649-e843-43ff-95e7-a21a072714be_0"],["pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_0","pin-type-component_edb09e16-b982-4564-8c59-d0c31b14f784_0"],["pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2","pin-type-component_515f6f7f-721f-439a-b2db-7f6c6ca7ad1f_0"],["pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_0","pin-type-component_0b4ba5d8-bcb4-4816-8dfe-3fa4ce9ed019_0"],["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2","pin-type-component_1b0f4904-14bf-429f-937d-c99b5c2da67c_0"],["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_0","pin-type-component_b2f3a979-ce1b-444a-a7e4-6ef67b25f077_0"],["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2","pin-type-component_fc486c6a-efa6-4e32-a1f3-0451662788c4_0"],["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_0","pin-type-component_3b6d34de-cd89-4ef4-9473-da4b3ae907df_0"],["pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_1","pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_1"],["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1"],["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1"],["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1"],["pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0","pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0"],["pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0"],["pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15"],["pin-type-component_a1044649-e843-43ff-95e7-a21a072714be_0","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15"],["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1"],["pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_1","pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_1"],["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1"],["pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_0"],["pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14"],["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_1","pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_1"],["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_1","pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_1"],["pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_0","pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0"],["pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13"],["pin-type-component_7419eacb-81ea-40c7-af9f-438e4f0521b0_0","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14"],["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_1","pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_1"],["pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_1","pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_1"],["pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_0","pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0"],["pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12"],["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_1","pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_1"],["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_1","pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_1"],["pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0","pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_0"],["pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_1","pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_1"],["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_1","pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_1"],["pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_0","pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0"],["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_1","pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_1"],["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_1","pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_1"],["pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0","pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_0"],["pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_1","pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_1"],["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_1","pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_1"],["pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_0","pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0"],["pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11"],["pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10"],["pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9"],["pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8"],["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_1","pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_1"],["pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_1","pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_1"],["pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_0","pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0"],["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_1","pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_1"],["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_1","pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_1"],["pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0","pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_0"],["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_1","pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_1"],["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_1","pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_1"],["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2","pin-type-component_a3ab8da7-d370-48c7-aed7-0afc87949c1f_0"],["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1","pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_1"],["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_1","pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_1"],["pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0","pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_0"],["pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0","pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_0"],["pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7"],["pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6"],["pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5"],["pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4"],["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_1","pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_1"],["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_1","pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_1"],["pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_0","pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0"],["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_1","pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_1"],["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_1","pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_1"],["pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_0","pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0"],["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_1","pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_1"],["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_1","pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_1"],["pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_0","pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0"],["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_1","pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_1"],["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_1","pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_1"],["pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_0","pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0"],["pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3"],["pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2"],["pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1"],["pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0"],["pin-type-component_77f3714c-986d-44d0-96fc-d08c3926bdf3_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"],["pin-type-component_77f3714c-986d-44d0-96fc-d08c3926bdf3_1","pin-type-component_6c05b0a4-5167-4fc7-aa40-154354a323db_0"],["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2"],["pin-type-component_6c05b0a4-5167-4fc7-aa40-154354a323db_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"],["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1","pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0"],["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2"],["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15"],["pin-type-component_2026dadb-8316-442a-8bdd-67cd7b7c35b5_0","pin-type-component_6af167c7-0fd0-4ca2-b611-5ff73a7d20c6_0"],["pin-type-component_6af167c7-0fd0-4ca2-b611-5ff73a7d20c6_1","pin-type-component_65174c61-423b-440d-87cd-92d054e20fb1_0"],["pin-type-component_65174c61-423b-440d-87cd-92d054e20fb1_1","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2"],["pin-type-component_65174c61-423b-440d-87cd-92d054e20fb1_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14"],["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1","pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2"],["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1"],["pin-type-component_4c09ece5-1761-45a0-a275-3834e713bd96_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0"],["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13"],["pin-type-component_643580bd-b866-47c4-b5fe-63ae91e7cd50_1","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2"],["pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_1","pin-type-component_643580bd-b866-47c4-b5fe-63ae91e7cd50_0"],["pin-type-component_4c09ece5-1761-45a0-a275-3834e713bd96_0","pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_0"],["pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0"],["pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0","pin-type-component_2026dadb-8316-442a-8bdd-67cd7b7c35b5_0"],["pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_0","pin-type-component_6af167c7-0fd0-4ca2-b611-5ff73a7d20c6_0"],["pin-type-component_6af167c7-0fd0-4ca2-b611-5ff73a7d20c6_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"],["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1","pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2"],["pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0"],["pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1","pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0"],["pin-type-component_566c9339-cfa0-4791-a41c-f6f6cc110bfa_1","pin-type-component_fcd5d325-6008-4d5c-8522-dfa7deaae9d5_0"],["pin-type-component_fcd5d325-6008-4d5c-8522-dfa7deaae9d5_1","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2"],["pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0","pin-type-component_566c9339-cfa0-4791-a41c-f6f6cc110bfa_0"],["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1","pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2"],["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0"],["pin-type-component_566c9339-cfa0-4791-a41c-f6f6cc110bfa_0","pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0"],["pin-type-component_08fc44c3-171b-463f-a521-c64edfef133b_1","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2"],["pin-type-component_08fc44c3-171b-463f-a521-c64edfef133b_0","pin-type-component_796f060b-5c39-4bf7-8a4c-fd057b19eb84_1"],["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_796f060b-5c39-4bf7-8a4c-fd057b19eb84_0"],["pin-type-component_643580bd-b866-47c4-b5fe-63ae91e7cd50_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12"],["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11"],["pin-type-component_fcd5d325-6008-4d5c-8522-dfa7deaae9d5_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10"],["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"],["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0"],["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2"],["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2"],["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1"],["pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0"],["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2"],["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2"],["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2"],["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0"],["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2"],["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1"],["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0"],["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14"],["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13"],["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12"],["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2","pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2"],["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2","pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2"],["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2","pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2"],["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2","pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2"],["pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_1","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_0"],["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1"],["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0","pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0"],["pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_1","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_0"],["pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0","pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0"],["pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0","pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0"],["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1"],["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1"],["pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0"],["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1"],["pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11"],["pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10"],["pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9"],["pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8"],["pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_1","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_0"],["pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_1","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_0"],["pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_1","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_0"],["pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_1","pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_0"],["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0"],["pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0","pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0"],["pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0","pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0"],["pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0","pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_0"],["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2","pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2"],["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2","pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2"],["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2"],["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2","pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2"],["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2","pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1"],["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1"],["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1"],["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1"],["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15"],["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14"],["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13"],["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12"],["pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_1","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_0"],["pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_1","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_0"],["pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11"],["pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10"],["pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9"],["pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8"],["pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_7"],["pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_6"],["pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_5"],["pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_4"],["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2"],["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2","pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2"],["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2","pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2"],["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2","pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2"],["pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1","pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_0"],["pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1","pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_0"],["pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1","pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_0"],["pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_1","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0"],["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0"],["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0"],["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0"],["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2","pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0"],["pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_0"],["pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_1"],["pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_2"],["pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_3"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_1"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0","pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_1"],["pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_0","pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_0"],["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_18"],["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16","pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0"],["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_18"],["pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_6"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_19","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_27"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_20","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_26"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_21","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_25"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_22","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_24"],["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_23","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_23"],["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_19","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_8"],["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_20","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_9"],["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_21","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_10"],["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_22","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_11"],["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_23","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_12"],["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_3"],["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_9","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_5"],["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_11","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_22"],["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_12","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_29"],["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_1","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_21"],["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_2","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_20"],["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_3","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_19"],["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_4","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_18"],["pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_4","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_7"],["pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_3","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_17"],["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"],["pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0"],["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1"],["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1"],["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1"],["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0"],["pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0"],["pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0"],["pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0"],["pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0"],["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0"],["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0"],["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_3faaa76b-f816-4c9f-8694-a0742ce9c0ad_4","pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_0"]]],[[],[["pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_0","pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_1"]]],[[],[["pin-type-component_f02b596c-ca03-491a-812a-3b2807a017f7_0","pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_2"]]],[[],[["pin-type-component_3faaa76b-f816-4c9f-8694-a0742ce9c0ad_3","pin-type-component_b4abe5c3-7b62-43ba-bf50-bd199eacd8c2_0"]]],[[],[["pin-type-component_f02b596c-ca03-491a-812a-3b2807a017f7_2","pin-type-component_0a6a9ae8-6690-4443-a873-564e66f0e654_0"]]],[[],[["pin-type-component_b4abe5c3-7b62-43ba-bf50-bd199eacd8c2_0","pin-type-component_0a6a9ae8-6690-4443-a873-564e66f0e654_2"]]],[[["pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_2","pin-type-component_f02b596c-ca03-491a-812a-3b2807a017f7_0"]],[]],[[],[["pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_3","pin-type-component_f02b596c-ca03-491a-812a-3b2807a017f7_0"]]],[[],[["pin-type-component_b5689c0d-8629-43ce-b194-b79107695973_2","pin-type-component_eeae5c5f-f233-4302-8f22-1b93da80a79f_2"]]],[[],[["pin-type-component_b5689c0d-8629-43ce-b194-b79107695973_0","pin-type-component_eeae5c5f-f233-4302-8f22-1b93da80a79f_0"]]],[[["pin-type-component_b5689c0d-8629-43ce-b194-b79107695973_0","pin-type-component_eeae5c5f-f233-4302-8f22-1b93da80a79f_0"]],[]],[[["pin-type-component_b5689c0d-8629-43ce-b194-b79107695973_2","pin-type-component_eeae5c5f-f233-4302-8f22-1b93da80a79f_2"]],[]],[[["pin-type-component_3faaa76b-f816-4c9f-8694-a0742ce9c0ad_4","pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_0"],["pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_0","pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_1"]],[["pin-type-component_3faaa76b-f816-4c9f-8694-a0742ce9c0ad_4","pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_1"]]],[[["pin-type-component_3faaa76b-f816-4c9f-8694-a0742ce9c0ad_4","pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_1"]],[]],[[["pin-type-component_d675a4a5-df4a-424c-b7ff-fd583a688e45_3","pin-type-component_f02b596c-ca03-491a-812a-3b2807a017f7_0"]],[]],[[],[["pin-type-component_3faaa76b-f816-4c9f-8694-a0742ce9c0ad_4","pin-type-component_f02b596c-ca03-491a-812a-3b2807a017f7_0"]]],[[["pin-type-component_0a6a9ae8-6690-4443-a873-564e66f0e654_0","pin-type-component_f02b596c-ca03-491a-812a-3b2807a017f7_2"]],[]],[[["pin-type-component_0a6a9ae8-6690-4443-a873-564e66f0e654_2","pin-type-component_b4abe5c3-7b62-43ba-bf50-bd199eacd8c2_0"]],[]],[[["pin-type-component_3faaa76b-f816-4c9f-8694-a0742ce9c0ad_4","pin-type-component_f02b596c-ca03-491a-812a-3b2807a017f7_0"]],[]],[[["pin-type-component_3faaa76b-f816-4c9f-8694-a0742ce9c0ad_3","pin-type-component_b4abe5c3-7b62-43ba-bf50-bd199eacd8c2_0"]],[]],[[],[["pin-type-component_49daef8d-a90d-4340-b3ab-604980de60c8_0","pin-type-component_b5689c0d-8629-43ce-b194-b79107695973_2"]]],[[],[["pin-type-component_49daef8d-a90d-4340-b3ab-604980de60c8_0","pin-type-component_eeae5c5f-f233-4302-8f22-1b93da80a79f_2"]]],[[["pin-type-component_49daef8d-a90d-4340-b3ab-604980de60c8_0","pin-type-component_eeae5c5f-f233-4302-8f22-1b93da80a79f_2"]],[]],[[],[["pin-type-component_b5689c0d-8629-43ce-b194-b79107695973_0","pin-type-component_3e91a306-3718-4e98-bb6f-276d56c43eeb_0"]]],[[],[["pin-type-component_1fbed37a-0c4e-445a-8971-de508f74e50f_0","pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_0"]]],[[],[["pin-type-component_7f11caa5-aeda-4da1-b237-8ef8c0d2c752_0","pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_2"]]],[[["pin-type-component_1fbed37a-0c4e-445a-8971-de508f74e50f_0","pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_0"]],[]],[[],[["pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_0","pin-type-component_1fbed37a-0c4e-445a-8971-de508f74e50f_0"]]],[[["pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_2","pin-type-component_7f11caa5-aeda-4da1-b237-8ef8c0d2c752_0"]],[]],[[],[["pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_2","pin-type-component_7f11caa5-aeda-4da1-b237-8ef8c0d2c752_0"]]],[[],[["pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_1","pin-type-component_8bbfc184-10a5-446c-98f6-e71beffecd3f_0"]]],[[["pin-type-component_3e91a306-3718-4e98-bb6f-276d56c43eeb_0","pin-type-component_b5689c0d-8629-43ce-b194-b79107695973_0"]],[]],[[["pin-type-component_49daef8d-a90d-4340-b3ab-604980de60c8_0","pin-type-component_b5689c0d-8629-43ce-b194-b79107695973_2"]],[]],[[["pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_1","pin-type-component_8bbfc184-10a5-446c-98f6-e71beffecd3f_0"]],[]],[[],[["pin-type-component_c86c6707-62b1-454e-8905-5c025e70ffa2_0","pin-type-component_854d4d60-1858-4ccb-99b2-38a7ca382402_0"]]],[[],[["pin-type-component_c86c6707-62b1-454e-8905-5c025e70ffa2_2","pin-type-component_6798c1e2-77da-48bf-b876-2e22f65ef2a4_0"]]],[[],[["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_0","pin-type-component_7e9999e8-686e-4f02-b1e7-bee04a417b43_0"]]],[[],[["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2","pin-type-component_e03f3631-cb55-4d48-bf80-427e34299dc2_0"]]],[[],[["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_0","pin-type-component_4bfdc0b0-0087-4f19-b9da-fe77fe2030bb_0"]]],[[],[["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2","pin-type-component_ada6e844-1bae-4716-870a-c40960a3bb4b_0"]]],[[],[["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_0","pin-type-component_725c2e06-513a-456a-a054-9a1efd2410b5_0"]]],[[],[["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2","pin-type-component_c9571346-472b-4672-95d7-be31dc07bc93_0"]]],[[],[["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_0","pin-type-component_84e67de5-59f5-4375-8901-060561a64dc9_0"]]],[[],[["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2","pin-type-component_5836c999-695f-47a8-8e7c-f38290544271_0"]]],[[["pin-type-component_6798c1e2-77da-48bf-b876-2e22f65ef2a4_0","pin-type-component_c86c6707-62b1-454e-8905-5c025e70ffa2_2"]],[]],[[["pin-type-component_854d4d60-1858-4ccb-99b2-38a7ca382402_0","pin-type-component_c86c6707-62b1-454e-8905-5c025e70ffa2_0"]],[]],[[["pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_2","pin-type-component_7f11caa5-aeda-4da1-b237-8ef8c0d2c752_0"]],[]],[[["pin-type-component_1fbed37a-0c4e-445a-8971-de508f74e50f_0","pin-type-component_43916a4e-c7c4-43ca-b750-0c6b91dabb72_0"]],[]],[[],[["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2","pin-type-component_34e49cee-f08a-4772-a6d4-df82dbc6905c_0"]]],[[],[["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_0","pin-type-component_a4a81ac1-f999-4c5f-bf1d-d39d1364ba7e_0"]]],[[],[["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2","pin-type-component_e4ccca5e-2f92-4742-9f88-17c0acf9d0e5_0"]]],[[],[["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_0","pin-type-component_84525e3e-ef29-4e0c-a293-959707966b26_0"]]],[[],[["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2","pin-type-component_45b045d9-de2e-4c1e-9f03-8f59566339f3_0"]]],[[],[["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_0","pin-type-component_ad7b12e6-293b-4cf0-b5fc-2ad4811766ad_0"]]],[[],[["pin-type-component_6131d2d5-4418-42b6-aa69-5becc7f7d213_2","pin-type-component_1266203a-634e-499d-8c59-c240f96559a6_0"]]],[[],[["pin-type-component_6131d2d5-4418-42b6-aa69-5becc7f7d213_0","pin-type-component_222e7ad6-20c2-4c60-bcc8-d81940d5a2c1_0"]]],[[["pin-type-component_1266203a-634e-499d-8c59-c240f96559a6_0","pin-type-component_6131d2d5-4418-42b6-aa69-5becc7f7d213_2"]],[]],[[["pin-type-component_222e7ad6-20c2-4c60-bcc8-d81940d5a2c1_0","pin-type-component_6131d2d5-4418-42b6-aa69-5becc7f7d213_0"]],[]],[[],[["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2","pin-type-component_1321abdf-76d2-4961-8eed-5e802ce03515_0"]]],[[],[["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_0","pin-type-component_69b6c16b-f2c6-4ab0-b694-b43efd7d7efa_0"]]],[[],[["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2","pin-type-component_80364b7e-c592-40e4-9f27-3a46aba92f9c_0"]]],[[],[["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_0","pin-type-component_5278fc75-d95d-4e4c-a86e-2e83a862e607_0"]]],[[],[["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1","pin-type-component_a3ab8da7-d370-48c7-aed7-0afc87949c1f_0"]]],[[],[["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_0","pin-type-component_0af45fa8-24bc-42e4-9c24-d15187e9fbc3_0"]]],[[],[["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2","pin-type-component_a723fcb8-a29a-44f7-91e6-b934c414e1d5_0"]]],[[],[["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_0","pin-type-component_266aa6bb-5bae-4ff3-85db-bbd370178ae8_0"]]],[[],[["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2","pin-type-component_9fb789aa-23a4-4c02-856a-7e2a62a5687c_0"]]],[[],[["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_0","pin-type-component_7fc8671b-e701-4c33-a644-f42eace24307_0"]]],[[],[["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2","pin-type-component_02c2443e-51cb-49a5-b48e-828fe43ba847_0"]]],[[],[["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_0","pin-type-component_34445add-d974-48d4-81af-972f5dd7934b_0"]]],[[],[["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2","pin-type-component_20c4afac-aed7-47a4-b18b-1cd7a3325c34_0"]]],[[],[["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_0","pin-type-component_3d109b51-1504-4d24-a9e7-9e3fe3074724_0"]]],[[],[["pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2","pin-type-component_78dc7030-f822-4db6-b90c-1a871bd2febd_0"]]],[[],[["pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_0","pin-type-component_e7d36833-6d1a-490c-96e9-4f178d942f47_0"]]],[[],[["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2","pin-type-component_d23f20e3-e8e7-4a94-b362-814ae84c95f1_0"]]],[[],[["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_0","pin-type-component_903934ae-30da-4a37-93c9-c64660e9c617_0"]]],[[],[["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2","pin-type-component_7dc8ce5e-7fe0-4560-a90a-24f57026c2ce_0"]]],[[],[["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_0","pin-type-component_7f294ee1-7ea8-4e70-bb0a-8c8b6b15b6c9_0"]]],[[],[["pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_0","pin-type-component_4732636d-ea0d-4b19-877e-d2ff4ddb5e8d_0"]]],[[],[["pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2","pin-type-component_f4cc5271-6fed-4fbe-b520-d7f27ca6d761_0"]]],[[],[["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2","pin-type-component_756a3f47-cc5c-4c12-8a88-5902936d2980_0"]]],[[],[["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_0","pin-type-component_62a268f0-68fa-4016-91c7-d55a738d6b46_0"]]],[[],[["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2","pin-type-component_5cc5144a-e27c-4a8c-a3b8-dfdff02281da_0"]]],[[],[["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_0","pin-type-component_5bdd54e6-172a-4994-8b34-5d8687be61e2_0"]]],[[],[["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2","pin-type-component_cb28eb0e-db83-4b4e-b021-b939f7a83c54_0"]]],[[],[["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_0","pin-type-component_29f2dcbd-c66e-4d22-9415-91c6505cd16b_0"]]],[[],[["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2","pin-type-component_4e5aed25-a709-4dca-a8d1-34d4dd3bbcf9_0"]]],[[],[["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_0","pin-type-component_d1e6942e-6a34-4356-87fa-da19b68ae6b8_0"]]],[[],[["pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2","pin-type-component_6544f2c2-1808-475f-8a33-efd3517c4989_0"]]],[[],[["pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_0","pin-type-component_0c082f01-0561-48cc-887e-4e37deace687_0"]]],[[],[["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2","pin-type-component_565c607a-48b0-4de4-800e-47cbf9473dce_0"]]],[[],[["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_0","pin-type-component_6d57b374-4a97-4f2c-b0da-4d4ccbef4f5a_0"]]],[[],[]],[[],[["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2","pin-type-component_c5d490e1-2b79-451a-b5af-757c0e65aa93_0"]]],[[],[["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_0","pin-type-component_dd44450f-fd4f-4059-aab9-565428093e7b_0"]]],[[],[["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2","pin-type-component_e808b193-47e2-4e3e-801b-fce476c62302_0"]]],[[],[["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_0","pin-type-component_e84ff89e-b801-43e3-905a-a7004860c743_0"]]],[[],[["pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2","pin-type-component_26138f80-3acc-4ecb-b94a-9f0d8ab839a6_0"]]],[[],[["pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_0","pin-type-component_636bd670-72c8-425e-8740-11540fc72a9f_0"]]],[[],[["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2","pin-type-component_7419eacb-81ea-40c7-af9f-438e4f0521b0_0"]]],[[],[["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_0","pin-type-component_bb4a8fb4-80b5-4764-a9f6-b3d9cae671c4_0"]]],[[],[["pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2","pin-type-component_a1044649-e843-43ff-95e7-a21a072714be_0"]]],[[],[["pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_0","pin-type-component_edb09e16-b982-4564-8c59-d0c31b14f784_0"]]],[[],[["pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2","pin-type-component_515f6f7f-721f-439a-b2db-7f6c6ca7ad1f_0"]]],[[],[["pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_0","pin-type-component_0b4ba5d8-bcb4-4816-8dfe-3fa4ce9ed019_0"]]],[[],[["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2","pin-type-component_1b0f4904-14bf-429f-937d-c99b5c2da67c_0"]]],[[],[["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_0","pin-type-component_b2f3a979-ce1b-444a-a7e4-6ef67b25f077_0"]]],[[],[["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2","pin-type-component_fc486c6a-efa6-4e32-a1f3-0451662788c4_0"]]],[[],[["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_0","pin-type-component_3b6d34de-cd89-4ef4-9473-da4b3ae907df_0"]]],[[],[["pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_1","pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_1"]]],[[],[["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1"]]],[[["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1"]],[]],[[],[["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1"]]],[[["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1"]],[]],[[],[["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1"]]],[[],[["pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0","pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0"]]],[[["pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0"]],[]],[[],[["pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0"]]],[[],[["pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15"]]],[[],[["pin-type-component_a1044649-e843-43ff-95e7-a21a072714be_0","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15"]]],[[],[["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1"]]],[[],[["pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_1","pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_1"]]],[[["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1"]],[]],[[],[["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1"]]],[[],[["pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_0"]]],[[],[["pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14"]]],[[],[["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_1","pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_1"]]],[[],[["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_1","pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_1"]]],[[],[["pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_0","pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0"]]],[[],[["pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13"]]],[[],[["pin-type-component_7419eacb-81ea-40c7-af9f-438e4f0521b0_0","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14"]]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14","pin-type-component_7419eacb-81ea-40c7-af9f-438e4f0521b0_0"]],[]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15","pin-type-component_a1044649-e843-43ff-95e7-a21a072714be_0"]],[]],[[],[["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_1","pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_1"]]],[[],[["pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_1","pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_1"]]],[[],[["pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_0","pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0"]]],[[],[["pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12"]]],[[],[["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_1","pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_1"]]],[[],[["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_1","pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_1"]]],[[],[["pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0","pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_0"]]],[[],[["pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_1","pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_1"]]],[[],[["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_1","pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_1"]]],[[],[["pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_0","pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0"]]],[[],[["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_1","pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_1"]]],[[],[["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_1","pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_1"]]],[[],[["pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0","pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_0"]]],[[],[["pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_1","pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_1"]]],[[],[["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_1","pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_1"]]],[[],[["pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_0","pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0"]]],[[],[["pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11"]]],[[],[["pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10"]]],[[],[["pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9"]]],[[],[["pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8"]]],[[],[["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_1","pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_1"]]],[[],[["pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_1","pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_1"]]],[[],[["pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_0","pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0"]]],[[],[["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_1","pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_1"]]],[[],[["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_1","pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_1"]]],[[],[["pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0","pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_0"]]],[[],[["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_1","pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_1"]]],[[],[["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_1","pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_1"]]],[[["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1","pin-type-component_a3ab8da7-d370-48c7-aed7-0afc87949c1f_0"]],[]],[[],[["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2","pin-type-component_a3ab8da7-d370-48c7-aed7-0afc87949c1f_0"]]],[[],[["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1","pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_1"]]],[[],[["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_1","pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_1"]]],[[],[["pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0","pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_0"]]],[[],[["pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0","pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_0"]]],[[],[["pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7"]]],[[],[["pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6"]]],[[],[["pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5"]]],[[],[["pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4"]]],[[],[["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_1","pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_1"]]],[[],[["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_1","pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_1"]]],[[],[["pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_0","pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0"]]],[[],[["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_1","pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_1"]]],[[],[["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_1","pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_1"]]],[[],[["pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_0","pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0"]]],[[],[["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_1","pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_1"]]],[[],[["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_1","pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_1"]]],[[],[["pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_0","pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0"]]],[[],[["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_1","pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_1"]]],[[],[["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_1","pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_1"]]],[[],[["pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_0","pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0"]]],[[],[["pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3"]]],[[],[["pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2"]]],[[],[["pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1"]]],[[],[["pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0"]]],[[["pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2","pin-type-component_a1044649-e843-43ff-95e7-a21a072714be_0"]],[]],[[["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2","pin-type-component_7419eacb-81ea-40c7-af9f-438e4f0521b0_0"]],[]],[[["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2","pin-type-component_e808b193-47e2-4e3e-801b-fce476c62302_0"]],[]],[[["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2","pin-type-component_c5d490e1-2b79-451a-b5af-757c0e65aa93_0"]],[]],[[["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2","pin-type-component_565c607a-48b0-4de4-800e-47cbf9473dce_0"]],[]],[[["pin-type-component_6544f2c2-1808-475f-8a33-efd3517c4989_0","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2"]],[]],[[["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2","pin-type-component_4e5aed25-a709-4dca-a8d1-34d4dd3bbcf9_0"]],[]],[[],[["pin-type-component_77f3714c-986d-44d0-96fc-d08c3926bdf3_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"]]],[[],[["pin-type-component_77f3714c-986d-44d0-96fc-d08c3926bdf3_1","pin-type-component_6c05b0a4-5167-4fc7-aa40-154354a323db_0"]]],[[],[["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2"]]],[[["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0","pin-type-component_77f3714c-986d-44d0-96fc-d08c3926bdf3_0"]],[]],[[["pin-type-component_6c05b0a4-5167-4fc7-aa40-154354a323db_0","pin-type-component_77f3714c-986d-44d0-96fc-d08c3926bdf3_1"]],[]],[[["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1"]],[]],[[],[["pin-type-component_6c05b0a4-5167-4fc7-aa40-154354a323db_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"]]],[[],[["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1","pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0"]]],[[],[["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2"]]],[[],[["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15"]]],[[],[["pin-type-component_2026dadb-8316-442a-8bdd-67cd7b7c35b5_0","pin-type-component_6af167c7-0fd0-4ca2-b611-5ff73a7d20c6_0"]]],[[],[["pin-type-component_6af167c7-0fd0-4ca2-b611-5ff73a7d20c6_1","pin-type-component_65174c61-423b-440d-87cd-92d054e20fb1_0"]]],[[],[["pin-type-component_65174c61-423b-440d-87cd-92d054e20fb1_1","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2"]]],[[],[["pin-type-component_65174c61-423b-440d-87cd-92d054e20fb1_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14"]]],[[],[["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1","pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2"]]],[[],[["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1"]]],[[],[["pin-type-component_4c09ece5-1761-45a0-a275-3834e713bd96_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0"]]],[[],[["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13"]]],[[],[["pin-type-component_643580bd-b866-47c4-b5fe-63ae91e7cd50_1","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2"]]],[[],[["pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_1","pin-type-component_643580bd-b866-47c4-b5fe-63ae91e7cd50_0"]]],[[],[["pin-type-component_4c09ece5-1761-45a0-a275-3834e713bd96_0","pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_0"]]],[[["pin-type-component_4c09ece5-1761-45a0-a275-3834e713bd96_0","pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_0"],["pin-type-component_4c09ece5-1761-45a0-a275-3834e713bd96_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0"]],[["pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0"]]],[[],[["pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0","pin-type-component_2026dadb-8316-442a-8bdd-67cd7b7c35b5_0"]]],[[["pin-type-component_2026dadb-8316-442a-8bdd-67cd7b7c35b5_0","pin-type-component_6af167c7-0fd0-4ca2-b611-5ff73a7d20c6_0"],["pin-type-component_2026dadb-8316-442a-8bdd-67cd7b7c35b5_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0"]],[["pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_0","pin-type-component_6af167c7-0fd0-4ca2-b611-5ff73a7d20c6_0"]]],[[],[["pin-type-component_6af167c7-0fd0-4ca2-b611-5ff73a7d20c6_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"]]],[[],[["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1","pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2"]]],[[],[["pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0"]]],[[],[["pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1","pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0"]]],[[["pin-type-component_26138f80-3acc-4ecb-b94a-9f0d8ab839a6_0","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2"]],[]],[[],[["pin-type-component_566c9339-cfa0-4791-a41c-f6f6cc110bfa_1","pin-type-component_fcd5d325-6008-4d5c-8522-dfa7deaae9d5_0"]]],[[],[["pin-type-component_fcd5d325-6008-4d5c-8522-dfa7deaae9d5_1","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2"]]],[[],[["pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0","pin-type-component_566c9339-cfa0-4791-a41c-f6f6cc110bfa_0"]]],[[],[["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1","pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2"]]],[[],[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0"]]],[[],[["pin-type-component_566c9339-cfa0-4791-a41c-f6f6cc110bfa_0","pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0"]]],[[],[["pin-type-component_08fc44c3-171b-463f-a521-c64edfef133b_1","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2"]]],[[],[["pin-type-component_08fc44c3-171b-463f-a521-c64edfef133b_0","pin-type-component_796f060b-5c39-4bf7-8a4c-fd057b19eb84_1"]]],[[],[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_796f060b-5c39-4bf7-8a4c-fd057b19eb84_0"]]],[[],[["pin-type-component_643580bd-b866-47c4-b5fe-63ae91e7cd50_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12"]]],[[],[["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11"]]],[[],[["pin-type-component_fcd5d325-6008-4d5c-8522-dfa7deaae9d5_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10"]]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14","pin-type-component_65174c61-423b-440d-87cd-92d054e20fb1_1"]],[]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12","pin-type-component_643580bd-b866-47c4-b5fe-63ae91e7cd50_1"]],[]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1"]],[]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11","pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1"]],[]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10","pin-type-component_fcd5d325-6008-4d5c-8522-dfa7deaae9d5_1"]],[]],[[["pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_0","pin-type-component_6af167c7-0fd0-4ca2-b611-5ff73a7d20c6_0"],["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0","pin-type-component_6af167c7-0fd0-4ca2-b611-5ff73a7d20c6_0"]],[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"]]],[[["pin-type-component_65174c61-423b-440d-87cd-92d054e20fb1_0","pin-type-component_6af167c7-0fd0-4ca2-b611-5ff73a7d20c6_1"]],[]],[[["pin-type-component_65174c61-423b-440d-87cd-92d054e20fb1_1","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2"]],[]],[[["pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_1","pin-type-component_643580bd-b866-47c4-b5fe-63ae91e7cd50_0"]],[]],[[["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2","pin-type-component_643580bd-b866-47c4-b5fe-63ae91e7cd50_1"]],[]],[[["pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0"],["pin-type-component_5fe70d92-e0f3-4ab0-90e2-f9cd6e3e1a0d_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0"]],[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0"]]],[[],[["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2"]]],[[],[["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2"]]],[[["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1","pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0"]],[]],[[],[["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1"]]],[[],[]],[[["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1"]],[]],[[["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0"]],[]],[[],[["pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0"]]],[[["pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2","pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0"]],[]],[[],[["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2"]]],[[],[["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2"]]],[[["pin-type-component_566c9339-cfa0-4791-a41c-f6f6cc110bfa_1","pin-type-component_fcd5d325-6008-4d5c-8522-dfa7deaae9d5_0"]],[]],[[["pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2","pin-type-component_fcd5d325-6008-4d5c-8522-dfa7deaae9d5_1"]],[]],[[],[["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2"]]],[[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_566c9339-cfa0-4791-a41c-f6f6cc110bfa_0"],["pin-type-component_566c9339-cfa0-4791-a41c-f6f6cc110bfa_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0"]],[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0"]]],[[["pin-type-component_08fc44c3-171b-463f-a521-c64edfef133b_0","pin-type-component_796f060b-5c39-4bf7-8a4c-fd057b19eb84_1"]],[]],[[["pin-type-component_08fc44c3-171b-463f-a521-c64edfef133b_1","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2"]],[]],[[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_796f060b-5c39-4bf7-8a4c-fd057b19eb84_0"]],[]],[[],[["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2"]]],[[["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1"]],[]],[[],[["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1"]]],[[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0"]],[]],[[],[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0"]]],[[],[["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14"]]],[[],[["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13"]]],[[],[["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12"]]],[[["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2","pin-type-component_fc486c6a-efa6-4e32-a1f3-0451662788c4_0"]],[]],[[["pin-type-component_1b0f4904-14bf-429f-937d-c99b5c2da67c_0","pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2"]],[]],[[["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2","pin-type-component_cb28eb0e-db83-4b4e-b021-b939f7a83c54_0"]],[]],[[["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2","pin-type-component_5cc5144a-e27c-4a8c-a3b8-dfdff02281da_0"]],[]],[[["pin-type-component_756a3f47-cc5c-4c12-8a88-5902936d2980_0","pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2"]],[]],[[["pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2","pin-type-component_f4cc5271-6fed-4fbe-b520-d7f27ca6d761_0"]],[]],[[["pin-type-component_515f6f7f-721f-439a-b2db-7f6c6ca7ad1f_0","pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2"]],[]],[[["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2","pin-type-component_7dc8ce5e-7fe0-4560-a90a-24f57026c2ce_0"]],[]],[[],[["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2","pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2"]]],[[],[["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2","pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2"]]],[[],[["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2","pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2"]]],[[],[["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2","pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2"]]],[[],[["pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_1","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_0"]]],[[],[["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1"]]],[[],[["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0","pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0"]]],[[],[["pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_1","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_0"]]],[[],[["pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0","pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0"]]],[[],[["pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0","pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0"]]],[[],[["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1"]]],[[],[["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1"]]],[[],[["pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0"]]],[[],[["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1"]]],[[],[["pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11"]]],[[],[["pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10"]]],[[],[["pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9"]]],[[],[["pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8"]]],[[],[["pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_1","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_0"]]],[[],[["pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_1","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_0"]]],[[],[["pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_1","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_0"]]],[[],[["pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_1","pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_0"]]],[[],[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0"]]],[[],[["pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0","pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0"]]],[[],[["pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0","pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0"]]],[[],[["pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0","pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_0"]]],[[["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2","pin-type-component_d23f20e3-e8e7-4a94-b362-814ae84c95f1_0"]],[]],[[["pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2","pin-type-component_78dc7030-f822-4db6-b90c-1a871bd2febd_0"]],[]],[[["pin-type-component_20c4afac-aed7-47a4-b18b-1cd7a3325c34_0","pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2"]],[]],[[["pin-type-component_02c2443e-51cb-49a5-b48e-828fe43ba847_0","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2"]],[]],[[["pin-type-component_9fb789aa-23a4-4c02-856a-7e2a62a5687c_0","pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2"]],[]],[[["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2","pin-type-component_a723fcb8-a29a-44f7-91e6-b934c414e1d5_0"]],[]],[[["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2","pin-type-component_a3ab8da7-d370-48c7-aed7-0afc87949c1f_0"]],[]],[[["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2","pin-type-component_80364b7e-c592-40e4-9f27-3a46aba92f9c_0"]],[]],[[],[["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2","pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2"]]],[[],[["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2","pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2"]]],[[],[["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2"]]],[[],[["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2","pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2"]]],[[],[["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2","pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1"]]],[[],[["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1"]]],[[],[["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1"]]],[[],[["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1"]]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15","pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1"]],[]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1"]],[]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13","pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1"]],[]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1"]],[]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1"]],[]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1"]],[]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1"]],[]],[[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1"]],[]],[[],[["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15"]]],[[],[["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14"]]],[[],[["pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13"]]],[[],[["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12"]]],[[],[["pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_1","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_0"]]],[[],[["pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_1","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_0"]]],[[],[["pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11"]]],[[],[["pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10"]]],[[],[["pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9"]]],[[],[["pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8"]]],[[],[["pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_7"]]],[[],[["pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_6"]]],[[],[["pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_5"]]],[[],[["pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_4"]]],[[["pin-type-component_1321abdf-76d2-4961-8eed-5e802ce03515_0","pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2"]],[]],[[["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2","pin-type-component_45b045d9-de2e-4c1e-9f03-8f59566339f3_0"]],[]],[[["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2","pin-type-component_e4ccca5e-2f92-4742-9f88-17c0acf9d0e5_0"]],[]],[[["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2","pin-type-component_34e49cee-f08a-4772-a6d4-df82dbc6905c_0"]],[]],[[["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2","pin-type-component_e03f3631-cb55-4d48-bf80-427e34299dc2_0"]],[]],[[["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2","pin-type-component_ada6e844-1bae-4716-870a-c40960a3bb4b_0"]],[]],[[["pin-type-component_5836c999-695f-47a8-8e7c-f38290544271_0","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2"]],[]],[[["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2","pin-type-component_c9571346-472b-4672-95d7-be31dc07bc93_0"]],[]],[[],[["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2"]]],[[],[["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2","pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2"]]],[[],[["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2","pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2"]]],[[],[["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2","pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2"]]],[[],[["pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1","pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_0"]]],[[],[["pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1","pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_0"]]],[[],[["pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1","pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_0"]]],[[],[["pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_1","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0"]]],[[],[["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0"]]],[[],[["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0"]]],[[],[["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0"]]],[[],[["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2","pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0"]]],[[],[["pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_0"]]],[[],[["pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_1"]]],[[],[["pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_2"]]],[[],[["pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_3"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1"]]],[[["pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12"]],[]],[[["pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11"]],[]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_1"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0","pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_1"]]],[[],[["pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_0","pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_0"]]],[[],[["pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_18"]]],[[],[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16","pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0"]]],[[],[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_18"]]],[[],[["pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_6"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_19","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_27"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_20","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_26"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_21","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_25"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_22","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_24"]]],[[],[["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_23","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_23"]]],[[],[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_19","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_8"]]],[[],[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_20","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_9"]]],[[],[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_21","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_10"]]],[[],[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_22","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_11"]]],[[],[["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_23","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_12"]]],[[],[["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_3"]]],[[],[["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_9","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_5"]]],[[],[["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_11","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_22"]]],[[],[["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_12","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_29"]]],[[],[["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_1","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_21"]]],[[],[["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_2","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_20"]]],[[],[["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_3","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_19"]]],[[],[["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_4","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_18"]]],[[],[["pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_4","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_7"]]],[[],[["pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_3","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_17"]]],[[],[["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"]]],[[["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0","pin-type-component_6c05b0a4-5167-4fc7-aa40-154354a323db_0"]],[]],[[["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"]],[]],[[],[["pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0"]]],[[["pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0"]],[]],[[["pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2"]],[]],[[],[["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1"]]],[[["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0"]],[]],[[],[["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1"]]],[[["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0"]],[]],[[],[["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1"]]],[[["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2","pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0"]],[]],[[],[["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0"]]],[[],[["pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0"]]],[[],[["pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0"]]],[[],[["pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0"]]],[[],[["pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0"]]],[[],[["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0"]]],[[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0"]],[]],[[],[]],[[],[]],[[],[["pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0"]]],[[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0"]],[]],[[],[["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0":"0000000000000066","pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_1":"0000000000000064","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0":"0000000000000102","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1":"0000000000000105","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2":"0000000000000108","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3":"0000000000000111","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4":"0000000000000098","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5":"0000000000000099","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6":"0000000000000093","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7":"0000000000000090","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8":"0000000000000087","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9":"0000000000000084","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10":"0000000000000081","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11":"0000000000000078","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12":"0000000000000075","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13":"0000000000000072","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14":"0000000000000069","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15":"0000000000000066","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16":"0000000000000116","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_17":"_","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_18":"0000000000000116","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_19":"0000000000000119","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_20":"0000000000000120","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_21":"0000000000000121","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_22":"0000000000000122","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_23":"0000000000000123","pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_0":"0000000000000004","pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_1":"0000000000000103","pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2":"0000000000000002","pin-type-component_7e9999e8-686e-4f02-b1e7-bee04a417b43_0":"0000000000000004","pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_0":"0000000000000006","pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_1":"0000000000000104","pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2":"0000000000000002","pin-type-component_4bfdc0b0-0087-4f19-b9da-fe77fe2030bb_0":"0000000000000006","pin-type-component_725c2e06-513a-456a-a054-9a1efd2410b5_0":"0000000000000008","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_0":"0000000000000010","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_1":"0000000000000101","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2":"0000000000000000","pin-type-component_84e67de5-59f5-4375-8901-060561a64dc9_0":"0000000000000010","pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_0":"0000000000000008","pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_1":"0000000000000100","pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2":"0000000000000000","pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_0":"0000000000000013","pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_1":"0000000000000110","pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2":"0000000000000007","pin-type-component_ad7b12e6-293b-4cf0-b5fc-2ad4811766ad_0":"0000000000000013","pin-type-component_84525e3e-ef29-4e0c-a293-959707966b26_0":"0000000000000003","pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_0":"0000000000000001","pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_1":"0000000000000107","pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2":"0000000000000005","pin-type-component_a4a81ac1-f999-4c5f-bf1d-d39d1364ba7e_0":"0000000000000001","pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_0":"0000000000000003","pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_1":"0000000000000106","pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2":"0000000000000005","pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_0":"0000000000000015","pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_1":"0000000000000109","pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2":"0000000000000007","pin-type-component_69b6c16b-f2c6-4ab0-b694-b43efd7d7efa_0":"0000000000000015","pin-type-component_7fc8671b-e701-4c33-a644-f42eace24307_0":"0000000000000023","pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_0":"0000000000000021","pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_1":"0000000000000095","pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2":"0000000000000018","pin-type-component_266aa6bb-5bae-4ff3-85db-bbd370178ae8_0":"0000000000000021","pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_0":"0000000000000023","pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_1":"0000000000000094","pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2":"0000000000000018","pin-type-component_0af45fa8-24bc-42e4-9c24-d15187e9fbc3_0":"0000000000000019","pin-type-component_5278fc75-d95d-4e4c-a86e-2e83a862e607_0":"0000000000000017","pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_0":"0000000000000019","pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1":"0000000000000096","pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2":"0000000000000016","pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_0":"0000000000000017","pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_1":"0000000000000097","pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2":"0000000000000016","pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_0":"0000000000000029","pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_1":"0000000000000089","pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2":"0000000000000022","pin-type-component_e7d36833-6d1a-490c-96e9-4f178d942f47_0":"0000000000000029","pin-type-component_3d109b51-1504-4d24-a9e7-9e3fe3074724_0":"0000000000000027","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_0":"0000000000000025","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_1":"0000000000000092","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2":"0000000000000020","pin-type-component_34445add-d974-48d4-81af-972f5dd7934b_0":"0000000000000025","pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_0":"0000000000000027","pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_1":"0000000000000091","pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2":"0000000000000020","pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_0":"0000000000000031","pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_1":"0000000000000088","pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2":"0000000000000022","pin-type-component_903934ae-30da-4a37-93c9-c64660e9c617_0":"0000000000000031","pin-type-component_5bdd54e6-172a-4994-8b34-5d8687be61e2_0":"0000000000000039","pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_0":"0000000000000037","pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_1":"0000000000000083","pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2":"0000000000000035","pin-type-component_62a268f0-68fa-4016-91c7-d55a738d6b46_0":"0000000000000037","pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_0":"0000000000000039","pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_1":"0000000000000082","pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2":"0000000000000035","pin-type-component_4732636d-ea0d-4b19-877e-d2ff4ddb5e8d_0":"0000000000000034","pin-type-component_7f294ee1-7ea8-4e70-bb0a-8c8b6b15b6c9_0":"0000000000000033","pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_0":"0000000000000034","pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_1":"0000000000000085","pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2":"0000000000000032","pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_0":"0000000000000033","pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_1":"0000000000000086","pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2":"0000000000000032","pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_0":"0000000000000061","pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_1":"0000000000000077","pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2":"0000000000000038","pin-type-component_b2f3a979-ce1b-444a-a7e4-6ef67b25f077_0":"0000000000000061","pin-type-component_0b4ba5d8-bcb4-4816-8dfe-3fa4ce9ed019_0":"0000000000000059","pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_0":"0000000000000041","pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_1":"0000000000000080","pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2":"0000000000000036","pin-type-component_29f2dcbd-c66e-4d22-9415-91c6505cd16b_0":"0000000000000041","pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_0":"0000000000000059","pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_1":"0000000000000079","pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2":"0000000000000036","pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_0":"0000000000000063","pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_1":"0000000000000076","pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2":"0000000000000038","pin-type-component_3b6d34de-cd89-4ef4-9473-da4b3ae907df_0":"0000000000000063","pin-type-component_dd44450f-fd4f-4059-aab9-565428093e7b_0":"0000000000000049","pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_0":"0000000000000047","pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_1":"0000000000000071","pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2":"0000000000000056","pin-type-component_6d57b374-4a97-4f2c-b0da-4d4ccbef4f5a_0":"0000000000000047","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_0":"0000000000000049","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_1":"0000000000000070","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2":"0000000000000056","pin-type-component_0c082f01-0561-48cc-887e-4e37deace687_0":"0000000000000045","pin-type-component_d1e6942e-6a34-4356-87fa-da19b68ae6b8_0":"0000000000000043","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_0":"0000000000000045","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_1":"0000000000000074","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2":"0000000000000046","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_0":"0000000000000043","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_1":"0000000000000073","pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2":"0000000000000046","pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_0":"0000000000000055","pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1":"0000000000000065","pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2":"0000000000000117","pin-type-component_bb4a8fb4-80b5-4764-a9f6-b3d9cae671c4_0":"0000000000000055","pin-type-component_636bd670-72c8-425e-8740-11540fc72a9f_0":"0000000000000053","pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_0":"0000000000000051","pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1":"0000000000000067","pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2":"0000000000000048","pin-type-component_e84ff89e-b801-43e3-905a-a7004860c743_0":"0000000000000051","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_0":"0000000000000053","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_1":"0000000000000068","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2":"0000000000000048","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_0":"0000000000000057","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_1":"0000000000000064","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2":"0000000000000117","pin-type-component_edb09e16-b982-4564-8c59-d0c31b14f784_0":"0000000000000057","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0":"0000000000000066","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1":"0000000000000065","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_0":"0000000000000028","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_1":"0000000000000030","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_2":"0000000000000114","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_3":"0000000000000115","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_4":"0000000000000016","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_5":"0000000000000018","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_6":"0000000000000020","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_7":"0000000000000022","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8":"0000000000000032","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9":"0000000000000035","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10":"0000000000000036","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11":"0000000000000038","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12":"0000000000000046","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13":"0000000000000056","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14":"0000000000000048","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15":"0000000000000117","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16":"0000000000000118","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_17":"_","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_18":"0000000000000118","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_19":"0000000000000124","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_20":"0000000000000125","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_21":"0000000000000126","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_22":"0000000000000127","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_23":"0000000000000128","pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0":"0000000000000069","pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_1":"0000000000000068","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_0":"0000000000000069","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1":"0000000000000067","pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0":"0000000000000072","pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_1":"0000000000000070","pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_0":"0000000000000072","pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_1":"0000000000000071","pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_0":"0000000000000075","pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_1":"0000000000000074","pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0":"0000000000000075","pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_1":"0000000000000073","pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_0":"0000000000000078","pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_1":"0000000000000076","pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0":"0000000000000078","pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_1":"0000000000000077","pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_0":"0000000000000081","pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_1":"0000000000000079","pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0":"0000000000000081","pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_1":"0000000000000080","pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_0":"0000000000000084","pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_1":"0000000000000082","pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0":"0000000000000084","pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_1":"0000000000000083","pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_0":"0000000000000087","pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_1":"0000000000000085","pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0":"0000000000000087","pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_1":"0000000000000086","pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_0":"0000000000000090","pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_1":"0000000000000088","pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0":"0000000000000090","pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_1":"0000000000000089","pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0":"0000000000000093","pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_1":"0000000000000091","pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_0":"0000000000000093","pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_1":"0000000000000092","pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0":"0000000000000099","pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_1":"0000000000000094","pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_0":"0000000000000099","pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_1":"0000000000000095","pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_0":"0000000000000098","pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_1":"0000000000000096","pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0":"0000000000000098","pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_1":"0000000000000097","pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_0":"0000000000000102","pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_1":"0000000000000100","pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0":"0000000000000102","pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_1":"0000000000000101","pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_0":"0000000000000105","pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_1":"0000000000000103","pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0":"0000000000000105","pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_1":"0000000000000104","pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_0":"0000000000000108","pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_1":"0000000000000106","pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0":"0000000000000108","pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_1":"0000000000000107","pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_0":"0000000000000111","pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_1":"0000000000000109","pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0":"0000000000000111","pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_1":"0000000000000110","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0":"0000000000000009","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1":"0000000000000044","pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0":"0000000000000044","pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1":"0000000000000046","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0":"0000000000000009","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1":"0000000000000050","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0":"0000000000000050","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1":"0000000000000056","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0":"0000000000000009","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1":"0000000000000052","pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0":"0000000000000052","pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1":"0000000000000048","pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0":"0000000000000009","pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1":"0000000000000054","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0":"0000000000000054","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1":"0000000000000117","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0":"0000000000000009","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_1":"0000000000000026","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_0":"0000000000000026","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1":"0000000000000038","pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0":"0000000000000009","pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_1":"0000000000000024","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_0":"0000000000000024","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1":"0000000000000036","pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0":"0000000000000009","pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_1":"0000000000000058","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_0":"0000000000000058","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1":"0000000000000035","pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0":"0000000000000009","pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_1":"0000000000000040","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_0":"0000000000000040","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1":"0000000000000032","pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0":"0000000000000009","pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_1":"0000000000000113","pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_0":"0000000000000113","pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1":"0000000000000022","pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0":"0000000000000009","pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_1":"0000000000000112","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_0":"0000000000000112","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1":"0000000000000020","pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0":"0000000000000009","pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_1":"0000000000000062","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_0":"0000000000000062","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1":"0000000000000018","pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_0":"0000000000000009","pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_1":"0000000000000060","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_0":"0000000000000060","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1":"0000000000000016","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0":"0000000000000009","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1":"0000000000000000","pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_0":"0000000000000000","pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_1":"0000000000000028","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0":"0000000000000009","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1":"0000000000000002","pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_0":"0000000000000002","pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_1":"0000000000000030","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0":"0000000000000009","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1":"0000000000000005","pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_0":"0000000000000005","pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_1":"0000000000000114","pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0":"0000000000000009","pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_1":"0000000000000007","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0":"0000000000000007","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_1":"0000000000000115","pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_0":"0000000000000116","pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_1":"0000000000000102","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_0":"0000000000000116","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_1":"0000000000000105","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_0":"0000000000000116","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_1":"0000000000000108","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_0":"0000000000000116","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_1":"0000000000000111","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_0":"0000000000000116","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_1":"0000000000000098","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_0":"0000000000000116","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_1":"0000000000000099","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_0":"0000000000000116","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_1":"0000000000000093","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_0":"0000000000000116","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_1":"0000000000000090","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_0":"0000000000000116","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_1":"0000000000000087","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_0":"0000000000000116","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_1":"0000000000000084","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_0":"0000000000000116","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_1":"0000000000000081","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_0":"0000000000000116","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_1":"0000000000000078","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_0":"0000000000000116","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1":"0000000000000075","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_0":"0000000000000116","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1":"0000000000000072","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_0":"0000000000000116","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_1":"0000000000000069","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_0":"0000000000000116","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_1":"0000000000000066","pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0":"0000000000000116","pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0":"0000000000000118","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_0":"_","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_1":"_","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_2":"_","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_3":"0000000000000009","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_4":"_","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_5":"0000000000000130","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_6":"0000000000000118","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_7":"0000000000000137","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_8":"0000000000000124","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_9":"0000000000000125","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_10":"0000000000000126","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_11":"0000000000000127","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_12":"0000000000000128","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_13":"_","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_14":"_","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_15":"_","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_16":"_","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_17":"0000000000000138","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_18":"0000000000000136","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_19":"0000000000000135","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_20":"0000000000000134","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_21":"0000000000000133","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_22":"0000000000000131","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_23":"0000000000000123","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_24":"0000000000000122","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_25":"0000000000000121","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_26":"0000000000000120","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_27":"0000000000000119","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_28":"_","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_29":"0000000000000132","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_30":"_","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_31":"_","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_0":"_","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_1":"0000000000000133","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_2":"0000000000000134","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_3":"0000000000000135","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_4":"0000000000000136","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_5":"_","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_6":"_","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_7":"_","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_8":"_","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_9":"0000000000000130","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10":"0000000000000009","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_11":"0000000000000131","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_12":"0000000000000132","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_13":"_","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_14":"_","pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_15":"_","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_0":"_","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_1":"_","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_2":"_","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_3":"0000000000000138","pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_4":"0000000000000137"},"component_id_to_pins":{"082451f0-7869-4209-aa80-c752e3204afe":["0","1"],"d448436c-9798-4335-8304-00153efa0c0f":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23"],"9e058603-a403-435e-a7b3-472988f8f796":["0","1","2"],"7e9999e8-686e-4f02-b1e7-bee04a417b43":["0"],"0fa29099-f06c-42e6-8abb-d829c961012c":["0","1","2"],"4bfdc0b0-0087-4f19-b9da-fe77fe2030bb":["0"],"725c2e06-513a-456a-a054-9a1efd2410b5":["0"],"f2a03157-3d3b-4891-9a96-ef7378eef59a":["0","1","2"],"84e67de5-59f5-4375-8901-060561a64dc9":["0"],"39ea5961-b6e7-49a0-8a1a-4a54142db333":["0","1","2"],"0ad2680b-02ba-49a2-a3e9-a96381a7d26e":["0","1","2"],"ad7b12e6-293b-4cf0-b5fc-2ad4811766ad":["0"],"84525e3e-ef29-4e0c-a293-959707966b26":["0"],"19cbe39d-a790-4e2e-bde4-0d5ef7c61da2":["0","1","2"],"a4a81ac1-f999-4c5f-bf1d-d39d1364ba7e":["0"],"548ad9b0-6450-4235-a7be-ccb79cd6080d":["0","1","2"],"d7dc068c-4b59-400e-ae50-562c7ccbc1ad":["0","1","2"],"69b6c16b-f2c6-4ab0-b694-b43efd7d7efa":["0"],"7fc8671b-e701-4c33-a644-f42eace24307":["0"],"8a57da25-4acd-4f0c-b8e8-8e9646645470":["0","1","2"],"266aa6bb-5bae-4ff3-85db-bbd370178ae8":["0"],"a42f6e75-c6ce-4431-8ab7-a546cadc6910":["0","1","2"],"0af45fa8-24bc-42e4-9c24-d15187e9fbc3":["0"],"5278fc75-d95d-4e4c-a86e-2e83a862e607":["0"],"8d75e431-ab93-4f28-a072-73fa2a9add70":["0","1","2"],"6fba6b65-b569-4c04-b286-0556b7aca02c":["0","1","2"],"458ace7d-db58-47fe-9e9e-81463f1cb31c":["0","1","2"],"e7d36833-6d1a-490c-96e9-4f178d942f47":["0"],"3d109b51-1504-4d24-a9e7-9e3fe3074724":["0"],"ddf014d2-e81b-4ce5-802e-4329eb48f7e0":["0","1","2"],"34445add-d974-48d4-81af-972f5dd7934b":["0"],"274be705-445b-40a5-9ab8-ea55a1873ac7":["0","1","2"],"8ac7020a-2504-45c9-b517-84bd506cb24c":["0","1","2"],"903934ae-30da-4a37-93c9-c64660e9c617":["0"],"5bdd54e6-172a-4994-8b34-5d8687be61e2":["0"],"a28b7076-045f-481a-8987-e6c379c85461":["0","1","2"],"62a268f0-68fa-4016-91c7-d55a738d6b46":["0"],"3cc0d351-6a54-4350-a5dc-29ea6ac8f53f":["0","1","2"],"4732636d-ea0d-4b19-877e-d2ff4ddb5e8d":["0"],"7f294ee1-7ea8-4e70-bb0a-8c8b6b15b6c9":["0"],"3569e0a5-063e-4474-b7f3-fd780070bcdd":["0","1","2"],"01ef38d5-a6be-49e6-b75b-fe4690ca3d8a":["0","1","2"],"b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99":["0","1","2"],"b2f3a979-ce1b-444a-a7e4-6ef67b25f077":["0"],"0b4ba5d8-bcb4-4816-8dfe-3fa4ce9ed019":["0"],"8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b":["0","1","2"],"29f2dcbd-c66e-4d22-9415-91c6505cd16b":["0"],"549bec3f-89a4-4854-8eed-2d9171821a2f":["0","1","2"],"1b855ccb-49a4-427a-9563-e1bcdb16e638":["0","1","2"],"3b6d34de-cd89-4ef4-9473-da4b3ae907df":["0"],"dd44450f-fd4f-4059-aab9-565428093e7b":["0"],"3a88c66b-feb0-48c3-be15-37e3d48518eb":["0","1","2"],"6d57b374-4a97-4f2c-b0da-4d4ccbef4f5a":["0"],"46f90c07-7d13-4392-a3bf-e813e3dabb36":["0","1","2"],"0c082f01-0561-48cc-887e-4e37deace687":["0"],"d1e6942e-6a34-4356-87fa-da19b68ae6b8":["0"],"83dcf7d9-214a-4ba8-8c4b-0198867c485d":["0","1","2"],"041b5070-e88a-4a6b-aa2c-a93c5f45650d":["0","1","2"],"67df4d37-3f2b-4d48-9904-dc3e640854f2":["0","1","2"],"bb4a8fb4-80b5-4764-a9f6-b3d9cae671c4":["0"],"636bd670-72c8-425e-8740-11540fc72a9f":["0"],"7cf5453a-9a65-47be-a0c1-a40e3c54981e":["0","1","2"],"e84ff89e-b801-43e3-905a-a7004860c743":["0"],"73ff6e4f-35de-4fa1-bb93-81012f621ef2":["0","1","2"],"8fd76732-6e42-40ac-b9ab-aae7428798a1":["0","1","2"],"edb09e16-b982-4564-8c59-d0c31b14f784":["0"],"eeac935f-c26f-4957-912d-5c92ef07716f":["0","1"],"11da4e6e-750e-4643-874f-89e7cea28441":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23"],"4505b10f-85e5-4973-b4b5-e3d656f3d0be":["0","1"],"b2e81b6c-d2d3-439c-82a2-c21100e871d6":["0","1"],"88c754f5-de3a-41e9-8e1a-6c44284e3b38":["0","1"],"ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1":["0","1"],"0077cc15-4d99-4651-a57e-536f288016fb":["0","1"],"dba2be22-3f32-4819-979e-cd2ac0c4cc6e":["0","1"],"7a6ab358-5837-431b-9348-a619c0d5eb4b":["0","1"],"8281ae65-4ada-4b48-aeec-e666f55d538a":["0","1"],"d121ccd5-ebd1-4e31-80c7-213974efb4b7":["0","1"],"c51e4057-62bf-4d4d-97d5-80d833dcecd9":["0","1"],"daff2923-49a4-426d-8290-92f3de68e4c8":["0","1"],"e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9":["0","1"],"c1ec2684-5203-484a-bb58-714d3d1ff689":["0","1"],"c2e4f40c-d3fa-4534-902a-b6ca784f2d33":["0","1"],"89080e17-209d-40ef-8155-edbb76fffbef":["0","1"],"dbc09422-6bd6-4f89-bf7e-49c71fb62af9":["0","1"],"9ab5a6ac-c827-4cf6-9b73-708335a1a9b0":["0","1"],"35a17054-5a08-4aee-9aa6-e124f96682e1":["0","1"],"d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c":["0","1"],"0152d242-8b4d-42db-8096-0f8dc98256f3":["0","1"],"35159cb3-cc74-4c90-b0f5-cff583f979a5":["0","1"],"2f031f22-1944-43ab-ae9c-f74e47cc4156":["0","1"],"625dbf85-54ff-48b2-a275-4089e5081167":["0","1"],"f86ac869-5086-4a06-8cd6-49f486548944":["0","1"],"0c68c6e3-0464-4e71-ab6a-9086b01a0e77":["0","1"],"709ba052-a0a0-4439-a40d-83aedf155550":["0","1"],"4b0e618a-0090-4173-a14d-dc77951515d3":["0","1"],"733ac60f-fd5b-4e01-bcd0-44ae417225ee":["0","1"],"114d5d14-5f5c-40e8-b182-5aaaa19436dd":["0","1"],"4f53b9c5-5f30-4a72-af1a-a8232ad99f6b":["0","1"],"621585ad-95ad-4cf3-9a10-1ca969371d4e":["0","1"],"995a17d1-5928-497f-b230-e981cff0c0da":["0","1"],"efd3f3bc-1ae1-45dd-a482-193032279b23":["0","1"],"81ae35b1-5b71-4716-a1af-fd111af3ac03":["0","1"],"a86bd662-6cba-44a0-8211-7ce5de8f1e54":["0","1"],"41446abf-3582-4e1a-bca9-cf131a5fba1c":["0","1"],"0d024f4d-e2f2-4b76-8f77-420b1168f36c":["0","1"],"3694689b-7dc6-49dc-a8fa-3e18614c7e29":["0","1"],"7807e964-3bc8-4b12-bb6c-44a1c1b24af9":["0","1"],"38df7453-f88c-4a99-82c0-fdb338cc7264":["0","1"],"4b269a77-3c6b-4832-bc03-819b3941bca2":["0","1"],"ca018356-08f3-4416-b12e-ca10c6c7bb67":["0","1"],"5712632d-8fa8-495b-a104-baf8f43c700a":["0","1"],"efcea04e-21d8-44a5-8f0d-74277474a2e0":["0","1"],"b69e0669-3879-4abd-9d7d-acc45f8eea74":["0","1"],"a8e515ed-cb32-4abf-ab34-4e8ba550aff5":["0","1"],"c90e906b-172f-43f0-a66d-c99371504fba":["0","1"],"15591579-4d1a-4075-aec4-52c43cc21020":["0","1"],"ee4052d6-2dbe-445a-8b8e-b1c8214d283a":["0","1"],"c58023a8-eade-4368-93d4-c18f7148e8e3":["0","1"],"ddbc596a-7cd5-4048-bdec-ae929062b39f":["0","1"],"e7200013-28f8-4ff6-9dbe-a2239e215492":["0","1"],"0b992200-29a8-47ae-9e2d-5041f24e3da4":["0","1"],"c107267e-960a-414d-898a-9b8f86844804":["0","1"],"3c883d29-f62b-49cf-a092-2c8c9f097c17":["0","1"],"f7984d9c-52aa-415e-b39c-e5fb625b93c2":["0","1"],"c525269a-6029-466e-8297-23d196a50c50":["0","1"],"c94229bb-b925-4416-b768-559f9d5d84b6":["0","1"],"42b98079-caa9-47e9-bd5d-65893e0dce4d":["0","1"],"662aa0ec-65ba-4d5d-a487-5ed33ea6d988":["0","1"],"5008935e-c93f-4fb4-a087-0abedc96eefb":["0","1"],"b45ca744-aa2b-4e0a-b23d-32ff2cca7a14":["0","1"],"fe152afb-21b1-47d5-b9c6-bd2b619f0439":["0","1"],"13bb41c2-0891-49e2-a36d-a0e52211de2b":["0","1"],"5d50f226-59dc-49dd-a79a-abbf5e3cb510":["0","1"],"58089c3e-bb30-4b9d-87df-71065baedba4":["0","1"],"824c2884-8b95-4bf2-9b1d-fc37145bfe37":["0","1"],"e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00":["0","1"],"a72804f7-e18d-407a-8183-98f8e53fe3d0":["0","1"],"bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1":["0","1"],"07965d4a-3c19-478e-9e88-2147d6a70aba":["0","1"],"b7e27884-48f5-44d6-9ad2-56da1f22ae1e":["0","1"],"b68f3984-33e3-4099-9fd0-2bf2992dd7c5":["0","1"],"ed5c99e1-3753-4905-b880-1ffcf976d135":["0","1"],"1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf":["0","1"],"6b9ac4cf-8b15-40e0-9908-87be89d7dd12":["0","1"],"6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88":["0","1"],"0e24347f-56a1-4fe8-a3eb-00f61ef717e3":["0","1"],"2d2c1fc2-9459-4e52-81e7-c39a9a7813f6":["0"],"935ec2c0-76f9-4c06-a88a-d876d661b1e8":["0"],"9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"],"0a8678a1-8b77-47ac-8524-d596b3cedd6d":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15"],"6fe13b46-5e6b-4103-adfc-cce8f32c36a7":["0","1","2","3","4"]},"uid_to_net":{"_":[],"0000000000000004":["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_0","pin-type-component_7e9999e8-686e-4f02-b1e7-bee04a417b43_0"],"0000000000000006":["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_0","pin-type-component_4bfdc0b0-0087-4f19-b9da-fe77fe2030bb_0"],"0000000000000008":["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_0","pin-type-component_725c2e06-513a-456a-a054-9a1efd2410b5_0"],"0000000000000010":["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_0","pin-type-component_84e67de5-59f5-4375-8901-060561a64dc9_0"],"0000000000000001":["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_0","pin-type-component_a4a81ac1-f999-4c5f-bf1d-d39d1364ba7e_0"],"0000000000000003":["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_0","pin-type-component_84525e3e-ef29-4e0c-a293-959707966b26_0"],"0000000000000013":["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_0","pin-type-component_ad7b12e6-293b-4cf0-b5fc-2ad4811766ad_0"],"0000000000000015":["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_0","pin-type-component_69b6c16b-f2c6-4ab0-b694-b43efd7d7efa_0"],"0000000000000017":["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_0","pin-type-component_5278fc75-d95d-4e4c-a86e-2e83a862e607_0"],"0000000000000019":["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_0","pin-type-component_0af45fa8-24bc-42e4-9c24-d15187e9fbc3_0"],"0000000000000021":["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_0","pin-type-component_266aa6bb-5bae-4ff3-85db-bbd370178ae8_0"],"0000000000000023":["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_0","pin-type-component_7fc8671b-e701-4c33-a644-f42eace24307_0"],"0000000000000025":["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_0","pin-type-component_34445add-d974-48d4-81af-972f5dd7934b_0"],"0000000000000027":["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_0","pin-type-component_3d109b51-1504-4d24-a9e7-9e3fe3074724_0"],"0000000000000029":["pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_0","pin-type-component_e7d36833-6d1a-490c-96e9-4f178d942f47_0"],"0000000000000031":["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_0","pin-type-component_903934ae-30da-4a37-93c9-c64660e9c617_0"],"0000000000000033":["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_0","pin-type-component_7f294ee1-7ea8-4e70-bb0a-8c8b6b15b6c9_0"],"0000000000000034":["pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_0","pin-type-component_4732636d-ea0d-4b19-877e-d2ff4ddb5e8d_0"],"0000000000000037":["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_0","pin-type-component_62a268f0-68fa-4016-91c7-d55a738d6b46_0"],"0000000000000039":["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_0","pin-type-component_5bdd54e6-172a-4994-8b34-5d8687be61e2_0"],"0000000000000041":["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_0","pin-type-component_29f2dcbd-c66e-4d22-9415-91c6505cd16b_0"],"0000000000000043":["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_0","pin-type-component_d1e6942e-6a34-4356-87fa-da19b68ae6b8_0"],"0000000000000045":["pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_0","pin-type-component_0c082f01-0561-48cc-887e-4e37deace687_0"],"0000000000000047":["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_0","pin-type-component_6d57b374-4a97-4f2c-b0da-4d4ccbef4f5a_0"],"0000000000000049":["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_0","pin-type-component_dd44450f-fd4f-4059-aab9-565428093e7b_0"],"0000000000000051":["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_0","pin-type-component_e84ff89e-b801-43e3-905a-a7004860c743_0"],"0000000000000053":["pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_0","pin-type-component_636bd670-72c8-425e-8740-11540fc72a9f_0"],"0000000000000055":["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_0","pin-type-component_bb4a8fb4-80b5-4764-a9f6-b3d9cae671c4_0"],"0000000000000057":["pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_0","pin-type-component_edb09e16-b982-4564-8c59-d0c31b14f784_0"],"0000000000000059":["pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_0","pin-type-component_0b4ba5d8-bcb4-4816-8dfe-3fa4ce9ed019_0"],"0000000000000061":["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_0","pin-type-component_b2f3a979-ce1b-444a-a7e4-6ef67b25f077_0"],"0000000000000063":["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_0","pin-type-component_3b6d34de-cd89-4ef4-9473-da4b3ae907df_0"],"0000000000000064":["pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_1","pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_1"],"0000000000000065":["pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1"],"0000000000000066":["pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15","pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_1"],"0000000000000068":["pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_1","pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_1"],"0000000000000067":["pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1"],"0000000000000069":["pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0","pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_1"],"0000000000000070":["pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_1","pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_1"],"0000000000000071":["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_1","pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_1"],"0000000000000072":["pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0","pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1"],"0000000000000073":["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_1","pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_1"],"0000000000000074":["pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_1","pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_1"],"0000000000000075":["pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12","pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1"],"0000000000000076":["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_1","pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_1"],"0000000000000077":["pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_1","pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_1"],"0000000000000078":["pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_0","pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_1"],"0000000000000079":["pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_1","pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_1"],"0000000000000080":["pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_1","pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_1"],"0000000000000081":["pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0","pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_1"],"0000000000000082":["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_1","pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_1"],"0000000000000083":["pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_1","pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_1"],"0000000000000084":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9","pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_0","pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_1"],"0000000000000085":["pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_1","pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_1"],"0000000000000086":["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_1","pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_1"],"0000000000000087":["pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_0","pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8","pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_1"],"0000000000000088":["pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_1","pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_1"],"0000000000000089":["pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_1","pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_1"],"0000000000000090":["pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7","pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_1"],"0000000000000091":["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_1","pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_1"],"0000000000000092":["pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_1","pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_1"],"0000000000000093":["pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_0","pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_1"],"0000000000000094":["pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_1","pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_1"],"0000000000000095":["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_1","pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_1"],"0000000000000096":["pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1","pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_1"],"0000000000000097":["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_1","pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_1"],"0000000000000098":["pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0","pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_1"],"0000000000000099":["pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5","pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_1"],"0000000000000100":["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_1","pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_1"],"0000000000000101":["pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_1","pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_1"],"0000000000000102":["pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0","pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0","pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_1"],"0000000000000103":["pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_1","pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_1"],"0000000000000104":["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_1","pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_1"],"0000000000000105":["pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_0","pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_1"],"0000000000000106":["pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_1","pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_1"],"0000000000000107":["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_1","pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_1"],"0000000000000108":["pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_0","pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_1"],"0000000000000109":["pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_1","pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_1"],"0000000000000110":["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_1","pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_1"],"0000000000000111":["pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_0","pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_1"],"0000000000000044":["pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1"],"0000000000000046":["pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2","pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2","pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12"],"0000000000000056":["pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2","pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13"],"0000000000000048":["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1","pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2","pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14"],"0000000000000117":["pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1","pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2","pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15"],"0000000000000050":["pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1","pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0"],"0000000000000052":["pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1"],"0000000000000054":["pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1","pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0"],"0000000000000032":["pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2","pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8"],"0000000000000035":["pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2","pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9"],"0000000000000036":["pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2","pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10"],"0000000000000038":["pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1","pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11"],"0000000000000040":["pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_1","pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_0"],"0000000000000058":["pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_1","pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_0"],"0000000000000060":["pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_1","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_0"],"0000000000000062":["pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_1","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_0"],"0000000000000112":["pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_1","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_0"],"0000000000000113":["pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_1","pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_0"],"0000000000000016":["pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2","pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2","pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_4"],"0000000000000018":["pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2","pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2","pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_5"],"0000000000000020":["pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2","pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1","pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_6"],"0000000000000022":["pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1","pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2","pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_7"],"0000000000000024":["pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_1","pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_0"],"0000000000000026":["pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_1","pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_0"],"0000000000000000":["pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1","pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2","pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_0"],"0000000000000002":["pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2","pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1","pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_0"],"0000000000000005":["pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1","pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2","pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_0"],"0000000000000007":["pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2","pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_1","pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0","pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2"],"0000000000000028":["pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_0"],"0000000000000030":["pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_1"],"0000000000000114":["pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_2"],"0000000000000115":["pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_1","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_3"],"0000000000000116":["pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_0","pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_0","pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_0","pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_0","pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0","pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_0","pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_0","pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_0","pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_0","pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_0","pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_0","pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_0","pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_0","pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16","pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_0","pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_0","pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_0","pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_18"],"0000000000000118":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16","pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_18","pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_6"],"0000000000000119":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_19","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_27"],"0000000000000120":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_20","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_26"],"0000000000000121":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_21","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_25"],"0000000000000122":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_22","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_24"],"0000000000000123":["pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_23","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_23"],"0000000000000124":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_19","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_8"],"0000000000000125":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_20","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_9"],"0000000000000126":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_21","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_10"],"0000000000000127":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_22","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_11"],"0000000000000128":["pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_23","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_12"],"0000000000000130":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_9","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_5"],"0000000000000131":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_11","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_22"],"0000000000000132":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_12","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_29"],"0000000000000133":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_1","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_21"],"0000000000000134":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_2","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_20"],"0000000000000135":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_3","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_19"],"0000000000000136":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_4","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_18"],"0000000000000137":["pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_4","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_7"],"0000000000000138":["pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_3","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_17"],"0000000000000009":["pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10","pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_0","pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0","pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0","pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0","pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0","pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0","pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0","pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0","pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0","pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_3","pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0","pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0","pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0","pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0","pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0","pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0","pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0"]},"uid_to_text_label":{"0000000000000004":"Net 4","0000000000000006":"Net 6","0000000000000008":"Net 8","0000000000000010":"Net 10","0000000000000001":"Net 1","0000000000000003":"Net 3","0000000000000013":"Net 13","0000000000000015":"Net 15","0000000000000017":"Net 17","0000000000000019":"Net 19","0000000000000021":"Net 21","0000000000000023":"Net 23","0000000000000025":"Net 25","0000000000000027":"Net 27","0000000000000029":"Net 29","0000000000000031":"Net 31","0000000000000033":"Net 33","0000000000000034":"Net 34","0000000000000037":"Net 37","0000000000000039":"Net 39","0000000000000041":"Net 41","0000000000000043":"Net 43","0000000000000045":"Net 45","0000000000000047":"Net 47","0000000000000049":"Net 49","0000000000000051":"Net 51","0000000000000053":"Net 53","0000000000000055":"Net 55","0000000000000057":"Net 57","0000000000000059":"Net 59","0000000000000061":"Net 61","0000000000000063":"Net 63","0000000000000064":"Net 64","0000000000000065":"Net 65","0000000000000066":"Net 66","0000000000000068":"Net 68","0000000000000067":"Net 67","0000000000000069":"Net 69","0000000000000070":"Net 70","0000000000000071":"Net 71","0000000000000072":"Net 72","0000000000000073":"Net 73","0000000000000074":"Net 74","0000000000000075":"Net 75","0000000000000076":"Net 76","0000000000000077":"Net 77","0000000000000078":"Net 78","0000000000000079":"Net 79","0000000000000080":"Net 80","0000000000000081":"Net 81","0000000000000082":"Net 82","0000000000000083":"Net 83","0000000000000084":"Net 84","0000000000000085":"Net 85","0000000000000086":"Net 86","0000000000000087":"Net 87","0000000000000088":"Net 88","0000000000000089":"Net 89","0000000000000090":"Net 90","0000000000000091":"Net 91","0000000000000092":"Net 92","0000000000000093":"Net 93","0000000000000094":"Net 94","0000000000000095":"Net 95","0000000000000096":"Net 96","0000000000000097":"Net 97","0000000000000098":"Net 98","0000000000000099":"Net 99","0000000000000100":"Net 100","0000000000000101":"Net 101","0000000000000102":"Net 102","0000000000000103":"Net 103","0000000000000104":"Net 104","0000000000000105":"Net 105","0000000000000106":"Net 106","0000000000000107":"Net 107","0000000000000108":"Net 108","0000000000000109":"Net 109","0000000000000110":"Net 110","0000000000000111":"Net 111","0000000000000044":"Net 44","0000000000000046":"Net 46","0000000000000056":"Net 56","0000000000000048":"Net 48","0000000000000117":"Net 117","0000000000000050":"Net 50","0000000000000052":"Net 52","0000000000000054":"Net 54","0000000000000032":"Net 32","0000000000000035":"Net 35","0000000000000036":"Net 36","0000000000000038":"Net 38","0000000000000040":"Net 40","0000000000000058":"Net 58","0000000000000060":"Net 60","0000000000000062":"Net 62","0000000000000112":"Net 112","0000000000000113":"Net 113","0000000000000016":"Net 16","0000000000000018":"Net 18","0000000000000020":"Net 20","0000000000000022":"Net 22","0000000000000024":"Net 24","0000000000000026":"Net 26","0000000000000000":"Net 0","0000000000000002":"Net 2","0000000000000005":"Net 5","0000000000000007":"Net 7","0000000000000028":"Net 28","0000000000000030":"Net 30","0000000000000114":"Net 114","0000000000000115":"Net 115","0000000000000116":"Net 116","0000000000000118":"Net 118","0000000000000119":"Net 119","0000000000000120":"Net 120","0000000000000121":"Net 121","0000000000000122":"Net 122","0000000000000123":"Net 123","0000000000000124":"Net 124","0000000000000125":"Net 125","0000000000000126":"Net 126","0000000000000127":"Net 127","0000000000000128":"Net 128","0000000000000130":"Net 130","0000000000000131":"Net 131","0000000000000132":"Net 132","0000000000000133":"Net 133","0000000000000134":"Net 134","0000000000000135":"Net 135","0000000000000136":"Net 136","0000000000000137":"Net 137","0000000000000138":"Net 138","0000000000000009":"Net 9"},"all_breadboard_info_list":[],"breadboard_info_list":[],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1707.5625005000006,-666.7614504999999],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"082451f0-7869-4209-aa80-c752e3204afe","orientation":"left","circleData":[[-1707.5,-640],[-1707.5,-695.7041515000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-372.5,-572.5000000000001],"typeId":"b7d4df28-c430-b8ca-f42b-be40986a361e","componentVersion":1,"instanceId":"d448436c-9798-4335-8304-00153efa0c0f","orientation":"up","circleData":[[-417.5,-460],[-417.5,-475.0000000000001],[-417.5,-490.0000000000001],[-417.5,-505],[-417.5,-520.0000000000001],[-417.5,-535.0000000000001],[-417.5,-550.0000000000001],[-417.5,-565.0000000000001],[-417.5,-580.0000000000001],[-417.5,-595.0000000000001],[-417.5,-610.0000000000001],[-417.5,-625.0000000000001],[-417.5,-640.0000000000003],[-417.5,-655.0000000000001],[-417.5,-670.0000000000003],[-417.5,-685.0000000000003],[-327.49999999999994,-520.0000000000001],[-327.49999999999994,-535.0000000000001],[-327.49999999999994,-550.0000000000001],[-327.49999999999994,-565.0000000000001],[-327.49999999999994,-580.0000000000001],[-327.49999999999994,-595.0000000000001],[-327.49999999999994,-610.0000000000001],[-327.49999999999994,-625.0000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1004.0648299999981,-189.85064199999965],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"7e9999e8-686e-4f02-b1e7-bee04a417b43","orientation":"left","circleData":[[-1032.499999999999,-189.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1087.4999749999997,-52.49997549999989],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"0fa29099-f06c-42e6-8abb-d829c961012c","orientation":"right","circleData":[[-1062.4999999999995,-69.99999999999982],[-1062.4999999999995,-54.99999999999976],[-1062.4999999999995,-39.99999999999976]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1004.0648299999988,-84.85064199999931],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"4bfdc0b0-0087-4f19-b9da-fe77fe2030bb","orientation":"left","circleData":[[-1032.499999999999,-84.99999999999982]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1087.4999750000002,-157.49997550000012],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"9e058603-a403-435e-a7b3-472988f8f796","orientation":"right","circleData":[[-1062.4999999999995,-175.00000000000006],[-1062.4999999999995,-159.9999999999999],[-1062.4999999999995,-144.9999999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1004.0648299999984,35.14935800000012],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"725c2e06-513a-456a-a054-9a1efd2410b5","orientation":"left","circleData":[[-1032.4999999999998,34.999999999999886]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1004.064829999999,140.14935800000057],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"84e67de5-59f5-4375-8901-060561a64dc9","orientation":"left","circleData":[[-1032.5,139.99999999999986]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1087.4999750000006,67.50002449999965],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"39ea5961-b6e7-49a0-8a1a-4a54142db333","orientation":"right","circleData":[[-1062.4999999999998,49.999999999999716],[-1062.4999999999998,64.99999999999989],[-1062.4999999999998,79.99999999999989]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1087.4999750000009,-577.4999755000001],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"0ad2680b-02ba-49a2-a3e9-a96381a7d26e","orientation":"right","circleData":[[-1062.5,-595],[-1062.5,-579.9999999999998],[-1062.5,-564.9999999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1004.0648299999991,-609.8506419999999],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"ad7b12e6-293b-4cf0-b5fc-2ad4811766ad","orientation":"left","circleData":[[-1032.4999999999995,-610.0000000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1004.0648299999987,-489.8506419999993],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"84525e3e-ef29-4e0c-a293-959707966b26","orientation":"left","circleData":[[-1032.5000000000002,-489.9999999999996]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1087.4999750000006,-352.4999754999999],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"19cbe39d-a790-4e2e-bde4-0d5ef7c61da2","orientation":"right","circleData":[[-1062.5000000000005,-369.99999999999955],[-1062.5000000000005,-354.9999999999995],[-1062.5000000000005,-339.99999999999955]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1004.0648299999995,-384.8506419999991],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"a4a81ac1-f999-4c5f-bf1d-d39d1364ba7e","orientation":"left","circleData":[[-1032.5000000000005,-384.99999999999955]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1087.499975000001,-457.49997549999966],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"548ad9b0-6450-4235-a7be-ccb79cd6080d","orientation":"right","circleData":[[-1062.5000000000002,-474.9999999999997],[-1062.5000000000002,-459.99999999999955],[-1062.5000000000002,-444.99999999999955]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1087.4999750000009,-697.4999755000001],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"d7dc068c-4b59-400e-ae50-562c7ccbc1ad","orientation":"right","circleData":[[-1062.5,-715.0000000000001],[-1062.5,-699.9999999999999],[-1062.5,-684.9999999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1004.0648299999991,-729.8506419999999],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"69b6c16b-f2c6-4ab0-b694-b43efd7d7efa","orientation":"left","circleData":[[-1032.4999999999995,-730.0000000000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1274.064829999999,-189.85064199999965],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"7fc8671b-e701-4c33-a644-f42eace24307","orientation":"left","circleData":[[-1302.4999999999993,-189.99999999999983]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1357.4999749999997,-52.49997549999989],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"8a57da25-4acd-4f0c-b8e8-8e9646645470","orientation":"right","circleData":[[-1332.4999999999995,-69.99999999999972],[-1332.4999999999995,-54.99999999999966],[-1332.4999999999995,-39.999999999999645]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1274.0648299999984,-84.8506419999992],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"266aa6bb-5bae-4ff3-85db-bbd370178ae8","orientation":"left","circleData":[[-1302.499999999999,-84.9999999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1357.4999750000002,-157.4999754999999],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"a42f6e75-c6ce-4431-8ab7-a546cadc6910","orientation":"right","circleData":[[-1332.4999999999995,-174.99999999999994],[-1332.4999999999995,-159.99999999999977],[-1332.4999999999995,-144.99999999999977]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1274.064829999999,35.14935800000012],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"0af45fa8-24bc-42e4-9c24-d15187e9fbc3","orientation":"left","circleData":[[-1302.4999999999998,34.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1274.0648299999993,140.14935800000035],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"5278fc75-d95d-4e4c-a86e-2e83a862e607","orientation":"left","circleData":[[-1302.5000000000002,139.99999999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1357.4999750000006,67.50002449999988],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"8d75e431-ab93-4f28-a072-73fa2a9add70","orientation":"right","circleData":[[-1332.4999999999998,49.99999999999984],[-1332.4999999999998,65],[-1332.4999999999998,80]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1357.4999750000002,172.50002449999965],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"6fba6b65-b569-4c04-b286-0556b7aca02c","orientation":"right","circleData":[[-1332.5,155],[-1332.5,170.00000000000006],[-1332.5,185.00000000000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1357.4999750000002,-577.4999755],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"458ace7d-db58-47fe-9e9e-81463f1cb31c","orientation":"right","circleData":[[-1332.5,-594.9999999999999],[-1332.5,-579.9999999999997],[-1332.5,-564.9999999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1274.0648299999991,-609.8506419999998],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"e7d36833-6d1a-490c-96e9-4f178d942f47","orientation":"left","circleData":[[-1302.4999999999995,-610.0000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1274.064829999999,-489.8506419999991],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"3d109b51-1504-4d24-a9e7-9e3fe3074724","orientation":"left","circleData":[[-1302.5000000000002,-489.99999999999955]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1357.4999750000009,-352.4999754999998],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"ddf014d2-e81b-4ce5-802e-4329eb48f7e0","orientation":"right","circleData":[[-1332.5000000000005,-369.99999999999943],[-1332.5000000000005,-354.9999999999994],[-1332.5000000000005,-339.99999999999943]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1274.0648300000007,-384.85064199999886],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"34445add-d974-48d4-81af-972f5dd7934b","orientation":"left","circleData":[[-1302.5000000000002,-384.99999999999943]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1357.499975000001,-457.49997549999955],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"274be705-445b-40a5-9ab8-ea55a1873ac7","orientation":"right","circleData":[[-1332.5000000000002,-474.99999999999955],[-1332.5000000000002,-459.99999999999943],[-1332.5000000000002,-444.99999999999943]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1357.4999750000006,-697.4999755],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"8ac7020a-2504-45c9-b517-84bd506cb24c","orientation":"right","circleData":[[-1332.5,-715],[-1332.5,-699.9999999999998],[-1332.5,-684.9999999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1274.0648299999991,-729.8506419999998],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"903934ae-30da-4a37-93c9-c64660e9c617","orientation":"left","circleData":[[-1302.4999999999995,-730.0000000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1529.064829999998,-204.85064200000033],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"5bdd54e6-172a-4994-8b34-5d8687be61e2","orientation":"left","circleData":[[-1557.4999999999986,-205.00000000000063]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1612.4999749999997,-172.4999755000008],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"3cc0d351-6a54-4350-a5dc-29ea6ac8f53f","orientation":"right","circleData":[[-1587.499999999999,-190.00000000000074],[-1587.499999999999,-175.00000000000057],[-1587.499999999999,-160.00000000000057]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1529.0648299999984,125.14935799999967],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"7f294ee1-7ea8-4e70-bb0a-8c8b6b15b6c9","orientation":"left","circleData":[[-1557.4999999999995,124.99999999999918]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1612.4999750000002,52.5000244999992],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"3569e0a5-063e-4474-b7f3-fd780070bcdd","orientation":"right","circleData":[[-1587.4999999999993,34.99999999999903],[-1587.4999999999993,49.9999999999992],[-1587.4999999999993,64.9999999999992]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1612.4999749999997,157.50002449999897],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"01ef38d5-a6be-49e6-b75b-fe4690ca3d8a","orientation":"right","circleData":[[-1587.4999999999995,139.9999999999992],[-1587.4999999999995,154.99999999999926],[-1587.4999999999995,169.9999999999992]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1612.499975,-592.4999755000008],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99","orientation":"right","circleData":[[-1587.4999999999995,-610.0000000000007],[-1587.4999999999995,-595.0000000000005],[-1587.4999999999995,-580.0000000000005]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1529.064829999999,-624.8506420000008],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"b2f3a979-ce1b-444a-a7e4-6ef67b25f077","orientation":"left","circleData":[[-1557.499999999999,-625.0000000000011]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1529.064829999999,-504.85064200000033],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"0b4ba5d8-bcb4-4816-8dfe-3fa4ce9ed019","orientation":"left","circleData":[[-1557.5,-505.0000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1612.4999750000002,-367.49997550000035],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b","orientation":"right","circleData":[[-1587.5,-385.00000000000006],[-1587.5,-370],[-1587.5,-355.00000000000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1529.0648299999993,-399.8506420000001],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"29f2dcbd-c66e-4d22-9415-91c6505cd16b","orientation":"left","circleData":[[-1557.5,-400.00000000000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1612.4999750000013,-472.4999755000001],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"549bec3f-89a4-4854-8eed-2d9171821a2f","orientation":"right","circleData":[[-1587.4999999999998,-490.0000000000002],[-1587.4999999999998,-475.00000000000006],[-1587.4999999999998,-460.00000000000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1612.4999750000004,-712.499975500001],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"1b855ccb-49a4-427a-9563-e1bcdb16e638","orientation":"right","circleData":[[-1587.4999999999995,-730.000000000001],[-1587.4999999999995,-715.0000000000008],[-1587.4999999999995,-700.0000000000008]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1529.064829999999,-744.8506420000008],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"3b6d34de-cd89-4ef4-9473-da4b3ae907df","orientation":"left","circleData":[[-1557.499999999999,-745.0000000000013]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1799.0648299999984,-204.85064200000056],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"dd44450f-fd4f-4059-aab9-565428093e7b","orientation":"left","circleData":[[-1827.4999999999989,-205.00000000000028]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1799.064829999999,125.14935799999944],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"d1e6942e-6a34-4356-87fa-da19b68ae6b8","orientation":"left","circleData":[[-1827.4999999999998,124.99999999999952]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1882.499974999999,-592.4999755000006],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"67df4d37-3f2b-4d48-9904-dc3e640854f2","orientation":"right","circleData":[[-1857.4999999999995,-610.0000000000005],[-1857.4999999999995,-595.0000000000002],[-1857.4999999999995,-580.0000000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1799.0648299999993,-624.8506420000006],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"bb4a8fb4-80b5-4764-a9f6-b3d9cae671c4","orientation":"left","circleData":[[-1827.499999999999,-625.0000000000009]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1799.0648299999984,-504.85064199999965],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"636bd670-72c8-425e-8740-11540fc72a9f","orientation":"left","circleData":[[-1827.4999999999998,-505.00000000000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1882.4999750000002,-367.49997550000035],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"7cf5453a-9a65-47be-a0c1-a40e3c54981e","orientation":"right","circleData":[[-1857.5,-384.99999999999994],[-1857.5,-369.9999999999999],[-1857.5,-354.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1799.0648299999993,-399.8506419999994],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"e84ff89e-b801-43e3-905a-a7004860c743","orientation":"left","circleData":[[-1827.4999999999998,-399.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1882.4999750000004,-472.4999755000001],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"73ff6e4f-35de-4fa1-bb93-81012f621ef2","orientation":"right","circleData":[[-1857.4999999999998,-490.00000000000006],[-1857.4999999999998,-474.99999999999994],[-1857.4999999999998,-459.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1882.499975,-712.4999755000008],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"8fd76732-6e42-40ac-b9ab-aae7428798a1","orientation":"right","circleData":[[-1857.4999999999995,-730.0000000000008],[-1857.4999999999995,-715.0000000000006],[-1857.4999999999995,-700.0000000000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1799.0648299999993,-744.8506420000006],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"edb09e16-b982-4564-8c59-d0c31b14f784","orientation":"left","circleData":[[-1827.499999999999,-745.000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1707.4374994999994,-598.2385495000005],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"eeac935f-c26f-4957-912d-5c92ef07716f","orientation":"right","circleData":[[-1707.5,-625],[-1707.5,-569.2958484999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1722.5625005000006,-456.7614504999999],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"4505b10f-85e5-4973-b4b5-e3d656f3d0be","orientation":"left","circleData":[[-1722.4999999999998,-429.99999999999994],[-1722.4999999999998,-485.70415149999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1722.4374994999994,-388.23854950000054],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"b2e81b6c-d2d3-439c-82a2-c21100e871d6","orientation":"right","circleData":[[-1722.4999999999998,-415.0000000000001],[-1722.4999999999998,-359.29584850000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1722.562500500001,-156.76145049999957],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"88c754f5-de3a-41e9-8e1a-6c44284e3b38","orientation":"left","circleData":[[-1722.4999999999995,-130],[-1722.4999999999995,-185.70415150000005]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1722.4374994999994,-88.23854950000054],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1","orientation":"right","circleData":[[-1722.4999999999995,-115.00000000000018],[-1722.4999999999995,-59.29584850000009]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-372.5,-182.5000000000001],"typeId":"b7d4df28-c430-b8ca-f42b-be40986a361e","componentVersion":1,"instanceId":"11da4e6e-750e-4643-874f-89e7cea28441","orientation":"up","circleData":[[-417.5,-69.99999999999997],[-417.5,-85.00000000000009],[-417.5,-100.00000000000009],[-417.5,-114.99999999999997],[-417.5,-130.00000000000009],[-417.5,-145.00000000000009],[-417.5,-160.00000000000009],[-417.5,-175.00000000000009],[-417.5,-190.0000000000001],[-417.5,-205.0000000000001],[-417.5,-220.0000000000001],[-417.5,-235.0000000000001],[-417.5,-250.00000000000037],[-417.5,-265],[-417.5,-280.0000000000002],[-417.5,-295.0000000000002],[-327.5,-130.00000000000009],[-327.5,-145.00000000000009],[-327.5,-160.00000000000009],[-327.5,-175.00000000000009],[-327.5,-190.0000000000001],[-327.5,-205.0000000000001],[-327.5,-220.0000000000001],[-327.5,-235.0000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1722.562500500001,68.23854949999986],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"0077cc15-4d99-4651-a57e-536f288016fb","orientation":"left","circleData":[[-1722.4999999999995,94.99999999999994],[-1722.4999999999995,39.29584849999989]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1722.4374994999994,136.76145049999923],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"dba2be22-3f32-4819-979e-cd2ac0c4cc6e","orientation":"right","circleData":[[-1722.4999999999995,109.99999999999976],[-1722.4999999999995,165.70415149999982]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1467.4374994999994,-613.2385495000004],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"8281ae65-4ada-4b48-aeec-e666f55d538a","orientation":"right","circleData":[[-1467.5,-639.9999999999999],[-1467.5,-584.2958484999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1087.4999750000002,172.50002449999965],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"f2a03157-3d3b-4891-9a96-ef7378eef59a","orientation":"right","circleData":[[-1062.5,154.9999999999999],[-1062.5,169.99999999999994],[-1062.5,184.99999999999991]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1612.4999749999993,-67.49997550000057],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"a28b7076-045f-481a-8987-e6c379c85461","orientation":"right","circleData":[[-1587.499999999999,-85.00000000000051],[-1587.499999999999,-70.00000000000044],[-1587.499999999999,-55.00000000000044]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1529.0648299999984,-99.85064200000011],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"62a268f0-68fa-4016-91c7-d55a738d6b46","orientation":"left","circleData":[[-1557.4999999999986,-100.00000000000051]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1467.562500500002,-681.7614504999995],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"7a6ab358-5837-431b-9348-a619c0d5eb4b","orientation":"left","circleData":[[-1467.5,-655],[-1467.5,-710.7041515000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1452.562500500001,-456.7614504999998],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"d121ccd5-ebd1-4e31-80c7-213974efb4b7","orientation":"left","circleData":[[-1452.5,-430.00000000000006],[-1452.5,-485.7041515000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1452.4374994999998,-388.2385495000008],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"c51e4057-62bf-4d4d-97d5-80d833dcecd9","orientation":"right","circleData":[[-1452.5,-415.0000000000002],[-1452.5,-359.29584850000015]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1467.562500500001,-156.76145050000036],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"daff2923-49a4-426d-8290-92f3de68e4c8","orientation":"left","circleData":[[-1467.5,-130.00000000000006],[-1467.5,-185.70415150000014]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1467.4374994999994,-88.23854950000054],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9","orientation":"right","circleData":[[-1467.5,-115.00000000000023],[-1467.5,-59.29584850000015]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1452.5625005000009,68.23854949999986],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"c1ec2684-5203-484a-bb58-714d3d1ff689","orientation":"left","circleData":[[-1452.5,94.99999999999999],[-1452.5,39.295848499999956]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1452.4374994999994,136.76145049999946],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"c2e4f40c-d3fa-4534-902a-b6ca784f2d33","orientation":"right","circleData":[[-1452.5,109.99999999999983],[-1452.5,165.7041514999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1197.5625005000009,-666.7614505],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"89080e17-209d-40ef-8155-edbb76fffbef","orientation":"left","circleData":[[-1197.5,-639.9999999999999],[-1197.5,-695.7041514999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1197.4374994999994,-598.2385495000005],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"dbc09422-6bd6-4f89-bf7e-49c71fb62af9","orientation":"right","circleData":[[-1197.5,-625],[-1197.5,-569.2958485]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1529.064829999998,20.149357999999438],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"4732636d-ea0d-4b19-877e-d2ff4ddb5e8d","orientation":"left","circleData":[[-1557.499999999999,19.999999999999147]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1799.064829999998,-99.85064200000033],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"6d57b374-4a97-4f2c-b0da-4d4ccbef4f5a","orientation":"left","circleData":[[-1827.4999999999986,-100.00000000000017]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1799.0648299999987,20.149357999999665],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"0c082f01-0561-48cc-887e-4e37deace687","orientation":"left","circleData":[[-1827.499999999999,19.99999999999949]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1197.562500500001,-441.76145050000014],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"9ab5a6ac-c827-4cf6-9b73-708335a1a9b0","orientation":"left","circleData":[[-1197.5,-415],[-1197.5,-470.7041515]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1197.4374994999994,-373.23854950000054],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"35a17054-5a08-4aee-9aa6-e124f96682e1","orientation":"right","circleData":[[-1197.5,-400.00000000000017],[-1197.5,-344.2958485000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1197.562500500001,-141.76145050000014],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c","orientation":"left","circleData":[[-1197.5,-115],[-1197.5,-170.70415150000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1197.4374994999994,-73.23854950000054],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"0152d242-8b4d-42db-8096-0f8dc98256f3","orientation":"right","circleData":[[-1197.5,-100.00000000000017],[-1197.5,-44.29584850000009]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1197.5625005000009,83.23854950000009],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"35159cb3-cc74-4c90-b0f5-cff583f979a5","orientation":"left","circleData":[[-1197.5,110.00000000000003],[-1197.5,54.295848500000005]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-1197.4374994999994,151.76145049999946],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"2f031f22-1944-43ab-ae9c-f74e47cc4156","orientation":"right","circleData":[[-1197.5,125],[-1197.5,180.7041514999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-942.5625005000006,83.23854949999986],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"625dbf85-54ff-48b2-a275-4089e5081167","orientation":"left","circleData":[[-942.4999999999999,110.00000000000001],[-942.4999999999999,54.29584850000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-942.4374994999991,151.76145049999946],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"f86ac869-5086-4a06-8cd6-49f486548944","orientation":"right","circleData":[[-942.4999999999999,124.99999999999989],[-942.4999999999999,180.70415149999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-927.5625005000013,-141.76145050000002],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"0c68c6e3-0464-4e71-ab6a-9086b01a0e77","orientation":"left","circleData":[[-927.5000000000001,-115.00000000000006],[-927.5000000000001,-170.70415150000008]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-927.4374994999994,-73.23854950000066],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"709ba052-a0a0-4439-a40d-83aedf155550","orientation":"right","circleData":[[-927.5000000000001,-100.00000000000023],[-927.5000000000001,-44.29584850000015]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-927.5625005000009,-441.7614505],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"4b0e618a-0090-4173-a14d-dc77951515d3","orientation":"left","circleData":[[-927.5,-415.00000000000006],[-927.5,-470.7041515000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-927.4374994999994,-373.2385495000008],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"733ac60f-fd5b-4e01-bcd0-44ae417225ee","orientation":"right","circleData":[[-927.5,-400.0000000000003],[-927.5,-344.2958485000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-912.5625005000007,-666.7614505],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"114d5d14-5f5c-40e8-b182-5aaaa19436dd","orientation":"left","circleData":[[-912.5,-640],[-912.5,-695.7041515000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1N4001-TP","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"MCC","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[-912.4374994999996,-598.2385495000005],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"4f53b9c5-5f30-4a72-af1a-a8232ad99f6b","orientation":"right","circleData":[[-912.5,-625.0000000000002],[-912.5,-569.2958485000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-2222.6758564999973,-361.19385550000004],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"621585ad-95ad-4cf3-9a10-1ca969371d4e","orientation":"up","circleData":[[-2292.5,-355.00000000000006],[-2154.3319999999976,-354.0745000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1882.4999749999984,157.5000244999992],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"041b5070-e88a-4a6b-aa2c-a93c5f45650d","orientation":"right","circleData":[[-1857.4999999999986,139.9999999999995],[-1857.4999999999986,154.99999999999955],[-1857.4999999999986,169.9999999999995]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1954.4657915,229.551062],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"995a17d1-5928-497f-b230-e981cff0c0da","orientation":"up","circleData":[[-1977.5,230],[-1932.5,230]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-2207.675856499998,-421.1938554999999],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"efd3f3bc-1ae1-45dd-a482-193032279b23","orientation":"up","circleData":[[-2277.5,-414.99999999999994],[-2139.3319999999985,-414.0745]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1954.4657915000003,-25.448938],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"81ae35b1-5b71-4716-a1af-fd111af3ac03","orientation":"up","circleData":[[-1977.5000000000002,-24.999999999999993],[-1932.5000000000002,-24.999999999999993]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1882.4999749999993,-172.49997550000035],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"46f90c07-7d13-4392-a3bf-e813e3dabb36","orientation":"right","circleData":[[-1857.499999999999,-190.0000000000004],[-1857.499999999999,-175.00000000000023],[-1857.499999999999,-160.00000000000023]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-2221.2502703637383,-486.41782413982327],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"a86bd662-6cba-44a0-8211-7ce5de8f1e54","orientation":"up","circleData":[[-2291.07441386374,-480.2239686398233],[-2152.9064138637377,-479.29846863982334]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1954.4657914999996,-295.44893799999994],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"41446abf-3582-4e1a-bca9-cf131a5fba1c","orientation":"up","circleData":[[-1977.4999999999998,-294.99999999999994],[-1932.4999999999998,-294.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-2207.675856499999,-541.1938555],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"0d024f4d-e2f2-4b76-8f77-420b1168f36c","orientation":"up","circleData":[[-2277.5,-535],[-2139.3319999999994,-534.0745000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1882.4999750000002,52.50002450000011],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"83dcf7d9-214a-4ba8-8c4b-0198867c485d","orientation":"right","circleData":[[-1857.5,34.99999999999999],[-1857.5,50.00000000000016],[-1857.5,65.0000000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1882.4999749999997,-97.49997550000012],"typeId":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"instanceId":"3a88c66b-feb0-48c3-be15-37e3d48518eb","orientation":"right","circleData":[[-1857.5,-115],[-1857.5,-99.99999999999994],[-1857.5,-84.99999999999993]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1547.675856499997,523.8061444999998],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"7807e964-3bc8-4b12-bb6c-44a1c1b24af9","orientation":"up","circleData":[[-1617.5,530],[-1479.3319999999974,530.9254999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1429.4657914999993,529.5510619999998],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"38df7453-f88c-4a99-82c0-fdb338cc7264","orientation":"up","circleData":[[-1452.4999999999995,529.9999999999998],[-1407.4999999999995,529.9999999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1547.6758564999977,448.80614449999985],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"4b269a77-3c6b-4832-bc03-819b3941bca2","orientation":"up","circleData":[[-1617.4999999999998,455],[-1479.331999999998,455.92549999999983]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1429.4657914999993,454.5510619999998],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"ca018356-08f3-4416-b12e-ca10c6c7bb67","orientation":"up","circleData":[[-1452.4999999999995,454.9999999999998],[-1407.4999999999995,454.9999999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1547.6758564999977,373.8061445000001],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"5712632d-8fa8-495b-a104-baf8f43c700a","orientation":"up","circleData":[[-1617.4999999999998,380],[-1479.3319999999972,380.92550000000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1429.4657914999993,379.5510619999998],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"efcea04e-21d8-44a5-8f0d-74277474a2e0","orientation":"up","circleData":[[-1452.4999999999995,379.9999999999998],[-1407.4999999999995,379.9999999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1547.6758564999984,298.80614449999996],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"b69e0669-3879-4abd-9d7d-acc45f8eea74","orientation":"up","circleData":[[-1617.5,305],[-1479.3319999999987,305.92549999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1444.4657914999996,304.55106199999994],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"a8e515ed-cb32-4abf-ab34-4e8ba550aff5","orientation":"up","circleData":[[-1467.4999999999993,304.99999999999994],[-1422.4999999999998,304.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1322.675856499997,-1021.1938555000004],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"c90e906b-172f-43f0-a66d-c99371504fba","orientation":"up","circleData":[[-1392.4999999999998,-1015.0000000000002],[-1254.3319999999974,-1014.0745000000004]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1219.4657914999996,-1015.448938],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"15591579-4d1a-4075-aec4-52c43cc21020","orientation":"up","circleData":[[-1242.4999999999998,-1015],[-1197.4999999999998,-1015]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1322.6758564999977,-1096.1938555000002],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"ee4052d6-2dbe-445a-8b8e-b1c8214d283a","orientation":"up","circleData":[[-1392.5,-1090],[-1254.331999999998,-1089.0745000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1219.4657914999996,-1090.4489380000002],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"c58023a8-eade-4368-93d4-c18f7148e8e3","orientation":"up","circleData":[[-1242.4999999999998,-1090.0000000000002],[-1197.4999999999998,-1090.0000000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1322.6758564999975,-1171.1938554999997],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"ddbc596a-7cd5-4048-bdec-ae929062b39f","orientation":"up","circleData":[[-1392.4999999999998,-1164.9999999999998],[-1254.331999999997,-1164.0744999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1219.4657914999996,-1165.4489380000002],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"e7200013-28f8-4ff6-9dbe-a2239e215492","orientation":"up","circleData":[[-1242.4999999999998,-1165.0000000000002],[-1197.4999999999998,-1165.0000000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1322.6758564999986,-1246.1938555000002],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"0b992200-29a8-47ae-9e2d-5041f24e3da4","orientation":"up","circleData":[[-1392.5,-1240],[-1254.331999999999,-1239.0745000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1234.4657914999998,-1240.448938],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"c107267e-960a-414d-898a-9b8f86844804","orientation":"up","circleData":[[-1257.4999999999995,-1240],[-1212.5,-1240]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-233.67163710292286,451.80051863723395],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"3c883d29-f62b-49cf-a092-2c8c9f097c17","orientation":"up","circleData":[[-303.4957806029257,457.99437413723405],[-165.32778060292313,458.9198741372339]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-115.46157210292509,457.5454361372339],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"f7984d9c-52aa-415e-b39c-e5fb625b93c2","orientation":"up","circleData":[[-138.4957806029253,457.9943741372339],[-93.4957806029253,457.9943741372338]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-233.67163710292354,376.80051863723395],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"c525269a-6029-466e-8297-23d196a50c50","orientation":"up","circleData":[[-303.4957806029255,382.9943741372341],[-165.3277806029238,383.9198741372339]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-115.46157210292509,382.5454361372339],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"c94229bb-b925-4416-b768-559f9d5d84b6","orientation":"up","circleData":[[-138.4957806029253,382.9943741372339],[-93.4957806029253,382.9943741372339]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-233.67163710292354,301.8005186372344],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"42b98079-caa9-47e9-bd5d-65893e0dce4d","orientation":"up","circleData":[[-303.4957806029255,307.99437413723433],[-165.3277806029229,308.9198741372344]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-115.46157210292509,307.545436137234],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"662aa0ec-65ba-4d5d-a487-5ed33ea6d988","orientation":"up","circleData":[[-138.4957806029253,307.99437413723405],[-93.4957806029253,307.99437413723405]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-233.67163710292422,226.80051863723406],"typeId":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"instanceId":"5008935e-c93f-4fb4-a087-0abedc96eefb","orientation":"up","circleData":[[-303.4957806029257,232.9943741372342],[-165.3277806029245,233.91987413723402]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-115.46157210292594,232.5454361372342],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"b45ca744-aa2b-4e0a-b23d-32ff2cca7a14","orientation":"up","circleData":[[-138.4957806029257,232.9943741372342],[-93.49578060292615,232.9943741372342]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-290.44893799999994,-849.6062409999997],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"fe152afb-21b1-47d5-b9c6-bd2b619f0439","orientation":"up","circleData":[[-267.49999999999994,-849.9999999999998],[-312.49999999999994,-849.9999999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-290.44893799999994,-819.606241],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"13bb41c2-0891-49e2-a36d-a0e52211de2b","orientation":"up","circleData":[[-267.49999999999994,-820],[-312.49999999999994,-820]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-290.44893799999994,-789.6062409999997],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"5d50f226-59dc-49dd-a79a-abbf5e3cb510","orientation":"up","circleData":[[-267.49999999999994,-789.9999999999998],[-312.49999999999994,-789.9999999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-290.44893799999994,-759.606241],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"58089c3e-bb30-4b9d-87df-71065baedba4","orientation":"up","circleData":[[-267.49999999999994,-760],[-312.49999999999994,-760]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-410.44893800000006,-849.606241],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"824c2884-8b95-4bf2-9b1d-fc37145bfe37","orientation":"up","circleData":[[-387.50000000000006,-850],[-432.50000000000006,-850]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-410.44893800000006,-819.6062410000002],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00","orientation":"up","circleData":[[-387.50000000000006,-820.0000000000002],[-432.50000000000006,-820.0000000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-410.44893800000006,-789.606241],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"a72804f7-e18d-407a-8183-98f8e53fe3d0","orientation":"up","circleData":[[-387.50000000000006,-790],[-432.50000000000006,-790]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-410.44893800000006,-759.6062410000002],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1","orientation":"up","circleData":[[-387.50000000000006,-760.0000000000002],[-432.50000000000006,-760.0000000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-545.448938,-849.6062409999998],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"07965d4a-3c19-478e-9e88-2147d6a70aba","orientation":"up","circleData":[[-522.5,-849.9999999999999],[-567.4999999999999,-849.9999999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-545.448938,-819.6062410000001],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"b7e27884-48f5-44d6-9ad2-56da1f22ae1e","orientation":"up","circleData":[[-522.5,-820.0000000000001],[-567.4999999999999,-820.0000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-545.448938,-789.6062409999998],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"b68f3984-33e3-4099-9fd0-2bf2992dd7c5","orientation":"up","circleData":[[-522.5,-789.9999999999999],[-567.4999999999999,-789.9999999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-545.448938,-759.6062410000001],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"ed5c99e1-3753-4905-b880-1ffcf976d135","orientation":"up","circleData":[[-522.5,-760.0000000000001],[-567.4999999999999,-760.0000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-665.448938,-849.606241],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf","orientation":"up","circleData":[[-642.5,-850],[-687.5,-850]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-665.448938,-819.6062410000002],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"6b9ac4cf-8b15-40e0-9908-87be89d7dd12","orientation":"up","circleData":[[-642.5,-820.0000000000002],[-687.5,-820.0000000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-665.448938,-789.606241],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88","orientation":"up","circleData":[[-642.5,-790],[-687.5,-790]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-665.448938,-759.6062410000002],"typeId":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"instanceId":"0e24347f-56a1-4fe8-a3eb-00f61ef717e3","orientation":"up","circleData":[[-642.5,-760.0000000000002],[-687.5,-760.0000000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-237.64935799999995,-671.5648299999999],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"2d2c1fc2-9459-4e52-81e7-c39a9a7813f6","orientation":"up","circleData":[[-237.49999999999997,-699.9999999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-222.64935799999992,-56.56483000000006],"typeId":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"instanceId":"935ec2c0-76f9-4c06-a88a-d876d661b1e8","orientation":"up","circleData":[[-222.49999999999994,-85]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"A000066","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Arduino","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[475,-501.25],"typeId":"23db5403-7550-740c-a02b-8b3755757442","componentVersion":1,"instanceId":"9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9","orientation":"right","circleData":[[332.5,-520],[332.5,-505],[332.5,-489.99999999999994],[332.5,-474.99999999999994],[332.5,-459.99999999999994],[332.5,-444.99999999999994],[332.5,-429.99999999999994],[332.5,-414.99999999999994],[332.5,-384.99999999999994],[332.5,-369.99999999999994],[332.5,-354.99999999999994],[332.5,-339.99999999999994],[332.5,-324.99999999999994],[332.5,-309.99999999999994],[617.5,-574],[617.5,-559],[617.5,-544],[617.5,-529],[617.5,-514],[617.5,-498.99999999999994],[617.5,-483.99999999999994],[617.5,-468.99999999999994],[617.5,-453.99999999999994],[617.5,-438.99999999999994],[617.5,-414.99999999999994],[617.5,-399.99999999999994],[617.5,-384.99999999999994],[617.5,-369.99999999999994],[617.5,-354.99999999999994],[617.5,-339.99999999999994],[617.5,-324.99999999999994],[617.5,-309.99999999999994]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"3a131a8a-799f-4763-ae9a-239860e7fa69\",\"explorerHtmlId\":\"ab7cdf34-f697-426a-bfe2-9de296e7f305\",\"nameHtmlId\":\"f6ec2471-315e-4968-b4e9-952a8dc2b7f2\",\"nameInputHtmlId\":\"be67a1a7-2817-4026-8c14-c0f0e76bd489\",\"explorerChildHtmlId\":\"2fd886e0-3231-43ee-8812-0c0debeb79fd\",\"explorerCarrotOpenHtmlId\":\"f0950f6e-4c24-48fd-9562-195c2fc6937a\",\"explorerCarrotClosedHtmlId\":\"cb37000b-415d-4b99-ba9d-acddd9152eca\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"d9103522-dc6c-4fb0-b6f6-8e6df09f7e8f\",\"explorerHtmlId\":\"ad64e1a0-2190-4869-9474-c4b55151bdcc\",\"nameHtmlId\":\"0a48bb7e-9e4d-4adb-9e71-616fc2b801a6\",\"nameInputHtmlId\":\"5abd8455-f67f-40cd-b1ad-8bf710ebb5dd\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"5915c6f4-6b83-4681-ba37-91ff2ff0039a\",\"explorerHtmlId\":\"f4b9b936-dd23-49ec-b392-9273e8c29a69\",\"nameHtmlId\":\"c4019432-91c8-4aa1-9298-c80f002b62c4\",\"nameInputHtmlId\":\"afe10960-a093-453c-8be6-53a66813410b\",\"code\":\"\"},0,","codeLabelPosition":[475,-658.75],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[494.3179315,-99.91661949999997],"typeId":"ea67bc39-2543-48d1-915c-5686eed5bac4","componentVersion":1,"instanceId":"0a8678a1-8b77-47ac-8524-d596b3cedd6d","orientation":"up","circleData":[[542.5,-99.99999999999999],[542.6500000000001,-89.49999999999999],[542.5,-79.59999999999997],[542.95,-68.94999999999996],[542.95,-58.599999999999966],[542.8,-47.79999999999997],[542.05,-27.09999999999998],[542.3499999999999,-38.34999999999998],[439.44999999999993,-99.69999999999997],[439.44999999999993,-89.64999999999996],[439.44999999999993,-79.59999999999997],[439.44999999999993,-69.09999999999997],[439.44999999999993,-58.29999999999997],[439.44999999999993,-48.39999999999996],[439.44999999999993,-37.59999999999998],[439.44999999999993,-26.949999999999974]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[488.4687385,-1050.618421],"typeId":"646c8823-36b2-4192-89ce-6ec44eb47b6e","componentVersion":1,"instanceId":"6fe13b46-5e6b-4103-adfc-cce8f32c36a7","orientation":"up","circleData":[[437.5,-940.0000000000001],[459.99999999999994,-940.0000000000001],[482.49999999999994,-940.0000000000001],[504.99999999999994,-940.0000000000001],[527.5000000000001,-940.0000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-1954.4657915000003,-535.448938],"typeId":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"instanceId":"3694689b-7dc6-49dc-a8fa-3e18614c7e29","orientation":"up","circleData":[[-1977.5,-535],[-1932.5000000000005,-535]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-1278.61541","left":"-2306.50000","width":"2949.00000","height":"1834.84310","x":"-2306.50000","y":"-1278.61541"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#FF74A3\",\"startPinId\":\"pin-type-component_7e9999e8-686e-4f02-b1e7-bee04a417b43_0\",\"endPinId\":\"pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_0\",\"rawStartPinId\":\"pin-type-component_7e9999e8-686e-4f02-b1e7-bee04a417b43_0\",\"rawEndPinId\":\"pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1032.5000000000_-190.0000000000\\\",\\\"-1047.5000000000_-190.0000000000\\\",\\\"-1047.5000000000_-175.0000000000\\\",\\\"-1062.5000000000_-175.0000000000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_0\",\"endPinId\":\"pin-type-component_4bfdc0b0-0087-4f19-b9da-fe77fe2030bb_0\",\"rawStartPinId\":\"pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_0\",\"rawEndPinId\":\"pin-type-component_4bfdc0b0-0087-4f19-b9da-fe77fe2030bb_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-70.0000000000\\\",\\\"-1047.5000000000_-70.0000000000\\\",\\\"-1047.5000000000_-85.0000000000\\\",\\\"-1032.5000000000_-85.0000000000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_0\",\"endPinId\":\"pin-type-component_725c2e06-513a-456a-a054-9a1efd2410b5_0\",\"rawStartPinId\":\"pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_0\",\"rawEndPinId\":\"pin-type-component_725c2e06-513a-456a-a054-9a1efd2410b5_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_50.0000000000\\\",\\\"-1047.5000000000_50.0000000000\\\",\\\"-1047.5000000000_35.0000000000\\\",\\\"-1032.5000000000_35.0000000000\\\"]}\"}","{\"color\":\"#BDC6FF\",\"startPinId\":\"pin-type-component_84e67de5-59f5-4375-8901-060561a64dc9_0\",\"endPinId\":\"pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_0\",\"rawStartPinId\":\"pin-type-component_84e67de5-59f5-4375-8901-060561a64dc9_0\",\"rawEndPinId\":\"pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1032.5000000000_140.0000000000\\\",\\\"-1047.5000000000_140.0000000000\\\",\\\"-1047.5000000000_155.0000000000\\\",\\\"-1062.5000000000_155.0000000000\\\"]}\"}","{\"color\":\"#A5FFD2\",\"startPinId\":\"pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_0\",\"endPinId\":\"pin-type-component_a4a81ac1-f999-4c5f-bf1d-d39d1364ba7e_0\",\"rawStartPinId\":\"pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_0\",\"rawEndPinId\":\"pin-type-component_a4a81ac1-f999-4c5f-bf1d-d39d1364ba7e_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-370.0000000000\\\",\\\"-1047.5000000000_-370.0000000000\\\",\\\"-1047.5000000000_-385.0000000000\\\",\\\"-1032.5000000000_-385.0000000000\\\"]}\"}","{\"color\":\"#774D00\",\"startPinId\":\"pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_0\",\"endPinId\":\"pin-type-component_84525e3e-ef29-4e0c-a293-959707966b26_0\",\"rawStartPinId\":\"pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_0\",\"rawEndPinId\":\"pin-type-component_84525e3e-ef29-4e0c-a293-959707966b26_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-475.0000000000\\\",\\\"-1047.5000000000_-475.0000000000\\\",\\\"-1047.5000000000_-490.0000000000\\\",\\\"-1032.5000000000_-490.0000000000\\\"]}\"}","{\"color\":\"#004754\",\"startPinId\":\"pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_0\",\"endPinId\":\"pin-type-component_ad7b12e6-293b-4cf0-b5fc-2ad4811766ad_0\",\"rawStartPinId\":\"pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_0\",\"rawEndPinId\":\"pin-type-component_ad7b12e6-293b-4cf0-b5fc-2ad4811766ad_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-595.0000000000\\\",\\\"-1047.5000000000_-595.0000000000\\\",\\\"-1047.5000000000_-610.0000000000\\\",\\\"-1032.5000000000_-610.0000000000\\\"]}\"}","{\"color\":\"#90FB92\",\"startPinId\":\"pin-type-component_69b6c16b-f2c6-4ab0-b694-b43efd7d7efa_0\",\"endPinId\":\"pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_0\",\"rawStartPinId\":\"pin-type-component_69b6c16b-f2c6-4ab0-b694-b43efd7d7efa_0\",\"rawEndPinId\":\"pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1032.5000000000_-730.0000000000\\\",\\\"-1047.5000000000_-730.0000000000\\\",\\\"-1047.5000000000_-715.0000000000\\\",\\\"-1062.5000000000_-715.0000000000\\\"]}\"}","{\"color\":\"#BDD393\",\"startPinId\":\"pin-type-component_5278fc75-d95d-4e4c-a86e-2e83a862e607_0\",\"endPinId\":\"pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_0\",\"rawStartPinId\":\"pin-type-component_5278fc75-d95d-4e4c-a86e-2e83a862e607_0\",\"rawEndPinId\":\"pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1302.5000000000_140.0000000000\\\",\\\"-1317.5000000000_140.0000000000\\\",\\\"-1317.5000000000_155.0000000000\\\",\\\"-1332.5000000000_155.0000000000\\\"]}\"}","{\"color\":\"#00FF78\",\"startPinId\":\"pin-type-component_0af45fa8-24bc-42e4-9c24-d15187e9fbc3_0\",\"endPinId\":\"pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_0\",\"rawStartPinId\":\"pin-type-component_0af45fa8-24bc-42e4-9c24-d15187e9fbc3_0\",\"rawEndPinId\":\"pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1302.5000000000_35.0000000000\\\",\\\"-1317.5000000000_35.0000000000\\\",\\\"-1317.5000000000_50.0000000000\\\",\\\"-1332.5000000000_50.0000000000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_266aa6bb-5bae-4ff3-85db-bbd370178ae8_0\",\"endPinId\":\"pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_0\",\"rawStartPinId\":\"pin-type-component_266aa6bb-5bae-4ff3-85db-bbd370178ae8_0\",\"rawEndPinId\":\"pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1302.5000000000_-85.0000000000\\\",\\\"-1317.5000000000_-85.0000000000\\\",\\\"-1317.5000000000_-70.0000000000\\\",\\\"-1332.5000000000_-70.0000000000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_7fc8671b-e701-4c33-a644-f42eace24307_0\",\"endPinId\":\"pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_0\",\"rawStartPinId\":\"pin-type-component_7fc8671b-e701-4c33-a644-f42eace24307_0\",\"rawEndPinId\":\"pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1302.5000000000_-190.0000000000\\\",\\\"-1317.5000000000_-190.0000000000\\\",\\\"-1317.5000000000_-175.0000000000\\\",\\\"-1332.5000000000_-175.0000000000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_34445add-d974-48d4-81af-972f5dd7934b_0\",\"endPinId\":\"pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_0\",\"rawStartPinId\":\"pin-type-component_34445add-d974-48d4-81af-972f5dd7934b_0\",\"rawEndPinId\":\"pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1302.5000000000_-385.0000000000\\\",\\\"-1317.5000000000_-385.0000000000\\\",\\\"-1317.5000000000_-370.0000000000\\\",\\\"-1332.5000000000_-370.0000000000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_0\",\"endPinId\":\"pin-type-component_3d109b51-1504-4d24-a9e7-9e3fe3074724_0\",\"rawStartPinId\":\"pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_0\",\"rawEndPinId\":\"pin-type-component_3d109b51-1504-4d24-a9e7-9e3fe3074724_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1332.5000000000_-475.0000000000\\\",\\\"-1317.5000000000_-475.0000000000\\\",\\\"-1317.5000000000_-490.0000000000\\\",\\\"-1302.5000000000_-490.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_0\",\"endPinId\":\"pin-type-component_e7d36833-6d1a-490c-96e9-4f178d942f47_0\",\"rawStartPinId\":\"pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_0\",\"rawEndPinId\":\"pin-type-component_e7d36833-6d1a-490c-96e9-4f178d942f47_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1332.5000000000_-595.0000000000\\\",\\\"-1317.5000000000_-595.0000000000\\\",\\\"-1317.5000000000_-610.0000000000\\\",\\\"-1302.5000000000_-610.0000000000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_0\",\"endPinId\":\"pin-type-component_903934ae-30da-4a37-93c9-c64660e9c617_0\",\"rawStartPinId\":\"pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_0\",\"rawEndPinId\":\"pin-type-component_903934ae-30da-4a37-93c9-c64660e9c617_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1332.5000000000_-715.0000000000\\\",\\\"-1317.5000000000_-715.0000000000\\\",\\\"-1317.5000000000_-730.0000000000\\\",\\\"-1302.5000000000_-730.0000000000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_0\",\"endPinId\":\"pin-type-component_7f294ee1-7ea8-4e70-bb0a-8c8b6b15b6c9_0\",\"rawStartPinId\":\"pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_0\",\"rawEndPinId\":\"pin-type-component_7f294ee1-7ea8-4e70-bb0a-8c8b6b15b6c9_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_140.0000000000\\\",\\\"-1572.5000000000_140.0000000000\\\",\\\"-1572.5000000000_125.0000000000\\\",\\\"-1557.5000000000_125.0000000000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_0\",\"endPinId\":\"pin-type-component_4732636d-ea0d-4b19-877e-d2ff4ddb5e8d_0\",\"rawStartPinId\":\"pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_0\",\"rawEndPinId\":\"pin-type-component_4732636d-ea0d-4b19-877e-d2ff4ddb5e8d_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_35.0000000000\\\",\\\"-1572.5000000000_35.0000000000\\\",\\\"-1572.5000000000_20.0000000000\\\",\\\"-1557.5000000000_20.0000000000\\\"]}\"}","{\"color\":\"#C28C9F\",\"startPinId\":\"pin-type-component_62a268f0-68fa-4016-91c7-d55a738d6b46_0\",\"endPinId\":\"pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_0\",\"rawStartPinId\":\"pin-type-component_62a268f0-68fa-4016-91c7-d55a738d6b46_0\",\"rawEndPinId\":\"pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1557.5000000000_-100.0000000000\\\",\\\"-1572.5000000000_-100.0000000000\\\",\\\"-1572.5000000000_-85.0000000000\\\",\\\"-1587.5000000000_-85.0000000000\\\"]}\"}","{\"color\":\"#5FAD4E\",\"startPinId\":\"pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_0\",\"endPinId\":\"pin-type-component_5bdd54e6-172a-4994-8b34-5d8687be61e2_0\",\"rawStartPinId\":\"pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_0\",\"rawEndPinId\":\"pin-type-component_5bdd54e6-172a-4994-8b34-5d8687be61e2_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_-190.0000000000\\\",\\\"-1572.5000000000_-190.0000000000\\\",\\\"-1572.5000000000_-205.0000000000\\\",\\\"-1557.5000000000_-205.0000000000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-component_29f2dcbd-c66e-4d22-9415-91c6505cd16b_0\",\"endPinId\":\"pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_0\",\"rawStartPinId\":\"pin-type-component_29f2dcbd-c66e-4d22-9415-91c6505cd16b_0\",\"rawEndPinId\":\"pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1557.5000000000_-400.0000000000\\\",\\\"-1572.5000000000_-400.0000000000\\\",\\\"-1572.5000000000_-385.0000000000\\\",\\\"-1587.5000000000_-385.0000000000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_0\",\"endPinId\":\"pin-type-component_d1e6942e-6a34-4356-87fa-da19b68ae6b8_0\",\"rawStartPinId\":\"pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_0\",\"rawEndPinId\":\"pin-type-component_d1e6942e-6a34-4356-87fa-da19b68ae6b8_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_140.0000000000\\\",\\\"-1842.5000000000_140.0000000000\\\",\\\"-1842.5000000000_125.0000000000\\\",\\\"-1827.5000000000_125.0000000000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-component_0c082f01-0561-48cc-887e-4e37deace687_0\",\"endPinId\":\"pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_0\",\"rawStartPinId\":\"pin-type-component_0c082f01-0561-48cc-887e-4e37deace687_0\",\"rawEndPinId\":\"pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1827.5000000000_20.0000000000\\\",\\\"-1857.5000000000_20.0000000000\\\",\\\"-1857.5000000000_35.0000000000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_0\",\"endPinId\":\"pin-type-component_6d57b374-4a97-4f2c-b0da-4d4ccbef4f5a_0\",\"rawStartPinId\":\"pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_0\",\"rawEndPinId\":\"pin-type-component_6d57b374-4a97-4f2c-b0da-4d4ccbef4f5a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_-115.0000000000\\\",\\\"-1842.5000000000_-115.0000000000\\\",\\\"-1842.5000000000_-100.0000000000\\\",\\\"-1827.5000000000_-100.0000000000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_0\",\"endPinId\":\"pin-type-component_dd44450f-fd4f-4059-aab9-565428093e7b_0\",\"rawStartPinId\":\"pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_0\",\"rawEndPinId\":\"pin-type-component_dd44450f-fd4f-4059-aab9-565428093e7b_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_-190.0000000000\\\",\\\"-1842.5000000000_-190.0000000000\\\",\\\"-1842.5000000000_-205.0000000000\\\",\\\"-1827.5000000000_-205.0000000000\\\"]}\"}","{\"color\":\"#A5FFD2\",\"startPinId\":\"pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_0\",\"endPinId\":\"pin-type-component_e84ff89e-b801-43e3-905a-a7004860c743_0\",\"rawStartPinId\":\"pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_0\",\"rawEndPinId\":\"pin-type-component_e84ff89e-b801-43e3-905a-a7004860c743_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_-385.0000000000\\\",\\\"-1842.5000000000_-385.0000000000\\\",\\\"-1842.5000000000_-400.0000000000\\\",\\\"-1827.5000000000_-400.0000000000\\\"]}\"}","{\"color\":\"#774D00\",\"startPinId\":\"pin-type-component_636bd670-72c8-425e-8740-11540fc72a9f_0\",\"endPinId\":\"pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_0\",\"rawStartPinId\":\"pin-type-component_636bd670-72c8-425e-8740-11540fc72a9f_0\",\"rawEndPinId\":\"pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1827.5000000000_-505.0000000000\\\",\\\"-1842.5000000000_-505.0000000000\\\",\\\"-1842.5000000000_-490.0000000000\\\",\\\"-1857.5000000000_-490.0000000000\\\"]}\"}","{\"color\":\"#004754\",\"startPinId\":\"pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_0\",\"endPinId\":\"pin-type-component_bb4a8fb4-80b5-4764-a9f6-b3d9cae671c4_0\",\"rawStartPinId\":\"pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_0\",\"rawEndPinId\":\"pin-type-component_bb4a8fb4-80b5-4764-a9f6-b3d9cae671c4_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_-610.0000000000\\\",\\\"-1842.5000000000_-610.0000000000\\\",\\\"-1842.5000000000_-625.0000000000\\\",\\\"-1827.5000000000_-625.0000000000\\\"]}\"}","{\"color\":\"#66ffa8\",\"startPinId\":\"pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_0\",\"endPinId\":\"pin-type-component_edb09e16-b982-4564-8c59-d0c31b14f784_0\",\"rawStartPinId\":\"pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_0\",\"rawEndPinId\":\"pin-type-component_edb09e16-b982-4564-8c59-d0c31b14f784_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_-730.0000000000\\\",\\\"-1842.5000000000_-730.0000000000\\\",\\\"-1842.5000000000_-745.0000000000\\\",\\\"-1827.5000000000_-745.0000000000\\\"]}\"}","{\"color\":\"#90FB92\",\"startPinId\":\"pin-type-component_0b4ba5d8-bcb4-4816-8dfe-3fa4ce9ed019_0\",\"endPinId\":\"pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_0\",\"rawStartPinId\":\"pin-type-component_0b4ba5d8-bcb4-4816-8dfe-3fa4ce9ed019_0\",\"rawEndPinId\":\"pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1557.5000000000_-505.0000000000\\\",\\\"-1572.5000000000_-505.0000000000\\\",\\\"-1572.5000000000_-490.0000000000\\\",\\\"-1587.5000000000_-490.0000000000\\\"]}\"}","{\"color\":\"#BDD393\",\"startPinId\":\"pin-type-component_b2f3a979-ce1b-444a-a7e4-6ef67b25f077_0\",\"endPinId\":\"pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_0\",\"rawStartPinId\":\"pin-type-component_b2f3a979-ce1b-444a-a7e4-6ef67b25f077_0\",\"rawEndPinId\":\"pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1557.5000000000_-625.0000000000\\\",\\\"-1572.5000000000_-625.0000000000\\\",\\\"-1572.5000000000_-610.0000000000\\\",\\\"-1587.5000000000_-610.0000000000\\\"]}\"}","{\"color\":\"#00FF78\",\"startPinId\":\"pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_0\",\"endPinId\":\"pin-type-component_3b6d34de-cd89-4ef4-9473-da4b3ae907df_0\",\"rawStartPinId\":\"pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_0\",\"rawEndPinId\":\"pin-type-component_3b6d34de-cd89-4ef4-9473-da4b3ae907df_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_-730.0000000000\\\",\\\"-1572.5000000000_-730.0000000000\\\",\\\"-1572.5000000000_-745.0000000000\\\",\\\"-1557.5000000000_-745.0000000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_1\",\"endPinId\":\"pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_1\",\"rawStartPinId\":\"pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_1\",\"rawEndPinId\":\"pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1707.5000000000_-695.7041515000\\\",\\\"-1707.5000000000_-715.0000000000\\\",\\\"-1857.5000000000_-715.0000000000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1\",\"endPinId\":\"pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1\",\"rawStartPinId\":\"pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_1\",\"rawEndPinId\":\"pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_-595.0000000000\\\",\\\"-1730.0000000000_-595.0000000000\\\",\\\"-1730.0000000000_-569.2958485000\\\",\\\"-1707.5000000000_-569.2958485000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0\",\"endPinId\":\"pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0\",\"rawStartPinId\":\"pin-type-component_082451f0-7869-4209-aa80-c752e3204afe_0\",\"rawEndPinId\":\"pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1707.5000000000_-640.0000000000\\\",\\\"-1707.5000000000_-625.0000000000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15\",\"endPinId\":\"pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0\",\"rawStartPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15\",\"rawEndPinId\":\"pin-type-component_eeac935f-c26f-4957-912d-5c92ef07716f_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-685.0000000000\\\",\\\"-747.5000000000_-685.0000000000\\\",\\\"-747.5000000000_-857.5000000000\\\",\\\"-1692.5000000000_-857.5000000000\\\",\\\"-1692.5000000000_-625.0000000000\\\",\\\"-1707.5000000000_-625.0000000000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15\",\"rawStartPinId\":\"pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_15\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-687.5000000000_-760.0000000000\\\",\\\"-687.5000000000_-685.0000000000\\\",\\\"-417.5000000000_-685.0000000000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_1\",\"endPinId\":\"pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_1\",\"rawStartPinId\":\"pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_1\",\"rawEndPinId\":\"pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1722.5000000000_-485.7041515000\\\",\\\"-1722.5000000000_-490.0000000000\\\",\\\"-1752.5000000000_-490.0000000000\\\",\\\"-1752.5000000000_-475.0000000000\\\",\\\"-1857.5000000000_-475.0000000000\\\"]}\"}","{\"color\":\"#00ff88\",\"startPinId\":\"pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1\",\"endPinId\":\"pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1\",\"rawStartPinId\":\"pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_1\",\"rawEndPinId\":\"pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_-370.0000000000\\\",\\\"-1745.0000000000_-370.0000000000\\\",\\\"-1745.0000000000_-355.0000000000\\\",\\\"-1722.5000000000_-355.0000000000\\\",\\\"-1722.5000000000_-359.2958485000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0\",\"endPinId\":\"pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_0\",\"rawStartPinId\":\"pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0\",\"rawEndPinId\":\"pin-type-component_b2e81b6c-d2d3-439c-82a2-c21100e871d6_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1722.5000000000_-430.0000000000\\\",\\\"-1722.5000000000_-415.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14\",\"rawStartPinId\":\"pin-type-component_4505b10f-85e5-4973-b4b5-e3d656f3d0be_0\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1722.5000000000_-430.0000000000\\\",\\\"-1722.5000000000_-415.0000000000\\\",\\\"-1677.5000000000_-415.0000000000\\\",\\\"-1677.5000000000_-835.0000000000\\\",\\\"-770.0000000000_-835.0000000000\\\",\\\"-770.0000000000_-670.0000000000\\\",\\\"-417.5000000000_-670.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14\",\"rawStartPinId\":\"pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_14\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-687.5000000000_-790.0000000000\\\",\\\"-695.0000000000_-790.0000000000\\\",\\\"-695.0000000000_-670.0000000000\\\",\\\"-417.5000000000_-670.0000000000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_1\",\"endPinId\":\"pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_1\",\"rawStartPinId\":\"pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_1\",\"rawEndPinId\":\"pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_-175.0000000000\\\",\\\"-1737.5000000000_-175.0000000000\\\",\\\"-1737.5000000000_-197.5000000000\\\",\\\"-1722.5000000000_-197.5000000000\\\",\\\"-1722.5000000000_-185.7041515000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_1\",\"endPinId\":\"pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_1\",\"rawStartPinId\":\"pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_1\",\"rawEndPinId\":\"pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_-100.0000000000\\\",\\\"-1737.5000000000_-100.0000000000\\\",\\\"-1737.5000000000_-40.0000000000\\\",\\\"-1722.5000000000_-40.0000000000\\\",\\\"-1722.5000000000_-59.2958485000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0\",\"endPinId\":\"pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_0\",\"rawStartPinId\":\"pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0\",\"rawEndPinId\":\"pin-type-component_ad0770a6-65b9-4ba6-ae56-ecc5dd50d5a1_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1722.5000000000_-130.0000000000\\\",\\\"-1722.5000000000_-115.0000000000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13\",\"rawStartPinId\":\"pin-type-component_88c754f5-de3a-41e9-8e1a-6c44284e3b38_0\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1722.5000000000_-130.0000000000\\\",\\\"-1722.5000000000_-160.0000000000\\\",\\\"-1662.5000000000_-160.0000000000\\\",\\\"-1662.5000000000_-805.0000000000\\\",\\\"-792.5000000000_-805.0000000000\\\",\\\"-792.5000000000_-655.0000000000\\\",\\\"-417.5000000000_-655.0000000000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13\",\"rawStartPinId\":\"pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_13\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-687.5000000000_-820.0000000000\\\",\\\"-702.5000000000_-820.0000000000\\\",\\\"-702.5000000000_-655.0000000000\\\",\\\"-417.5000000000_-655.0000000000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_1\",\"endPinId\":\"pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_1\",\"rawStartPinId\":\"pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_1\",\"rawEndPinId\":\"pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_155.0000000000\\\",\\\"-1745.0000000000_155.0000000000\\\",\\\"-1745.0000000000_170.0000000000\\\",\\\"-1722.5000000000_170.0000000000\\\",\\\"-1722.5000000000_165.7041515000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_1\",\"endPinId\":\"pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_1\",\"rawStartPinId\":\"pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_1\",\"rawEndPinId\":\"pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1722.5000000000_39.2958485000\\\",\\\"-1722.5000000000_27.5000000000\\\",\\\"-1745.0000000000_27.5000000000\\\",\\\"-1745.0000000000_50.0000000000\\\",\\\"-1857.5000000000_50.0000000000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_0\",\"endPinId\":\"pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0\",\"rawStartPinId\":\"pin-type-component_0077cc15-4d99-4651-a57e-536f288016fb_0\",\"rawEndPinId\":\"pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1722.5000000000_95.0000000000\\\",\\\"-1722.5000000000_110.0000000000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12\",\"endPinId\":\"pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0\",\"rawStartPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12\",\"rawEndPinId\":\"pin-type-component_dba2be22-3f32-4819-979e-cd2ac0c4cc6e_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-640.0000000000\\\",\\\"-807.5000000000_-640.0000000000\\\",\\\"-807.5000000000_-782.5000000000\\\",\\\"-1647.5000000000_-782.5000000000\\\",\\\"-1647.5000000000_110.0000000000\\\",\\\"-1722.5000000000_110.0000000000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12\",\"rawStartPinId\":\"pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_12\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-687.5000000000_-850.0000000000\\\",\\\"-710.0000000000_-850.0000000000\\\",\\\"-710.0000000000_-640.0000000000\\\",\\\"-417.5000000000_-640.0000000000\\\"]}\"}","{\"color\":\"#00AE7E\",\"startPinId\":\"pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_1\",\"endPinId\":\"pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_1\",\"rawStartPinId\":\"pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_1\",\"rawEndPinId\":\"pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_-715.0000000000\\\",\\\"-1467.5000000000_-715.0000000000\\\",\\\"-1467.5000000000_-710.7041515000\\\"]}\"}","{\"color\":\"#C28C9F\",\"startPinId\":\"pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_1\",\"endPinId\":\"pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_1\",\"rawStartPinId\":\"pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_1\",\"rawEndPinId\":\"pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1467.5000000000_-584.2958485000\\\",\\\"-1467.5000000000_-580.0000000000\\\",\\\"-1490.0000000000_-580.0000000000\\\",\\\"-1490.0000000000_-595.0000000000\\\",\\\"-1587.5000000000_-595.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_0\",\"endPinId\":\"pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0\",\"rawStartPinId\":\"pin-type-component_7a6ab358-5837-431b-9348-a619c0d5eb4b_0\",\"rawEndPinId\":\"pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1467.5000000000_-655.0000000000\\\",\\\"-1467.5000000000_-640.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11\",\"rawStartPinId\":\"pin-type-component_8281ae65-4ada-4b48-aeec-e666f55d538a_0\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1467.5000000000_-640.0000000000\\\",\\\"-1400.0000000000_-640.0000000000\\\",\\\"-1400.0000000000_-302.5000000000\\\",\\\"-822.5000000000_-302.5000000000\\\",\\\"-822.5000000000_-625.0000000000\\\",\\\"-417.5000000000_-625.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11\",\"endPinId\":\"pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_1\",\"rawStartPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_11\",\"rawEndPinId\":\"pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-625.0000000000\\\",\\\"-567.5000000000_-625.0000000000\\\",\\\"-567.5000000000_-760.0000000000\\\"]}\"}","{\"color\":\"#5FAD4E\",\"startPinId\":\"pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_1\",\"endPinId\":\"pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_1\",\"rawStartPinId\":\"pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_1\",\"rawEndPinId\":\"pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_-475.0000000000\\\",\\\"-1482.5000000000_-475.0000000000\\\",\\\"-1482.5000000000_-497.5000000000\\\",\\\"-1452.5000000000_-497.5000000000\\\",\\\"-1452.5000000000_-485.7041515000\\\"]}\"}","{\"color\":\"#FF029D\",\"startPinId\":\"pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_1\",\"endPinId\":\"pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_1\",\"rawStartPinId\":\"pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_1\",\"rawEndPinId\":\"pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_-370.0000000000\\\",\\\"-1475.0000000000_-370.0000000000\\\",\\\"-1475.0000000000_-340.0000000000\\\",\\\"-1452.5000000000_-340.0000000000\\\",\\\"-1452.5000000000_-359.2958485000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0\",\"endPinId\":\"pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_0\",\"rawStartPinId\":\"pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0\",\"rawEndPinId\":\"pin-type-component_d121ccd5-ebd1-4e31-80c7-213974efb4b7_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1452.5000000000_-415.0000000000\\\",\\\"-1452.5000000000_-430.0000000000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10\",\"rawStartPinId\":\"pin-type-component_c51e4057-62bf-4d4d-97d5-80d833dcecd9_0\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1452.5000000000_-415.0000000000\\\",\\\"-1415.0000000000_-415.0000000000\\\",\\\"-1415.0000000000_-295.0000000000\\\",\\\"-807.5000000000_-295.0000000000\\\",\\\"-807.5000000000_-610.0000000000\\\",\\\"-417.5000000000_-610.0000000000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10\",\"rawStartPinId\":\"pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_10\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-567.5000000000_-790.0000000000\\\",\\\"-575.0000000000_-790.0000000000\\\",\\\"-575.0000000000_-610.0000000000\\\",\\\"-417.5000000000_-610.0000000000\\\"]}\"}","{\"color\":\"#FF74A3\",\"startPinId\":\"pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_1\",\"endPinId\":\"pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_1\",\"rawStartPinId\":\"pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_1\",\"rawEndPinId\":\"pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_-175.0000000000\\\",\\\"-1482.5000000000_-175.0000000000\\\",\\\"-1482.5000000000_-190.0000000000\\\",\\\"-1467.5000000000_-190.0000000000\\\",\\\"-1467.5000000000_-185.7041515000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_1\",\"endPinId\":\"pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_1\",\"rawStartPinId\":\"pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_1\",\"rawEndPinId\":\"pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_-70.0000000000\\\",\\\"-1482.5000000000_-70.0000000000\\\",\\\"-1482.5000000000_-62.5000000000\\\",\\\"-1467.5000000000_-62.5000000000\\\",\\\"-1467.5000000000_-59.2958485000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_0\",\"endPinId\":\"pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0\",\"rawStartPinId\":\"pin-type-component_daff2923-49a4-426d-8290-92f3de68e4c8_0\",\"rawEndPinId\":\"pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1467.5000000000_-130.0000000000\\\",\\\"-1467.5000000000_-115.0000000000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9\",\"endPinId\":\"pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0\",\"rawStartPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9\",\"rawEndPinId\":\"pin-type-component_e16687ab-42e5-4e99-9d84-e9c8ffa4d6e9_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-595.0000000000\\\",\\\"-792.5000000000_-595.0000000000\\\",\\\"-792.5000000000_-287.5000000000\\\",\\\"-1415.0000000000_-287.5000000000\\\",\\\"-1415.0000000000_-115.0000000000\\\",\\\"-1467.5000000000_-115.0000000000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9\",\"rawStartPinId\":\"pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-567.5000000000_-820.0000000000\\\",\\\"-582.5000000000_-820.0000000000\\\",\\\"-582.5000000000_-595.0000000000\\\",\\\"-417.5000000000_-595.0000000000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_1\",\"endPinId\":\"pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_1\",\"rawStartPinId\":\"pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_1\",\"rawEndPinId\":\"pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_50.0000000000\\\",\\\"-1475.0000000000_50.0000000000\\\",\\\"-1475.0000000000_27.5000000000\\\",\\\"-1452.5000000000_27.5000000000\\\",\\\"-1452.5000000000_39.2958485000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_1\",\"endPinId\":\"pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_1\",\"rawStartPinId\":\"pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_1\",\"rawEndPinId\":\"pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_155.0000000000\\\",\\\"-1475.0000000000_155.0000000000\\\",\\\"-1475.0000000000_177.5000000000\\\",\\\"-1452.5000000000_177.5000000000\\\",\\\"-1452.5000000000_165.7041515000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_0\",\"endPinId\":\"pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0\",\"rawStartPinId\":\"pin-type-component_c1ec2684-5203-484a-bb58-714d3d1ff689_0\",\"rawEndPinId\":\"pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1452.5000000000_95.0000000000\\\",\\\"-1452.5000000000_110.0000000000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8\",\"rawStartPinId\":\"pin-type-component_c2e4f40c-d3fa-4534-902a-b6ca784f2d33_0\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1452.5000000000_110.0000000000\\\",\\\"-1400.0000000000_110.0000000000\\\",\\\"-1400.0000000000_-280.0000000000\\\",\\\"-777.5000000000_-280.0000000000\\\",\\\"-777.5000000000_-580.0000000000\\\",\\\"-417.5000000000_-580.0000000000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8\",\"rawStartPinId\":\"pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_8\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-567.5000000000_-850.0000000000\\\",\\\"-590.0000000000_-850.0000000000\\\",\\\"-590.0000000000_-580.0000000000\\\",\\\"-417.5000000000_-580.0000000000\\\"]}\"}","{\"color\":\"#BDC6FF\",\"startPinId\":\"pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_1\",\"endPinId\":\"pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_1\",\"rawStartPinId\":\"pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_1\",\"rawEndPinId\":\"pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_-695.7041515000\\\",\\\"-1197.5000000000_-700.0000000000\\\",\\\"-1332.5000000000_-700.0000000000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_1\",\"endPinId\":\"pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_1\",\"rawStartPinId\":\"pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_1\",\"rawEndPinId\":\"pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1332.5000000000_-580.0000000000\\\",\\\"-1212.5000000000_-580.0000000000\\\",\\\"-1212.5000000000_-550.0000000000\\\",\\\"-1197.5000000000_-550.0000000000\\\",\\\"-1197.5000000000_-569.2958485000\\\"]}\"}","{\"color\":\"#7544B1\",\"startPinId\":\"pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_0\",\"endPinId\":\"pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0\",\"rawStartPinId\":\"pin-type-component_89080e17-209d-40ef-8155-edbb76fffbef_0\",\"rawEndPinId\":\"pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_-640.0000000000\\\",\\\"-1197.5000000000_-625.0000000000\\\"]}\"}","{\"color\":\"#7544B1\",\"startPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7\",\"endPinId\":\"pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0\",\"rawStartPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7\",\"rawEndPinId\":\"pin-type-component_dbc09422-6bd6-4f89-bf7e-49c71fb62af9_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-565.0000000000\\\",\\\"-762.5000000000_-565.0000000000\\\",\\\"-762.5000000000_-265.0000000000\\\",\\\"-1160.0000000000_-265.0000000000\\\",\\\"-1160.0000000000_-625.0000000000\\\",\\\"-1197.5000000000_-625.0000000000\\\"]}\"}","{\"color\":\"#7544B1\",\"startPinId\":\"pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7\",\"rawStartPinId\":\"pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-432.5000000000_-760.0000000000\\\",\\\"-462.5000000000_-760.0000000000\\\",\\\"-462.5000000000_-565.0000000000\\\",\\\"-417.5000000000_-565.0000000000\\\"]}\"}","{\"color\":\"#A5FFD2\",\"startPinId\":\"pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_1\",\"endPinId\":\"pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_1\",\"rawStartPinId\":\"pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_1\",\"rawEndPinId\":\"pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1332.5000000000_-460.0000000000\\\",\\\"-1197.5000000000_-460.0000000000\\\",\\\"-1197.5000000000_-470.7041515000\\\"]}\"}","{\"color\":\"#FFA6FE\",\"startPinId\":\"pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_1\",\"endPinId\":\"pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_1\",\"rawStartPinId\":\"pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_1\",\"rawEndPinId\":\"pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_-344.2958485000\\\",\\\"-1197.5000000000_-340.0000000000\\\",\\\"-1220.0000000000_-340.0000000000\\\",\\\"-1220.0000000000_-355.0000000000\\\",\\\"-1332.5000000000_-355.0000000000\\\"]}\"}","{\"color\":\"#774D00\",\"startPinId\":\"pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_0\",\"endPinId\":\"pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0\",\"rawStartPinId\":\"pin-type-component_35a17054-5a08-4aee-9aa6-e124f96682e1_0\",\"rawEndPinId\":\"pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_-400.0000000000\\\",\\\"-1197.5000000000_-415.0000000000\\\"]}\"}","{\"color\":\"#774D00\",\"startPinId\":\"pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6\",\"rawStartPinId\":\"pin-type-component_9ab5a6ac-c827-4cf6-9b73-708335a1a9b0_0\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_-415.0000000000\\\",\\\"-1197.5000000000_-400.0000000000\\\",\\\"-1175.0000000000_-400.0000000000\\\",\\\"-1175.0000000000_-257.5000000000\\\",\\\"-747.5000000000_-257.5000000000\\\",\\\"-747.5000000000_-550.0000000000\\\",\\\"-417.5000000000_-550.0000000000\\\"]}\"}","{\"color\":\"#774D00\",\"startPinId\":\"pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6\",\"rawStartPinId\":\"pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-432.5000000000_-790.0000000000\\\",\\\"-470.0000000000_-790.0000000000\\\",\\\"-470.0000000000_-550.0000000000\\\",\\\"-417.5000000000_-550.0000000000\\\"]}\"}","{\"color\":\"#7A4782\",\"startPinId\":\"pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_1\",\"endPinId\":\"pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_1\",\"rawStartPinId\":\"pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_1\",\"rawEndPinId\":\"pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1332.5000000000_-160.0000000000\\\",\\\"-1220.0000000000_-160.0000000000\\\",\\\"-1220.0000000000_-175.0000000000\\\",\\\"-1197.5000000000_-175.0000000000\\\",\\\"-1197.5000000000_-170.7041515000\\\"]}\"}","{\"color\":\"#004754\",\"startPinId\":\"pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_1\",\"endPinId\":\"pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_1\",\"rawStartPinId\":\"pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_1\",\"rawEndPinId\":\"pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_-44.2958485000\\\",\\\"-1197.5000000000_-25.0000000000\\\",\\\"-1220.0000000000_-25.0000000000\\\",\\\"-1220.0000000000_-55.0000000000\\\",\\\"-1332.5000000000_-55.0000000000\\\"]}\"}","{\"color\":\"#FFB167\",\"startPinId\":\"pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_1\",\"endPinId\":\"pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1\",\"rawStartPinId\":\"pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_1\",\"rawEndPinId\":\"pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_54.2958485000\\\",\\\"-1197.5000000000_50.0000000000\\\",\\\"-1220.0000000000_50.0000000000\\\",\\\"-1220.0000000000_65.0000000000\\\",\\\"-1332.5000000000_65.0000000000\\\"]}\"}","{\"color\":\"#6685ff\",\"startPinId\":\"pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_1\",\"endPinId\":\"pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_1\",\"rawStartPinId\":\"pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_1\",\"rawEndPinId\":\"pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_180.7041515000\\\",\\\"-1197.5000000000_192.5000000000\\\",\\\"-1220.0000000000_192.5000000000\\\",\\\"-1220.0000000000_170.0000000000\\\",\\\"-1332.5000000000_170.0000000000\\\"]}\"}","{\"color\":\"#90FB92\",\"startPinId\":\"pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0\",\"endPinId\":\"pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_0\",\"rawStartPinId\":\"pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0\",\"rawEndPinId\":\"pin-type-component_35159cb3-cc74-4c90-b0f5-cff583f979a5_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_125.0000000000\\\",\\\"-1197.5000000000_110.0000000000\\\"]}\"}","{\"color\":\"#90FB92\",\"startPinId\":\"pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4\",\"rawStartPinId\":\"pin-type-component_2f031f22-1944-43ab-ae9c-f74e47cc4156_0\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_125.0000000000\\\",\\\"-1160.0000000000_125.0000000000\\\",\\\"-1160.0000000000_-242.5000000000\\\",\\\"-725.0000000000_-242.5000000000\\\",\\\"-725.0000000000_-520.0000000000\\\",\\\"-417.5000000000_-520.0000000000\\\"]}\"}","{\"color\":\"#90FB92\",\"startPinId\":\"pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4\",\"rawStartPinId\":\"pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-432.5000000000_-850.0000000000\\\",\\\"-485.0000000000_-850.0000000000\\\",\\\"-485.0000000000_-520.0000000000\\\",\\\"-417.5000000000_-520.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_0\",\"endPinId\":\"pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0\",\"rawStartPinId\":\"pin-type-component_0152d242-8b4d-42db-8096-0f8dc98256f3_0\",\"rawEndPinId\":\"pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_-100.0000000000\\\",\\\"-1197.5000000000_-115.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5\",\"endPinId\":\"pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0\",\"rawStartPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5\",\"rawEndPinId\":\"pin-type-component_d6e5c84b-c20b-48f5-a42a-5c5a8ecfc61c_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-535.0000000000\\\",\\\"-740.0000000000_-535.0000000000\\\",\\\"-740.0000000000_-250.0000000000\\\",\\\"-1175.0000000000_-250.0000000000\\\",\\\"-1175.0000000000_-100.0000000000\\\",\\\"-1197.5000000000_-100.0000000000\\\",\\\"-1197.5000000000_-115.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5\",\"endPinId\":\"pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_1\",\"rawStartPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_5\",\"rawEndPinId\":\"pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-535.0000000000\\\",\\\"-477.5000000000_-535.0000000000\\\",\\\"-477.5000000000_-820.0000000000\\\",\\\"-432.5000000000_-820.0000000000\\\"]}\"}","{\"color\":\"#BDD393\",\"startPinId\":\"pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_1\",\"endPinId\":\"pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_1\",\"rawStartPinId\":\"pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_1\",\"rawEndPinId\":\"pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_65.0000000000\\\",\\\"-957.5000000000_65.0000000000\\\",\\\"-957.5000000000_42.5000000000\\\",\\\"-942.5000000000_42.5000000000\\\",\\\"-942.5000000000_54.2958485000\\\"]}\"}","{\"color\":\"#E56FFE\",\"startPinId\":\"pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_1\",\"endPinId\":\"pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_1\",\"rawStartPinId\":\"pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_1\",\"rawEndPinId\":\"pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_170.0000000000\\\",\\\"-957.5000000000_170.0000000000\\\",\\\"-957.5000000000_192.5000000000\\\",\\\"-942.5000000000_192.5000000000\\\",\\\"-942.5000000000_180.7041515000\\\"]}\"}","{\"color\":\"#001eff\",\"startPinId\":\"pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_0\",\"endPinId\":\"pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0\",\"rawStartPinId\":\"pin-type-component_625dbf85-54ff-48b2-a275-4089e5081167_0\",\"rawEndPinId\":\"pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-942.5000000000_110.0000000000\\\",\\\"-942.5000000000_125.0000000000\\\"]}\"}","{\"color\":\"#001eff\",\"startPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0\",\"endPinId\":\"pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0\",\"rawStartPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0\",\"rawEndPinId\":\"pin-type-component_f86ac869-5086-4a06-8cd6-49f486548944_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-460.0000000000\\\",\\\"-665.0000000000_-460.0000000000\\\",\\\"-665.0000000000_125.0000000000\\\",\\\"-942.5000000000_125.0000000000\\\"]}\"}","{\"color\":\"#001eff\",\"startPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0\",\"endPinId\":\"pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_1\",\"rawStartPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_0\",\"rawEndPinId\":\"pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-460.0000000000\\\",\\\"-455.0000000000_-460.0000000000\\\",\\\"-455.0000000000_-737.5000000000\\\",\\\"-350.0000000000_-737.5000000000\\\",\\\"-350.0000000000_-850.0000000000\\\",\\\"-312.5000000000_-850.0000000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_1\",\"endPinId\":\"pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_1\",\"rawStartPinId\":\"pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_1\",\"rawEndPinId\":\"pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-927.5000000000_-170.7041515000\\\",\\\"-927.5000000000_-190.0000000000\\\",\\\"-950.0000000000_-190.0000000000\\\",\\\"-950.0000000000_-160.0000000000\\\",\\\"-1062.5000000000_-160.0000000000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_1\",\"endPinId\":\"pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_1\",\"rawStartPinId\":\"pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_1\",\"rawEndPinId\":\"pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-55.0000000000\\\",\\\"-950.0000000000_-55.0000000000\\\",\\\"-950.0000000000_-32.5000000000\\\",\\\"-927.5000000000_-32.5000000000\\\",\\\"-927.5000000000_-44.2958485000\\\"]}\"}","{\"color\":\"#00FFC6\",\"startPinId\":\"pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_0\",\"endPinId\":\"pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0\",\"rawStartPinId\":\"pin-type-component_0c68c6e3-0464-4e71-ab6a-9086b01a0e77_0\",\"rawEndPinId\":\"pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-927.5000000000_-115.0000000000\\\",\\\"-927.5000000000_-100.0000000000\\\"]}\"}","{\"color\":\"#00FFC6\",\"startPinId\":\"pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1\",\"rawStartPinId\":\"pin-type-component_709ba052-a0a0-4439-a40d-83aedf155550_0\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-927.5000000000_-100.0000000000\\\",\\\"-680.0000000000_-100.0000000000\\\",\\\"-680.0000000000_-475.0000000000\\\",\\\"-417.5000000000_-475.0000000000\\\"]}\"}","{\"color\":\"#00FFC6\",\"startPinId\":\"pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1\",\"rawStartPinId\":\"pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-312.5000000000_-820.0000000000\\\",\\\"-342.5000000000_-820.0000000000\\\",\\\"-342.5000000000_-730.0000000000\\\",\\\"-447.5000000000_-730.0000000000\\\",\\\"-447.5000000000_-475.0000000000\\\",\\\"-417.5000000000_-475.0000000000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_1\",\"endPinId\":\"pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_1\",\"rawStartPinId\":\"pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_1\",\"rawEndPinId\":\"pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-927.5000000000_-470.7041515000\\\",\\\"-927.5000000000_-490.0000000000\\\",\\\"-957.5000000000_-490.0000000000\\\",\\\"-957.5000000000_-460.0000000000\\\",\\\"-1062.5000000000_-460.0000000000\\\"]}\"}","{\"color\":\"#E85EBE\",\"startPinId\":\"pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_1\",\"endPinId\":\"pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_1\",\"rawStartPinId\":\"pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_1\",\"rawEndPinId\":\"pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-355.0000000000\\\",\\\"-942.5000000000_-355.0000000000\\\",\\\"-942.5000000000_-325.0000000000\\\",\\\"-927.5000000000_-325.0000000000\\\",\\\"-927.5000000000_-344.2958485000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_0\",\"endPinId\":\"pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0\",\"rawStartPinId\":\"pin-type-component_4b0e618a-0090-4173-a14d-dc77951515d3_0\",\"rawEndPinId\":\"pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-927.5000000000_-415.0000000000\\\",\\\"-927.5000000000_-400.0000000000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2\",\"rawStartPinId\":\"pin-type-component_733ac60f-fd5b-4e01-bcd0-44ae417225ee_0\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-927.5000000000_-400.0000000000\\\",\\\"-867.5000000000_-400.0000000000\\\",\\\"-867.5000000000_-205.0000000000\\\",\\\"-695.0000000000_-205.0000000000\\\",\\\"-695.0000000000_-490.0000000000\\\",\\\"-417.5000000000_-490.0000000000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2\",\"rawStartPinId\":\"pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-312.5000000000_-790.0000000000\\\",\\\"-327.5000000000_-790.0000000000\\\",\\\"-327.5000000000_-722.5000000000\\\",\\\"-440.0000000000_-722.5000000000\\\",\\\"-440.0000000000_-490.0000000000\\\",\\\"-417.5000000000_-490.0000000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_1\",\"endPinId\":\"pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_1\",\"rawStartPinId\":\"pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_1\",\"rawEndPinId\":\"pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-912.5000000000_-695.7041515000\\\",\\\"-912.5000000000_-700.0000000000\\\",\\\"-1062.5000000000_-700.0000000000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_1\",\"endPinId\":\"pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_1\",\"rawStartPinId\":\"pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_1\",\"rawEndPinId\":\"pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-580.0000000000\\\",\\\"-935.0000000000_-580.0000000000\\\",\\\"-935.0000000000_-542.5000000000\\\",\\\"-912.5000000000_-542.5000000000\\\",\\\"-912.5000000000_-569.2958485000\\\"]}\"}","{\"color\":\"#ff0066\",\"startPinId\":\"pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_0\",\"endPinId\":\"pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0\",\"rawStartPinId\":\"pin-type-component_114d5d14-5f5c-40e8-b182-5aaaa19436dd_0\",\"rawEndPinId\":\"pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-912.5000000000_-640.0000000000\\\",\\\"-912.5000000000_-625.0000000000\\\"]}\"}","{\"color\":\"#ff0066\",\"startPinId\":\"pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3\",\"rawStartPinId\":\"pin-type-component_4f53b9c5-5f30-4a72-af1a-a8232ad99f6b_0\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-912.5000000000_-625.0000000000\\\",\\\"-845.0000000000_-625.0000000000\\\",\\\"-845.0000000000_-227.5000000000\\\",\\\"-710.0000000000_-227.5000000000\\\",\\\"-710.0000000000_-505.0000000000\\\",\\\"-417.5000000000_-505.0000000000\\\"]}\"}","{\"color\":\"#ff0066\",\"startPinId\":\"pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_1\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3\",\"rawStartPinId\":\"pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_1\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-312.5000000000_-760.0000000000\\\",\\\"-312.5000000000_-707.5000000000\\\",\\\"-432.5000000000_-707.5000000000\\\",\\\"-432.5000000000_-505.0000000000\\\",\\\"-417.5000000000_-505.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0\",\"endPinId\":\"pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0\",\"rawStartPinId\":\"pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0\",\"rawEndPinId\":\"pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-2277.5000000000_-535.0000000000\\\",\\\"-2307.5000000000_-535.0000000000\\\",\\\"-2307.5000000000_-415.0000000000\\\",\\\"-2277.5000000000_-415.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0\",\"endPinId\":\"pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0\",\"rawStartPinId\":\"pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0\",\"rawEndPinId\":\"pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-2277.5000000000_-535.0000000000\\\",\\\"-2307.5000000000_-535.0000000000\\\",\\\"-2307.5000000000_-1015.0000000000\\\",\\\"-1392.5000000000_-1015.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0\",\"endPinId\":\"pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0\",\"rawStartPinId\":\"pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_0\",\"rawEndPinId\":\"pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1392.5000000000_-1015.0000000000\\\",\\\"-1407.5000000000_-1015.0000000000\\\",\\\"-1407.5000000000_-1090.0000000000\\\",\\\"-1392.5000000000_-1090.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0\",\"endPinId\":\"pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0\",\"rawStartPinId\":\"pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0\",\"rawEndPinId\":\"pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1392.5000000000_-1165.0000000000\\\",\\\"-1407.5000000000_-1165.0000000000\\\",\\\"-1407.5000000000_-1090.0000000000\\\",\\\"-1392.5000000000_-1090.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_0\",\"endPinId\":\"pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0\",\"rawStartPinId\":\"pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_0\",\"rawEndPinId\":\"pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1392.5000000000_-1240.0000000000\\\",\\\"-1407.5000000000_-1240.0000000000\\\",\\\"-1407.5000000000_-1165.0000000000\\\",\\\"-1392.5000000000_-1165.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0\",\"endPinId\":\"pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0\",\"rawStartPinId\":\"pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0\",\"rawEndPinId\":\"pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-2292.5000000000_-355.0000000000\\\",\\\"-2307.5000000000_-355.0000000000\\\",\\\"-2307.5000000000_305.0000000000\\\",\\\"-1617.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0\",\"endPinId\":\"pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0\",\"rawStartPinId\":\"pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0\",\"rawEndPinId\":\"pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1617.5000000000_380.0000000000\\\",\\\"-1632.5000000000_380.0000000000\\\",\\\"-1632.5000000000_305.0000000000\\\",\\\"-1617.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0\",\"endPinId\":\"pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0\",\"rawStartPinId\":\"pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0\",\"rawEndPinId\":\"pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1617.5000000000_455.0000000000\\\",\\\"-1632.5000000000_455.0000000000\\\",\\\"-1632.5000000000_380.0000000000\\\",\\\"-1617.5000000000_380.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0\",\"endPinId\":\"pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0\",\"rawStartPinId\":\"pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_0\",\"rawEndPinId\":\"pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1617.5000000000_455.0000000000\\\",\\\"-1632.5000000000_455.0000000000\\\",\\\"-1632.5000000000_530.0000000000\\\",\\\"-1617.5000000000_530.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0\",\"endPinId\":\"pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0\",\"rawStartPinId\":\"pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0\",\"rawEndPinId\":\"pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-303.4957806029_307.9943741372\\\",\\\"-327.5000000000_307.9943741372\\\",\\\"-327.5000000000_232.9943741372\\\",\\\"-303.4957806029_232.9943741372\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0\",\"endPinId\":\"pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0\",\"rawStartPinId\":\"pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_0\",\"rawEndPinId\":\"pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-303.4957806029_307.9943741372\\\",\\\"-327.5000000000_307.9943741372\\\",\\\"-327.5000000000_382.9943741372\\\",\\\"-303.4957806029_382.9943741372\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0\",\"endPinId\":\"pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0\",\"rawStartPinId\":\"pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0\",\"rawEndPinId\":\"pin-type-component_c525269a-6029-466e-8297-23d196a50c50_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-303.4957806029_457.9943741372\\\",\\\"-327.5000000000_457.9943741372\\\",\\\"-327.5000000000_382.9943741372\\\",\\\"-303.4957806029_382.9943741372\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0\",\"endPinId\":\"pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0\",\"rawStartPinId\":\"pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0\",\"rawEndPinId\":\"pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-303.4957806029_457.9943741372\\\",\\\"-303.4957806029_590.0000000000\\\",\\\"-1632.5000000000_590.0000000000\\\",\\\"-1632.5000000000_530.0000000000\\\",\\\"-1617.5000000000_530.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_3\",\"rawStartPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"439.4500000000_-79.6000000000\\\",\\\"302.5000000000_-79.6000000000\\\",\\\"302.5000000000_-475.0000000000\\\",\\\"332.5000000000_-475.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10\",\"endPinId\":\"pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0\",\"rawStartPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_10\",\"rawEndPinId\":\"pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"439.4500000000_-79.6000000000\\\",\\\"439.4500000000_590.0000000000\\\",\\\"-305.0000000000_590.0000000000\\\",\\\"-305.0000000000_457.9943741372\\\",\\\"-303.4957806029_457.9943741372\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0\",\"endPinId\":\"pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0\",\"rawStartPinId\":\"pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_0\",\"rawEndPinId\":\"pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-2292.5000000000_-355.0000000000\\\",\\\"-2307.5000000000_-355.0000000000\\\",\\\"-2307.5000000000_-415.0000000000\\\",\\\"-2277.5000000000_-415.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0\",\"endPinId\":\"pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0\",\"rawStartPinId\":\"pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_0\",\"rawEndPinId\":\"pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-2277.5000000000_-535.0000000000\\\",\\\"-2307.5000000000_-535.0000000000\\\",\\\"-2307.5000000000_-480.2239686398\\\",\\\"-2291.0744138637_-480.2239686398\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1\",\"endPinId\":\"pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0\",\"rawStartPinId\":\"pin-type-component_621585ad-95ad-4cf3-9a10-1ca969371d4e_1\",\"rawEndPinId\":\"pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-2154.3320000000_-354.0745000000\\\",\\\"-2142.5000000000_-354.0745000000\\\",\\\"-2142.5000000000_230.0000000000\\\",\\\"-1977.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2\",\"endPinId\":\"pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1\",\"rawStartPinId\":\"pin-type-component_041b5070-e88a-4a6b-aa2c-a93c5f45650d_2\",\"rawEndPinId\":\"pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_170.0000000000\\\",\\\"-1827.5000000000_170.0000000000\\\",\\\"-1827.5000000000_230.0000000000\\\",\\\"-1932.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2\",\"endPinId\":\"pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1\",\"rawStartPinId\":\"pin-type-component_83dcf7d9-214a-4ba8-8c4b-0198867c485d_2\",\"rawEndPinId\":\"pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_65.0000000000\\\",\\\"-1857.5000000000_110.0000000000\\\",\\\"-1932.5000000000_110.0000000000\\\",\\\"-1932.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12\",\"endPinId\":\"pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_12\",\"rawEndPinId\":\"pin-type-component_995a17d1-5928-497f-b230-e981cff0c0da_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-250.0000000000\\\",\\\"-507.5000000000_-250.0000000000\\\",\\\"-507.5000000000_-347.5000000000\\\",\\\"-125.0000000000_-347.5000000000\\\",\\\"-125.0000000000_-880.0000000000\\\",\\\"-2112.5000000000_-880.0000000000\\\",\\\"-2112.5000000000_230.0000000000\\\",\\\"-1932.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2\",\"endPinId\":\"pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1\",\"rawStartPinId\":\"pin-type-component_3a88c66b-feb0-48c3-be15-37e3d48518eb_2\",\"rawEndPinId\":\"pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_-85.0000000000\\\",\\\"-1812.5000000000_-85.0000000000\\\",\\\"-1812.5000000000_-25.0000000000\\\",\\\"-1932.5000000000_-25.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2\",\"endPinId\":\"pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1\",\"rawStartPinId\":\"pin-type-component_46f90c07-7d13-4392-a3bf-e813e3dabb36_2\",\"rawEndPinId\":\"pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1857.5000000000_-160.0000000000\\\",\\\"-1857.5000000000_-137.5000000000\\\",\\\"-1932.5000000000_-137.5000000000\\\",\\\"-1932.5000000000_-25.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13\",\"endPinId\":\"pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_13\",\"rawEndPinId\":\"pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-265.0000000000\\\",\\\"-492.5000000000_-265.0000000000\\\",\\\"-492.5000000000_-362.5000000000\\\",\\\"-147.5000000000_-362.5000000000\\\",\\\"-147.5000000000_-910.0000000000\\\",\\\"-2037.5000000000_-910.0000000000\\\",\\\"-2037.5000000000_-25.0000000000\\\",\\\"-1932.5000000000_-25.0000000000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1\",\"endPinId\":\"pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2\",\"rawStartPinId\":\"pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1\",\"rawEndPinId\":\"pin-type-component_7cf5453a-9a65-47be-a0c1-a40e3c54981e_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1932.5000000000_-295.0000000000\\\",\\\"-1812.5000000000_-295.0000000000\\\",\\\"-1812.5000000000_-355.0000000000\\\",\\\"-1857.5000000000_-355.0000000000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1\",\"endPinId\":\"pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2\",\"rawStartPinId\":\"pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1\",\"rawEndPinId\":\"pin-type-component_73ff6e4f-35de-4fa1-bb93-81012f621ef2_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1932.5000000000_-295.0000000000\\\",\\\"-1925.0000000000_-295.0000000000\\\",\\\"-1925.0000000000_-422.5000000000\\\",\\\"-1857.5000000000_-422.5000000000\\\",\\\"-1857.5000000000_-460.0000000000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14\",\"endPinId\":\"pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_14\",\"rawEndPinId\":\"pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-280.0000000000\\\",\\\"-470.0000000000_-280.0000000000\\\",\\\"-470.0000000000_-385.0000000000\\\",\\\"-170.0000000000_-385.0000000000\\\",\\\"-170.0000000000_-970.0000000000\\\",\\\"-1992.5000000000_-970.0000000000\\\",\\\"-1992.5000000000_-295.0000000000\\\",\\\"-1932.5000000000_-295.0000000000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1\",\"endPinId\":\"pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2\",\"rawStartPinId\":\"pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1\",\"rawEndPinId\":\"pin-type-component_67df4d37-3f2b-4d48-9904-dc3e640854f2_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1932.5000000000_-535.0000000000\\\",\\\"-1812.5000000000_-535.0000000000\\\",\\\"-1812.5000000000_-580.0000000000\\\",\\\"-1857.5000000000_-580.0000000000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1\",\"endPinId\":\"pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2\",\"rawStartPinId\":\"pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1\",\"rawEndPinId\":\"pin-type-component_8fd76732-6e42-40ac-b9ab-aae7428798a1_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1932.5000000000_-535.0000000000\\\",\\\"-1932.5000000000_-655.0000000000\\\",\\\"-1857.5000000000_-655.0000000000\\\",\\\"-1857.5000000000_-700.0000000000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15\",\"endPinId\":\"pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_15\",\"rawEndPinId\":\"pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-295.0000000000\\\",\\\"-440.0000000000_-295.0000000000\\\",\\\"-440.0000000000_-407.5000000000\\\",\\\"-192.5000000000_-407.5000000000\\\",\\\"-192.5000000000_-940.0000000000\\\",\\\"-1932.5000000000_-940.0000000000\\\",\\\"-1932.5000000000_-535.0000000000\\\"]}\"}","{\"color\":\"#A5FFD2\",\"startPinId\":\"pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0\",\"endPinId\":\"pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1\",\"rawStartPinId\":\"pin-type-component_81ae35b1-5b71-4716-a1af-fd111af3ac03_0\",\"rawEndPinId\":\"pin-type-component_efd3f3bc-1ae1-45dd-a482-193032279b23_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1977.5000000000_-25.0000000000\\\",\\\"-2022.5000000000_-25.0000000000\\\",\\\"-2022.5000000000_-414.0745000000\\\",\\\"-2139.3320000000_-414.0745000000\\\"]}\"}","{\"color\":\"#FFA6FE\",\"startPinId\":\"pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0\",\"endPinId\":\"pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1\",\"rawStartPinId\":\"pin-type-component_41446abf-3582-4e1a-bca9-cf131a5fba1c_0\",\"rawEndPinId\":\"pin-type-component_a86bd662-6cba-44a0-8211-7ce5de8f1e54_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1977.5000000000_-295.0000000000\\\",\\\"-2007.5000000000_-295.0000000000\\\",\\\"-2007.5000000000_-479.2984686398\\\",\\\"-2152.9064138637_-479.2984686398\\\"]}\"}","{\"color\":\"#774D00\",\"startPinId\":\"pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1\",\"endPinId\":\"pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0\",\"rawStartPinId\":\"pin-type-component_0d024f4d-e2f2-4b76-8f77-420b1168f36c_1\",\"rawEndPinId\":\"pin-type-component_3694689b-7dc6-49dc-a8fa-3e18614c7e29_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-2139.3320000000_-534.0745000000\\\",\\\"-1983.4160000000_-534.0745000000\\\",\\\"-1983.4160000000_-535.0000000000\\\",\\\"-1977.5000000000_-535.0000000000\\\"]}\"}","{\"color\":\"#7A4782\",\"startPinId\":\"pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2\",\"endPinId\":\"pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2\",\"rawStartPinId\":\"pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2\",\"rawEndPinId\":\"pin-type-component_3569e0a5-063e-4474-b7f3-fd780070bcdd_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_170.0000000000\\\",\\\"-1542.5000000000_170.0000000000\\\",\\\"-1542.5000000000_65.0000000000\\\",\\\"-1587.5000000000_65.0000000000\\\"]}\"}","{\"color\":\"#7A4782\",\"startPinId\":\"pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2\",\"endPinId\":\"pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1\",\"rawStartPinId\":\"pin-type-component_01ef38d5-a6be-49e6-b75b-fe4690ca3d8a_2\",\"rawEndPinId\":\"pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_170.0000000000\\\",\\\"-1542.5000000000_170.0000000000\\\",\\\"-1542.5000000000_305.0000000000\\\",\\\"-1422.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#7A4782\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8\",\"endPinId\":\"pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_8\",\"rawEndPinId\":\"pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-190.0000000000\\\",\\\"-515.0000000000_-190.0000000000\\\",\\\"-515.0000000000_305.0000000000\\\",\\\"-1422.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#004754\",\"startPinId\":\"pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2\",\"endPinId\":\"pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2\",\"rawStartPinId\":\"pin-type-component_3cc0d351-6a54-4350-a5dc-29ea6ac8f53f_2\",\"rawEndPinId\":\"pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_-160.0000000000\\\",\\\"-1542.5000000000_-160.0000000000\\\",\\\"-1542.5000000000_-55.0000000000\\\",\\\"-1587.5000000000_-55.0000000000\\\"]}\"}","{\"color\":\"#004754\",\"startPinId\":\"pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2\",\"endPinId\":\"pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1\",\"rawStartPinId\":\"pin-type-component_a28b7076-045f-481a-8987-e6c379c85461_2\",\"rawEndPinId\":\"pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_-55.0000000000\\\",\\\"-1497.5000000000_-55.0000000000\\\",\\\"-1497.5000000000_380.0000000000\\\",\\\"-1407.5000000000_380.0000000000\\\"]}\"}","{\"color\":\"#004754\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9\",\"endPinId\":\"pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_9\",\"rawEndPinId\":\"pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-205.0000000000\\\",\\\"-537.5000000000_-205.0000000000\\\",\\\"-537.5000000000_380.0000000000\\\",\\\"-1407.5000000000_380.0000000000\\\"]}\"}","{\"color\":\"#B500FF\",\"startPinId\":\"pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2\",\"endPinId\":\"pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2\",\"rawStartPinId\":\"pin-type-component_549bec3f-89a4-4854-8eed-2d9171821a2f_2\",\"rawEndPinId\":\"pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_-460.0000000000\\\",\\\"-1542.5000000000_-460.0000000000\\\",\\\"-1542.5000000000_-355.0000000000\\\",\\\"-1587.5000000000_-355.0000000000\\\"]}\"}","{\"color\":\"#B500FF\",\"startPinId\":\"pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2\",\"endPinId\":\"pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1\",\"rawStartPinId\":\"pin-type-component_8649ae8f-4a7d-41ac-b7cc-e72e54b8f55b_2\",\"rawEndPinId\":\"pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_-355.0000000000\\\",\\\"-1587.5000000000_-257.5000000000\\\",\\\"-1490.0000000000_-257.5000000000\\\",\\\"-1490.0000000000_455.0000000000\\\",\\\"-1407.5000000000_455.0000000000\\\"]}\"}","{\"color\":\"#B500FF\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10\",\"endPinId\":\"pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_10\",\"rawEndPinId\":\"pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-220.0000000000\\\",\\\"-560.0000000000_-220.0000000000\\\",\\\"-560.0000000000_455.0000000000\\\",\\\"-1407.5000000000_455.0000000000\\\"]}\"}","{\"color\":\"#f50a0a\",\"startPinId\":\"pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2\",\"endPinId\":\"pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2\",\"rawStartPinId\":\"pin-type-component_1b855ccb-49a4-427a-9563-e1bcdb16e638_2\",\"rawEndPinId\":\"pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1587.5000000000_-700.0000000000\\\",\\\"-1542.5000000000_-700.0000000000\\\",\\\"-1542.5000000000_-580.0000000000\\\",\\\"-1587.5000000000_-580.0000000000\\\"]}\"}","{\"color\":\"#f50a0a\",\"startPinId\":\"pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1\",\"endPinId\":\"pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2\",\"rawStartPinId\":\"pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1\",\"rawEndPinId\":\"pin-type-component_b3ed5ea8-d9ad-4aa4-b08b-9e6ddb1d9e99_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1407.5000000000_530.0000000000\\\",\\\"-1415.0000000000_530.0000000000\\\",\\\"-1415.0000000000_-550.0000000000\\\",\\\"-1587.5000000000_-550.0000000000\\\",\\\"-1587.5000000000_-580.0000000000\\\"]}\"}","{\"color\":\"#f50a0a\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11\",\"endPinId\":\"pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_11\",\"rawEndPinId\":\"pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-235.0000000000\\\",\\\"-590.0000000000_-235.0000000000\\\",\\\"-590.0000000000_530.0000000000\\\",\\\"-1407.5000000000_530.0000000000\\\"]}\"}","{\"color\":\"#FFDB66\",\"startPinId\":\"pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_0\",\"endPinId\":\"pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_1\",\"rawStartPinId\":\"pin-type-component_a8e515ed-cb32-4abf-ab34-4e8ba550aff5_0\",\"rawEndPinId\":\"pin-type-component_b69e0669-3879-4abd-9d7d-acc45f8eea74_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1467.5000000000_305.0000000000\\\",\\\"-1473.4160000000_305.0000000000\\\",\\\"-1473.4160000000_305.9255000000\\\",\\\"-1479.3320000000_305.9255000000\\\"]}\"}","{\"color\":\"#90FB92\",\"startPinId\":\"pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_1\",\"endPinId\":\"pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_0\",\"rawStartPinId\":\"pin-type-component_5712632d-8fa8-495b-a104-baf8f43c700a_1\",\"rawEndPinId\":\"pin-type-component_efcea04e-21d8-44a5-8f0d-74277474a2e0_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1479.3320000000_380.9255000000\\\",\\\"-1458.4160000000_380.9255000000\\\",\\\"-1458.4160000000_380.0000000000\\\",\\\"-1452.5000000000_380.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_1\",\"endPinId\":\"pin-type-component_c107267e-960a-414d-898a-9b8f86844804_0\",\"rawStartPinId\":\"pin-type-component_0b992200-29a8-47ae-9e2d-5041f24e3da4_1\",\"rawEndPinId\":\"pin-type-component_c107267e-960a-414d-898a-9b8f86844804_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1254.3320000000_-1239.0745000000\\\",\\\"-1263.4160000000_-1239.0745000000\\\",\\\"-1263.4160000000_-1240.0000000000\\\",\\\"-1257.5000000000_-1240.0000000000\\\"]}\"}","{\"color\":\"#BDD393\",\"startPinId\":\"pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_1\",\"endPinId\":\"pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_0\",\"rawStartPinId\":\"pin-type-component_ddbc596a-7cd5-4048-bdec-ae929062b39f_1\",\"rawEndPinId\":\"pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1254.3320000000_-1164.0745000000\\\",\\\"-1248.4160000000_-1164.0745000000\\\",\\\"-1248.4160000000_-1165.0000000000\\\",\\\"-1242.5000000000_-1165.0000000000\\\"]}\"}","{\"color\":\"#E56FFE\",\"startPinId\":\"pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_0\",\"endPinId\":\"pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_1\",\"rawStartPinId\":\"pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_0\",\"rawEndPinId\":\"pin-type-component_ee4052d6-2dbe-445a-8b8e-b1c8214d283a_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1242.5000000000_-1090.0000000000\\\",\\\"-1248.4160000000_-1090.0000000000\\\",\\\"-1248.4160000000_-1089.0745000000\\\",\\\"-1254.3320000000_-1089.0745000000\\\"]}\"}","{\"color\":\"#00FF78\",\"startPinId\":\"pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_0\",\"endPinId\":\"pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_1\",\"rawStartPinId\":\"pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_0\",\"rawEndPinId\":\"pin-type-component_c90e906b-172f-43f0-a66d-c99371504fba_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1242.5000000000_-1015.0000000000\\\",\\\"-1248.4160000000_-1015.0000000000\\\",\\\"-1248.4160000000_-1014.0745000000\\\",\\\"-1254.3320000000_-1014.0745000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2\",\"endPinId\":\"pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2\",\"rawStartPinId\":\"pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2\",\"rawEndPinId\":\"pin-type-component_8d75e431-ab93-4f28-a072-73fa2a9add70_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1332.5000000000_185.0000000000\\\",\\\"-1287.5000000000_185.0000000000\\\",\\\"-1287.5000000000_80.0000000000\\\",\\\"-1332.5000000000_80.0000000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2\",\"endPinId\":\"pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1\",\"rawStartPinId\":\"pin-type-component_6fba6b65-b569-4c04-b286-0556b7aca02c_2\",\"rawEndPinId\":\"pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1332.5000000000_185.0000000000\\\",\\\"-1332.5000000000_200.0000000000\\\",\\\"-1122.5000000000_200.0000000000\\\",\\\"-1122.5000000000_-1240.0000000000\\\",\\\"-1212.5000000000_-1240.0000000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_4\",\"endPinId\":\"pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_4\",\"rawEndPinId\":\"pin-type-component_c107267e-960a-414d-898a-9b8f86844804_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-130.0000000000\\\",\\\"-455.0000000000_-130.0000000000\\\",\\\"-455.0000000000_20.0000000000\\\",\\\"122.5000000000_20.0000000000\\\",\\\"122.5000000000_-1240.0000000000\\\",\\\"-1212.5000000000_-1240.0000000000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2\",\"endPinId\":\"pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2\",\"rawStartPinId\":\"pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2\",\"rawEndPinId\":\"pin-type-component_a42f6e75-c6ce-4431-8ab7-a546cadc6910_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1332.5000000000_-40.0000000000\\\",\\\"-1287.5000000000_-40.0000000000\\\",\\\"-1287.5000000000_-145.0000000000\\\",\\\"-1332.5000000000_-145.0000000000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2\",\"endPinId\":\"pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1\",\"rawStartPinId\":\"pin-type-component_8a57da25-4acd-4f0c-b8e8-8e9646645470_2\",\"rawEndPinId\":\"pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1332.5000000000_-40.0000000000\\\",\\\"-1332.5000000000_-10.0000000000\\\",\\\"-1137.5000000000_-10.0000000000\\\",\\\"-1137.5000000000_-1165.0000000000\\\",\\\"-1197.5000000000_-1165.0000000000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_5\",\"endPinId\":\"pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_5\",\"rawEndPinId\":\"pin-type-component_e7200013-28f8-4ff6-9dbe-a2239e215492_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-145.0000000000\\\",\\\"-470.0000000000_-145.0000000000\\\",\\\"-470.0000000000_42.5000000000\\\",\\\"92.5000000000_42.5000000000\\\",\\\"92.5000000000_-1165.0000000000\\\",\\\"-1197.5000000000_-1165.0000000000\\\"]}\"}","{\"color\":\"#00FFC6\",\"startPinId\":\"pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2\",\"endPinId\":\"pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2\",\"rawStartPinId\":\"pin-type-component_274be705-445b-40a5-9ab8-ea55a1873ac7_2\",\"rawEndPinId\":\"pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1332.5000000000_-445.0000000000\\\",\\\"-1287.5000000000_-445.0000000000\\\",\\\"-1287.5000000000_-340.0000000000\\\",\\\"-1332.5000000000_-340.0000000000\\\"]}\"}","{\"color\":\"#00FFC6\",\"startPinId\":\"pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1\",\"endPinId\":\"pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2\",\"rawStartPinId\":\"pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1\",\"rawEndPinId\":\"pin-type-component_ddf014d2-e81b-4ce5-802e-4329eb48f7e0_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_-1090.0000000000\\\",\\\"-1145.0000000000_-1090.0000000000\\\",\\\"-1145.0000000000_-332.5000000000\\\",\\\"-1332.5000000000_-332.5000000000\\\",\\\"-1332.5000000000_-340.0000000000\\\"]}\"}","{\"color\":\"#00FFC6\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_6\",\"endPinId\":\"pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_6\",\"rawEndPinId\":\"pin-type-component_c58023a8-eade-4368-93d4-c18f7148e8e3_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-160.0000000000\\\",\\\"-485.0000000000_-160.0000000000\\\",\\\"-485.0000000000_72.5000000000\\\",\\\"70.0000000000_72.5000000000\\\",\\\"70.0000000000_-1090.0000000000\\\",\\\"-1197.5000000000_-1090.0000000000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2\",\"endPinId\":\"pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2\",\"rawStartPinId\":\"pin-type-component_458ace7d-db58-47fe-9e9e-81463f1cb31c_2\",\"rawEndPinId\":\"pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1332.5000000000_-565.0000000000\\\",\\\"-1287.5000000000_-565.0000000000\\\",\\\"-1287.5000000000_-685.0000000000\\\",\\\"-1332.5000000000_-685.0000000000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1\",\"endPinId\":\"pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2\",\"rawStartPinId\":\"pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1\",\"rawEndPinId\":\"pin-type-component_8ac7020a-2504-45c9-b517-84bd506cb24c_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1197.5000000000_-1015.0000000000\\\",\\\"-1160.0000000000_-1015.0000000000\\\",\\\"-1160.0000000000_-685.0000000000\\\",\\\"-1332.5000000000_-685.0000000000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_7\",\"endPinId\":\"pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_7\",\"rawEndPinId\":\"pin-type-component_15591579-4d1a-4075-aec4-52c43cc21020_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-175.0000000000\\\",\\\"-500.0000000000_-175.0000000000\\\",\\\"-500.0000000000_87.5000000000\\\",\\\"40.0000000000_87.5000000000\\\",\\\"40.0000000000_-1015.0000000000\\\",\\\"-1197.5000000000_-1015.0000000000\\\"]}\"}","{\"color\":\"#E85EBE\",\"startPinId\":\"pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_1\",\"endPinId\":\"pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_0\",\"rawStartPinId\":\"pin-type-component_4b269a77-3c6b-4832-bc03-819b3941bca2_1\",\"rawEndPinId\":\"pin-type-component_ca018356-08f3-4416-b12e-ca10c6c7bb67_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1479.3320000000_455.9255000000\\\",\\\"-1465.9160000000_455.9255000000\\\",\\\"-1465.9160000000_455.0000000000\\\",\\\"-1452.5000000000_455.0000000000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_0\",\"endPinId\":\"pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_1\",\"rawStartPinId\":\"pin-type-component_38df7453-f88c-4a99-82c0-fdb338cc7264_0\",\"rawEndPinId\":\"pin-type-component_7807e964-3bc8-4b12-bb6c-44a1c1b24af9_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1452.5000000000_530.0000000000\\\",\\\"-1465.9160000000_530.0000000000\\\",\\\"-1465.9160000000_530.9255000000\\\",\\\"-1479.3320000000_530.9255000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2\",\"endPinId\":\"pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2\",\"rawStartPinId\":\"pin-type-component_39ea5961-b6e7-49a0-8a1a-4a54142db333_2\",\"rawEndPinId\":\"pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_80.0000000000\\\",\\\"-1017.5000000000_80.0000000000\\\",\\\"-1017.5000000000_185.0000000000\\\",\\\"-1062.5000000000_185.0000000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1\",\"endPinId\":\"pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_0\",\"rawStartPinId\":\"pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1\",\"rawEndPinId\":\"pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-165.3277806029_458.9198741372\\\",\\\"-151.9117806029_458.9198741372\\\",\\\"-151.9117806029_457.9943741372\\\",\\\"-138.4957806029_457.9943741372\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1\",\"endPinId\":\"pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2\",\"rawStartPinId\":\"pin-type-component_3c883d29-f62b-49cf-a092-2c8c9f097c17_1\",\"rawEndPinId\":\"pin-type-component_f2a03157-3d3b-4891-9a96-ef7378eef59a_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-165.3277806029_458.9198741372\\\",\\\"-147.5000000000_458.9198741372\\\",\\\"-147.5000000000_492.5000000000\\\",\\\"-1062.5000000000_492.5000000000\\\",\\\"-1062.5000000000_185.0000000000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2\",\"endPinId\":\"pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2\",\"rawStartPinId\":\"pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2\",\"rawEndPinId\":\"pin-type-component_9e058603-a403-435e-a7b3-472988f8f796_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-40.0000000000\\\",\\\"-1017.5000000000_-40.0000000000\\\",\\\"-1017.5000000000_-145.0000000000\\\",\\\"-1062.5000000000_-145.0000000000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1\",\"endPinId\":\"pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_0\",\"rawStartPinId\":\"pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1\",\"rawEndPinId\":\"pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-165.3277806029_383.9198741372\\\",\\\"-151.9117806029_383.9198741372\\\",\\\"-151.9117806029_382.9943741372\\\",\\\"-138.4957806029_382.9943741372\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2\",\"endPinId\":\"pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1\",\"rawStartPinId\":\"pin-type-component_0fa29099-f06c-42e6-8abb-d829c961012c_2\",\"rawEndPinId\":\"pin-type-component_c525269a-6029-466e-8297-23d196a50c50_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-40.0000000000\\\",\\\"-1062.5000000000_-2.5000000000\\\",\\\"-882.5000000000_-2.5000000000\\\",\\\"-882.5000000000_417.5000000000\\\",\\\"-147.5000000000_417.5000000000\\\",\\\"-147.5000000000_383.9198741372\\\",\\\"-165.3277806029_383.9198741372\\\"]}\"}","{\"color\":\"#ff1100\",\"startPinId\":\"pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2\",\"endPinId\":\"pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2\",\"rawStartPinId\":\"pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2\",\"rawEndPinId\":\"pin-type-component_548ad9b0-6450-4235-a7be-ccb79cd6080d_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-340.0000000000\\\",\\\"-1017.5000000000_-340.0000000000\\\",\\\"-1017.5000000000_-445.0000000000\\\",\\\"-1062.5000000000_-445.0000000000\\\"]}\"}","{\"color\":\"#ff1100\",\"startPinId\":\"pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1\",\"endPinId\":\"pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_0\",\"rawStartPinId\":\"pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1\",\"rawEndPinId\":\"pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-165.3277806029_308.9198741372\\\",\\\"-151.9117806029_308.9198741372\\\",\\\"-151.9117806029_307.9943741372\\\",\\\"-138.4957806029_307.9943741372\\\"]}\"}","{\"color\":\"#ff1100\",\"startPinId\":\"pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2\",\"endPinId\":\"pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1\",\"rawStartPinId\":\"pin-type-component_19cbe39d-a790-4e2e-bde4-0d5ef7c61da2_2\",\"rawEndPinId\":\"pin-type-component_42b98079-caa9-47e9-bd5d-65893e0dce4d_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-340.0000000000\\\",\\\"-1062.5000000000_-317.5000000000\\\",\\\"-620.0000000000_-317.5000000000\\\",\\\"-620.0000000000_342.5000000000\\\",\\\"-165.3277806029_342.5000000000\\\",\\\"-165.3277806029_308.9198741372\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2\",\"endPinId\":\"pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2\",\"rawStartPinId\":\"pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2\",\"rawEndPinId\":\"pin-type-component_d7dc068c-4b59-400e-ae50-562c7ccbc1ad_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-565.0000000000\\\",\\\"-1017.5000000000_-565.0000000000\\\",\\\"-1017.5000000000_-685.0000000000\\\",\\\"-1062.5000000000_-685.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_1\",\"endPinId\":\"pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0\",\"rawStartPinId\":\"pin-type-component_5008935e-c93f-4fb4-a087-0abedc96eefb_1\",\"rawEndPinId\":\"pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-165.3277806029_233.9198741372\\\",\\\"-159.4117806029_233.9198741372\\\",\\\"-159.4117806029_232.9943741372\\\",\\\"-138.4957806029_232.9943741372\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2\",\"endPinId\":\"pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0\",\"rawStartPinId\":\"pin-type-component_0ad2680b-02ba-49a2-a3e9-a96381a7d26e_2\",\"rawEndPinId\":\"pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-1062.5000000000_-565.0000000000\\\",\\\"-1062.5000000000_-527.5000000000\\\",\\\"-860.0000000000_-527.5000000000\\\",\\\"-860.0000000000_-430.0000000000\\\",\\\"-605.0000000000_-430.0000000000\\\",\\\"-605.0000000000_192.5000000000\\\",\\\"-138.4957806029_192.5000000000\\\",\\\"-138.4957806029_232.9943741372\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_0\",\"endPinId\":\"pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_0\",\"rawEndPinId\":\"pin-type-component_f7984d9c-52aa-415e-b39c-e5fb625b93c2_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-70.0000000000\\\",\\\"-417.5000000000_515.0000000000\\\",\\\"-87.5000000000_515.0000000000\\\",\\\"-87.5000000000_457.9943741372\\\",\\\"-93.4957806029_457.9943741372\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_1\",\"endPinId\":\"pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_1\",\"rawEndPinId\":\"pin-type-component_c94229bb-b925-4416-b768-559f9d5d84b6_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-85.0000000000\\\",\\\"-440.0000000000_-85.0000000000\\\",\\\"-440.0000000000_537.5000000000\\\",\\\"-57.5000000000_537.5000000000\\\",\\\"-57.5000000000_382.9943741372\\\",\\\"-93.4957806029_382.9943741372\\\"]}\"}","{\"color\":\"#00AE7E\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_2\",\"endPinId\":\"pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_2\",\"rawEndPinId\":\"pin-type-component_662aa0ec-65ba-4d5d-a487-5ed33ea6d988_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-100.0000000000\\\",\\\"-447.5000000000_-100.0000000000\\\",\\\"-447.5000000000_110.0000000000\\\",\\\"-12.5000000000_110.0000000000\\\",\\\"-12.5000000000_307.9943741372\\\",\\\"-93.4957806029_307.9943741372\\\"]}\"}","{\"color\":\"#C28C9F\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_3\",\"endPinId\":\"pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_1\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_3\",\"rawEndPinId\":\"pin-type-component_b45ca744-aa2b-4e0a-b23d-32ff2cca7a14_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-417.5000000000_-115.0000000000\\\",\\\"-432.5000000000_-115.0000000000\\\",\\\"-432.5000000000_170.0000000000\\\",\\\"-50.0000000000_170.0000000000\\\",\\\"-50.0000000000_232.9943741372\\\",\\\"-93.4957806029_232.9943741372\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_0\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_fe152afb-21b1-47d5-b9c6-bd2b619f0439_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-850.0000000000\\\",\\\"-267.5000000000_-850.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_0\",\"endPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawStartPinId\":\"pin-type-component_13bb41c2-0891-49e2-a36d-a0e52211de2b_0\",\"rawEndPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-267.5000000000_-820.0000000000\\\",\\\"-237.5000000000_-820.0000000000\\\",\\\"-237.5000000000_-700.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_0\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_5d50f226-59dc-49dd-a79a-abbf5e3cb510_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-790.0000000000\\\",\\\"-267.5000000000_-790.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_0\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_58089c3e-bb30-4b9d-87df-71065baedba4_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-760.0000000000\\\",\\\"-267.5000000000_-760.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_0\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_824c2884-8b95-4bf2-9b1d-fc37145bfe37_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-865.0000000000\\\",\\\"-387.5000000000_-865.0000000000\\\",\\\"-387.5000000000_-850.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_0\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_e12ba4ec-e1ec-4be3-a465-c2fc7f1b0f00_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-865.0000000000\\\",\\\"-387.5000000000_-865.0000000000\\\",\\\"-387.5000000000_-820.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_0\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_a72804f7-e18d-407a-8183-98f8e53fe3d0_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-865.0000000000\\\",\\\"-387.5000000000_-865.0000000000\\\",\\\"-387.5000000000_-790.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_0\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_bf3dc0fb-dd6e-4c59-903b-6bbbab3fccf1_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-865.0000000000\\\",\\\"-387.5000000000_-865.0000000000\\\",\\\"-387.5000000000_-760.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_0\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_ed5c99e1-3753-4905-b880-1ffcf976d135_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-865.0000000000\\\",\\\"-522.5000000000_-865.0000000000\\\",\\\"-522.5000000000_-760.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_0\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_b68f3984-33e3-4099-9fd0-2bf2992dd7c5_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-865.0000000000\\\",\\\"-522.5000000000_-865.0000000000\\\",\\\"-522.5000000000_-790.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_0\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_b7e27884-48f5-44d6-9ad2-56da1f22ae1e_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-865.0000000000\\\",\\\"-522.5000000000_-865.0000000000\\\",\\\"-522.5000000000_-820.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_0\",\"endPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawStartPinId\":\"pin-type-component_07965d4a-3c19-478e-9e88-2147d6a70aba_0\",\"rawEndPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-522.5000000000_-850.0000000000\\\",\\\"-522.5000000000_-865.0000000000\\\",\\\"-237.5000000000_-865.0000000000\\\",\\\"-237.5000000000_-700.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_0\",\"endPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawStartPinId\":\"pin-type-component_1d1c2d9f-e2bf-4916-b8b3-7bed2f551ddf_0\",\"rawEndPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-642.5000000000_-850.0000000000\\\",\\\"-642.5000000000_-865.0000000000\\\",\\\"-237.5000000000_-865.0000000000\\\",\\\"-237.5000000000_-700.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_0\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_6b9ac4cf-8b15-40e0-9908-87be89d7dd12_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-865.0000000000\\\",\\\"-642.5000000000_-865.0000000000\\\",\\\"-642.5000000000_-820.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_0\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_6d10b9b7-629d-43f1-9a8c-9eb4ed2f0e88_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-865.0000000000\\\",\\\"-642.5000000000_-865.0000000000\\\",\\\"-642.5000000000_-790.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_0\",\"endPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawStartPinId\":\"pin-type-component_0e24347f-56a1-4fe8-a3eb-00f61ef717e3_0\",\"rawEndPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-642.5000000000_-760.0000000000\\\",\\\"-642.5000000000_-865.0000000000\\\",\\\"-237.5000000000_-865.0000000000\\\",\\\"-237.5000000000_-700.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16\",\"rawStartPinId\":\"pin-type-component_2d2c1fc2-9459-4e52-81e7-c39a9a7813f6_0\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-237.5000000000_-700.0000000000\\\",\\\"-237.5000000000_-715.0000000000\\\",\\\"-275.0000000000_-715.0000000000\\\",\\\"-275.0000000000_-520.0000000000\\\",\\\"-327.5000000000_-520.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_18\",\"rawStartPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_16\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_18\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-327.5000000000_-520.0000000000\\\",\\\"-297.5000000000_-520.0000000000\\\",\\\"-297.5000000000_-550.0000000000\\\",\\\"-327.5000000000_-550.0000000000\\\"]}\"}","{\"color\":\"#5FAD4E\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16\",\"endPinId\":\"pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16\",\"rawEndPinId\":\"pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-327.5000000000_-130.0000000000\\\",\\\"-222.5000000000_-130.0000000000\\\",\\\"-222.5000000000_-85.0000000000\\\"]}\"}","{\"color\":\"#5FAD4E\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16\",\"endPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_18\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_16\",\"rawEndPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_18\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-327.5000000000_-130.0000000000\\\",\\\"-297.5000000000_-130.0000000000\\\",\\\"-297.5000000000_-160.0000000000\\\",\\\"-327.5000000000_-160.0000000000\\\"]}\"}","{\"color\":\"#5FAD4E\",\"startPinId\":\"pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_6\",\"rawStartPinId\":\"pin-type-component_935ec2c0-76f9-4c06-a88a-d876d661b1e8_0\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-222.5000000000_-85.0000000000\\\",\\\"-222.5000000000_-130.0000000000\\\",\\\"152.5000000000_-130.0000000000\\\",\\\"152.5000000000_-430.0000000000\\\",\\\"332.5000000000_-430.0000000000\\\"]}\"}","{\"color\":\"#FF029D\",\"startPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_27\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_19\",\"rawStartPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_27\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_19\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"617.5000000000_-370.0000000000\\\",\\\"790.0000000000_-370.0000000000\\\",\\\"790.0000000000_-565.0000000000\\\",\\\"-327.5000000000_-565.0000000000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_26\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_20\",\"rawStartPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_26\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_20\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"617.5000000000_-385.0000000000\\\",\\\"775.0000000000_-385.0000000000\\\",\\\"775.0000000000_-580.0000000000\\\",\\\"-327.5000000000_-580.0000000000\\\"]}\"}","{\"color\":\"#FF74A3\",\"startPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_25\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_21\",\"rawStartPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_25\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_21\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"617.5000000000_-400.0000000000\\\",\\\"760.0000000000_-400.0000000000\\\",\\\"760.0000000000_-595.0000000000\\\",\\\"-327.5000000000_-595.0000000000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_24\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_22\",\"rawStartPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_24\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_22\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"617.5000000000_-415.0000000000\\\",\\\"745.0000000000_-415.0000000000\\\",\\\"745.0000000000_-610.0000000000\\\",\\\"-327.5000000000_-610.0000000000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_23\",\"endPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_23\",\"rawStartPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_23\",\"rawEndPinId\":\"pin-type-component_d448436c-9798-4335-8304-00153efa0c0f_23\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"617.5000000000_-439.0000000000\\\",\\\"730.0000000000_-439.0000000000\\\",\\\"730.0000000000_-625.0000000000\\\",\\\"-327.5000000000_-625.0000000000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_19\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_8\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_19\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_8\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-327.5000000000_-175.0000000000\\\",\\\"182.5000000000_-175.0000000000\\\",\\\"182.5000000000_-385.0000000000\\\",\\\"332.5000000000_-385.0000000000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_20\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_9\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_20\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-327.5000000000_-190.0000000000\\\",\\\"205.0000000000_-190.0000000000\\\",\\\"205.0000000000_-370.0000000000\\\",\\\"332.5000000000_-370.0000000000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_21\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_10\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_21\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_10\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-327.5000000000_-205.0000000000\\\",\\\"227.5000000000_-205.0000000000\\\",\\\"227.5000000000_-355.0000000000\\\",\\\"332.5000000000_-355.0000000000\\\"]}\"}","{\"color\":\"#BDC6FF\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_22\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_11\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_22\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_11\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-327.5000000000_-220.0000000000\\\",\\\"250.0000000000_-220.0000000000\\\",\\\"250.0000000000_-340.0000000000\\\",\\\"332.5000000000_-340.0000000000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_23\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_12\",\"rawStartPinId\":\"pin-type-component_11da4e6e-750e-4643-874f-89e7cea28441_23\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_12\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-327.5000000000_-235.0000000000\\\",\\\"272.5000000000_-235.0000000000\\\",\\\"272.5000000000_-325.0000000000\\\",\\\"332.5000000000_-325.0000000000\\\"]}\"}","{\"color\":\"#A5FFD2\",\"startPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_9\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_5\",\"rawStartPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_9\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"439.4500000000_-89.6500000000\\\",\\\"287.5000000000_-89.6500000000\\\",\\\"287.5000000000_-445.0000000000\\\",\\\"332.5000000000_-445.0000000000\\\"]}\"}","{\"color\":\"#08d46a\",\"startPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_11\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_22\",\"rawStartPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_11\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_22\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"439.4500000000_-69.1000000000\\\",\\\"422.5000000000_-69.1000000000\\\",\\\"422.5000000000_-10.0000000000\\\",\\\"715.0000000000_-10.0000000000\\\",\\\"715.0000000000_-454.0000000000\\\",\\\"617.5000000000_-454.0000000000\\\"]}\"}","{\"color\":\"#774D00\",\"startPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_12\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_29\",\"rawStartPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_12\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_29\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"439.4500000000_-58.3000000000\\\",\\\"407.5000000000_-58.3000000000\\\",\\\"407.5000000000_-2.5000000000\\\",\\\"730.0000000000_-2.5000000000\\\",\\\"730.0000000000_-340.0000000000\\\",\\\"617.5000000000_-340.0000000000\\\"]}\"}","{\"color\":\"#e11934\",\"startPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_1\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_21\",\"rawStartPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_1\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_21\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"542.6500000000_-89.5000000000\\\",\\\"655.0000000000_-89.5000000000\\\",\\\"655.0000000000_-469.0000000000\\\",\\\"617.5000000000_-469.0000000000\\\"]}\"}","{\"color\":\"#004754\",\"startPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_2\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_20\",\"rawStartPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_2\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_20\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"542.5000000000_-79.6000000000\\\",\\\"670.0000000000_-79.6000000000\\\",\\\"670.0000000000_-484.0000000000\\\",\\\"617.5000000000_-484.0000000000\\\"]}\"}","{\"color\":\"#B500FF\",\"startPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_3\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_19\",\"rawStartPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_3\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_19\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"542.9500000000_-68.9500000000\\\",\\\"685.0000000000_-68.9500000000\\\",\\\"685.0000000000_-499.0000000000\\\",\\\"617.5000000000_-499.0000000000\\\"]}\"}","{\"color\":\"#FFB167\",\"startPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_4\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_18\",\"rawStartPinId\":\"pin-type-component_0a8678a1-8b77-47ac-8524-d596b3cedd6d_4\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_18\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"542.9500000000_-58.6000000000\\\",\\\"700.0000000000_-58.6000000000\\\",\\\"700.0000000000_-514.0000000000\\\",\\\"617.5000000000_-514.0000000000\\\"]}\"}","{\"color\":\"#f73302\",\"startPinId\":\"pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_4\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_7\",\"rawStartPinId\":\"pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_4\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"527.5000000000_-940.0000000000\\\",\\\"527.5000000000_-857.5000000000\\\",\\\"227.5000000000_-857.5000000000\\\",\\\"227.5000000000_-415.0000000000\\\",\\\"332.5000000000_-415.0000000000\\\"]}\"}","{\"color\":\"#06f40a\",\"startPinId\":\"pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_3\",\"endPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_17\",\"rawStartPinId\":\"pin-type-component_6fe13b46-5e6b-4103-adfc-cce8f32c36a7_3\",\"rawEndPinId\":\"pin-type-component_9e84bb7d-bdbc-45f5-a0ed-5a200d52e2b9_17\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"505.0000000000_-940.0000000000\\\",\\\"505.0000000000_-842.5000000000\\\",\\\"647.5000000000_-842.5000000000\\\",\\\"647.5000000000_-529.0000000000\\\",\\\"617.5000000000_-529.0000000000\\\"]}\"}"],"projectDescription":""}PK
     ��Z               jsons/PK
     ��Z����� ��    jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"16 - Channel Analog Multiplexer","category":["User Defined"],"userDefined":true,"id":"b7d4df28-c430-b8ca-f42b-be40986a361e","subtypeDescription":"","subtypePic":"793ea4e6-6f4c-45cd-8a04-0920ddad3581.png","iconPic":"627c2b90-5d53-4228-8b10-5ea0a126027c.png","imageLocation":"local_cache","componentVersion":1,"pinInfo":{"numDisplayCols":"7.00000","numDisplayRows":"16.00000","pins":[{"uniquePinIdString":"0","positionMil":"50.00000,50.00000","isAnchorPin":true,"label":"C0"},{"uniquePinIdString":"1","positionMil":"50.00000,150.00000","isAnchorPin":false,"label":"C1"},{"uniquePinIdString":"2","positionMil":"50.00000,250.00000","isAnchorPin":false,"label":"C2"},{"uniquePinIdString":"3","positionMil":"50.00000,350.00000","isAnchorPin":false,"label":"C3"},{"uniquePinIdString":"4","positionMil":"50.00000,450.00000","isAnchorPin":false,"label":"C4"},{"uniquePinIdString":"5","positionMil":"50.00000,550.00000","isAnchorPin":false,"label":"C5"},{"uniquePinIdString":"6","positionMil":"50.00000,650.00000","isAnchorPin":false,"label":"C6"},{"uniquePinIdString":"7","positionMil":"50.00000,750.00000","isAnchorPin":false,"label":"C7"},{"uniquePinIdString":"8","positionMil":"50.00000,850.00000","isAnchorPin":false,"label":"C8"},{"uniquePinIdString":"9","positionMil":"50.00000,950.00000","isAnchorPin":false,"label":"C9"},{"uniquePinIdString":"10","positionMil":"50.00000,1050.00000","isAnchorPin":false,"label":"C10"},{"uniquePinIdString":"11","positionMil":"50.00000,1150.00000","isAnchorPin":false,"label":"C11"},{"uniquePinIdString":"12","positionMil":"50.00000,1250.00000","isAnchorPin":false,"label":"C12"},{"uniquePinIdString":"13","positionMil":"50.00000,1350.00000","isAnchorPin":false,"label":"C13"},{"uniquePinIdString":"14","positionMil":"50.00000,1450.00000","isAnchorPin":false,"label":"C14"},{"uniquePinIdString":"15","positionMil":"50.00000,1550.00000","isAnchorPin":false,"label":"C15"},{"uniquePinIdString":"16","positionMil":"650.00000,450.00000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"17","positionMil":"650.00000,550.00000","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"18","positionMil":"650.00000,650.00000","isAnchorPin":false,"label":"EN"},{"uniquePinIdString":"19","positionMil":"650.00000,750.00000","isAnchorPin":false,"label":"S0"},{"uniquePinIdString":"20","positionMil":"650.00000,850.00000","isAnchorPin":false,"label":"S1"},{"uniquePinIdString":"21","positionMil":"650.00000,950.00000","isAnchorPin":false,"label":"S2"},{"uniquePinIdString":"22","positionMil":"650.00000,1050.00000","isAnchorPin":false,"label":"S3"},{"uniquePinIdString":"23","positionMil":"650.00000,1150.00000","isAnchorPin":false,"label":"SIG"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"16 - Channel Analog Multiplexer","category":["User Defined"],"userDefined":true,"id":"b7d4df28-c430-b8ca-f42b-be40986a361e","subtypeDescription":"","subtypePic":"793ea4e6-6f4c-45cd-8a04-0920ddad3581.png","iconPic":"627c2b90-5d53-4228-8b10-5ea0a126027c.png","imageLocation":"local_cache","componentVersion":1,"pinInfo":{"numDisplayCols":"7.00000","numDisplayRows":"16.00000","pins":[{"uniquePinIdString":"0","positionMil":"50.00000,50.00000","isAnchorPin":true,"label":"C0"},{"uniquePinIdString":"1","positionMil":"50.00000,150.00000","isAnchorPin":false,"label":"C1"},{"uniquePinIdString":"2","positionMil":"50.00000,250.00000","isAnchorPin":false,"label":"C2"},{"uniquePinIdString":"3","positionMil":"50.00000,350.00000","isAnchorPin":false,"label":"C3"},{"uniquePinIdString":"4","positionMil":"50.00000,450.00000","isAnchorPin":false,"label":"C4"},{"uniquePinIdString":"5","positionMil":"50.00000,550.00000","isAnchorPin":false,"label":"C5"},{"uniquePinIdString":"6","positionMil":"50.00000,650.00000","isAnchorPin":false,"label":"C6"},{"uniquePinIdString":"7","positionMil":"50.00000,750.00000","isAnchorPin":false,"label":"C7"},{"uniquePinIdString":"8","positionMil":"50.00000,850.00000","isAnchorPin":false,"label":"C8"},{"uniquePinIdString":"9","positionMil":"50.00000,950.00000","isAnchorPin":false,"label":"C9"},{"uniquePinIdString":"10","positionMil":"50.00000,1050.00000","isAnchorPin":false,"label":"C10"},{"uniquePinIdString":"11","positionMil":"50.00000,1150.00000","isAnchorPin":false,"label":"C11"},{"uniquePinIdString":"12","positionMil":"50.00000,1250.00000","isAnchorPin":false,"label":"C12"},{"uniquePinIdString":"13","positionMil":"50.00000,1350.00000","isAnchorPin":false,"label":"C13"},{"uniquePinIdString":"14","positionMil":"50.00000,1450.00000","isAnchorPin":false,"label":"C14"},{"uniquePinIdString":"15","positionMil":"50.00000,1550.00000","isAnchorPin":false,"label":"C15"},{"uniquePinIdString":"16","positionMil":"650.00000,450.00000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"17","positionMil":"650.00000,550.00000","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"18","positionMil":"650.00000,650.00000","isAnchorPin":false,"label":"EN"},{"uniquePinIdString":"19","positionMil":"650.00000,750.00000","isAnchorPin":false,"label":"S0"},{"uniquePinIdString":"20","positionMil":"650.00000,850.00000","isAnchorPin":false,"label":"S1"},{"uniquePinIdString":"21","positionMil":"650.00000,950.00000","isAnchorPin":false,"label":"S2"},{"uniquePinIdString":"22","positionMil":"650.00000,1050.00000","isAnchorPin":false,"label":"S3"},{"uniquePinIdString":"23","positionMil":"650.00000,1150.00000","isAnchorPin":false,"label":"SIG"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Touch Sensor TTP233","category":["User Defined"],"id":"7529b28e-1847-4d84-acce-e52ea11a6606","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1c06f444-5387-4cb2-91f2-17a999ad4bd8.png","iconPic":"995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.66667","pins":[{"uniquePinIdString":"0","positionMil":"216.66667,500.00000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"316.66667,500.00000","isAnchorPin":false,"label":"I/O"},{"uniquePinIdString":"2","positionMil":"416.66667,500.00000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Switch Symbol SPST","category":["User Defined"],"id":"2d44b201-0eba-4542-b8d6-a72ddb6878af","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"6bfc6843-1883-4a57-a768-11efac5c5eb3.png","iconPic":"9d204b9c-624e-42df-9128-467635275a1c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.44065","numDisplayRows":"2.98954","pins":[{"uniquePinIdString":"0","positionMil":"6.53821,108.18463","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"927.65821,102.01463","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"LED_RED","category":["User Defined"],"id":"820a18f0-1f12-49e5-aa5e-d4450deb7c7d","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"3d3e563e-9ba6-48b4-a3f8-79399330dfef.png","iconPic":"89208456-78cc-4fe1-a1e6-da24e243623e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"302.99292,52.62506","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"2.99292,52.62506","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"GND","category":["User Defined"],"id":"d9393c8d-28d0-481b-9226-0c2455840b61","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"7260fbed-8271-43c5-b1e8-f8e9900a221b.png","iconPic":"e3aa425b-adcd-4ef1-9309-97e806748a2c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.35393","numDisplayRows":"5.10062","pins":[{"uniquePinIdString":"0","positionMil":"168.69222,444.59880","isAnchorPin":true,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Arduino UNO","category":["Microcontroller"],"userDefined":false,"id":"23db5403-7550-740c-a02b-8b3755757442","subtypeDescription":"","subtypePic":"0b351edc-7875-4477-b820-546ce15be531.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"LoRa Ra-02 SX1278","category":["User Defined"],"id":"ea67bc39-2543-48d1-915c-5686eed5bac4","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"ae1d0bb1-db79-4eca-b526-eb1d648f9ad0.png","iconPic":"1348d1eb-e6ae-43d4-937f-d455f2ad4bcd.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.31437","numDisplayRows":"12.64394","pins":[{"uniquePinIdString":"0","positionMil":"786.93229,632.75287","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"787.93229,562.75287","isAnchorPin":false,"label":"NSS"},{"uniquePinIdString":"2","positionMil":"786.93229,496.75287","isAnchorPin":false,"label":"MOSI"},{"uniquePinIdString":"3","positionMil":"789.93229,425.75287","isAnchorPin":false,"label":"MISO"},{"uniquePinIdString":"4","positionMil":"789.93229,356.75287","isAnchorPin":false,"label":"SCK"},{"uniquePinIdString":"5","positionMil":"788.93229,284.75287","isAnchorPin":false,"label":"D105"},{"uniquePinIdString":"6","positionMil":"783.93229,146.75287","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"785.93229,221.75287","isAnchorPin":false,"label":"DI04"},{"uniquePinIdString":"8","positionMil":"99.93229,630.75287","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"9","positionMil":"99.93229,563.75287","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"10","positionMil":"99.93229,496.75287","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"11","positionMil":"99.93229,426.75287","isAnchorPin":false,"label":"RST"},{"uniquePinIdString":"12","positionMil":"99.93229,354.75287","isAnchorPin":false,"label":"DI00"},{"uniquePinIdString":"13","positionMil":"99.93229,288.75287","isAnchorPin":false,"label":"DI01"},{"uniquePinIdString":"14","positionMil":"99.93229,216.75287","isAnchorPin":false,"label":"D102"},{"uniquePinIdString":"15","positionMil":"99.93229,145.75287","isAnchorPin":false,"label":"DI03"}],"pinType":"wired"},"properties":[]},{"subtypeName":"POWER SUPPLY 5V 5AMP","category":["User Defined"],"id":"646c8823-36b2-4192-89ce-6ec44eb47b6e","userDefined":true,"subtypeDescription":"","subtypePic":"483af35d-09f4-402a-a8a9-75c28eb4643f.png","pinInfo":{"numDisplayCols":"13.51513","numDisplayRows":"18.87938","pins":[{"uniquePinIdString":"0","positionMil":"335.96491,206.51286","isAnchorPin":true,"label":"220V Positive Pole (AC)"},{"uniquePinIdString":"1","positionMil":"485.96491,206.51286","isAnchorPin":false,"label":"220V Negative Pole (AC)"},{"uniquePinIdString":"2","positionMil":"635.96491,206.51286","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"3","positionMil":"785.96491,206.51286","isAnchorPin":false,"label":"GND (DC)"},{"uniquePinIdString":"4","positionMil":"935.96491,206.51286","isAnchorPin":false,"label":"12V-24V Output (DC)"}],"pinType":"wired"},"properties":[],"iconPic":"0a03a94b-1490-4d51-a356-eaee23e4f5f0.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"LED_GREEN","category":["User Defined"],"id":"6daab273-1bed-42a8-91c6-8d14a3f51d8d","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png","iconPic":"f39c2bb7-8598-4025-b62d-e677fac223ba.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"1.00000","pins":[{"uniquePinIdString":"0","positionMil":"-3.56139,47.00708","isAnchorPin":true,"label":"Anode"},{"uniquePinIdString":"1","positionMil":"296.43861,47.00708","isAnchorPin":false,"label":"Cathode"}],"pinType":"wired"},"properties":[]}]}PK
     ��Z               images/PK
     ��Z
�8b  8b  /   images/a7e3301e-fb46-458d-916f-a05c0bde95f4.png�PNG

   IHDR  �  �   ��O3   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���]l��}����%R�(��(�"mY�-?(˃���S�$]Ңht�:l��u����C�m�i˴�Л]�z�a7	$C
�hs5�r��b9�]�ReZ�����"��8�BQ<�����z��s>�o��/S  �laa�G�"⹈8Px� ����N�*=Z�7�7�^(=   ��.Eę��}��� "6K ��T�  ���=�"�E�gC�     t�LD|:���^8z��J ��� xU�s���C      �ӓ9�?>z��ϖ  M� ��������K�      �!�9��>??���C  `��  <P>�R���w      찱�����=Uz  �� �I�."z��      �TUU���8Qz  �� ��ѣG�^D�.�     `�����ߔ  �"p �����8�s���w      4�_=z���G  �0� x �u��#��;      ��9/�  � p �A�"⟖     РO�����  �iw  :onn�q��     �&���Xz  �4�;  ��R�g�7      𩹹��,=  v�� �N;r��#)�ϖ�     PBUU���  �Iw  :������     Fק���*=  v� �NK)���      JJ)���  `�� 謥����;      JJ)�Å��=�w  �N� �Yu]���      Z�@���K�  �� p ��r���     �6H)���  `'� 褣G�.F��K�      h��.--�(=  �� �N�9��     �6?_z  �/�;  ��s�L�      -��  ��� �E���'K�      h�g���N�  �C� @�,,,<ӥw      ��`0���  �~� �ϔ      �R�Pz   ��;  ]���      Z�������#  `��  tʣ�>�;"�)�     ��R]�~.  �%p �Snܸ�LD���     �bw  :K� @�|��      ������  �!p �k�      wwpaa�åG  �v� ���     ��L�  �w  :c~~���8\z     @��?[z  l�� ��H)=Wz     @���9v�؁�;  �^	� �ӥ      tD������#  �^	� ��;     ��?^z  �+�;  ]ы��Rz     @�|��   �W��  `+���zO�[UUU���݆Q��������p'ccc�k׮�3    �j}}��az�ȑ#�o�����C  `�7  tB]ק�z�~����1111>>����v�~����cccQUU�z=A;���<fggKπV���?O>�d�    [���q�֭�y�f���ō7�ڵkq�ڵ�~�z\�v-rΥ�ދ�~��\D|��  �*  ]�����XLOO���t�߿?���SSS�gOg�     ;dll,���bϞ=q���;>���o��V���ƛo��.]�˗/G]��ݺ���C� @�� ���LLL���|������LLMM��.     `D���8t�P:t�����|�r\�x1.]�/^��7o\�#>Qz   ��;  ]PE�������Ǐ�������     �]�^/>�~�sׯ_�.�믿���zlll\��7B�%G  �V	� h����G��ޭ>_UU;v,�񘙙�4     �199'N��'ND]ױ�����Z���q�����,..>�ꫯ�m�� `;�  ��`08���RJq�ĉ8u�T�ݻ�     `h����������ӧOǕ+W��^�������J#��pD� ��;  ��Rz_����8p �}����      m355SSS��OƵk��ܹs���/�[o�5���9�DD�ǡ�  � �;  ��s~�n__ZZ��~������     莽{�ƩS��ԩSq���x饗��_����}��҇w� `���  `��^_8~�x|���     �6==�>�l|��}�C199��/�����=;��  0,w  Z����c�؝�v�Сx��g#���*     ��ؽ{w<��S��}.>�āv�e����x!  6g. h�7�x㉈�u���>}:z�^Ë      ����8~�x?~<^y�8s�L\�zuۯ�s���x~� �p� h�������gggcvv��9      �{��cii)���ę3gb}}��_#���� ��� �vO��sssM�      (���x�������g�Ɵ�ٟE��^^���  ;�*=   ~�������ɦw      �{��x�gⓟ�dLLL��o=y�ر�a� ��"p ��N�      �6�����?��1;;���ҿu�����  ;A� @���x�N_�r�J�S      �eϞ=�O}*�����|J��C�  �M� @k-...Dľ;}mee��5      �������x���o�q�;  �'p ��r�'��k/^����&�      �RUU�},&''����  t�� �6{��="��_lj     @��޽;������9��GDjf  l�� �6�k�~�ܹXYYij     @�;v,�����ȁ������  �!p ���q<��󱶶��     �V��*:t�gRJw?�  �	� h����������矏����     �j9���SM�  ��� �VUD<������<������-     �k0ĥK���L��Ɇ�  ���K  �;YXXX���[}��W^����|�#����5     �����o����]�I)�� @��� @+UUu�^�+��_���bmmm�      Z���_�o~�[y��� �b�Y ��꺾��="bee%���/����NO     h��^z)����G]�[y|����C��  �%p ��rΏl��޸q#��կ�ٳg���      �s�ʕ��?����7�qO'�����,  �/��  �NRJۺ�~[]���o~3Ο?�=�\LOO��4     ���_���ַ⥗^�ֱ������/��2  �w  ����._�_��W�G�~��111�/     Ш�s\�p!�����������>�S�  `�	� h�	�#������w������O�O<�w�ީ�     �����p�B���k�ꫯ����N��� ��� �:���;��q�������'O���'O��     ����f\�|9.^�.\�����x����  ��  �N��{h�����/��b|�[ߊ�z(N�<��[     ����㭷ފ���������t�R\�|9�n������YYYy��7 �{!p �u��Zl�}꺎s��Źs�b߾}q�ĉ8v�X�ݻ���     F���f\�v-�^�������o��V\�r��������c!p �u�  ��R�ox���8s�L�9s&<KKK�����R�s     ��X[[��7o�͛7�ƍq��ոv�Z\�~=�]�kkk�'���"���  �&p �����^�|��x��7�^�]�v���\������L8p �}�F    �����X__�[�n��������vȾ��7n܈����W��GJ��  �N�9  �Q��������{��^|�{ߋ����bjj*���SSS�o߾����ݻw���x���^     �����9G�9666""b0�����u]���f�����ǃ� ����3d���,�?�Qu]� h%�;  m�Tz�{��:VWWcuu�=���z���\���c����X��J_��W��ٳ�g    r;Dg�\p ���  �Qk.�o���/�hx�(��ݾ~   @+=)"r�!  �NU�  p���     ���\\\\(=  �M� @����싈��;      F�c�  ��	� h�~��z;     @��� ��� �*UU-��      0
RJ���   �&p �m\p     h�#�  ��	� h�;     @3�  ��� ��Y,=      `D/=   �M� @��     �1}�����G  �;	� h���      Fŭ[����   �$p �m\p     hH����  ���  ����̾��*�     `T���  ��� �������      0J\p �m�  �FJi��     �s��   x'�;  ��RZ*�     `ĸ� @�� h���      F̱�H�G  �mw  �d��      ����ѣӥG  �mw  Z#�t��     ��Tz   �&p �5rγ�7      ����  �6�;  m�;     @��  ��� �6�     4��룥7  �mw  Z�رc�1Uz     ��I)�� @k� h������      F�� ��� �
u])�     `D-�   �	� h�^��;     @.� �w  Z!��;     @�=����#   B� @{��     PH]׮� �
w  Z!�,p     (dssS� @+� h��ґ�      FUJI� @+� h�     
� �w  ��w     �r�  ��� ��p�     ��;  � p ���8Tz     �� �
w  �;r��LD�K�      aK�  @�� �v�-=      `�훞��*=  �  ������      0�v�ڵXz  � (.��;     @aUU	� (N� @q9g�     �[*=   �  WU��      �� @qw  ��9.�     �8Zz   � h�;     @y�  �� �6�.=      `��gKo   �;  m p     (,�t��  � �w     ��\p �8�;  mp��       bbfff_�  �6�;  E9rd2"�K�       b||�H�  �6�;  E�z���      ����gKo  `�	� (*�$p     h����  %p �4�;     @KTU%p �(�;  E�u-p     h���l�  �6�;  E����      ���  %p �4�     Z"�|��  F�� ��\p     h����  %p �����      ��;  E	� (��k�;     @{�� @Qw  �r�     �U<�裻K�  `t	� (M�     ���͛�K�  `t	� (M�     �"9���  ]w  J�     �H]�GJo  `t	� (�駟�{K�      �/�z=� (F� @1+++��     �L��w  �� PL���     ���  #p �����      -�Rr� �b�  �$p     h����  #p �����     �}\p ��;  %	�     ��w  �� PL��@�      ����H�G  0��  �R�*�     �16==���  F�� �br�w     �;Tz  �I� @1.�     �SUUӥ7  0��  �s�_z      ?*�$p ��;  ��]p     h'�;  E� (&�$p     h!� (E� @Iw     �v� P�� ���      -T׵� �"�  �ҋ���#      �Q)%�;  E� (�رc�""��     �	� (B� @�n��_z      �I� @w  ���zS�7      ��  !p �����      �%p ��;  E�     Z�PD��#  =w  ���J�     �^c333{K�  `�� ("�,p     h������  =w  �p�     ��RJw  'p ��     �M� @	w  �H)	�     �M� @��  �;     @��u-p �qw  ��     �ޡ�  =w  �H)	�     Z,�t��  F�� �R��      �]M�  ��� P��      �&p �qw  J�     ��� ��	� (E�     �b)%�;  �� PB{K�      ����  ��� и����J�      ��  ��� и��I��     �o��G�]z  �E� @�rΓ�7      ��]�vm��  F�� ��	�     �allL� @��  4N�     ���@� @��  � p     耪����  �h� �8�     ���k� h�� ��      �s� �(�;  %�     : ����  F�� ��UU%p     � � h�� ��      �R� �(�;  ��9�     �A� @��  � p     ���  0Z�  � p     �� h�� ��      �R� �(�;  %�     : 缿�  F�� ����      ��;  M� и���      �s� �(�;  �s�     �3��  �h� P��     ��'J�  `t� (A�     ����S�7  0:�  � p     �]�v	� h�� ��U1^z      [3���  ��� ШÇTz      [SU��  4F� @�RJ��7      �u9g�;  �� �(�;     @������  ��� Ш��1�;     @��� @��  4*�,p     萔�� ��� h��     �C\p �Iw  �;     @�� h�� ���)=      ��K)�/� ��!p �i�      pO��^  #p �Q)���      �'w  #p �iw     �n� ��;  ���Z�     �-w  #p �Q)%�;     @����  4F� @��      �s� ��;  M�     t�� ��� hTJI�     �-{""� �h� Ш���      �R-..�;  !p �Q)���      �7u]O��  �h� �4�=      :&�,p �w  �&p     ��;  M� �4�;     @�� h�� �F���      ������  �h� Ш���     �{\p �w  �6Qz       �&�,p �w  ��;     @�� h�� ��	�     �G� @#�  4M�     �=w  !p �iw     ���9� h�� �&��      �"p �w  3333Qz      ���*�;  �� И~�?^z      �.�,p �w  SU��     ���  4B� @c�      �%p �w  �$p     �&�;  �� И��M�;     @7	� h�� �Ƥ�&Jo      `[�  4B� @cRJ.�     t�� �F� h��     ����  �h� И����      ؖ=�  0�  4��k�;     @7�N�>=Vz  >�;  �I)�*�     ��y�W�Ko  ��'p �1w     �����w  �N� @cr�~l%     @GUU%p `��  4�w     ��J)M��  ��O� @c��     tTJ�w  �N� @c\p     �4�;  C'p �19��      ؞�` p `��  4�w     ��J)	� :�;  �I)��     �]w  �N� @cr�.�     t��  4A� @��      �%p `��  4�w     ���Z� ��	� hLJI�     �Q)%�;  C'p �1)���      �6�;  C'p �19g�     �K� ��	� h��     ��RJ�Ko  ��'p �Iw  ��ha    IDAT   �����w  �N� @��      �R�(� ��� ����Jo      `�\p `��  4&��;     @w	� :�;  M�     t�� ��� �$�;     @G���  �� �&	�     :*�,p `��  4i��       �M� ��	� h��      �%p `��  4I�     �]w  �N� @��      �%p `��  4i��       �M� ��	� hJ?|�	     �ew  ��_z��Z^^���z����ґ�����@UU�1Q����R*��-�@D��Ǜ)�A�y="�kq3���s^����N (f}}�������g      �MUUM-//���; �aUJi<�<����kWD�RJ�rν��w5"���=�9窪V#�f]�k?��r���^�wq0\��_��K�w�"��}�K_ZJ)=]����HD����"b|0DDD�9""RJ?�1�u���V?       �v9�^���Z 5��~x�c�1��v����v㻼���"���nD�\U՟���W~�W�7�yT�w�o��o���깈x6">�r��  �w�      �)�9g��Q2O�������:""���W#�ň��񍺮������_����6����Ω�ҧ"��\D�� �j���     ���ATUUz @������^UU,//�DğD���9��~��^,����[�{��{677&��3񩈘+�	 �K�d     ��s� �f#��"��RJ���|!"��s�r����������:A�~��[�����?�s��`0�k)��қ  ��v     t�`0(= �K�"�SJ�86�����R�������7~�7^/=�������9��9����l���G  ;@�     �}�� `��"�r�?���������?�9��]�v��_��_�Rz\���#"眖��2��Ku]����(�	 �A�s����}�eg]�߳ϝ	I�$Pe����ش�VQ���"(-��ը���ҁ{�3#Jr@��9�d���j��"�6`*��,|c�l�4�,�$& M($s3q^�~�G��I2/����}���]k��������^��]:      [d�; �XT9��F�s�9r�`0�����f�d3�������������L)}M�<  ��4     ���� 0vgG�����8~�����ѣ���׼����2��<��녈�ќ�9��  ��     ��w ���g)���:�+���[��:����ҡ�6S����_\U՞�h�҈�� 0K�     �Ϟ ���~�h4z�`0xw]�����sK�\M���{����)�+"��J� �E�y      ��= �Fu"�������`����~fqq��5iS]pEľ�����
�       �V��t �Y�����}0�^J銥����4)SYp_�Rzm������\  �0��      �g� ��/�9�`0��N��waa�s�C��T�{������WD��s��� �?��	     �~�Ѩt  "���l4����:�������C�KU:�������*"���v �m&�\:      [d� ��rnJ�ʺ�?9_T:̸�~����r4��/+� �S��	     �~&� lKO�9�w0�nJ駖����t��h���s���F���v �mN�     ����  lk/�9|8�"�J�٬V��������9�_���K� ��rΥ#      �E&� l{��i8~`8>�t��h]�}8^RUխ���Y  X?�<      �Ϟ @k<?����`𓥃l�\� 뵲�����9����Y  �8�     ��w �V9?"���F?�w�ރ��G+&���:��M�� �R�y      ��= �VzY�ӹy����*d=�}�}m,��qQ�,  l��N     ���� �Z�����u�����N�����ڵ�@�����  �u9��      آ�hT:  �����~0����՟��zGJ:�m9���o|����@� `z��     �~�|  ��ڵ돮��'�r2ۮ������s�Λ#�y��  0>&�     ��	�  �!���cǎ}���?�t�G�V�~���)�E�SJg `�L�      h?{>  S�))�?ۿ�w�r�mSp����>����8�t  ��w     ��3� `��WU��~����A���~��;���xL�,  L�i      �g� `*�L)�z���]:H�6(��=)�k�C  &�b'     @��� �ZUJ���`pE� %/����F�J�  4#�\:      [4�JG  `�^7�*�X�}0�.�T�? ���     �~�|  �_�y�`0(6ļH�����"���z  �c�;     @��� 03��u��x����2�te�� �,�<      ��P# �ّR�r0,5}�F��ಔҵM^ ���b'     @�;v�t  ��?��+�����6yM  �w     ���� 0sRD��.x#)��߿���;#����  �~,v     ��= ��ԩ��7����k�b/����\PU�{"b~�� `���	     �~u]��  @9�s������I_k�����]�N���I^        �<C�  f�W��ͽweee�$/2��{�9u:�_��gL�  ���N        h�g��ͽ#�&u��������dR� �]�     گ���  (,����p�<��O������-��I�        (C� �5o�9���ྲ�rAD�fD̍��  ��	�      �g� �5U��k���x�'��zU��y{J���</  �g�     ����  p\J��UU���덵�>֓���w#���<'        �=�u]:  �HJ�[�=�ܥq�sl��`����q� ��b�     @��� ��RJoX뒏�X
��]w�Y����9�� 0},v       �T�����3�����~�ȑ+"�_��\        ��T�u�  lO_}����8N���p8|fD,�!  S�w     ��Sp �TRJ{����z�-ܯ���9�GĎ� `�)�       �T���_�����-�R�}uu�?F�3�r        �Lp ��y���Wn��.�_s�5O�9_��� 0;Lp     h?w  ��u+++l��M܏;֏��7{<  �E�     ����  ����z�f�T�}���ύ���E          �N)���:����{UU�#"m�X        ���. �vHUU]�s�p�|���`��ƍ �l��	     �~�|  ؀��n�m��~�7t"��7z           fKJ�M�^on#�l��~�w�<".�P*  ���s�      l�	�  l�����d#���6�}�F @��;     �4Pp `~f#S��]p��;~0"���H  �<w     ���� �&<u׮]�a�_^W�}mz��l:  3/�T:      [�� �f�_��I?�u�o����o)  3��*     �O� �Mz�Z'���UpO)-n-        0�� ؤ��|���p�����-� `�Y�     ��}  ،�ҿ���g쥟���s�=�H  �2�      ���  �UU���-����\/["  f��N     ��P�u�  �T������)���>77���1�T        @k)� �;:�Ώ���,��S���          ��X�9���S�8���D        Z�w  �����N��)�u]�|2y           �a�쪟�����/�X           f�K����O��I�v�zaD�h$        �urΥ#  �~�u]��d����s�d�y           �a'�?�����Ή�N<           3)��=�~��G���������1�H*           fN������G����{J�I        �Nιt  �DUU/x�{�|#���<  lUJ�t        `�9� ���b��
����9���          �z�`0���xX�����l           f�N|Q=��om.           �,��-'�~��~�7tRJ��|$  fAJ�t        `�y�7��9�⡂�w��8�H$           f�y��v�3���N����          `���겟Xp��Y           �a)������g� ��H)��      ��KG  `�\|�UD�u�]w^D��bq           �UO�ꪫΏX+�>|��0R          ����;w>+b���*          �6��6b���R��e�  0�R��      �i�s. ����k�����f `�)�        ��Rzz�?LpWp          ���+++�"�+
� `�yT%        p_y�uםW���=�t        �6 `R>�UU]�O* ��R*        �ƪ�zR�Rzb�         @;�� ���u��*"�          (�UD\P:           �-���*"�Q�   L��R�        �6�s~\�+        h��s�  L����;           ��㪈xl�           ̼�V9�sK�  `���JG      `��  0A�V)��S  0�,t        g��J)�,� ���        ���*�l�;        �. 0A;���+� ��g�     `:�� `�vTq�t
  �_UU�#      0
�  L��*�t�t
  ���N     ��`� �	:Z圏�N ����	        ���*�l�;  ��     0��  0AG���j�  L?�      ӡ���  �^�W��)  �~
�      ���  ��R�b_, ��g�     `:�� `Rr�_4� �FX�        N'���*"�_�   L?w     ��`� �II)}���ϖ ����	     0��  0)9绪���t  ���N     ��`� �	��J)�Y:  ��B'     �t�� �����4� �FX�        N'�|Wu����J `�)�     L�>  L�h4��ڷo߽�w��  0�,t     �_Jɾ  ��}���[���T�(  L=�      �g� �I�9*"���H)�U�8  L;��        ���W9�O�� ������_     `[3� �	�ˈ�����Y  �v;     �Ϟ  ��s�h�Z���ѣ�DD.� ��f�     ����  0!ynn�ck�}����.	 ��f�     ����  0!���𥈵���[
� `X�        N����P�=���2Y        �60� �	���?N,��L  fAUUg�      ۚ=  &�.�Cw���w��"�`�8  L=�<      �Ϟ  ������_<Tp��z�RJ.�	 �ig�     ����  0�����g����<  ���        �I�ɉ/Vp����� ��Pp     h?{>  �[J��'�~X�}yy�/"�F 0,v     ��=  ��s������7VpO)���F# 0��:�      ��� �����:�9Y����        ���;  �s~�#�{T�}uu��#��F 03:�N�      l��� 0.)�C9�?x�������z��w  ��b'     @�j ���߻������j�k�y  �1
�      �R* �)�R:ig��-�����E��D 0S�     ��w  �!�t����?�g'm�z�C��&�
 ����     �~&� 0u]�{yy���}vʖQJ魓� ��Qp     h?{>  ��)�ꧼ�\\\�����$�  0{L�      h?w  ��o�����Mp�)��O&  ���锎      �)� 0oI)�S}x�;Δ�["���# 0sLp     h?w  ��hUUo=�N{ǹ��xWD�8�H  �$�     �O� �-�����)��3�|���  0�,v     ���F  lEJ���3�����?>�D  ̬�R�      l�=  ��楥�������Ѽf�a  �q�y      ���� ���|i]w�^x��-� `���     �~
�  lҧWWWߵ�/����K/��V��	 �Yf�     ����  �9�_��z����u�q��Ͽ#"n�l(  f��N     ����^  6*�t����������[F�_~�є�U�� ��Sp     h�N�S:  ���^�wd�_�P���O~�/�?��L  �:w     ��3� ������[6r��ZF�^z�(�t��2 ����<     ��P#  6"����/���F���g��}wD|x�� 0��     گ�锎  @{�����=h�R�/"�&� `F)�     ���  �)G�rJiÝ�Mܻ��"�77s,  ��D     �v����� `���~c�s�a����z1"����  �=      �M� �u8�Rڳك7}ǹgϞ��9�a�� 0{Lp     h7w  �$�����Ż6{���8�;�k"��[9  ��w     �vSp �>>??�VN��;��/��hJ�#��V� �l��	     �n�{  8�c�c�_~����[��\ZZ�hJ�ꭞ ����tJG      `<� ��t����Փ��O*w��qeD|b� `zY�     h7�  8�������8�X
�w�>�s�ш��8y  ��O     �v���ԍ  �.Gs�?�����8N6�;���古�^7�� 0}Lp     h7w  N������q�l�w�|SD��8�	 ��0�     ��� x�]x�+�<�X�8{�^=�~8"�0�� 0Lp     h7�=  �����.����8O:�?�ܻw�9�E�X� �~&z      ��'� ��������{�O<������SJWN��  ��O     �v�� ���v���O�������Ɯ�oM��  ��O     �v��^  "�w����4��O�3���:���['u  �ł'     @���͕�  @Y��ܹ�R��&�0ڽ{�}�N�E��I^ �v0�     ����  ̴{�~��ݻ��E&>BsaaᶈxaD�?�k ����     �n�� 0�H)}��={>=�5r���vo����Q� `{��	     �n ̤QD�����MM\���Q�۽1"~,"rS� `{��J     �v�� 0srD��Z�����v�o�9���k �}X�     h7�=  3g_��}s�l�����|]����.  �UU㷟      ����\�  4��nw�-�0Z^^����ĵ (�D     �v�� 0r΃n����.6Bsyyy9"^_��  4ς'     @�yb/ �Lؿ��.��g�۽2缯d  ���     �^UUEJ�t  &(����v���P�O*���WRJ��Kg `��     ��^ �T�)�奥���ˋ�#"���)������  09Y	     �^
�  S�X��'�����Dl��{D���ү��^��� �dX�     h/{=  S��������_)�mSp��XZZ�ú��w�� ��Y�     h�����  �;���n����AN��
�{��e�ΝGćJg `��     ګ��]� �ͻ���|ݞ={n)䑶�]��ݻ�޹s�wD��Jg `|�     ��^ �������maa�s���̶}n��ݻG������)�AD�H\�    IDATU:  [c�     ����m� ��9�s�.//�b� ��-'��hyy���ƈ�t�,  l��V     ��aF  �R�#���۽�т�{DĞ={n9v�س#���Y  �<��      �e� @k�x���g,--�T:�z��A���7"�w8^�s�>"W:  ��     �^ss�� ��"b���t��hݟU.--�+"�6"��t  6F�     ����  �������m+�G�����vo_]]}~D�:"VK� `}<�     ��� Za5"^����M���]:�f���A�^���kWVV���t������ ��yl%     @{)� l{���v�����o�ݻ��q�`0xID\O*	 �S0�     ��� ��;#�U�n���A�ajF�n����է��E���y  x4��      �e� `{I)J)��F�����1�O���E���W_�ku]_?ST� h;��      �e� `����,,,�V:̸MU�����Ż"��~���RJWD�K#"� 0���     ���; ��������vo.dR���~�������K���3s�?��� 0�����     `�)� ����~vqq��K���h---�E<XtND��9�8"� hXUU�R��s�(      l��; @���{"b����M��4e&
�ǭ��}Ɂ�Z���r�?g�� 0K����hT:      �i�  �9����iaaᓥ�4m&�:>�:p������҈xUD\T8 �L���Sp     h!� &��9��r�Yg�e���w�S�L܏[XX�RD������9�����.��F�Y�� L-�      �d�; �D��߫���C�}���ե��3"�~>8p��c�����e���ʦ �.
�      �� 0V7G�;v����Y��~2�:am���Fį��D�Kr�/N)����� �"�      �d� `KF9���RzOD���vo/h�r�yk�8"��`0��ҋr���_V6 @;Y�     h'�<  ��������rο���|O�@m�s����=�x[�׫�9�g���=�������xlр  -��x(     @�ر�t ���K������СC��zu�Pm��	k�h����s��k��꺮����礔.���"�ܢA �!�=      ��> �����9�RU�MUU}�կ~�_��r�`m�s�~?��󶈈^�W���_u�ر����RJO�������'� �L2�     ��<� �AG#�o#�o"�orΟ��O���}��{����Jd�:
��������<⳹��?��ǎ{|J�	)�'�u��qVUU��9?&"Ύ��a
�vw,"��.�9?����D�h���	?D�߯� 3�ȑ#�O*�     ���9�N<8� fI'"��:�:᧳��s�{;"b5">Q #�s(�r�联���u�ň8\U�=9���??77w����{w��;V �LSp/`��sk?  3�.xgD|�      l�[��֟���?�K�  `�U�  0s(      �����P�  L?w  ����      �qw�}�}  &N� �F�-|     �ϑ�8V:  �O� ��=P:       f� �F(� Ш��Lp     h�C�  0� hT�Y�     �eRJ&� �w  �f�     �er��x  h��;  M3�     �eRJ�Jg  `6(� Ш���;     @˘� @S� h��O     ��1� �F(� ШN�c�;     @�b @#� h��W     ��=  �� @�Lp     h�C�  0� h��      �c� �F(� Ш��	�      �c�;  �Pp �Q9g�=      ��  �Pp �Q���w     ��Qp �
�  4j~~^�     �}� h��;  �:��-~     �ϡ�  �
�  4��[o=��9      �C�  h��;  %.      �1� �F(� P�	      -�s�� @#� (�(     @��� �
�  �`     �ERJ��3  0� (���      X?w  ��� @	�J      `������  �lPp ��     Z����7� �F(� P��;     @{�{���  �Pp ��C�      �n�"�. �٠� @	&|      ����  �
�  4.�d�;     @{��  ��Pp ��     �C� ��(� P�	�      �� @c� h\]�&�     �DJ�`�  �w  J0�     �%r�&� �w  J0�     �=� h��;  %��     �K  `v(� и��	�      -�R2� ��(� P��;     @K�u�� @c� (�P�       ��	�  4I� �ƥ�Lp     hw  �� @	&�     �DJ�`�  �w  ��tLp     h���Mp �1
�  4n׮]
�      -�RRp �1
�  4��[o=�J�      ��RJKg  `v(� Pʡ�      8���Lp �1
�  �r�       ���Ç� h��;  ���     �sssKg  `v(� P�	�      �_���~���!  �
�  �b�;  ��ۻ�9ӳ������n�7Yd��,k,Y���@H��D�!eI@BBd�a�r��d�'$�x�v������~� ��C���y��kg�]��޼���.   �w��ҲG  �>�  dq�     �w�  �^�  d�     ��N�   ֋� �,��      �J.� �Tw  ���     й�� �Tw  Rx3     �����  ��;  )�q���     ����;  K%p  ED�     :�Z��� ��"p  ��     ��5� X*�;  )�q�     t."�  ,�� �.�     L���  ��;  )�      �s� �e� �b�ϲ7      �r�5�;  K%p  ��      ������  �z� �b�;     @��qt� ��� ����w     ���� �R	� H�����2f�      ��Ο?�;  K%p  �XJ��=     �:���z�= ��"p  ӝ�      ����  ��;  �>�      �d  `�� ��;     @�"B� ��	� �$p     �Tk�v�  ֏� �Lw     �N��\p `��  d�     t*"\p `��  �i�	�     ��;  K'p  MD�     :w  �N� @�;     @�Zk��7  �~�  ����      <��  d� ��w     �~�� @�;  i�      ���w  �N� @�q�      ��A� ��	� H�;     @����ogo  `�� HSk�     tjcc�w  �N� @�Ǐ�     �Ԯ^��Y�  ֏� �4��̛�      }�[J9� ��� �f{{���Ҳw      �7�  ���  d:*���     �� H!p  ���      |�� �w  �d      ��  �� ��w     ��� H!p  ��     �?w  R� �&p     �� �w  �	�     �#p  �� �T�5�;     @gZkw  R� H�      ��;  )�  �r�     �?�8
� H!p  U�U�     ЙǏ� H!p  ��      �y|�֭;�#  XOw  R��(p     �˭RJ� �z� �j6�	�     �r3{   �K� @���#�;     @_�  �� ��_���     �/w  �� Hu���ǥ���;      �w  �� �+�      �� �F� @�      �� �F� @�      �� �F� @�֚�     �w  �� Hw     �N���  �� ��;     @'�  d� ��w     �~��(p  �� �t����      �֗����do  `}	� H�Zs�     ��.]z�= ��%p  ]�U�     Ё���� ��&p  ]k�V�      Ji����  �z� ��@      ���  �z� ��;     @�  �� ����X�     Ё֚� �Tw  �-�{���;      �]D� H%p ���      ������  �z� Ћ��      ��8�.� �J� @/�      �j�w  R	� ��~�      �u���)p  �� �.��\p     �������#  Xow  z!p     ��z;  ��  t��*p     H�Z� �N� @/�      �"b/{  � �BD�go      Xs.� �N� @/\p     H�Z� �N� @/�      �"B� @:�;  ]��
�     	� �� �.\�z�v)�({     ���q/{  � �E+��&{     ������ @:�;  =��=      `]mnn
� H'p �'w     �/_�|�=  �  �d?{      ��r� �.� ��      	Zkw  � p �'w     �!p �w  z"p     ȱ�=   J� ��;     @�֚�  tA� @O��      ���� ��;  ���)     @�k�  ��;  9::�     $h�ͳ7  @)w  �"p     H0���  tA� @7�ŽR���      k�p�X��  �� �+�      Kۥ���  J� ��;     �r]�   �� ��;     �����  �sw  ��Z�     ,��  tC� @W"B�     �\.� ��;  ]�     ,�� �n� ��8�w     �庖=   >'p �+���     `��� @7�  te�     ��p�X��  �� Е�
�     �g^Ji�#  �sw  �r�ƍ���{�;      �AD̳7  ���  ��z�      �u�Z� ��;  =Zd      Xײ  ���  �h/{      ��p� ��� �Nk�w     ��� ��;  ݉�;     �r\�   O� �#�;     ��� @W�  t��&p     8{����F�  x�� ��D��     ���K)-{  <M� @wj�w     �3��  �,�;  ��q;{     ��k�meo  �g	� ������Rʭ�      +���  �,�;  ��      g("�  tG� @�Zkw     �3�Z���  �%p �Wײ      ��Z��  tG� @�j���      V��|>��  �� Х��<{     �
�*���#  �Yw  z%p     8;�f  ��� Ыk�      V�� �.	� �����     ��� �� �.-�{����;      VQk�r�  x�;  ݊�y�     �UTk�u�  x�;  �j�	�     ����� �.	� �ٵ�      +ho�N�  x�;  =��      ��~�=   ^d�=   ^b�Z+��� /t���rpp�=���ѣ2�c�    �Rk-E� @��  t��6?<<�]������׳g@��Ey��a�    ��/}��R>��  /R�  ���֮eo      X5�V� �� �n	�     N�� �n	� ������Z���      �""������  �"w  z��      �
"��Rv����do �� е����      �
��d�  ��� е��V�     �U�����  �2w  �VkuE     �<��.p �kw  ����     `DD��;  ]� е�l�MV     �S�$p�8{  ��� ��=z��'_�	     �[���������  /#p �k7nܸ�;      V�/J)-{  ��� �)pI     �-DD��^��  �"p �{�֭�      S�����  �*w  ��Z�${     ���ZK)���  �*w  �7�k"      o��Zj�>s �{w  �7�k"      o!"������;  �U�  tocc�W�=     `�"�J)c�  x�;  ݻr��^��a�     ������  pw  ��E�N�     �)�����G�;  �$�  L�V�      �)� 0%w  &�����      Smss�g�;  �$�  L�0���      0E����u;{  ��� ���yDdo      ��Z�G�  ��  L�0��     ���(�0|��  NJ� �$���Ok���w      LI����x1{  ��� ��8��ne�      ��Zk���d�  ��� 0�q�     �)�����ٹ��  NJ� �d��Q�     �)q� ��� 0%��     �$"��Z��  ^�: �ɨ�
�     N���*�w  ��P 0��엵�1{     ��Z˹s�~��  ^�� �����zW�w      LA�u�ʕ+��;  �u� ��a~��     `
�a�Q�  x]w  �惈��      еZk)��w�  x]w  &����'o�     ���w  &G �������     ��axx���w  ��R 0)����Z���      =����ҥK��w  ��� 05���Q�     �^ED��~/{  �	�;  �DD�     �.�P"���;  �M� ����Ok�(     �<�0���d�  �7�
 `���     <_D\��緲w  ��P 09���G�0<��     Л�(����  oJ� ��\�x�q����      ����R���  oJ� �$E�k�8     �ak����  oJ �$��~$p     �]�0|o>�?��  oJ �$���'_�	     @)��g'���  oC� �$]�v�r�u?{     @/�a(�n�  xw  ��E�k�H     PJ)�ֽ���f�  ��� `���     �����RJ��  oC �d�����0d�      H7��J)�;�;  �m	� ������#� {     @�Z��W����w  ��� 0e���Z=�     ��Z�a�ǋ/>��  oK	 ��E�{�0d�      H�䳒�d�  �� p `�Zk��;     ��f���Rʻ�;  �4(�  ����݋�0lg�      �Pk-�͝����[  �4� ��VJ��'_�	     �Vf�Y���g�  ��"p `���     XG�0�r{{��;  �� X��� {     �2=������o� �� p `�vvv�R��V��     ��������7�w  �iR  �*�9�Ͳ7      ,E����wׯ__do ��$p `%Dķ�a���     `f��8���d�  ��&p `%���܏����#.     ��"��f�o���}��  N�� ��Qk��l6˞     p�666Jk�w  �Y� �2���{��̥     `eED���������-  p�  ���Z�+W�    �U���qw�?��  gE� �J�����l6�u�     ����c�  �IDAT6C��/���v�  8+w  V�q��/�a��     p�Ν;�㝝����  gI� ��������s��-{     �i����Mk�OJ)��[  �,	� XE-"�l6���     �f��݈���b�i�  8kw  V����s���iq�     ���l�����{{{?��  � p `e���~kss�K)7��      ��Z��l������������{  `Yf�  �,-�*�|�TJ���X=<x��͛���:�[Jy�=  ���ZJN�Ν���͎�����f��8����儍Gk���x*��g�M�^��~ "�k��[��Q)�=��G���q)�w��a~�5#�?���Xk�=����s�  �v���R�y�L    IEND�B`�PK
     ��Z'�Y��  �  /   images/4bf63cb1-3675-4452-8ab6-1403298522d5.png�PNG

   IHDR   d      X�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  SIDATx���KA�_�&�Ҕj�PZL-1����?�7O=x��[�ދ'�{�xl=x#"�P"�ɖ�T�[b�&���ݢv��xa��o�;o�f&
I ��ё��v��F��5�M������Yj�ۧ�����ZZZ��v�����$��\�v�T�)�Q�Z���?�;r�V�B�x�1E����� &M6���������FM�0��UUu���[�;<<$��K�Z�L���B�@�LF/_7Ft�o}<YB��.��Ȉ�8��p�\�b�hY��|>D�A=�\����l!�>����=�����y�ϐ!v�[V�������ѓ�=��a��ò���;�\��)�mr.�&�277'�A,C�d�����ƉpF��F)�uI�
f�`���(_���X��N�ǐ�v�����4�q$����"�q�	T���.�[�$�F���E��:MdW���a��n��4�'�b�to���f�����<��.�1L� �=�%n ���r�F�I�wQR�V!��{�G"[��Zbh_+���Ol3$����%��;�'���������(Ϥ'�0�j�����U�99��Xf{Ƕk�Cv�8����
�����v� ;;;����W��t)�x�D�ֱLmll ��PX���ښ^����.�P̂(p$mP!��/eqqQh��!Fk�\��jX� 8.1�d�"��{�n��Il�~�&#��r���>�t�z�JE���>��-��ޞ^�n�a<I��+nDE#E������O�[V�0��T*u�pZl�k'���UV�R1�n�y0q�<��>���$���I�"�t}�4���������J�u�    IEND�B`�PK
     ��Zgm=� � /   images/793ea4e6-6f4c-45cd-8a04-0920ddad3581.png�PNG

   IHDR  �  �   z�P   	pHYs  \F  \F�CA  ��IDATx���	xT��w23��,Y'�d�$�	��� ��J�Z�r�^�Z�*��ڽ�^�j�ֺ�V\ZmŵT��m�Jdq!��	��}���d���$�$�3�$���y��$99s&�y�}�;��j��n�2���" ���"���"���"���"���"�_��/N����*=^(�\�	|$"�����p�����G�	Δxxuq}���V+t�-0�4B��
��("��J���E[q:&��m����@P��#'Ms��iG�'�H�S+��(��-���X4Ξ�����Cڗ���Eh)�,�RZ�>ĸ� "���@��~~�4:
'l-�'�2!�#��DD��H"0敢m�x'�N���gÖ} �@0)�~Qtt �)��E��aN�HӁ��x侹J�DD=H"�|�NS"F��l����0��r�Q	9��4ݡ�sG%�z8S�px�<�[W��;"�(r �kF�LF�)��-��|��h�)�,r�}C(ڊ
`�mB|W��u�ɧQF$��z����54�P:���t�6�����6U�4W�f�WwY��4�cЅ<b;2���F^O""�d��Qիӄ��N�/�@�S��ڕ�����;[7{��nY��e��>[nƊP�ITyh�9�w����.Y'~Db�u(�55�ˬ/?�V�����{Q���]Sv�Ք�%L�r_K�*Jݾ_*�JDDc��@j+*����f���Q�_�t�3��K0�E��[��ٲ��*Z���e�B��#���0�Άڔ
�^��W�aX�}�G��+ojP����b(TG���߂���s��@i07Z��DD�"x ) J�K��HƮW�T��F�/��%kg?�^Rm�I�5Rj�����=���JLB�+�q嵈��_���ڌ��W�ȟ���r����㑲�"�π!�P��|���sK�n�z,y?���IA���x�:��DD�#h 9�M��v�kF�&k�r����5K�8��5^�.�����#-�ƶ�^G7q
&�z�̬ޯ������l6i��W mN�2Y7}iK�B�����t�B���c��$[N��%�{\�5#9.[������i�V�\������I�j�W�
�1^��c�z�<t/l����m^>�/�
�W|J������n���~޶sL^��1-�\�Ͼ��N�GH��jՉ��-;[nE���*WX;�˼��$��l��_�R���_�Fu���t�=��<t ����<��_?p���_y��,M��H�w.��H����L6B����˶n��@��t���x�ը����� {��C_t���}���щ�M�w�U�|�k� ހ��W��m;�yj������A�8V�Z�O�KX�W]�����{e�Q/?���ۀ�䍋��#��^�a��87��P���AI,�6�̔�wU}��݈4
u,g�J׮b4x;�a�x���zDDcQ���J>��>�Xk�^���b�P�F_<]��$�vEfq֔�*=>϶{j�-:��/���IXZ�7�ϯ��bS��t�� ��v(�q@L���aZ	��Z��G��?�"�h1` ɹ�ß��� oj-D��䩲�u_W��?���k�!�X?؈��W���N8k�g�Fsb�μ�$�@�@Ί��ؿmo�"�h0` ��ܐ����a
$WR�<Yv����O,��P�/�4�ꧧ|���E��-��7��� ���J_7�2��(Z!y�
7Y+�D���{0|:ͥr�S�UΨ�g9^�Gu�>������8�\�<Q\~!�
&H3��ƺ�א��V�d��g�Ғ������7Vj�S���V�f�������'`L��F˿^�Iu�HD��������;=�T�܇��7!����y�q����u-��i߷~g`4����t�4m��t-��ij�}�c#<"��$CM#����YG�y��k��-$�\r^VSA��r���5Bq�cS��@@mJC��R���B�v��Eި��(�!5�"�j�;>x�oQo�Ӕ���2���w�(��M�ȧ�7:����*����I'�XȽ��l~O*�*���hI��������(R��H�_-�0��37�����j�'�d �^ȼ��n��3��
�����h{�$��X�3�U��������$�����nl�?ᦊO8����e^s�%���6�4�p5�����c��T��t�쮱�����޺k�f�:}���/���N�bϑF1^/�wW"TU?�q�0�_��/-B���n��h���i9�EC����3�^���g��:�U��W(��E'}Mt��t�Bx;���VF7'����/����W^B玊��0�
�����_�W/��K���EY��r�����w,:�:�uk�Ů�3�^T�h��f�����e^/w��G��*���/���������Ie_�$���������>{�T�N�lꭔ X��pʾD�ى>��k��y�I�y�Q�jE$��\<z�v"�N$���{�n� DD�Bv頴�}蘘o�ry��֒IW+;s�|qe�N����(���t���5g���|��Sΐ���7`�i����P��ƥҽ=���̳�b�����������'�A�Q�UW0Q�� �Fb%`���A��}�� "�&�)��F��Yxv�/�3��N�83afްCV��`D�X�#��b��S�k:�.܍pT}
_��ߟ��mxrƐ��e�?����њ:5]���w9�nn�#B��Q4
��jBe-l��>5� ��*��E8��N���h����@<��N!W�6o�wb<�fF��H327� E��I��#�͍8xQ��Iq-�c����[���Š�!)]�]���#��P8���#qDD=ݠOT�����疠�� #A\3�tE�!u��w��m��6�~~��6�!Z`����DD9���<����F4Ϝ����U��.Fa)�Q���(K���(r�'9p��R��]Hݾ�Ņh������}Q[�H�_-�L""{�H=�].�mك��=p�%Ö�GV*\I������Sۺ�i�H��D	�jw�R��h�{ �
���Mz�XiQ�ի�¯>��1n/T]N�x�Ns<""�H}�#z+}ވQHDDHDDHDDHDDHDDHDDHDDHDDHDDHDDHDDHDDF4�D�	_��c�'���?It�%"�����p�����G�	Δxxu}7�S9��m�BW�C�h���}DD����7N���tL΃�(���*�x䤣iNb;�H���{�a�E���_���S�>5_�;"Țf��t�Ji��r����WX�R����%��(�D��L�˄\dl܎��ZQtR ��h�W����1�<:-j�[������ADD�eЁ$����9#EL����F(]Q�T �0:�28M�iv�	/*����JDDQ$�@�t���0��LM��E�0n]9��Dȁ$��3Mmb�T?���m "��/�@�L���h+*���	�U\}GD4��$�F���E�6�W�мC�p�C���h�Zv۽~4��\��y>�����k�Ǡy�vd~	�����DD4�� q��W�	m�_ڧ|��+/yo_w��w�q��ee�����l�+B	&Q�y�dl�""�d��E�%ס��4Ԙ,����[Mr�_P^�E9n[wMٽ����%��D������B�DD46�
����+k�]�������z@>S�нy/z/�b�ϖ5G�W��Z\��-{0J�	gχ�t6ԦT(�z��v�jú�CX�|�n���AMV�S��P���~�s�Ǧ7 q��������`���E�@R@*�*��P���]���(=�z_2d�K��~^��-']�H�}R�*��J�*!Y7|K�E����G��f4��G��'x��������E�8}��:�����[
wC=+�w �������}w��?��(Z$G�Iv�nq���d-]P�!78��fi�lg���k��y��p�%C�����&N�����9��k�8>���&����
��ɓB&�� m�U��[|�~��[���~��p�\�_~5���Y�@����Y���^3������\���i���lo�N)����P��U(������8�н��<��&m^~ �B�߀�`�s~��}����W/Eҹ�c(b�t�����VH�~C�Q�
>BʔW�N,�n��r+�LW���i^�5%9�&`���*�*L���aT���8��{������H�d��<������_y���n��kL����P�Q����kx�/$"�ZAəl�q�;�m����?R�zaE�.�Qt��+9A�~�.����y{�;�щ�t޾���u���f�1�W]'-����vĦ���(ZH~��߶㟧��_�0Qwu�}$O�X�jb<�/a�}���~#+�z���~^�F��_Fb118��Ҫ:E��+{GZ���$�ùAֆ
���Hby��d�����3���F��^�}č/��p5j��;E� #$��|��}&����r��Ū����x�tI�튼⬆�񙯽Iz~����%"��",-̇���W�s'N}��jIj5
�~P
��W_�V��$9�bz��S6b(�����|]�2����݆H�}�w�{���8t� ":]H�.7�r���c�ɕ7Oֆ݁�q?���(��K"7ݤ�R���7����DD�� #$T�.Y+�ڸ���0�)�l���Q��r����}H�ML���:��6J�uDD���א��V�dR��4��%Sc�i31ho�,�4��N�����9\�����O@$H��U�}Qb�v��_��bu`�mTǦ}�좯DD�*h ��[`�	~���a�2�>�	a��(|�k��5���k��O��=�;�����t�4m��t-ذ�Mϔ>*TjL{�͠��������mo�"��,h j�4�H��:����]Sv�h!�0���
�dW��5��N�&:6�#��@mJ��:��DD4z����Zk���ⷨ7�iJ��n�Z�{	���|����Zl�c�_XUԤ�$���sX6�'G�C��W}©ṧ����G9ƒY����}��:�����ƺ��!u�����rt�f�c�؝�vP�������T�s��r&��C!�B�~�mo����CW8	X��n�Y��H��_��;�����N��z�1uR�I����m;EY7�&�BK�d�]c-��3�W/�^wM��P���^�%�s�I[�9��(��E��J��꧷!.F�DO�����P��!���o�_�nBT��Xz�g����V�b�\���N����#�܅�v��n��>%+�T��P�>Q��m9���$Cݚe����U�ھ↙�jE�íy��˝�둲�
*g��D�׏�����Ie_�$���������_�U
#U`dr��J��O-�':�N|��~_+��{O�\L=�@""�%�tPZ�>tL̅7N��}Lkɤ���9W���h���|EcqnTw���&�Qs�+A;�g�^�+=�9�aOy�.������On\�Ĺ��|ݷ`�y�Ti[t�=�yw�tP�ߞD��""
/ف�r#s�v�,<;��uJ�Q7#�t�̼a��rA�tlZ/=�HG?����>���8�>�FL���mxr�S��w��5��FKH�U*ka�>������W!�@-�IT���Q""Y!W�6o�wb<�]�(�iF� "��r )�~侹/*�35	�!��#p����V""�ꇤty��v=_p���B�$FF"��1Q�t�>QU;/0R��[����q�HL�qdDD}��1VLߙ˷A_ۄ��%��T�h�a~oG�0Q�K�Zj�<s
ڊ�W��3���FE�>�p,�&"�������J�w!u�~��}R<2
��Em�#i�Th0��h�	[ �Pv���e�*����[v:Y�p%�ã�{JOm낦�"�3-$���!J%"��/��+(��6�c�}DqV�N����Ƹ�Pu9���xDD4��/�� �G�V"��Dzc�l�Sӡ���im����۷��P�h3��DD�ӿ�d^����~�sVW����h��s�Z:@HD"~�٘��G���v\�rV~�O�B�#���7�&�D���D��u�W�~R߭`D���jΘ��/�o�
����D4�
���/�):����{ѹ�����(z0��FQ��)�Z���?�6����h��&LF���eo/V�U��}�E-�(ɸ�Z(Tj��7FG��1Q�b ������]U��(�1��FA�F�XSZH?W0Dь�D41!�Hڥ_G�����h�@""T�͍�Mː�3�T䬸���e�m3�݄���u�Dc�h�����LP(���G�~4�}i���g�������n�����X�@"%�����YRuq#m�=A����U�Z��7�Si�Ǥ?�տ�)�{D�nDI����i�;�~B��J��DgX�Ӎ��}8��?!����` �rn�!�眃���*��HW8I���i ������>��rE��$E�\Z
l��pd��L��W�w�>���V+t�-0Ԉ}�l�G���G~���K!�����hx�)tlZ����3���A�;ޭY���î��2\��A��H�8-ڊ�19n���"�l⑓��9E��#�j$�
��D���v��G�F��#��J�Y7}GzD���	�=����(���ڣ��@�kb�8{*ڧ�K�a�BY��"��N�B)�bb\nE#��;Q��CȾ�{��:��_����A��H����/�FG�$��e�DX&�"c�v$Tւ(�<�;�!_�ז���|��$�XC
$�J�6u<��G�E�³a�> s �^?���ߏ������,��]�g��s�"͠IL�U/:s*F��t'�#�͍P�< �&���g߽���)��I��H�H"�|�NS"F��l����0��r�E<�)���D��ub�V+<m-p����}��G$9|r�2L}������cJ8s�"Qȁ$��-�;*a�Ù��Ë�aܺrN�Q�Q(����"���|�UW���?W}���S�/ZL���������;ӎ/@L���,(�H⚑=ӄ�&FJ�sK`.��EQATR��:P������N��񴶠�g�u�a?Fq_��p"l�w�(��H�	9þ�!mE0�6!����h��h����Ң���QQ�Ͼ+{֊��a!FHD�Fv �4�������9����J����F�ײ[|ݦJ��J���j�.�2��{��GlG�@_���I4�����~�Hh{�͐�7�m&b4�E�(d��Qիӄ��N�/�@�S��ڕ�����;[7{��nY��e��>[nƊP�ITyh�9�w�h��#��+���r��ϸ�.�A Q��u�A$�\�B_�Pcj����o5��~Ay��m�5e�ZM�[��-��D������B�D�A�B��M����ay��*HpC�@�H$+�ڊ
C*d���vEës/��]�LyC��{�{�k~��9B�J���B�mك�)�Ϛ'�X�MM;��a����[?�u���ʛԘ����j��y����w��9p"KfIw�61��]�fk�b�m�vP�5�ʾt����E����g��m��+����7Ȣ
��<��
�ʥ?T$c׫g*�C�ޗY�����W/����)�O�CZŞAU	Kk�n�62�.C�6���<-M��j���1x��������EI��������m=�����Q����B���Ώй}�~z��F��gk�r0�P��o�Y]��6��d�Zw���B�> �H4��&�U��5#S��tA9���H�Қ�s�I��Atx��Ñ�]c[H���8E�3^�hz��Ҏ�{�ڠ4��ˇ6'O
��o݆�˯B��i'�'鼅Ƚ��
�J�F���L�
p�}��L�}�BbW������9]���\�fג�G�^�Fͮ�Z���&w�!���R���$n��BE���d�I�\	��{�H��Vo���r�_ڦ.���-;=�@�NEϮ�*>A�\L�~��>˪h� }�R�_�@H���?�ݾo���bZ�t�%H:�|���w�P�؃��TU�2=(�s���A�쳠NNA�~��+���PDL㚾z�������z�h�!e���O,�n�����tq�+���e^c�Q��l��ۯ�������0�{�a��=���S,����<������_y���n���B�,y�����}�at�W��_���)���8-�����H4���FY;�khޱl�ְ����J�+�wY���\�	����p1�ӥ����F'��ݰ����Uf8�r/b�V�ŗKi��MR	"�����"р�����k;�yj������A�8V�Z�O�KX�W]����߄�E�?���z�3�iOk3��+=���oE��+{GZ���Dcqn����ic��X�m(9ZI���3����X�N1�8c��\,E׭��)|v�"Q���J>��>�Xk�^���b�P�F_<]��$�vE~qV��N��p�|dݰR��%�7�kZD�hy}-�"UXZ�7�ϯ���ɽG�.K�����)_�&Z�x��m������`����"Հ�$�ZL�rj�����)�����|]�2��M��16}��r���]1��ǡ������6` ���_�p���c�ɕ'��ew l�������7L$Ks�^{��<F�Flf6�%3�{�DO�og�%��aQY
N����"]��G�p���N��|�����\*g;u�X��|��eT�xD"q�Ȳ����&�5��WLy�y�:Ҥ?�;�g�O�X�y��;A�^CҶZa�H���KK����fb��XY�iHO�4m��?��/.ƒ��y�w��;�«�_��/�D��y���2���D#!h ��[`�I�#��He�}�{¨�Q���'k^M_�"k��}{��g����t�4m7�J����o)�Qȕ�D�i��:�
	�X4�5�h�S$kg����)�S��@�s�yYMYW��^_�(k;qIԋK��R����о�m�'6zS���BI������M�D�(����V;���+~�zs��ԭ�!o����@�\n�G>���Q��8V��U���HB��~&]��{���*�r=�i%���G@�ybj���JU�Ɗ�^��J�_-�0��37�����j�'�d �^ȼ��n��3��
����Mh{�Mi��h� 
�~v���T�@���
��q7�Ο�p>�g���x�������7���?�>��\�Bc�����=Uh)�,�k�%?{�h��١N߭��K�粓��s�Q�׋�ݡ7����w�+�(���T��{�[�����I5�#睋���I����-*?$��褯�F=��]o����IQ�\:���ͯ����z��k]��w�������?�бi�T>�H�A�����>x>�dD#NV ����4}���N��$Cݚe����U�ھ↙�jE�íy��˝�둲�
*g���hd��1��?!��I��������ik��^�0R%��t���So���j��D����'}~��Gq�s��%R.����!�O���<�jJ����jT�p��M�h��}E<�b:&�����s�A�Z2�jegΕ/�,ک�;_�R՝.�nN�Qs�+A;�g�^�+=�9�aOy�.�����%�c(q�������BLl����N���R5<�԰��o|�Ҕa�Y�z[�>�D1�ƿ������Ktz��*��/���dR�ˍ��Q���_�g�)-F݌��3���ӱ�]�!�@?�X�ȪJH�.
���U���;�����3�t�o�&=Dis�#6-��4��������'R?&:�yZ�����*/���/N�Q�i�pBe-l��>5� ��*��E8��hO{�i:>�A��D�Z�A��'}�����mk�����O����R�7��7n�;1v�.|�4#s��ebʭ��H
��on�����LM�h�k��&(|�۹�h(�տ�E��"��Ѡn�W�<�_��/8GVY�p##F��ƪ�?܏�����t�QU;/0R��[����q�HL�qdDc��~����lH������|��M��_"�M�`���v�}�HkX�g�Q?�R�3����F4Ϝ�����T�S��R�"q�Q8�v����^��_�DԷ����t26�B���h-.D��<xdd��jG��j��`*0EQ�I����t3Q�޻@��Bږ=H��GZ2l��pd����)=���v���H����v�6����'7_��tDA_3�@��ۤ����Y�:-��/��B��D�w�4�#
����������"؈vw�#z+�|�N�'�����v�D�@:ݿ�Z�*;��@"
��nT��VX�� "���Df���%Z��DQ�>UG��#�(t$�0i��:��� ��a ���eT��[x�+�0������&X?��_����D4D��=���"���"���"���"���"�h;���w������'�ΰDDtz�@R ���r���0�����}*G��V��[`��Z٠���4�@��i�V\���yp�0Ae��t4�)Bl���T#yOU �x�!�� l���Ģq�T�O͗:�����Eh)�,�RZ�>ĸ� "���@��~~�4:
'l-�'�2!�#���7���ՐIFüR�M����iQ��lز�&��,���͠IL�U/:s*F��t'�#�͍P�< "��1�@at�kep�1��f^T��3����Hȁ$��-�;*a�Ù��Ë�aܺrN�E��I\3�g�0��H�~n	���@DDc_H�d��3�B�VT Cm⫸���h��H>�:0")ԋ�;^]c�vU�s����������[W�e�����]��L)�t!�؎�/����ד���8� nT��4����K8P�T���˶n�+16{��ݲ2U�d�}�܌�����<s
26��]�N�"�Ē�P�kjL�Y_~��&9�/(/�������^�)uK ��徖(U��}�T�����&Y��VTR9 cU��+�מ�x�P��g���`܋ދ�X�e��U*�"m��R�G�Y�`,����4����w�ᬫAg��V|�n���A�9�)�P������߂��������>�i���4K��v�þg7��~��E�����T(U.12l��d�g������zI�-']�H�}R�*��J�*!YׯD�U�"F��v��&4���y^���is�!傋`�>��CmJ;��[�-���~�㈟}�o�	s�bb��f�O���C����G"�� h 9�M��v�m���J��X��a�3�X�5��<�z8Ғ�kl�ut&c�g�Mws#���g�Ai0@��mN�2�ߺ�_����N�O�y_F�w��H���H��z8DׁJ��
�
&H�������������aQtH��4�_U���kFr\�zC�ߗ���6�p���m��!���~���s��r�<�[t��i�<�Ҏ+�R�_qM ����_��������vn���K�t������/=��7��Ys��%�S�	�=
u�	��/F�%_GӚ�AD���2�ժ����-�"�tq�+���e^c�Q��l��ۯB�V��Q������>%�z8��p�w���'Pp��O�~�+/�a���P�8��?��~x�>N$��[�C���ހiK�2��(j$g�Q֎��w���{H?R�zaE�.�Qt��+9A�~�.��x��������D��z���S��t`���>��XX��/M5�'MQ�0��bu�.r���W0LT��>$O�X�jb<ޠ�̼���5�FV���6bŝ$0�#�����(BH޸X�;����&�s���f�66h ��݆����Ϥ�>c��j�˟ =���aDDQ#�I~%e�w�I��}��m}�j��l�/�.�����KRMZ� ������EXZ�7�ϯ���M�=\��1Vh�s��=�so{�DD�b�@�s-��?A)��˛Z�21Y��{�;��
e��^N^�c���0�w�Ai���a}���uZAD-$U�[�����@r%�̓݁�q?�+(��K"�F�zR�!��W�x� "�&AFH��M�J;�6���{0|:ͥr�S�UΨ�g9^�Ge�G$�	#Q	B���8��?��(����m��&#��̦�/-�{��{��dxce��!=udдY ���xC��k���a���+���/@D���������;=�T�܇��7!����y�q����u�`�����%R5�Β��}C.�V
�|�0Z���k�Q�
H��F4�)����|��uה�)ZH ��伬�����n��k�����Ա��_�@*��8�׿�H!�5�����	G�hE 4�/2!"k����Zk���ⷨ7�iJ��n��cHg��%P>���O/otk��U~aՆ�>�{�����`���ny����,���0,bbPpσH��ҧ#":]��H�_-�0��37����sۆB����T�s��r&��C!�B�|�	mo���/-��B���~�4�7Qe{��`���;���R/��S��Nd����
-��ew���g����]�4;�黵W|��\v�{��0��z�������w�+�(���T����B��}RWV�ހ�y�"��N�~ש���4[���N��&+��yҹ��8>��:X%�\:Q�w����Wz.�P����>?�cû���{���"+�T��P�>Q��E�Wg��nͲ��q��׋��m_q�Lu�"��ּ���N��H�]�3��}�����c��B�Γ*!�
�������R�>�R��Ԑ`���ۭb�ZiB����Ϗ<�(}.��Jz��0��?}�/��@"�� �tPZ�>tL̅7N+{�^�>��d���Μ+_\Y�Siw�"
��;]���=F���<�A{���3�t�=�ػ`�:�2z"���pe`� �k�㬳����T�ѫ�[��kx�)i�����Kv Ÿ��ܰ5��E|F��bԉ23f�;d�
�c��C,�O)�FE��D�v���U�_
���Q���3�t{��? ":]�T\5����h���H��q��"�Ģ���[@DD#+�j����N���l�h�iF� "��r )�~侹/*�35	�!��#p���jQ�T?$�˃���q��sd�
'12a$�����Ǡ��y��R���`$�kFb��##"��3���b��\���&��/�զb0D�{;¾����"GXZ�'T��Pۈ�S�V\ �*<���(,%0*��ci7E��$�^W�ؼ����������Q��/j�I���r@���@DDcO����˅�-{�V���dز���J�+)}�Szj[4����h!!U��P*�}a�^�@�5�I+�#��zuZ��G_6�텪ˉod5�#"��7|��<����h ���DDD��DDD��DDD��DDD��DDD��DDD��DDD��DDD��DDD��DDD��DDD��DDDaDI����i�;�~B��J��DgX""=�p~�@R ���r���0�����}*G��V��[`��Z٠��h�D��9��Ӣ�� ���6�ka.~6��IGӜ"�vڑ�I5��T~.��E��9l���Ģq�T�O͗:���E5�.BK�d�M�U�C��""
�X9?�%�,�9��_"�o8�_\��L�E���H���7���C
$q@�J�6u<��G�E�³a�> s��+�~Q����yЁ$��Ջ΁Ü��"����x侹J�DDt��z~T �7{�kep�1��f^T��3���>g,��C$1<�x���$^4�֕s���蘱~~9�Ĝ�=ӄ�&��~n	���@DDc��R Y&���P��Pۄ�*��#��[4��e�O�$^�Lmsxu�;��?4���e���W@�8͕����i.��t�A�����ky=��N[�r~���F(�N���:���O�:kW^��޾�z����w��T-����r3V����]��3� c�.��F���Z�}�:>�F�Q'���P�ϲN�⍊%}���4Ԙ,����[Mr�_P^�E9n[wMٽ����%��D)�����B�DD��<?߲f��_�2Ҷ؆��,+�ڊ
C*7a���vEës/Ç]�LyC���x�5?[�ԯR���i[�`(b�tH8k�����&}�s�᪫A��a���^yCOM࿗~�4(�j����o��t�t<
�q7� ��>��"�#y~�l��z��칸�Z�]"�gB9?$�B|r�����Ꙋ���l�K~Q�K��~^��-']V�O�CZŞAU�U%$"���ȸ�Z�h�����҄Ɨ�E�ӫ�ZN��6wR.���3`8�4h�'}빥p7�=��Yg"�_�g&�ӡ�z�笮��HDt�蝟g=��s�@r��dW�s��&k�r���x�k�6�v&k���s��x=i��5���:�	�1yճИ�{��nnD�g�B�
U|| l�C���)�7�_�s���������Ce��$-X"�`���4�l9i�2�@��r�$��ÿ/���mZ�r9�۲�C
$1�)Z�j t��-��Q��oѹk[ �O�r1m��d)ү�JC|����x`߻[�y��m0]x	��=��uZa۽�;���W����D�}~^s����3&\'g{9���#�Ly�������-�"�tq�+���erVv8�&`�����3X�Fu�?�ÿ��� ��u�
�~{�yw����7��"�����U�!TU?�����g��Kډ��JJ��+� ~�Y���!F����-�o��#��ܾ�7�����ϛ��9p.����-�\��b4$�=	�!.��dS�kZx-�ҵf��;���;��b$���9NWu��3��:?$g�Qށ54�X�uk�Ϝ��t���x�ը����� {���/������F'r7�c��W��u��� �SQp��܀��~��u߂��\}tr���q���O�G�w~���XX+>8�bb��� ��[����&�s`��e���B�
�=� �׿��m��ɯV������v�+&�.��o�8V�^N�����2k���0��g�<��d��f�}���ϭ[ޗ�#�"sg�@�쳠P��2�c���QW�}�"���~���"����>���$h��#~�Y����X2�{{����:w8D��y�@����>(��^�a��� kC���$���X:Kz�U��t݇��q=5g���ގv|�oHSs}S�_[�&��F{FF|�_8O��Ys���%Z�~��?LE�_��V�@
����� #$��"��}&����r��Ū���aZ	ʣ�M, ��#��/I'~����F��=��oO������F��о�WH!�q�a�?^@�kk�Q��=|7�G��9,-̇���W�s'�#�=";�����:b�y���s��޺|�0:����n�C�J�/������<` ɹ�ß�����@��<U��������/�y�6�r�4�p�����N9�����k�Ut�$��'9v
���y�@Ru�!�#^7��]Iq�dm�x����|b�������ჽ�3�y#:6�����Yg�>o{�MD�P��]F�0��AFH�]�Vrx�q�>܃a ʟ��N8V95�N(�3��7D4����o��]�roQ{r�>D���Y����YC����{v"҄r~>v�� ���א��V�d��.�i�KK���S�|��XY�iHO�4m�!n���?D4v��^��}��8)6ӌ�o�&}�����}R1dQ��c�z�k�!n�=�O����H��Y�3�码��o�-'=�f=�T�܇��7!����y�q����u-��i߷��/,��[L��Z"yͯ�]>C��ۑ8A�Y�oY?�Xz�{��ށ_� ���L>Q�쉨�?��/-��ϳ��U?�.�K(�g�1�����p�~���A�Pӈ�9Er^����)�S��@�s�yYMYW��^_�(k;qɲ�=� ��(�8�\�Z�b�'7]-ݔ*Zƈ*��3ϔ*����HF�����������k!�]LL���0��S�?az��}ta8�r~��g]8?�"����GHM�����^QV�3�4�n}�yC�(۽��rS>���o��8V��U�y\
$!���KA�X�n �ב��D4��R��w�#=1�!FM9���T�_��
�yX�_IN���Z;��@qϓ(/�������=񇓾f����Q�p���s��X7���Zj�+Ggn�9�{��ik� Jz���}!�
{n�Y��$~z(�^H�7��I�@���~�>��-A��5���q�Ο"�<��p�[oHM1��Y#՘���?KQ���e�GL��&]�W8�ߊ.�]ۥǉ2�q��R���e�ƒ�T��t�쮄���ϫ�T���iv��õW|��\v�{��7��"yw%BU���@���R�4%��Q��!i��U�C4��zbN:~���N��Z�ϗ|��������}�t�B�
qQر���E�F��'}My�xdL�8R.��I�u�X���Tb)x�Ĕ'��>7L�u�uۖ���H�ſ�H-1M�gY��r��������Ж�L2ԭY�:�p�zQv��+n���V�?ܚ�y��a`���UP9C_<"*t���W0��?���IM�
~�;����A��`��O�k�]}��LԼ�O�������'š>I�5�o?���翷o���c#��/�Cz���/����Dט����ʣ%�"��r4��e�)�*��cb.�qZ��5�cZK&]��̹�ŕE;�v�+�s��ӵK|�cԜ�J������JO9CN��Sހ����/�$BI���d^v��Β���=wiK���i��g�B�ۑw��J�}�̐;ę1e���z���4\�ӫ��y~Nt�v�=^�h��eR�ˍ��Q��l��g�)-F݌��3���#ݳx���􁡽��;>['��M�Z����^܌��������E+ѐOi�G�˫�{��#f-rV���y_3���N$�9J��h����?JCjW3�y~���#�P��!]uK���-� ڧ�#$\���'qA�s�G ��$�X��_!��[Ѵ�9i�Bܓ�io��hk2���o��[�+�$���C��z�-����Q�ÕRwi��\�n�e������-�K�m��
���qR?��K.�]v�������s��@��Ý�hG;��G���i����}�:�T�a���c �}���s_Q�ĬŞ���?"n|�������������_�#i���C$�׏�77��Eep�&a4ĵt�a�Ȼ�HDë������$/XC�L) D����+]U�������'��n�g����4�M��&ܝ~AZ�j��R��:K�6<�E��~�6���g�*#m����P^�� �z��Ye+�I$�x����4!Y?�,=$11�d�����@(��Eb����3>o�by��r-����D�X�$�3�@�����h���A߹%�����~n	ڊ
0Ĝ�rdDD�%
&�X4y��pr75H�H4V��C��X��۠�mB��Ye�C�X7��#�����X<?���EBU-��h�9m���S2C�|J u�:�p,�&":݌��s؊-�9Ìͻ��}?Z��>)����ڑ��Z*71�
DDt�X9?�����˅�-{�V���dز���J�+)}�CF���v��/C�(���F�}gDDc^�����m��u�m��JG��^�~�ї�q{��r"���xDD#&B��#P�8��D�""�,�p~�@"""����"���"���"���"���"���"���"���"���"���"���"���"�(k���w������s�΃DD4z"��<|�� i)��Ña�3%�ߞ�'���
]}5�T+��=?�=��qZ�o{��<���Z�_�M<r��4���v$~R��=U�_�DD4t�~~[ �5�h�=�S�΃C!~QM���R:Yz�i��
o�v"���X9?�%�,�9��_"�o8�_\��L�E���H���7���C
$q@�J�6u<��G�E�³a�> s��+�~Q����yЁ$��Ջ΁Ü��"����x侹J�DDt��z~T �7{�kep�1��f^T��3���>g,��C$1<�x���$^4�֕s���蘱~~9�Ĝ�=ӄ�&��~n	���@DDc��R Y&���P��Pۄ�*��#��[4��e�O�$^�Lmsxu�;��?4���e���M�0͕�����]�e6M�t!�؎�/����ד������W@�8?���t�K��9?�~q#�W�	�`T�_ڧ|��+/yo_wNm8���ݲ2U�d�}�܌��qqq��)�ؼDD��a:?�w�q�8?�j��Ϻ�k�ɾ�6���x�bI_(�55�ˬ/?�V�����{Q���]Sv�Ք�%L�r_K��Hݾ_*HDt:���-k����+#-p~�̒�Z���eR[QaH�&��5ۮhxu��e���)o�^�q/z/�b�ϖ5��Th-.Dږ=
�N�����X:jS*�z=|v;\��a�����n����&+�)�P�����׿������#y�W�1�YW]��y��\�ADG���������=WX�K��L(������T�O.���#�^=SQ���}��/�{���ϫ�T�r�e���'�!�bϠ�Ъ��u�Jd\y-b�����6����8��?�k���=m�x�,���3`<�)'ߐ���R��e��`D�]�#e��N��8ζ�^G�O�{�1�if��ϳ��]r(p~�5R�{~H�t�쪰bN��d-]P�!7�oz�҆9�$c��|����#-�ƶ�^G7q
&�z�F���z8>�>�M%i�@��'�L�M�Aڒ�P1����$�����C�P�0��'�pN�����:�{'���_�b ��!���@�l��eK�w��,��j��ϳ�}~H��4��p��q�s�r���ߗ���6�p���m��!���~Jc��yǦ��y�^�vm?uۼ|�_~ү��4����]�ϋi5Ӆ� i�B�"c��0j^��4����G��~�i�d�y&��݂�?�Dtz����tO��1�:9��9?!eʫ�$���l�a���\a�4/����a6[��W�D&�~Uoխz���4�����.�?�8
~��)�o~�E4��3�=ǯ1%�;���h���U�)�~���0���ʟ�C�,iD���&�x|;�h���b�=�̹�̈*>^���&��ѹ}�[ޗ�+���:=g��8c�
& 6-S��wv��p֊������r��}~��Uݢ���f���Aəl�q�;�m����?R�zaE�.�Qt��+9A�~�.����y��������ƫN���ҁ�*��)���N��.�}
y߿#��%��ٻ𶪳�M[�{�+q��$ę�$(3�̆R!lH[�|-���-�Z �2Z6�P�4�E!v��xٚ��w��؉�+�ږ���<z,GWҽ�����{�{�t�ih��[`�E&�a�����U���4��
�n����S^{�¢>�K����$o��`�����d�FZ|0!t�~��=����:������#�{�}�u���}��Vf�������~^ҼӺ﷬����>|O$���pBb,2i�^����P���������cx���	}f6�SJ�I�:� ��^=�s�
���I�? �M��M�u"�r����Qw�%��O���+Z����V$>��|�읊�;J1H�l6�>�x}Є$��%3�}W�.�������'5�������{o�aGgrƱ��Z�Ǩ_�^$��ǃoz�?�O��J�(����x�z��G�环��S��1�V��˯¨����Bj���K���%���h����Yʈ�AZH�+EhZ|;0H���_��֯�Ad����o��9=����m����ԇ�-���Q�M�c��D���iPWyɈ��"6�O�;o������Y!�Y��/��dF��в棰�{$�gE�0ln@�����3���d�h��t��l�A���t�V���&�ccLL��b�,sTTھ�B$$Bs ����W4�I��<`B�s-�K QS,��׵"MRJ��mۃ_��q���#ZPw �Q=��].�S��@/��caP����������9�t�)\��go�~"b >���.��.�	�y��$���Pj$h������?УF��@%�)~�~94�1��=���]��7^���6(�Eׯ�\ �ӀǶMW(��e1����AZH^�&k$-!!����ʟ��N'����pɝ~G���)*h����6�OJ�}g��Cs����>+[ٞ��1����zѽ�k	ޅ�Q�R�D=K]z��f�u��EHsw�y{D�VB�χb�r%�s�S���V�e0�g���b}?e���β�����)r��k�W��S}��l(�hAׅDBJ�����y�C+���N����}V�`���}�u�F�f]��ńX�����{b$���[�=x����}�8��
1Z6Rr�3�g�9hB2V7���l3�FZK�����CA.g��>�AV���@���t��.���5˴�����v�AŸvW�rF��D1D�����U�|N9c��}�[/<y7�&jEvY�Z8Tq�n4�
,�]~'�oZ�J�C��S�<'%R(�Yc�{D���AAJ��	�\Y��ٓ�Z
�W�^<�w������r���\!w{�y�8(з�+E�w�1��*�57���H>�t�pL'��ms��Qi*3$��MdKn0�:Qy�]����v$L�ӔXJf"a����+ix���e>�耯Wvbg�T���\Q�ٺ�:��a���G|�(���s(��V��T�Ͽ�����T�}��	�+�R=�����GA�e;B�B~�~��쫷٥}��}Ee;(!���������ϥ:rtARi�s��,7�z���MH�߻��Ƙrh�*u�э�	b¬�{�mb�)��7hݰ���(9ry��G��|V<���"皛���{�5��s��\@�νb�\9��j��wd�
k(�����}a�#?�*�9I��i-��/֣��w���1Qm�+��g7>M���w.��yS���-�o��1����y��^�B��~(��c�>cl�P���kD����e��+�(��Z�R����Οa�{��|�EWE��FZ|�516e{�M��*��0w:-��zqݬP���.=��Bn�G���U�|H�����_�"��P�O9����)�xM�'�h�Ps�*wg-Z*Δ���I/S�8�ǿu]�!ɧ��=��P�q�<j�s  5�c�#Uȋ�zY$I�o&��,%ή��G�-c,B��˽�	I�U�9TT�N&Ū��eO���H�ϲ����<����]h�u'��\��`�sU�h��kg���2n,ȾFn3�K�
hݡ�&�W?X��{E���H�]����oS#��61�ã�S]�l�htt��=��{��O=~?���b���7h5��KKP�{�L���@��]j_zVMe���}�UQ���@�Ku�kG ��T#)>�.�Q�-���3��O�M�ƒ�Wh��.{y٤-��u*��k�l�ǽ���<��s�����f�'g��^�p!mc�e�()}s�"$�9֥7�2��ѥ��[7�CHM���M�L{��;8+�E޲�E�gdu?F�T��1t�16���СdB�#��V}�Z��V�V���9������T��e'$���k6���C�'�-F��b�.ݝ�Y�l�U.(����t�c�0ڔT1'�.p��ֈ�o뿤��a�'dA)u�� *S7���/�(i�Ֆ����HA,�f��ӏx�����zG�ﭟ���8�h��ppM5)����I��C	J��j('��Rq���*�sw��8:*L�|U����ׂ�K��F��2D�@�s9���a�Lm4!�'?G���e��?����^�QC�i��x��F�L�\��zVj^x����Bd��
4��R6���tBKUUⲭ0�/F�%W�
�V��{�yŎc$�琫}[�nB{R�4'��zd����ȡ7��)�+4�zC���R1I�hTA�zՍ�6���v\�C��~�z|9!�|俻{Λw�ДN?���EڇuP�g�V�ر���m��L1Җ��L�Sz/c��!&�R�a�k�G�[��讣U�-�g�*D�s�����WQ��+�2B6��sX�!i<^����>IV�
%Q楃�}`�1%8�o�.4�HjR�p:੩��+-�y���ō���\z*DZ���PT����}T��@���sJ�4i��IR3�[F���DS-�t�pI-*���[o(�j|�h�XjZK������Jd�A�X�~�Y��16R�b|Vd	�Ċ*��jQ?c"�&�A@�����S��K�ؕ��cǚX����:�-��oE���h�\�����(��]��;��r�T``�1vX��g�R�˃�ۑQ�Ό�s3��I�'9^S�MF�݅�f�X/�J����!Je�1\��g�R7i���M�C�#��������m��>h]n�}\y�1ƆL����KH}���;c�E�h��C��c���pBb�18!1��
��c�ENH�1Ƣ'$�cQ�c����	�1�XT���c,*pBb�18!1��
��c�ENH�1Ƣ&$*k�7��������s�ʃ�1ƆO4���KH*���
{~&�Yip�&���;����
cu̕� T#/��c�%J��	�g�붷L(@�E����-/u�'A��@�7{���B�cx�c,r��KH�8=jg���P�<	�C�͚��i�Ag��ڣ���1v�����HB��z^�ȾJ�?\��q���G��MH,�c�1�b)>G��h�j�NCS�h&�1�g�{�nX�W�`�1ֿX��a'$j�=�$8��*��lOJ@��k��x�c��X��a%$:���χ;-	C�aMÞ��c�����c�(��CNH�ܷ`ΰlwz2��3�V�r�c���9�D}���47���sJ`-��1�b?>���lc��Y(�&����	<��1vl	�YvB��餌7-��ٝ>cM�f������Z�϶����4œd��7�]$e��^�1���y%0U���$��1k��g�o@�|Ƹ�vF���'�����j�%�~��̩Oݖ<��a��^{~�͡8�"��1Y뷂1ƎEC���j�s��b�=�6��,+�ӁҐ�P�*k*�jl3�z��:9۟ZZ�C)nY�x��liie�����E�0�7�� c�X2������������`��,+!5M*
�܄����Kkޘ�z~��ϖ�t,D�˾6���j��Z4N.BƆ툄�hB��`�6��thL&�x���u��h��:|7=U-�N>��ρ>ˊ������Z�9��Ucc���|��k�E|�^P�:&�D�sB����
��\�}����q��4��~K�ձpլu���2ee����(�VZmbr��1�]u|��5����{�y|�1�Zm��L���{����V�W����P���^S������/ꕏ�A�33MvUX�L�k�vj)"^@�z墚Y�dK����қ`�3#�ڦ���8n"&<�O�Ys������ow�o��VR��1��+�.59��/Gٜ�=^'���u�z��ݾuھ�B�O�ZK���E������ե��gkc�Eb���	ɞ�!{'wxBn���<|�j��MS�����=73���?
��K��ݶ����[z���VO�%�#��Ac��x�~����(@��nA��/�@�����Q����0z
�編��a��Hw|^���L�qc���^N|�BʖW��6li�	f4����f]"gd�Ӛl���t�g܃Ot'�O<�����5����w�]�~�	�Y�`��2.�!�I��~͋��LFDz̓O?�H=�H�`!�{P\�b�E:�L=�<$�>I�h-���Dw=���m*C����5�G�I'�<u:�kh�f�l6�*�E�G�A�G�ï�*���Ɗ��m9W*��&$w�rj�7/ٸQ��@)��t�䭭c���Dٯ�r��&'�7�~8`2:}(w\��ǿ%�xr���7_�����^	��a�Y����?
�XtH;�B���qM�?��\!~6��
�n���c��)s��g_��MC��?�v�z=��;#���LH���em��s���A�s�赃�W�WZ^��ٗneV>���F�z�g��9|�ɽo�O�VV�����	��(���|���QѽN۷�e���< F�҈Y��b�:� ��z�]��JF���M���+v����&���&��ul���=bB�Fb|0!�z�;ow�b��[�kdm(}�����	��w�Kf����]p|�-��SK�.�����NG�}j�3Ɔ]����E2
x<���kE�Z��J�(������u�@�3+���7{\Ҙ�(��CH9�\��F�����E�H��AZH�+EhZ|;0H���_��֯�Ad�t�C�fľ5��^��5X<.;G|(����}_��mBb���cC�2�x1��Լ�T�Ɉ�.ԯz��ǚ?yo�s��ZJ�~v#J�^���|$�=E\{��4���#1>+���`s�*%_O�~xd��@eį��j+,S;[\������%3{�NP9!16�hJG�f���� '�P���w���z�X���Ѱ���B�����GR2>���\��H�K?�bh�R�eo����&��EK�t���wV!k�q?�����w��Бt)��.�y��c�L�K�?�:\��q��Gۅ��)�����<`BҺ�!�3�8�t��d�\YvH���G�����H�m���#�h�(]��!�m�6��f��Qw�^ttx�P���r�rƆ�{����T����W᷷����t^���p�.�uB��.���G}|�B�B�t���7\,����ʟ��N'����p7Y_�e�Q��Cc0�:v4Ҧ��W{m���z��׊�����n�e��r^��l
�0��b.�M��R���]jT'�*����pT0���C1t9���9�5���V�e�˚6�����~ʘ��eEq5��S C\���1���F
�B	����+������p����v���{+P���~z&>���7����A�?�(��2��YэN󐲯�N�h:�b(1���DI��@�ALc�L�$j�U�>�ˍϴ�Q,��	�X� {^f��5����������\΢�}��~5ӁY��ر]���!��i3E�]#cBA�A#p�(�J������A�~��Ֆ^�c����Zl����|���]dY�ƌ��D��P����)&ƆD��Y��53���ˈ�뺄�5��G��|�t|��̕���=I�����z����GKH@o-<-�nL�r�7���]CjYW���-.b&�;͟| EIgVG��K<a�8K"���1=h���o��p;���hdl����"B�b���C�i���dNl��Q�D���_�����PⳭ0g����9x���V����zFmi�?���H+�v,����/�&y�Wo�K�*��*դ��D�����@���,�5�T@H�e��U����_/�1}������FhR���{�m�')�ٯѺa=��6�b���"Բ�w���ב���C� �v�K��і�eU�.��#cUX@���������i�LI��i-$`@�R�X f]�}`���F]y����;�c㼩E�O~��Y'��tf�m�׽�^ti��ѭ7��ǐv�"�d]��wP���dԲ�#T��ce��GX|�516e{�M��*��0w����{W/��j�pե�[_�M��ȓ�j�)�B% R2�%!�9]���8��!4}����ۅ&�Ҭ�EK��rB�5i�պj��]8w|%����D�ߺ�$�v�؎�U��~0�bLG��rogB�-�*�5����#�y��^�P���,+!i��΃�:N�>Ѕ�\w����%���=�PU؁�/�v�n�*��Ƃ�k�6��n����4]���Pt�H�������P������ [�HF�����l�h��1�:���W�N�5ʮ���q����d�>��}���U*���n�+���,�NFa��f$�g٥�2�v�e\>|�x��3�ԍ%�д�]��I[4��q6�Z]�g+=���I���7�_�53�89+�: �i�/�DI�
&�9֥7�2�Ѳ�I�]���CHM�����ZW�=�P+��!G&#�S��38��#����MqTf�PE����/ҏ��.d^�X��d�E�����oqx}��ϲ��ӎ�5�Py扡����f1N��N�¬k6�*L�EL�i�0ڔT1"�.p����Y�h1���T���j4�!���`;��!ތE)�J�骟y\TO�����zG�ﭟ��M�m�F�����*%�s���j|��jby칻�\\�h��UvWAI�l�\��M��6x�GcJRM���/`]|��Cؼ�c��w��J�C�M'��xˡ�ԳB�Gʸ�R�\s��O=!Td9���|���>RO���C��m]�	�I	p�r���t�����d���^�EG^�UY���K{|"]�^	�j)���)��H�����@��k���p�'c8Z�}X����c��u��^|�ik�>[jM��ޭ�CL�m���b#դ<��ܕ�Bzo����z|k=$�ǋ�U�`��'�*[�$ʼt���1�Z��n]���bM��,]G����s_����X��a/�GU[�L\=�M��`(P�$5�e�L����b5>G�b,5��_�TU��y%�ʠ��J�[?ݬ� ��b1>+��ybE�U���1M�� �Ufet��R֥q�J�f��cM,�ge����Y�"}�N4N.B��x�[�[��@�ν��D8c�+�Y���E�� c�vd�m�3#��L8s��IN���w�Qgw!��&�ˠ�*l�Rc���Y��M�acm���P�*��3�#��|[u�Z�j_��1��)J���%�>Ё���1ƢK4��!MH�1�X8!1��
��c�ENH�1Ƣ'��|��ȸ�
x���
��#cǂ����s�+�D�'��NH1�z�2��+0ƂK9�,��8��#`��R�^չN��nG]]c}��Ȁ�l�NH��RQi:��.��bTUU�`�b���2�˅����?���ΰ���[1���F,��zQ]]�}���p8P[[����u��;�b'�p:��wtt�/���CRR;ֵ�������G~gX���Er�;��uզ�&���	i�/#u�1v��x<`��c���0�	�ʚ�q�*o������� c����y��
pf��	gVܩ	���Nk��7��X� s%- ���1��`����xB��ź�-
�n��D.�!�t��D��Iз9���^�l����7�cJ����XB
��Q;��Ņb��H��n�$4L� :�l�e�ng��cE��gE��(��JD�U�����ml>��nBbyc��K�9��D;T3w��Gc0y��<�D�sw�*�� c����b|;!Qp�9'�iM�P��f{R��]����0�X_b5>����`w�?/Y㰦a�y�1��RNJ�1v�X��!'$j�[0gX��;=�ϙ�Q�K���1����rB�>IGv�e��9%��~	�c��CJH��y�~�,M���\U��
}�;����,;!��tRƛ֎��N���~����W\�g��g�F�n�&N�$����.vYӦz�Ɛ[l��TU�דc�,���P!.I��ƹ~c�ER�kH��7��P>c\H;�ms�wW���V��W��k�ԚC�{>�?_�0�t�=?��P�f�Ϙ���[�cǢA�ϟ�-���X�P���|�왵��gY������TYS�Vc�y�s�������RJq�����Ԛ��AJL�rߋJa�o�)
2�رd��M+ͻۓ�!�����J|����&�Tn�R^��5o�V�
?B��gKk:b�˾6���j��Z4N.BƆ툄�hB�	sa�6���F��T�m��h��:|7=U-�杊��' �*�T��p8��f;�>x�cL)C�/~~M��^�^P�:&�D�sB����
��\�}����q��4��~K�ձpլu���2e���� �l{XUh��Iȹ���Z��xC��y�P���~�q�Zm�O<i>��}g":
MO��ߡ��b�=w"��1�"5|�y������,��$7>MH��4�Ua�O2��uک��x:蕋jf��-�>s�>Ko�	ΌkC[��8n"&<��I���Ν_�o�Cc6#���yХe ��[�y��(�3���$�<W<�N'~w�.G��2�m-��%��N�Z�G楋�ϲ�~$������s|��t|���y�w2q��'��I�A��׮6=�4��j9��s3CJH�R����*h������П`��{�|��1�\�HJ(?��TB��G����d$%�=�5j^xZj���?���H�ɧ���3�E�{��c����r�����.��������-�l���(�h(���ͺD���5�(�u�Z��Vt'�O<����o�Ž�����>�1���>#�Iǉ��e��湿�~��=�����������]NH�E�Ɍ�s�C��s�I��b���ަ��V�mSZ�X���sk�R�y�t�&H�F-�����p9����c�Mڶ�+���A�;�"o�j�7/ٸQ��@)��t�䭭c���Dٯ�r��'O��K?0���;�]���ti�?�����-���D2���c,z��{!F�y�H$������φ�_Ǯ�n���e�d^v��s�HhG�{�E�H��&��N�ﲶG�9�_� �:]��~=`����.��5�/?�ʬ|菡]�	����ml辯��?�S�;O$<5�`�E���c�}�J_R��ݱ}+Z�~O�A1�V���$�0W|�Z�����#���C����u.��"�y���3�e�T��Q�Ags�����Y���&$�m.�!�*v�������ZM�%G׉�?I^���gF���>��ag�?�������I�_���Z4�^���H=�{0����:�*��m�ж�Kطl��ꛥ����w��g}�{��e�� -$��"4-�$���!�_��.�6��SE��oU�8�Ժ���r�{`��W���`��˥$�W<L����0ꎻ��4������~��C����^����&#B�m�������y�~�ǿQ7�`��Y�%���P)�z4鵋RU��v8ȿ�W�(���6��ڠ��I)�v�����<��� c
�)]�d1"Q:�C��+C��d|0!ɹ�%��)�~��Z�&)�X������i_��9�P
}��}S:�J��^&4f��u?��hz�E/j2�"�Rwߥ���"���M�OD�������	�y��$���P:9Ѹ����T�%7b(,�Ŀ������4���MQE���|��v���@7j%������zt��K֢�P���<Q,��g��|2b >i!yi���������*.g;���r����e��DJ�Y�AJF�������Jа�{B�w/�hNC�_�clx�����j賲ŉ��7��D�/֣m��Z��B�χb����%�s�kH񍭰�8`Z�蕅��~ʘ��eEq5��S C\�rx�Oj3�E��O=S��#4���Q{҇��׷�a��-�s�M�&��� cl��w���0��Qtڤdd/�^����m��Qɥ���DUJ���3���4!�`���B���֒�0���P��Y���b�կf:� 9;��4��2m�趋d��q����.��n��+��O�Z7����e�l-�\x�n�)g�+z=�
��q�F=T`�%5��
� �����="���|��sЄd��E��Ir�-�֫W/��;ZB
xk�i9ucr�����@����%���-Z+4?�����O]Jj�}_Kˀ���Z��kL�"2������<EZ��|�4�Kf���TR�P�{���gd��=B�϶�R|�m4���-��F�[hO<��Q[Z�Ə� Ҋ��y!?��I^����Ҿ�/�Z�'EB"���Zj���d־е"O���߽G�1����|g�ϥ>���5�k�1Ɔu����D�MN�u"�n�M�Y"���e��}�f�����C� �v�K��і�eU�.��#cUX@���������V��I�v_Hk!�>_'�K9���F�V�숺�B���w.��yS��;uS���������s��b��Rh-���nt��NX�[o�}��2CP��u��ߡx��wnd�gYcS�W�a�٫�
s���z���
�y���ӭ/�&op��?X�χ�m�U�/
c�8Q�S�۟��������z��ގ�%�=Y��JgJ'���)j^�D\N�O;Ez���{ҭJ��Zcg����f^��3���� *�rogB���e]�t#)>�JHZ��󠧎�\�ҫ;�|`����k�*�@ۗ];C�W��pcA�5r��]R�U@�}���v����z�N>M$�»�������JF�����L�H�Xv�~��zY��At���K7}���T���U��1[���vVcP��6�+l:�FR|�]:(�lZ���g���#>�I�X2�
M[�e//��E�p�N�Rum�����w�'1~��������<�� .�m�L%��^&��N���`�y�(�H����[	҇��u�W�Ua�z��ȿ����D	��Z�Zo��\��>��g��19�1��С��u�Q%�s�ۿ�����#>�NHjO;��lB�'��O�[���8]�;
���,�\P0��F7j�&N#�h]��I<W�N����S��˖�9�b�5�3���--��]p�����247�F�U?󸘚��%ɿ����[?_�h�d|Vra�P�sH�U˫`�ݍ��BD���*��;�ʍ��A4;;4`�u�g`�E?�ф�����עn��hY�1\�v����V#�B��T�(k���L�����{��z�ۑךro��t�{��%%5���	�9�j�ֵ�О� -G;�L둽nx�\2�F�C���X�� n�Νˮ�1�Z��kn���T+���]-��s�	I� �ݵ�s�|�ӓ1-�>�����_���4�>�-<[�K4O�%ZCG^�::D֦���gV�����G�]�>����+w&W����C�x�(\�	��}���J��KK��cJ�	�GNr�n:ZFF�"�r�Ir�NRWަ3��p����}T��@���sJ�4i��IR3�[F���D����b5>G�b,5��_�TU��y%�ʠ��J�[?ݬ� ��b1>+��ybE�U���1M�� �Ufet��R֥q�J�f��cM,�ge����Y�"}�N4N.B��x«f�ku y�^Qn"�
�1�����XB�qy��a;2ʶÙ�{n&�9��$'�k�ɨ���l�eP�rQ6�B��1Ƃ����xB�&��I�p�t����u�������/���c��(J���%�>Ё���1ƢK4��!MH�1�X8!1��
��c�ENH�1Ƣ'$�cQ�c����	�1�XT���c,*pBb�18!1��
��c�ENH�1Ƣ'$�cQaH�5���?T�\����9h�A�c�'���%$��H�=?ά4�S�]ӝ�d�ol����JZ ���c�����Y��3ċu�[&��"o�\�C�閗��ٓ�os 雽H�^!�1<`�1�h�ϊ%�@�����\\(V����fMBô	�3�v@�Qv�v�;V�J|V$!ي�P=�Dd_%��a�8���#k�&$�W�1Ƙ|��#JH�C5s���x4����3O�=w7�ҁ�|0��_,��5��s��tjn�'% �ݵ�x�`�1�[�������Ý���氦a�y�1��RNJ�1v�X��!'$j�[0gX��;=�ϙ�Q�K���1����rB�>IGv�e��9%��~	�c��CJH��y�~�,M���\U��
}�;����,;!��tRƛ֎��N���~����W\�g��g���T�K��I2���.���T��r�����j�zc�i|6T�o�9ۥ��\��7~��T^K�dw�q��h�ؑ�z��byS��Yv��P>c\H;�ms�wW���V��W��k�ԧ�n�?�?_�X�P���B9p�E\?c"��oc��)>���a�ⳬ�DJC�Ba���L���<����lji�O:��V.�w�'+c�=?;G�{Q)��M;E!@�;����,+!5M*
�܄����Kkޘ�z~�����Tw,D����Z���yN@�E��"dl؎Hh�&$�0�i��Oπ�`D���@%��>Ck�����nzj���(=/�Vl�?c�Eb$���	IQ�O.Ӿ�Y[�8^U��v����X�j�����y��2q��d�m�
�61	9�,C��WAo�w;oCj_}�O?.Jè1�O����m���c,#,>MH��4�Ua�O2��uک��x:蕋jf��-�>s�>Ko�	Όk�Bz��	���9�Ys�����Ν_�o�Cc6#���yХe ��[�y��(�3�h-�/c,��W]z`���+��&${^��L�}�	�}�rP�p�R�3�Ǎ]*g{{nfH	)>&=��	��w��RT>�g�m�R��=Sy��
ʼd2/],%����m.�'d}���{Yf/�׽�c,��/xi���&˳R|�J��r�s�R��ZH4t�aK�O�0���&m[ΕrFv8�i�Fy���h1�������`���{%�.����P����A��0z,�g��m�6�U����1��z�yH�}���-�N>-���mj@{]���-C���9|nM��s�v�B���X���߲�u��_sh=9����|��+��&$w�Eގ��o^�q�Ⓛ<R�y���[[-Ơ��=)��_7��0O�*�7�~8`2:R{m5v\sB�~��,���u�X�I;�����r2�#���ױ���F�ף���~��{>P4�'͇u��u�M�G&R#->��:]���M�h�D�r�k=`����.��5�/?�X��e%�n���3Qk,�����aG�o�1=R����=�}��ؾ-�>�ZB��Z}�U���hZ����\����dD=!�Edk��d&���>t�i���3�j���}�5��	�g��ީx�#�t�}�{���ϒ?^4!��ns�q�>0���a0%�|���~�;o��t�1�E3�Ww�d�x����������`D��߃q̸>O�s
�/���O=/���*�����������gDR������3C;>�H��AZH�+�hZ|;0H���_��֯�Ad�t�C�b߶	�-��v߯[�"cу�R;��Ծ�t�Ɉ\NԿ�r����t��鷷���7w'�.����=��K���x
���UJ\���Y�%���P)�z]��ڏ�D��SN�]��ň<�X��)]"�~�3�Ťz����4��]�3+DB"�g�vB
���W4�I��<`B�s-�K QS,�X�A�IJ)��m{��v�����>��)���Pi;�	j_}��(�Rwߥ����Z]�j���PH'���}"&�0/��%>{S��y���u�C.g�����r��d���<������T��؆$�K;���E���1]���t��Zt�W�"��p�u%מ�������YٝC��m!�_(��e1����AZH^h�.Y#9|񆋥�`��r��I�*��o;\�GkI�`�Q5���i�G�����Xti�����A]n��"L�p��Nd�b��3�_����s��{��`e��EE�ɱ㫐�;��|(�.� P2>����
��vYӦ���X�O󰽳�(�&3]V���&��T��f(���c0�=b,*��Q��c£ϊQtT,9{���F#�h$n�_���1(����d�d�˾�Z[��Sy�pɍϴ�\,��	�X� {^f��@��i-�__��E��,Y�j��^ӱc;n�zi�6St�u�î5�'1<t���~{�AE&�1���k���3�w�mH9�\���-$�`���nTÒ�\���o����^��1t&�%���(�t�X�P�ƒ���������A���u�'�y?�Z�^�x���li����r���\!w{ӁZY��5��u�H����"fҼS���P�U�:c��׋�'<Ƙ��<خ��(�)R�/�q�D��e����2��{���gd��ӏ�x~�����\�N�oK���]��r�B�϶�R|�m4���-��F�[hO^Q�����o�x>
"�(۱��S���e_��.���P5�xR$$�ۯ��D}����O��������c��&����X܈JJ	�ND�M�uG.��7�b?-#�%�tv��&&��T�lE2Q~�����:���{��r��gYվ>��X�P�-��})��2G~�U�s����ZH��׉Y�)��#���B�tvtdS�/)g,��;���yS�݆��H8���}���`��&j��	+}����XgW�Z��^)%��voGX�h��"�~^}�GX|�516e{�M��*��0w����{W/��j�pե�[_�M��ȓ�j�)����_�Ƣqbi	JL%�KQ��!4ӈ��#>\Rs=i�)Ⱥ|�8S:z���D먫��J��؈��/�v_6O:���4���>#��o�})� .^�儧�`D�5�ⳬ��uz:z�8�e���u'��\��`�sU�h��kg���2n,ȾFn3�K�
hݡ��0�.Y �*R����|Q_
w�'�vh$��ѥ�v�"t�ԟ#�RAŦ��cldp���Y{N:�Tz�nsl��}��=��Y�Np�S:W�u4C,�|���e��(ہ�q���e��lR7���BӖw���&m�8ܯ���kumQ��k�;Γ?�o��hkf�qrV�u �6�_���Ҏk/�Z@��z���<A[��?]���CH�|5��]t���H����5�ץc�/����h���%Gk%�:G����{!�{��©T�z�OT���9������T��e'$���k6���C�'�-F��b�.ݝ�Y�l�U.(����4�4q�hѺ(t��>x��A���Oޗ�z,c,:P����~vnw�����[����U:A=�����֫o�a�Xd�p1j^x��6��ro�,�J����JE�A��\��C*��X^{�n4"�|U����Wnj��ٌ�c��h�&{������];Ee�V#*8�&LF��뺋���Z{%r��G����Ѩ_�AJ@��}���ٚa)��ѿ���^%��F�j$�琫}[�nB{R��02�G���`�����C�"�%7��@h���eW��X��1�n�͍?B�S��kEy�n��5�g5*�3���9䄤����Z�9o>�����i�A��b c�Q7���g�y�4!���5G׸��EX�>��X>b���}˗�rީȿ�W�5���P���g��ZM�{a���z|k=$�ǋ�U�`��'�*[�$ʼt���1���z�$W�­KI�J����B��!M`����n�^� �ѻ�xx��^�H���r|{�>��Z e��9%h�4C��$��-#��`j���HќE*�:�b5>G�b,5��_�TU��y%�ʠ��J�[?ݬ� ��b1>+��ybE�U���1M�� �Ufet��R֥q�J�f��cM,�ge����Y�"}�N4N.B��xe�닮Ձ�{E��p*00�;,V�b	����AƆ��(�gF
칙p�Ó� ���&���B\�M��A%�EUX��0��1-���	������&qá�T��g�G@����v�.7�>^+�1ƆL����KH}���;c�E�h��C��c���pB�f��1v����hj��b4�N��b�J�BZZ�ر,99Z�������Q��RQ���)eddpˈ�C,�j5jkי��aяR�Z�O��!++F��1փ�dBvv���]�MK8!Ő�O�\�r%ZZZ��[RR�����a��R9�ԣ(��oxc2�w��NH1����
׮o�~�%�����XO�܃�hB�����C���	)����d����c����	�1�XT���c,*pBb�1�4!QYs�!�C��5^�X��Vd�16|�!>^BRΌT��3��J�;5��5�iM���V�`���y�>�,Q�OH>C�X��eB�-�ȥ?��ny���=	�6��ً�����c�����XB
��Q;��Ņb��H��n�$4L� :�l�e�ng��cE��gE��(��JD�U�����ml>��nBbyc��K�9��D;T3w��Gc0y��<�D�sw�*�� c����b|;!Qp�9'�iM�P��f{R��]���c��j|+!���>>�iIjk��7��,��cG���rB�f�s��`��ӓ���������c�X��!'$�td�a�Q&��Sk�`�1��9��d�7��B�4i�UuH���w��c�H�ϲ�?N'e�ia혮��3��o�:=+�Z���>�6�/�B\�O�q��w��էz�Ɛ[l��TU�דcǬ��e�M���B�m�ӟ����[o^�qc_{�������6L0�k�Ϻ9��Y��3&"k�V0�رh(�scQ�C��s��Y��gֆ�e~:P�
SeMeZ�m�YϽ_'g�SKK}(�-����--�̑��#���F���� c�K�0>ߴrѼ�=Y��e%��IE!���TTm��z��W�G���liM�B��`Cka��6h@�E��"dl؎H�F$�0�i��O����xT�m��h-�>yMO�%ɧ��qӠKIC������ھ���f0�X��2>_���j������-��P�s����(�'e�p��-��v,\5�E��}��LY��y|2ʶ�U�V����k�!�򫠎7�������<��gV��j�{ߵ:X���7�"Z�::���޿�1���3_�+��&$gf�쪰:��G��H����E5��ɖJ�9x��7�gF
��M!��q�LX�⬹���^_׮o���
mB��G#.7����x+2p��L��Zj����O=����C-"j��F�=�`(-m��n�8d�����&${^��L�8��>I9�y��զ���]-g{{nfH	)>&=���t�����|��h���H&G2������y�bh�	}�ި_/�NF�e�a�on�kOE�m�Y�H[p!;c,��W.5>�x�إr���������B��۰��'P��P~sk�u���Nk�Q��4�}`Ew2:��#����^��%�}���>�1����e��Ȕ�oیW_����k���j|�Q0ƢG¬`)��s�?� �]������׊��mjD��|]j2.�T�oYW
���Bڇ��c�Mڶ�+���A�;�"o�j�7�3t0")��t�䭭c���Dٯ�r��'O��K?0���;���׿[��V�r*q�oo�31ƢS��S�s]h񺽾�WB�[v;4��1ӵ�m�6����,���kq�P���FZ|0!t�~��=����:����z�^i_i]x9k�g]~��Y��e%�n�������|JgW}�B�P1Ƣ�tڃ/8����/���1Fb|0!�z�;ow�b��[�kdm(5P����	�F�Y�u6�]�"N &����>���bW4�q��������M�>c,z�\v�[7E��=��0�D$�|Z>�J��9HI~�M�o����k����:�lc�R"}X:���D�L&w�w|��眇Q��=��=��6֣��C��O��"c�Ŕ�5�8�KMG�m�F��Oz��Dj$�gE�0ln@���Ѥ�.�����69��~���A�eW��Ԥ�!�t�>�t��?�R2�n���c#���'��}7�/Fڂа�_ö?�_�z$%��	Iε�.�DM��c-�&)�X������i��S`���r��"%��{��u�=/9���Ϗ����݋ж������j_��t��^��h��jYצ�
%>{S��y���u���9��0H�I6̕����иe���$��F�#г�����>������u����.����s�O���/�C��Tf��{1�޿".'/W�$4��처OF�� -$/�N����x��ҏ{0�����tҾ�9k��Z��k-	�T��<���M�{��>�����ֈ�]_2M>�-�� c�D������'p�d�^}0�k5��:�Ko�i�$��x�_Y�VB(��P]�A�d|z)��v첦M}ea���W�V�M*ygYQ\Mf���d�����2�E�|�ÅR]{�l�8��!�x��E���2�	ފ��E��h�|p9&�x^t�g_y�} J��i=�X��A������`���0�Z���
r9��Y���Ld��c�v�.QH��fSZ$ñ�,D���^W�}_��c,���{���x�X��	�/��Fy�*�P�ƒ���������A���u�'�y?�Z�^�x��h		(୅��ԍɹB�������vm�?E�ig���IsO�p9�9\V��|}�g���W1�16|���^���	m���A�K��1��s폱��;��PⳭ0g����9x���V��W��zFmi�?���SK�����м�����$/��mvi_�V�~�	��H��~�����O����ݕ��[Ø��5f���h|�}�7����S�k�.8�+�u��24}�.RN?Y�-A�sq#R#->���$��+�ȕ�-?˪�]�yGƪ��9��})��2G~�U�s����ZHԄn���H���b	���?.�QW�@���;���yS{�{���EM*]J*Ri��[+{=�V�I'����Gדcǆ��ߍ�S�U]ro�M��"6�ⳬ��)�+�0m��U	m���_�-ܻzqݬP���.=��Bn�G���U�|H�V�PU��0���h�P�)Y]������z��jLfѭG��H���z�sO��i�N���*��_��@Մ�,��B����c;��Ih��W�q��~���B�JI�YVB�:=�=u��}�m��d�K���{����m_v��^U�Í���mvI�V�;��#4�{�����EҼ��"|c~?p�}�65��4f�h�t%�*���FC����
?�R[-��#�%E��w��ЅF�4��cǖʇ���s/�:>y?���=R#)>�.�Q�-���3����٤n,��-ﲗ�Mڢq�_������<���k�;Γ?�o��hkf�qrV�u �6���EI�����d]r=,3O�t���&�f����~�/�/�:����Qw܅���-+�hs����{���r4��-0Ǝ=TI��ŧ�Xs�X̓�]+A�����oqx}��ϲ��ӎ�5�Py扡����f1N��N�¬k6�*C�7O�"mR2��61��sI���h�U�皧L-���)�'9�wr7cǸ+F��AcI@ε�yM%�s5�j|��jby칻�\\�h��UvWAI4����/"~_K�Hp��ؒ~�%b�P04()��"���M;Q�H��!W���݄��8�iN����^��1���EKdmGe��X��
d��J賲��X��!'$�/��w�b�y��NO�p04�H��*���0ƎM>�-�yAަ�^�F�ͨ�&1(j ����ǲ���6D*��sX�!i<^����>IV�
%Q楃�}`�1%|�Qq�Ԗ�O��m�k/���b9>��@Um-�2q��4M��@}���c��/V�sD+�R��Z�%LUu��W"�z8�ĺ��͊``���*�"K�'VT�\U���4yZeVF�,�*e]Ǯ��n�;��R|Vf���o��~+�7�D��"4�/�WF����ZH޹W���c���b%>+���h\dl؎���pf����	gN:<�	��n2��.�5��zT�\T�����1��h�ϊ'�n�k���JGP�?�1]�۪�}к�P��_�1�X��4>^B����c,�DC|҄�c���c����	�1�XT���c,*pBb�18!1��
��c�ENH�1Ƣ'$�cQ�c����	�1�XT���c,*pBb�1�4!QYs�!�C��5^�X��Vd�16|�!>^BRΌT��3��J�;5��5�iM���V�`���y�>�,Q�OH>C�X��eB�-�ȥ?��ny���=	�6��ً�����c�����XB
��Q;��Ņb��H��n�$4L� :�l�e�ng��cE��gE��(��JD�U�����ml>��nBbyc��K�9��D;T3w��Gc0y��<�D�sw�*�� c����b|;!Qp�9'�iM�P��f{R��]���c��j|+!���>>�iIjk��7��,��cG���rB�f�s��`��ӓ���������c�X��!'$�td�a�Q&�����2{�o��m���A[�E@�q�q�����?��踍�(.��;�n�����esd-�(m龥I��I���+	-M��6)�����饹���&�{�������yH���0��?>�$H��>A��#��/�Dd!W�1sl��gق�UK�7�G�6Y���J����z�*��a�ޤ�i�������ע�����]I�'1s����9��j���,�ϖU*S�V�éh�0�Zc��Z�����F�#�>/`�u|�- �ʮ��bT�GԞ���%�]�d���S+>�a�U�P�"SF�_��VW���5��0s,��9���A�kr6L��0�:>���RI�/�ˋ���|��J9�O�ϷKo���s�<b4į��)M��
#~�Na�0s,ч���-�=�[R�4>'��=�/�,A����D����f�2A����o䗷�Ā��3���dŠN�
5�9HX[�ޠ��u�dD��!J�����0��+����V���S7,a���������0��/���,�����[f�3f���y�/�wAR@��EWTv i�'�+�}��SJ�Q�3��W=s�)=QV�T7$	�
z�B���A���!��ֵ�FKM*�,Ɓ�� ����s���B�+e�o��sѸ�0��#7>�{W3�H�eEJr�g��dI4�v������8fj>z�@�������1�v���eK���Xh+|�<���a�Ko#�]�\Q��;�0�D�6 a�P��#��7 a�X71�0G�#9>/�UJ��~��^ɔ� �"����,7')
?�R�z��Y��)-�'A
���ş@)�]��G?�L�7t�73�]��Y�A�����UX?y4�a͑�g����R]�5�].g9��)Y��Vo��~F�{��1e���K�X/�
�
��|�-F�/=��O=,���cJk�-�eo���� �0}�B�F�_��B�@K]-*?|ǧ��G��	'���U?¼}k�硹���S��u�A�-������/�Q���p6�k�@7�1SOG��ܴ:&����K���Z�~�����	Gz|�^�jL���٫ Yc# ����֯��b���� w�1B���%���gL�n�(�]��݊Q{�+˱}��`�o����)��>������_�q��:a�xm��x�'n��ȸ�v�e���S%QI�=O�z�/���"�F��
MIC���aڹ@HH����� 1���~M>��]�&ߜ���ܭ 9��.������1��������n��������|����g�%Fn���0G�ʏ�m$i��?�"�����ׅ�e��#�r��wx^�Tb���#�ݸ�R[�ϫ`;P��ID7����ndUQ�H��&1����΁G���1��ס��!��a�i�z��mb��G 45M��"K=i*�'��_'�R�'X�guS�/�s��d�Ⱦ�0�9"���J֎
���*HTޭ�+��
�y��J'�g�H��PQ�gol@��]�����1Ӊگ��q�B�N�1S���|�f\�R*����y�d\bDK2�=z�?�P���h��d$Ͻ
I�̣/|����?��w���Z��?����:�K���ӧ!�7@;d�?�,㳦޺R֎2�g/�|'e�};��X�M��j/��rG��0a��_sV�!y_t�OJ-��(�5�r�a�㰘Q�ϐp�,Q��7��v�"����	Z�Q��������y׈m���΃u��.GU�E��/�(����=�[������.�EiȚ/?E��_ ���$m����g��04V�S�m�4�*S����f�B�"(�m������>�T��2���t����� ��]�U�hވ�s���>���P������nŨ=M{v�G{bN=��#�vݏ�t+F����@�P:~C����[A�3���.���Z�et�p��6{��SF�b7����
EU�������p��� )*�<q��a�n�0�c\����+�m���}�	�����.�"*�v�̣�Z���6-�hX��Wזx��v�O#��2>��j��(��$U���xK�v2�m1�d�(E�J��kno�C!�?(_����7�m���Vb��o D�A�98�ڿ�d)�0>��*EI ��[EA@�i�Q��#���"����y>_9a�{���zuY49�x�Mi�ƍ�H|��"�'#@�ssL�dY;���DH-T�&���~���! �6�|9���k�s��h8d��:�)�ԯ�e�}IXQ�D��1�a��
ү��m~輋���?���T̠yȎͼuS��)<{�{�ȴe#�/���1ta �î;O�~r�g�sHa5F�d����f�tac�c��.'�<1~��}Ck [١�$<k���/?�DЂ;�az���?�B�I'#�ē���5I	�Y�l����;W>ӢW�1+�{uM��\Y��@��lN>:�g���-��)=�끨��2"�Y`�|��&K΋��pYy5]i��c���u!a�3N�������T�G���W*?zO����t!J_~����S��m������Jݡ��N��Wף��N;�47��6>{$}q*'��s>4d�^�|�{����g3OM��N���J�ݕ�R��|���,Q�M!��h4�I�mZ�0Lϡ�m*�y���/F�+�vX�Ա��]O����P1�B#]��cٚ��!�<�\����=B����hFs�wGY�3j4į�a
2{�(�:�w2�~u�䩯��$]�|cU�#A"2n�KT��-Ŧ�ٔ2�3��޶�]��0��|����_ֶ&i�qh��f�F�-�\(��Z����9{��Cr_詧�8V���h��m|��I��޹O�ȕCcFR��>��քe�{� ����T�%�Xg�HL����]E>�B2��F��O�9���������=��x���ޔ~!z7�Bd�����m*Q���+0�;(mG�DPq�K�bN9��8�]E�Q�M*wA)>s��V۞h*���)�X}B?�e-��-(D�����R��w�3��ϭ�kxHa`Yf�ZSzb��ׄ��ݲ�Rx��Ĉ�
Ş6y��@�KϠ����R}ȥ��MDO:I��>Z�/���r����X�0|�������c�xR��?w��]���9dFJ�\�9�7}�=t��~&\p0]'	Q���w�zZ7�"�����f_o�UӾ=�;�<T"����4>�$�����G�{4іj�ї.��Y��{��v�?UkX�=_��2Wn�"nK!TVߋG(������Y��$*@hj:��_���$��Qxf�c�ziM�����\� �\�S��(y�I0�*?~���-�b�p��,�	OF��1��	��:�;w��ط�Nݠ}�ZI�^�@�I"��=�@ӟ�g��A	붣~p��a��]���2G՘q	Y���Mk�֕�j�hDb�Ӎ�EUT�^�d)��`�7`n�a}�m��÷c�l᠐r�5�{BBCE	g�2N
ũ̴�WQ�}�t[S�.��&_-�.F�
�����`�T�7�!��%H"&�X��*�*fpA)����D����"�������&5b�w��(_�R���DY��/��n��������u��
��d5dL�����Y� �ؚ��r��8��k�#�ȞܫE�����(�.��j���tCs���m��r6Y�\Q�$:]���
��9�!��k�E���2�(�d�P����? ��u���'<�z����7�aEDQ�]���yj{G��ٔ{AKmuA"s��gCƍ����o,Ŏ����y�Oroɼ��?yt�����>��F�.�)m�g!��Z��=��ߡCO-?�L�v�`����}!H����`	OF��p�����0��żO�eWI�:�o�&��l�%hmn��F�VDT�G���q8T~N�N�Y"7��D���>�eg��P���n^)�H�w�J�����g��U�	s�G݁*$��=�0�O�_��WC<�p#��,ǖ�Ġ�_@Ę�BH�ٽ�6Ef5����N'v�x5�vހԿ� � ��U��VQ1�X�����gAR؝��r��3��	«�kX��;�2�VDT��0��f{I�ܾ6�$����h�p�%�ꎊ:��a�e���EW�/�U/�>Is�D�tLQ
~X���j���5���o�J�]��s��!)m-�Z�#��u�,�
B�Ko���a�E�ӏ�Go�_�xPт&.^D]T��0��\V�S/���r���b7>J�^� i�G �����ȵ5SRⲉy�����('Ia GF��S�����ۭ���G��ܫ�����]I%�&�ɲA�	d���b���a�+G����Q�%ЗT�j�0��fé�OgtR�8Iu������0�G���+C[�2i�f�o؉����D��?O��f���'�&z���0��h��&H.�M6$�-@ºXbaJK�%5��H��<��jSB�D��(��>�2�0�	�����F�`mE�x�u��ٵap��N�l��Ɋ{���1�0	��9p��zcԻ�a�	.�a|�SAb�a��`Ab�a�$�a&(`Ab�a�$�a&(`Ab�a�$�a&(`Ab�a�$�a&(`Ab�a�$�a&(`Ab�a�$�a&(�SA"[sGx(�͕-vџ�:2�0�v�1�~=�3T����J�!�������=^�IX�`�H�%� k\d�=ݩ'{X�ڲj苩T7�c��[l$
/<G�~��ʺ.��� ���D�����h���"���D��DTNM��;�!��P+�a������A����%B��@BV9~�����n�:��w;�0\�E�r�Q69ODG����z�`4�@Ҫ��]�a��+A"�(�4��"��h�P|Ɖ0��A�$L
��0L��ǂD)�}�N�%%}���#���*(m-`�a�=$�=�N����Ɯb��s�`��,J�0����tE�'1ra����i�0`y>���a�	>���8�P�T61)���a�9��I�����jGdC_R��B��c�9ڑ-H�P�����Iԍ{xE�F�Ŷ4�޺Zoo�b�;�i��NrhCϗ���-z��ہ�yЕT�|�0L��9��j����Q�ٶ:\e��$��
�>צ��Ѕ�gI2�����+�O@U��P��hqD�)y�zS͂y��{R��2EU=T�Ȕ����7N.Uc�!i�f0�0�1>�x��@O�g��I�N$DTr����bCyø3���R��S����Ǎ��Ny��`Xg�HN�{.�*�߰S�2�0�ӗ�/���9>�E���U��x��l{���3���}�ZcV���S�BMn��7(�:D�8c�Cm��R���l��d?���q��h����9�t����X�TW¸�0�	�z|��0J�)oO߬���k[g.��zf�)=Q���Dº�������z�ߐ4�r�px���
�K��^��� ��q����'_v��~��� ]�a���H��r�*H�D�l�n��b�0�7o�c����֘�b�^�5<k����mE�O����/��Д4��+�aٵ�IDIa���	u\<R�zf^�us�[���\�a�#͑���U�L�	��/,}EnNR,^Y�ᕺ�kG�\)gSZ�O��1 ��?�2���UÚ|���6u^����ċ.E�ˠ�G�:��>(��u?~#�v�0G�#=>��{��,ϫ�ԷvS���3�����)���Uؒb ��;�B��4�����?���9�g-ڃ�E��썗���I�Ǐ9�L�x�e5b��`Ab� B����OB�IS�2��8��z�4ԣ���M�_�#�۶ty���P$_v������P���n�K7�qgL۴/��=���0L?��k�F��+��� �	�"�g9x$k��h ��jc���b���m�-��l��z�@��F�>n��!ҍ%����V��C��W��vUd��}Dl�r��+�0��p��H��f!�#f�Gqg�����e�Nx�YT-�pv�	C�����������`+-���ڜ���X~��I��2v8f�H�B�V��T-� -5��'�0>ˡ[Ar��]��t ��#uS����o�E�V�Z����c&_z�{���e��g��y���MB7�G��o@�+�0Q��x�C"���k���F#���!E)QN�m��<��ط���=~�F#	�-�}���r���{��:$n!:��EJ�5@���μ�n�]s#�-������X.�0>ު��}G�p��
olZ� �������p�i�
�w��Ɗ��߻�}%z�T$�w�(�s��m�ł�0~��QD���$�Y�qi��bN=��>W
�BB�=v��!�F��s.U�T��[*?|�Rtv8T�KKM�.���ӧ�9��OA��җ���x�#���%����K�$_������ź@c��&w_����t��>��i���Y�:=������W��C�0Lg����[�(M��/�v�kO�V���|��o�D���^�m�|��$�J7݁��@�Z���J��bΣ�n;���´e�x�_ֆ���ES�M�����Hw.���J�-w!49U�䅧�0L �n�(�%p:��M�����⃷��f+;��ů!��kEAR���Ѹ>�ک0��Ef���������.���_����s|�V���ŸpF)�K?V! (�c��޷����]��T�9�$$^|�����w8�,`��D�:�!mCB��E�A ��Z�E�R�����K�A_P�d1���Gx� D��ղ�sb����%V3�0>{єnI��,�<�Dj'#@o�9&l��[�7l�~��s̔'�-!a��~�qq�F2���a�3�Nto�~�e��c��ÁמGƍ�#�	��z�~�G����l)2n�M�3r��ɗM��q��g�/���*K��J;{X�ҏ� �ڰ��짖�UNT�h8�?V\����1��Z�{�^08t�G������_��+H��r�槹��߉��@cڸν�1��>!v�,j�#��m�����y�C
�1�$C��R�?�9\sђm��*|q]Nhyb�H9����󗳕�7�gBo�2��9m�K�B��;D����P��B�r?O���&0#Ul�{���o���{ɿ��
�����D$������dA�[�����n~ė�Y^I[VSz���@=2�����Ï4Yr^�G��ʫ�J�-&�U�$�j�3N��zzףNHt�����莨�N��_w�����.��G�κ�a1w�"�<����Z�*d�	Q�vʼ�b�-�|�L�Lrppq�nO���bʖ���WÏ�2>��� �+P9a���5d�^�|�{Ȣ~೙��Vf�ʮ�ԕV�ڏ��W�#�gAmH@�䩨��[0�8mV�6-^��VR)�p�)�'BT����x�������0'^2e�}	��}���
��٩�K���Gj|������͑���Ϩ����)Ȝ��	N�΄򝌸_:y�i0I�*�X�<�H������r�zDiwY��6mހ���������b�q�Z�}�N��R�_{�9�7Ի��Q]��XK�����:���.QY�����3���,����_/���Q��Q�Kӵ���Gr|���uH�@��}���3�R���&,�S�s�?L�^�u������U�S/$�k�B9ZM�@��x	��|��9Z,7��X?y��7}(��O�*�ݍ9���0L�X�����������������Ğ6�G�D�oE�?���y_��\~��y�B7b�{�,��ő��"kallA!����2�:	R��s+��RX��֔��,�5Tm�e7|���.�Q��l�A��|�����+ь�YyDO:I��@���q�t�9R4���i���w�����=�)PWi:���v����S�?����d	��bk�уe�:	Zc��K�i���^孺��5,M����J��k��*�d�����Y�<b��A�0�
���t�0g�Ĉ��ۯW�%�0G���V�Vd�E^s�O�;}E\#��O�a�]{�)��+�#���� 8D��������mG����� �^R�7d��1��(W��>��+�զ���9N7�UQ{y�adO:��M0��M�Ҏ��=��\q"ƞ |��;,=�H!{�ϫP�֫���+0sd�Er¦��>�����+���������z|ul��>�E�D�_�Ґ��g�2&D��v|�قbkF��(>�D�
�#�Ȟ�/=3ړ�r�,� o�	=��E74W�u�rKZ�@��,����'P��OC��0�(y�1ĝ6���T����O=,LTU�Ş>M�/L�j�_�I�6p���Ijˆ���j>"�㳯�d�����=���` vk!"��4U�	����VI3|P�ݮ���W�7�$�T��_׮��� �MI�:_���N�*��\��!��E�~��
���h���榩����u����w
6|v�NY��ё0S��#��@�Wo�0�&� s˅gbТ�}�Xs�y�=^_G�{��G��]���b���˅*z����w���W���OMC�	>���DƗ����)����H^]/]�j(=��a��"�-OG�ɧ"�Y�u_��f��SP
��7��ۯ��*	���Hl��=ose�p�?�b��<��P��u���Y� -�V��[a�֟�B�Fz��\f�����g�$�VȟPdDb��-�0���ߋ�cP�� $4N�Y,��֐� ��p���Iޕ¿�H�|9�N����v�)�M�C�l�4gDi:������������^u���]J�oЕT�lr��6=�Z`������a&x�K���K*P5vjs��T��3:EaqRTD��Q��0�/�Q��+%�ٌ�;Q����!�h�a��	�ь����PO�a���	�e�	k��� ��X��aI��-&-:�)=��	�u�������^�#�0�1��ɍ$(ڊZ��Ak2g�k��T��6��U��k[[�a�#��Fd/��o�s*C�E�AmE�J�!~,"�k��	�Hx���0�;h<����h�O�a�a���a�	
X��a����a�	
X��a����a�	
X��a����a�	
X��a����a�	
X��a����a�	
X��a���O��N8�C�8�~B�b���3,�0sl8AR ��8�2aI2�	��s�>��	a5Fh˪�/�}5ܠ�a���dCmn6�f�9B^s*=�Q9a4�fD�؇؂BI�l`�a�?~$g�㇣nx���H�*Ǐ@���B��mG���0L��/�Ԑ����y":�'$lգ�aP�Vm@��0�0��^		F��1�>��E��3N�)mR$aR����a�	z,H���7�$XR��WP:�9:_�����a���#A"1�s�X��k�)�=g
~�Ϣ�0ӏ�Y�(MW4}�#���6	��s��a��� ќ�9ـ#EJe���a����aPz�|�vD6�%��,��;�a��ق�UKɘ�D�h�k+�7���KÌ�U�֦���fExnS�v�#<�Kr\^�^�s�v`rt%<��0s�#[ h��]����&�]�^�S��f����=)�ꃏ��2EU=T�Ȕ���a"����Ð�f3�a��Y?	�\������P�0�̷�������|;�q��S1��J&�\dU�a�0je�a�Nd	R���"
K��*[v�b	�^��o䗷�Ā�3~m�J;N�k�*jrs��� �A��!�I�3����kᴘa--F��_`\�3Z�]�5��獃v�Ph�P����(�^�3�W�w�z�a�c�0J�EF=#�)�׶�\6�]��}��DY�RݐL$�+�K�**�W�I��!$,���Z�+Q�d1�^vcC�熿�Q'N��$W-@sy��w+�~��0LG�
�%� ۵��(M�1rA�X>�r�5&�Į�z�Z"u�$�B[Q��y���a�o!4��5WU��s&�z=�2���	�!i�܈ċ.ź�#;G-ETD��k�>4W�I�7B���aB�4I�����u�ը��s0�0��*H������"w�H�������kG�\)gSZ�O��1 #�^Ud��wÚ|���6u^�6 �3g#q�e�HEvz���Ѵ�?������9ul����s�P*�u�#����fv0g�q�=BJ��UG�Q����g��S��#�GI��^�qJ=�[�J_~��|H
q<����
Q��~���2�>���җ���\-�5�s�P�{��ψq'H��0L^�!�@��U�(��ӟ�m{o������EP��(�Ǎ=c:����v]�w݊Q{�+˱����	��}%��$&�a�9D���T��l;��@�G��U�Z�ku�Ui�{=f�W����~X��q��?O��n�� �0s�n���}��Ʀ��B��d� a��D�����b���w��mA�		A�g�M�c2m� �a�^"$�N>�z�v��n��}5�^���sH�is`�Y�2O7tR.���O�U�;��3�����y��:�
O�r�VZs��"��v�Y�ŵ%/>���߃a��H��$g.ƅ3J9\�!/��#�����m�^W��<���n6�/ �����	�0Lg�$U��u2�H-�D�l1�d��*����5���uA�f���b�H�fial�=�TDO<{��	�a�^"��,M�*��a�H?B phCϗ��Z�V9Q������*"���΁W����?��^s�&��n�0ӆ�9��#L2�)�0����5-��W��/��	-O�	���+��j��5}AKMv�zF}��(�H�����ƫ�0ô�U��e�0�'z=�0RF�?l�?�d�y�.+��+��uL��1�C�rcƉ�]����{2λU�R�&�B?�g��a�+^I_\��	#d�!+���s��Ct���<5�2;u���u����R��|���,Q�=y*�~�}�����A�:*
�a��Re4F3�#�;~��\�!~�S�95�K�<�:�w2�~u��EG��t��U��|E���
_9�f��P��+��",���GO^�0ӟ�~��
D��'Z�ˡ1#)Ea��kk²�=mC!	������)r_��ȧ^H��F�_"��i�*�V��Z�e��EGE	�'�v��Z�.tU(�y�RdԶl�~�`�a!+o[P��1Cew�5f��yW=�h���q���(MW��֔.�}4�nG����;n�6g�h-A��
����0A�"J}�'����W���c���ٗ#���P�d1���$:�RZP�VCm��n�H�u��br�.�50�0��%H*��M�F�}`IPR�1�ҥ�4���{�"�����j:KӠ�+�R��Mӹ��R����>�j�\4�{�'����td����[$�F��#1R��uX�䩬;b�X�pA��ɭ�ι�9�7ԃa�9����u�Q?8��0���u!5yC�3.yoA�f���c�ѺR_m�Jϛ�t#�c�&۵a�'F������`X�s=��W_"E@S���)
�h���7��B�(�����Q��;�e���.FU/�H����}1�0m��[3�Wn@�'�|*�6F�Q���k�SVn�e��U?�����.�T�@v?͕hڽ��y"s�f��ob��ڝk��E�r���F4�����=n[�0s,�S�q������nx��ح���SBE�����RE�e��0���ϋaRVm@st$��.��;P����0��|$�݉�/Wa�9S`���� ��^���P88�0�_�]��ւ�e?b�Y'ɲ�'��50�0���א�v�)�M�C�l�4gDi:���a��2T��]J�oЕT�lr��6=�Z`������a&x���gTa	�%�;���p��8���8)*�uF�(�f�a��YNӜNҚ͈߰5�9������P͈ٹO��ā�a�9��{e�	k��� ��X��aI��-&-:�)=��	�u������>�2�0G?�k�#	���V<p�ڇ�Y��08�m�i�C�dE�=����a��O�đ�Po%�a�9n[�0�,H�0LP���0�,H�0LP���0�,H�0LP���0�,H�0LP���0�,H�0LP���0�,H�0LP���0�}*H�v�
������D�a�a�c��	��$����K�ָHص���,M�1B[V}15��}�0�~${xjs�Q?4��Z��P�葞��	#�i4#z�>�Jbe�0��� 9C5�?uóDg��@BV9~�����n;Bl�`�a�/~���t�M�ё?!a�=�2��j�v��a���J�H0�'�A���$-�0�q"Li{�"	����0ӿ� Q�nߴ�`I�G_A����Hd|�
J[�a��C���hϹS`5D��1����)�i>��0L?�gA�4]��GD�\X�c��$X���;�a�~�ςDsF�d�4)�M�CJ�o`�a�~|��A�/`����ЗT"�����a�vd�#T-E$czt��bזWmTZ����V��[�v���#m��Im��R�5�E��9b;09��
�Ob�9ʑ- �Pծ����GԞ���%�]�d����+>�0e��&'�i������앵��P5v��l�0s�"K�H����t��ņ�qg��M������ۑ��[:{��������T��"���;�Q+�0st"K�jG��d����Y�LP,����`�ʲ֙�|�e�:cvZ���8U*��� amz�R�C�	�1f<4�		��i1�ZZ��u?ø��ڻN���!��1�8�Ȓ^.�����[�9�(T�n���&D���E:_�w����.P����������UL,2n�]l���,l%��/�Ia�*]Qف�͟���]�ܧ���u�q�jf��eEJuC2����G.᪨h�^u�.�\��.�k��DŒ�({�E؍�߇��!�o�@ܴs�9��y�]���K��h���=4�놏�^���q� ~o)܅��X�ӱH�fΆa���˅RG�Vip2mZ��������#ǟ����A���g�ntZ�TU�q�:ԯ���|��3�"q�қAs�$?���x��]��]� ǫ Y�]�i��Pi35�npD��tv�xkLD�]�}N�%RKB,��>�G;h(����8\4WU��s&�4x������L�	H��F�~)�M��?�	��qѡk���e�V8�f�J��s(�JĞ6M�����ˢ�$�)W.��[³r0�� <gp��+#"�8�Gn�_)45�<��'wz�����dI��$�� ��z��,��h�a���dJO�}��=�/˝3���^��oͨAW��ߔ�� �]��ş@%�ݰ&�O?��ͿuJ��Ȗ�h6g͕D*�ӱf�>~՟}��- ��a1��5F�ۀ������h�R�b�ln�e�v��B���8t1�����'�����"2���B%		�h5	I��f����;PǵYi��lD�M��,E�U"J#A��8��^���AH��o8���7ԃa9R�<�:*��T}=�L����T���SygI1 ��W�Ta�/�ň����\�e�ߺ�E�ޏ�7^A��';<Gi��N� {�g1��ߋ�W�Bޗ�ĀE�=��.�FLg�W|�ڟ`޶M���b��;�RG�?HH�zZ���ɂ��/���5�v���=�oo��А�^o#�Fd�#����W:}�(*6l�D�$^|)2�q/�9�WA��F�:Pxy��y���=�0��ݶ��n6Fh�.�����bϘ}�h�M���Ĩ=�e�~�%~g-.��:�/���$ϹR��S*ɴ�]&<Q��z}J�E�;Al����ȍ�w�S����N���a���n�ou�Q��aڼAD�r����lļS�o��.�y3��	N[�*Qi>��aj��1��'D�qM��C�`�:'[��'�$�4pv�v�p��� �MMtl���"]�S�BH��)��Ke��~ط/y���:�6�p���Ȧ����v��Ο%��v��~�i��w�~����m��+�Ō��A�Suy#D�e	3.FĘq� En�@������J��UDO7j��l��o���}{���f�8C̣T�S�ɇ(y�	��>���k�M7{�*M�r�ϻ�]�B�D�/�D��m�#|`6��]��SNs�XI�[��_E�W���t+H�p���a&s>��޺R֎
���*Ht���+�)%D���@;x��I�M{~�R�*݈��>�9�����SE�BT,y[�m��$ C��b�pV�_�g���
'����$0�:�4i�\$���i��&�җ4��r���p���v�E��8
)���7"49M���g{H�R��VD�[/=�-�%G���uuL������b~���{�2�,��T{��H�{52�q�H�tcG¬IHgzPݞ�o���?sD�!�w�Q�۷#@h�u����Ш�-��Iw����
� �r�L9MlY���)�{�����5o�(><㦝#Rk�v�tC�5_.�]�֫��YsAW�8�2�c(}�9Qa-)BXj:�\(�ul�4H߃��uz-���e���¸�gwCi���3���;E����Ħ��t�6p׃"����[�h�s�DAFڵ7!�̳EY~�%�MS���z��bP��#RT���B��<W��k�-���� E�n�_lSy��'��]S��)R�D��"EY�2e�^���<�XN�?�G�^]�źJ�z�E������� 8Bۙ|��c��$.��A�E*��~�%"�֣s�\�'�]-=<�'(�)�ㆶ���P���ߏ���k���Š|�\L��t�X�V�HBe��F-�^�EJ��q8T������	�����
a�?wf��������E�_z/�
��� r���:���Hù��w��Q�w�k�v�.��G��B�"�GŇ��Z���nI�\�g�r��c�2:v��}���U(#�r�{������!J���W�-�Z��Ak�\��>�R��
*��9*�����犻�a/-���N��$�*���h��u=�zt%U�| ��@ZG�pXd�I��C�a�O+�����4�[A�����}�V/�H��vȰ67�."��_�t�Ǘ����<Q{7��/q/T�
׮R���-�l��=^� i^�9:�V�TM�*�K��VD�l1�d�(}^�V���~�
�@B�"��R�d4X��MI��>��o��=����]7����:$]�!PIs�ч��
9x.?�]��)x��� Ԇ�e�{��F�4�ڭ�S�����Uw�
�6-&K-��Q���r����~/�u�h'H�ƴ��hO��pZ��b5��S��s��%Bj���$���~��# �-�����Z�V9Q���Н�*"���(��6}av�8�']� *ovoKw��tw]��=�;c��������D�U��<PY����nl[�Jw��A�
Z����Ci���!!b�%�/W����Z���u�ט��PըHGwu�����v���9m�(E>���A�ש<T��&�Lp�u)���AjJ1��`�pMm&z��儖'Ə�Bk�\le�� �Y�ڋU2�fN���	�(E�U	�ɩ_���}�y��w�a�^�@D���K�ȅA �@X� q>������J�)@�TVM7b��mK"�;��N�K�������-={/��EJ�F�t���Ps��U��e�0�'z=5�SEd<l�+�H�%�E{D������r0o/�@�iZ�A)F.��k/F��/�DL�о���HC<�J3I����t�W����O�:f���nÈ���M�zJ��S�bT��?�����X�COw��6�;Jz~^��E��zM��[��x$}q*'��u����+�ϝr��o��|6������9r�וV@t�X�:_��t�%��s���Ś	�-Fl�ڧ�BN�t\s�!Rmq�+p���BY��R��
��&�$�z$Hh�-����д;��2���H�\�8��GH�5��h����M~s����?LAfo�[gB�NFܯ���H�`��U�ڞ�7_q/:���?Ѱf�l*+���brq������A�u��E䄓�g�KA��ܶ�[��b���P�r��E�Z��{��z9МI�����<*��U��K1�x��v�k���$�$���L���:$��/z�>��\�I)!���&,�Q�>qJI��K>o�9#1E�k�w���Je�?Q[K���h�����:�{�t��!��<���)m�u�,FAB�� Q�-��<��𧅝-��)�X3��I£0g��Q_+�a�C��,��_�g��}�auQd�y�]~i�h*?xɗ]-R��q�����s䑵06���c���ې�vܻ���ϭ�k�n٬�R�I�YkN�/F!v;b�솯��C*��J$����(y�i�}�UJ�DO:EرК��*��4��'ŝ8�e���ۺ�+Ȯȓ��f�6�cu�����F���e��NQF���!�"Bʾ쇉�����lhh�RO�t9|StL��_� ￍ�%o�L��ATm�`��)�/�یJ��q�(�"������+Ϻ#%��(@7O���~�M{E3LZ�D뮆H�OѢu�ސ`E�=^�5�|��_�-2}�,ARYlm�4Z�$�)=1��/]:O�8\��*r��n�uW�U�S$>S��|��4���-�PY}O��d/�B��BT(����ǁ�CKm���Q4�#��!�ڡ1ڽ���<��}���XX�<�:��|��9�����"K�V7�š��?��eb����>�.���y	�DA���oݖ7��eADQ2�I���]N�(�C������ ������q�D�7�&�Y��N�%!E��k{h vȘU%}��P��6���������"K��Y��Д�`�^d[%�ێ�����A.v�.�&o�ec�%�_7b��l�8���J�h3�-��lQa����7'ƍ����07����6z$JdCs )�_��q'Q�<{{��˥/2<��?: �����w>("\*�v�f��}�h\��_�G4�z�u��	EA����uQ�$�B���	$���^��G��S�3������_%�-r��;�Q&�~�H�� �Z����z���Q�&�oK�� [�Bl�H^��g���IZeC������Ϥ��(�.�􁧇H	�Q-ȣ/qse���뮬eJ^xR<���ۯ�ihﻸ��?�m"?w�-ŉHƲkG@J���m�w
��A��2��5���Պ�QW��Oýg���Cw�?Tp���Y"]��+\��������w�xx�u9��5_|����'�|^�1�;
d��TPDVET=IBD��<�l]P$��x|2W��]S���B0���{z�j9��7nX�A&Ԉ�ϐ"j*n��ޡ���ZN�ȣ	[���e�ы�n�)�6�9:fj~��B��`�a�>���DƗ����)����H^]/]�j(ܾ�a��У~HJ[�����g�$�VȟPdDbD��0��zܠ�\�3�H�lbjGd�/�9#J�qd�0���U�XJߥ��]I%�&��jS��Fʊ�~/``�a���0�*,���Uc��67N�:�S'EE������0L���@ۼRҚ͈߰5�9����ȞY���f���'�z���0�}�M�\(�lHX[��u�$��Kj<l1�h�yN�MM�k�����p�fE�a�c
��IP��⁃�>d�j׆��n;mH��&+B��֛a�X'p����0��g�P��<��g���SAb��B�"�E�0o�ԥ�`02��u�ɨ\��w��x��	z�*��p��(~�Q�<���_� 1AO��v�Qۿg��ŧ�޺�a�#�(��)�\v@tB�F�Q�O����?� 1A������;o��^�*2
�R�Ă�0�$&���A��~Z���}�ċ.Eܙg�Fx�Fc��Տ���"uu�.�`'U���ס~��3iWP��:�j�:!����	[E��K`��R�]^�C�C���:Xv�����Z��ɧ"b��һ��\4��θi��aٵM{v�a�$&hQ�#܃hղ%���	'A�ξ�i�⃷�|}��"�Z�[6NCΣ�F�)�uڏ��^���Nυef!��O:��?�ݷ]������Ys�q��K��P��}��+�{W�F� �^@���F�7݁�����o"�$�?� J�<�	6X����0�\��kE4����/		E���$7!J~�5D�0	Ƶ?I�X'7��M�n�Hy�5l��ٝ
%TB���8EC��[ET�6$ b�8I�NG�ɧběcˬ?��辒��f�I���*?z��bh��p��ŜY���H�ǁW�����9�1��%"���҂�O?��Bz�Tnw��u�`�`��	Z���~]ہ�N�"JZ���oE��b0nڽ��ㄥgB#�ۯ��+���\ֽ���D?�8D?Q��CQώ��A݊�<V�����ב:�z}�	F����Mj��Wl�zvQ+{�e{��^3n���~b�F���G�bDk��͛	s�f��￉8I�?�"&�aAb���D�ۇ�������"E>!"%W���^�W����Ĉ(��H��(Tj1s� ����q���zο��xP��\H�HT��a�M�;EX4w�������+�� ����ڹ��)�(O��gu#5_|����$EJg�a�$&(��G�5_-�𜭬TT�E�8��\(��Ch�wߞ�z�G�\U[�~��FX��]k㺟�OJ텦��t�����׉��?�8�EX��Cݏ_A��4!��p�l���S��Uu��sRTɂ�;,HLСP�?c�خ����d�EI$H4�Cs8u����h��^_���r!H$]�5qg�I�7��ms[������$���"�#(��Ƶ?A�s��qGBT�GP����¼}&�aAb�����=�C�����4�ߝ ��u_�����sKqP�C�y9=��i�Ⱥve���ɪ�X�vWё[��ձ�Cǈl��k������^T 2L_ѧ�Dm'�pl?�l���I��a\��n���9�B�����.k���_kϛkeݷ�M��c�~�%j��M{~o�H������ðW����
E;�f��<�NJ�po��|];k%O�� �s�� I�KBL��$`���]��K��4!��mY5��Ԡ����P:,f���S��T�@sI^���B��t\���g����]��g_#{�!�rUL,���_ܯ��?�]ז��$&u����T0L��wA����67�C3�!��9	��鉨�0�F3�w�ClA�$V60�I H`������������CDG�&�߂���sGaU�,�z��������w�;��./W%ER��Ce�47D�}��(��"P;d8&�� 9C5�?uóDg��@BV9~�����n;Bl�`�?�t�yG��E���=�s��6g�Ӧ��v-!�a������k;�}���R��҂��\讞k���B�q�oJ���Ү�Ql';E�<��K����`�`�/�Ԑ����y":�'$lգ�aP�Vm@��0��d�����l��א+	A��OA����)�hٽ����q����Q�������_$��q�]���?;�y�=�����MhX����� �/�E�o��F2o�K,�e�`�W�D�Q>ij��l��\Z�a(>�D��� E&�����Gܑ�Ӊ���z�?7�."%������pZ�~��L�:vڂ[���g������.�\�dg1f|��Q��b�@\��\)��*?|G���$�"�K��{�IW�ŲN�(��ߑ��ra��u�c�@χi��������/�.��ؿ��'h��ǂD)�}�N�%%}���#���*(m-`�T^'	
AVA�e�K�Me�p�XGD�-���9��~˵��{PKb�2��hO�{oH�[��w>��I$��y�\z�eQ-=i�x-�}�u+iި`���y��6;%I@��:>�Q�S��a���0G�	�ўs��j�F_cN1`�9S0��|�~�&!��֓o�T-{_�G"ڷ����-5��.%j�����uz���7��)z��RC4�C-'*��Ƹ�Q�V�J�{6�HN����$Er�-=���(v̟-ZG�\�n�!�t2s�b2v�J�m�u�(��K���j�\U���W
�VWO)�.��0L0� Q��h��#"F.��1�?m,���]?���jL��zz-E��y�ri�k�h}�����y�r�bȁ��<���F��L��<_���ۦ�M`�`�gA�9#s�G���&�!%����!'�ԫ�&�)�km�0}�O��0(=��P;"��JDr�sl3�e({�eY-\$��#�?r��D�s��a�ق�UKɘ�D�h��WTmTYlKC뭫���-f�S��葶h�$�6�|)�ݢ�����]I�'1�4�c' r�	b���ֈ� �\�ڊ�gu���0G�@U��P��hqD�)y�zS͂y��{R��2EU=T�Ȕ���a"����Ð�f3�Xe��� b���uBBS��褐���U��_��~���I����t��ņ�qg��M������ۑ��ϝ�H���Μ!�|����7�F�s,R��+��捜�͢��-���9>�E���U��x�8�#g��_�:���g�5f���:U*��� amz���EZ䨉O���\�n\��(������1�B���F���`�a��Gb��	�0J�EF=#�)�׶�\6�]��"Sz��H�nH&���%\�ԫ�+ﻳ�'�1�e)��K����#�s��Y�h�;<���1^{�0��x$K�A�k��d�S��7b䂎�tv�xkLD�]����D�`I�����@�iC_z[ث����M��D�Ud�$6��!&�Ӯ�	������"Ĝz&2n��0L��*H����,,}E.X����+u�׎̹R����D�����?�v�L*��~T8*n�Bc	3g#q�\(��[]����u�z2�4�}bN9�0�w�GH���(:��T}=��6|�cc�<{��(ɒb ��;.95z�%�������請h��B=z?��x����|������D���S��{g�T���7��,M�tߡ-��(�!�>��q�Qtd\���FGg�yF�g�q)�����(m龤MҤM��=_I��&�iSH��=O��&7_n���|�9�a��G@A�����U�n���= f.+v�u��m�F}��)F����f
�/���K�b��~�wm��E;k昀LP�Ι!|��^|����Zc�׊������A�%W�x��ZN����$�Z���ᨭm���uk+�P�ڥcu�U�hw3庹]�e/>-K��p�ޠ��W���]�����>���濾R��z�q�r�`�?�W^/��"H�6I����`	R��S���t4��$�N#{ ��Z�AB�d_#kG��j
�s'M�t�H�>Lx�P(��u"��Y�e��x�
��R��!�l(�e���"풇�F��o�ay�����MΝ$4͍;���Ҩ��OԄ��E�FfLXB5_�$^z�^z�odJSS��
����l[��Fp�/!����V�r<�!��Ʉ'Mk�F�爔���N8}���C��s��w��
P�#�1Ӊ_A�����̗~�� ��5��޷-p^�2�;��i��	O(����j�A�" _������шv�֟��� �z�4�<X�4���N��ۃxoz\�lW�>ǉ��.TL��ݻi#��$Uk�b��O� 	�#Nw��;�/�=�1{��S�7��~�����]�}�����#j>x�x���ƿ�)ԦT����|��x�����hS.�1���c�+뾇�~�==�9��e�탠b�>.�C����S{�w��_q�Y�*^{	)W߀�kn��}��\$VP�@�rTcs��.�r����OK`��sF��c�+o 23[��{\-ͽƥ����~�qp۬�~W��F������I���t5�.0j����;�%*d ����v��>����#c��H�芮B���BūK�DH�P�Zee�9��˥�0P{
9���c�չ���T�h0�K×��+u�����^"��/<�(�Z}�ι��x�1�IJ�%���9u�E�����Cm�7o�^�oJ)��cm�N�dk��3a�_F�Ix�m;%|���w�:-[6 X��Y&� ұ�+E������.@�w�����xaƯ�H���ǟِ��~�]0�3Cl?��^b�p�e�}b�$�Z�;��)���إ[��3���[zyA�Z���IH��7?�=�_T��C�5$m}3,2�5-a�;��5W��!?���g�"��'@����&u9���/t���G"=:�z	Rҡd��o�gS#�&��MJ*&��������h8��z���+~u|�(ަ�}�\ȴ��1G>�H��I��^x��Vd#E���"���˗�ꍿ���^<L�$9��DO9U���PU�a�m[P��I���1!\�߮�����'#����ڏ�E�wz�<��g_�A��Tx�qI�(-���ȼ�Ai�s������"���5�l�P��?�V]-�}��~wkF>I_YKfr��@=�T�,)6�1!�Ֆ��Ө�5�f���5�ug���zJ��i�g_j�[�����S�DW�	].�k�}�6�����N�����KbD�%H')լ\!�s>/"��yw���\HD<�V{��k<�N�s�5"
����}�.;�GV ǜ<U�3⡅hټ��]"���D6��t/����cӔ_���:��M(��
�<���2]6�$�O	�~�>�@JT�����tU�}�ه��g�)��5'��5XSN�-�̙���@�x���5������PQ-k?ZC2�_-�@�n$��3�[�Pc9:9��wMR�g��u{}-�V��
���}��y�M��0O�+%^|%J�](;�<�Pq8���8}Aj��O ����p�xƎ�(�V�wa�_��pԒ��>kr�\"ֆ��w�;��ڟ����]˖,�!F�T���(b�K��)H-���!F��$p�TSM�mс��o�%!q��ӑ}V!���A�,(�̊��e�i��X�OWP�:	A���o�����C8*+�9�+����J�S��ti�t]�G�)��
����x���I�(J�f����$���vD�R����~E�y÷��\�*��+U��	��7�OǄw>I�e?N�ig��n��s|_H�ռa�$O1��cd�<�됤���]�Es9�d��E8/�_GҪ��ۆ����K7Z����>'vwiP����[��/�%\�K4��W��׿�a�G>���Ms��h%2�_,�SM�u�ĝٙ�M�uÙ@}�l{~�ڦu9�DS������B�;����0P1��G#�-���y�7��:��+ҍ8ԁZ��q����9���'EþpT3��Uk**Aݤ���ƚs2N��z��O��L	v�n��禽����)_�"�N��#X��E���Ў�BS�I!ʗ��Ư�-�3=P6M���-��U��З�������:y:��#8����m@q�C'e�wk;�L%饫nZ�'ۧ�S��m��~w��tm��*���#;���  <IDATq���Z���E^�������3��d9�Z�'Z
����Xf�#K�T6G�(M�X2�3�qQ�ݤY���7�\��������K�S�ɝ����*{��}�����è�^F촳E-�����P'���Rw=W�D���;J[�}�V�c=M8��JY����H��&�pȩ}P��!50� )�J]w���&kL� Z�j��?���^׷8�1��9/F<��f_�g������)����^�M��?����6�D��,8uZ��e��/s��%�ڷ��Ai�i��U�8Ĥr�1�xG��tW���m�������X[����W�$J�N�)��0N>E\���@�)�J�� )-���#�$Q�%]����t�}��|��s���P|��3!����k�G��==�%�k�'r�9� �)i12�'���{D鳽3�ڪ
��:��ܘ��!H�6��ق�>*��2�f��VPO@�I[�U�]P ��|%n�
N�u�G�|���ji�Ή����f𠌯��?�lـC�G������!�j}wB6�pr���;�B��D(��6Jq�e�szg#H�͊��ݲ�l����\$��@n�� ��Z�K	w��(��n�]��[�+�\h��1�ǟ R�&(s՘�rX2��1?���D��e���T��2�	Y�P=
�&3�x�H]�����3:�g���c���1ilo׆�@5=�_ѧ�e�Şڹ��O��6$K$�.�0Z�;�pU�4�ߋ�_��믈m��)�	g����aۥ�:-���̻�ٿyEs��w3<��;m���FÚvt+�k��n+�crc�#C�W�v54��q�}b��#Jt�'����=>M#�葥5Ƴl�,��H����gR��1%���'Et���g]����y�5��M'sZ�$��qr�x^(�z�Ճ2�(���k���˺D�fF/yU���%�X:��C����6�:�*~=�Y�ߐ
}�i�x������w��
Egg]I0����z)fx� )�nd}��.�{b���&��A��EN&8��),۷�+����N�7¶g�p���*y�WB�����-Gޢŉ�,}�����
�����[ɥ�^�_�o$��$`PA,%	�O�߀���Q#���gB��47J��R��Q�5e4���>]�h!B{~sg��T��u%���qǽ=��V�.
���?~՗pT�����F��U,fxӯ~HJG;rV}�3N�e+J(2"1�c`�`��O���H��@넞N�m��D5A�"^2�M����C��Y���ji���^�܅�	��m�L�/z4��4���5?G��;�:�fq�$�=����y]�p7�pwF8�3/FҬ�b��?�����bN=CD����ڑ�+K���[6�`��\��%�X��7��F�2Û~K�U;[��*��a\.��fD�t_hJg �!t���?�<t�׊4ʸ�����)%�@���:y:��{�����c���Ow�.!z)�!�z�MX�n�nT�{���*NS��//Q	e2��R�h?���s�?��J79:�&Il�&��C	E4�(���{�|{ �<N$^�c,Mߥn�����
d����#m�֐'00�6��a�u&˪A��r��j[�I�f�z2�	I�rD�W�����0>nUh:�S/EETg��n�a&|	�r�s])e�6$nم��yh��v��}�n�"n�~a��af�2A�lu iC�6��d�%#��D8��n�{JOmiEd�Y�3�µ���a�)B.H]H���n7��!sV�^���e#ڜP�����xs8�������f0̱��	R��Po%�a���G�0�GT��a�,H�0LX���0Ä,H�0LX���0Ä,H�0LX���0Ä,H�0LX���0Ä,H�0LX���0Ä,H�0LX���0ÄGT���K	ס��v��D�a�a�c��$`K��%+�������ݠOek�����:D�Q��zn��0s�rAr�h�����h3�kaNBe�[f2jNM��?퇩�D+�a��O���A��|4��ΰ���f�8�M+D)i�ND8��0�_B"H�LTN+�Q(!a��8�QYHY�1��`�a�'$���'�!$�v�e�
K�^�I¤p��0�/�-H4E����`KKđ���b����Z(�`�a��$��O�=!GkZ�]4#?*dQb�F-H4MW:s�Q#��8��t�������a�	A�YSp��H�rj�
7�a��%H�Q�����rU^��ξc���$W�Z�H&��E��S_U�Ui����X�4o��-��	�X�T�Nw�-5��=Jt�vpZ�ռ��03đ- T���G7x�����/���W���We�C����>]U7��%+��`��\jO<)뷁a���:�Q�u0ʪ��̓��5r�?��ЉB��ɜ��4'$n��)C�k�UQ�]¨�a�����qyA���6_]��I��p{@����cF��dCsN��9B�J���yH�P����s�4'M�:!J�.���h��=�����S���4$̼�Qc�ף��M�W�i�W���0s,X�F�r1�VL���Ɋ��Ũ�%%!똵j�?ճ�[2�eEJ�c�����_.��8�ߺ )�ތ�o����ZԬ\������>\��y���_C�R�x(庹��{�ö{'�a��$[r�l�nZ3J�i�tV!���D��U'��e�(}��=� [�	�ꆠ^G?�8�]�"Sӻ�k���m�OpY,"JҎȅ63��D�ϿI���Ʃ�{��!=�y��b��Ҍ�/>���ÄDO>��1��ۻ�~�"�b�a�	(H��$ك��xU._����[�7LȻE�����I�5�W|�1Z�޴����,۶��7;�W^��o�2���q��q�\�k�m��#v�r���<�\{#F>�4Ԧx�>�;�\�a���R�<�:J����.�����斴����Q�--�$o\�R��K�w�Q��q���������{Q��������,��xƝ��ho����#��Ϳ!������sĜ<�SNA���0�tP��&#䠫��zӦM!_������֝�5����Ο	ø��v�7��+F޴�Ta�m����D-n��b���~`_�ϭxu�$��X��a��+Hn��g���Q[�>� ����/�(H�ұ��*D�^�J�nn�v��gd�Q��y�(ԝI�u��|�u�v�UYx����0Ӎ_Ar�4��Z��$"����vT .�&� QzwT��b��d�����ӵm��?��e�f�K���	�!
.��0L�I�����9h�̚��r�ui�P��0~�XC",�nΪ�]4�nn�oWv�Bm���!�0�p!$-��˭�x���mGEـ��κs�����x_�z�0�*~I�Z�w�2_�!oj-H���|���ΫPFw'?8C0e��^gs�����e�u�!
�0L'~I���آ��0H��ӝ.k��$o|���=
�|K$�x%9(TJ��@
U�G��p�0�0̰!@��Nn�2�ZUz.� ��G^&g?�t�r�:����Gu�i xG=��X�٫|����,�6+�a�N�!i�a�!H�i	ߙ����f��|� /�*9q��}#̐������.g����*&V�*��{�����z�0̱D@A�W����h7P#�1s��6��V[�+N�Nּ���N֘֝Ep�[E�b�4YL�u����ֽ�]���`��}�#:;��t��t�a�N
RTY5jN'k0sN��O�L�ZH |<���������o������4�+��P'$!v�Y­���vug�GM(��������X0Yl��6C�0L'�#��zh��h���M~s-	������:~ŵ�ͬ��]yё�l��U��*yґ Y�=���p�ɛm$gpGeE������d!d:�BT���}>�t�Ϻ2����0L7��:��]�Es9�d��)��|ߑ�jJ�����J�d�5+9M�sbw������h��3�Λ)�B�Z�{�CL���t��a�#OaӴ�]�Q�S��*$_u���hLۛ����)+���w�0�t#�0�TT��Icew��N��T�*�dN��`��h��2;~�%39U�s"�N��#XJ~{���э̅��P��jT,_*R�뺻hPk��g"e�\���v�n�^��$^t"tz�=�{5����C!>���<��>�Ĉ,��a�nd	�������e,	J�=.�⽛4+tQ��k���)���:�嚜�9r��<�o/��|ru}���{�e�M?G���<�,r~��7��em�wjS�h-����^cQS�ݿ�c��U<g����G�Sy���.�"k�6�[��a��ȶJڸM����i!g�!��`�����k��������پ&���#=n�7Lh��Ns굗V�$L������"aS�m�H�~�m6b�������x�)����r"c�CG�HV���kh�"�����f_���,�!T�1�F�T`��8��)�[m`�az"[�"mH]�e��P�v�1��Gl!,ik�ʲ
u��[�V���P�⅘�x�UW�V�[D;�hٺ�.;O�=���AeuI-?lf!b��CP�1��d�Ec~�ӏ%��[�P�ۅ���qc�a���w��-h���5-G��Z���
�afx� )�nd}��.�{b���&��A�r�a�����ю�U�����d�
���H���a��C����v�)UN-@ø\	h͈��82b�~�c,Mߥn�����
d����#m�֐'00�0�CHZ�ǔ�#���'���p�B����x)*�:�P�v3�0�Kh���J)�!q�.ԏ�C�l��0d�u�q��;��800�0C��	�e�I�����$,ɰ�'��vC�SzjK+"͢�����A�2�0C��R������}Ȝթ�­�|و6'T�vD8���a�� �	�Vb�a��9���0�0�`Ab�a�$�a&,`Ab�a�$�a&,`Ab�a�N���n�S�    IEND�B`�PK
     ��ZĊ���4  �4  /   images/627c2b90-5d53-4228-8b10-5ea0a126027c.png�PNG

   IHDR   d   �   nR��   	pHYs  \F  \F�CA  4�IDATx��]x��>��d�{��ك@B #��вn�RF˺-��A�v mo[(�P���(a��2!��m�{�u�{~I�m9q�HF�y����K��������V��PW
H��3��B	�uz�B����3�ɝl��FC:��D��'3�v^�Xj�8��)�|Q!��I)�+){�v�w8(��P��T��q��D��O
���j��)��V�M%�-'C�MvN���}�j���DhĄ�;*�@��B;C���g���y���;��>��
{n&U�5��}�B}%����.#�oS���,��N}N���l�k~���\KPϤ�`3B;���)m�sZƖ��uͣK�H�y ¹��4�9�d�i"??�w��d.A~Lۚ��:TAE?�	�,��j^{��O�B7�A��Jj^���ׯf��)A=��6#(�g �X���ڴ�����7�:�3+���Ք2�L2�C����t���mm����!��Q�Ct�
�\������)�%��$����6�	[�s���+�e�K��(���3I��[(�v�bҐ���U���v�� �����Աu#e}�*�46P�s!Eo��L:�lvm]�K��E][5mҜ�O֐O�����9�d����}dli#bO�]SE��ϖ��zH�l%��U}4����z�d,.���}B� ] �ڦ�S'���6��x}�)���
���;�NKI�l?�L&j]���'O�����>��줎��)��+H����b�J?�2d�QˊOĨ'�rdR�:���u;�V�-?��F���]Vc���9]��b#i�^5��R��G�T\�1���S�xS�O<$^��� ?�3�G.�`��8:�6$�KJ�_A�gN����)xN�8�������*kYZ��pq��Y~P}��a��u�b��`\�ؿW}^�0轡0�`��[�9�Rɑ�&׌�i�k�$>	#���k"$m��'��iنrU��2�5�טɸ�H�E�#��M ��d�&5��F:_ѐ��p�(�K����NQྲ��t�Hrd��N1�uPڮ2J�[�f�;f@�p��wF���f�$xX�F��rd�Q��"J�~�
?YK�$�� �;�mDU�u����ݮ���ey�rLr1�!#�&��BU��l�U�H�V�H��� �cu��B<"�4	�w4ҁ�pgQ��'�¨3����8o�G�=i�#�泪:�,c�>2�tp\��3΢��fQ����%����r����YE͟,��n��\�mwK6�}�D��(�S~�W99�@�u{��J����G��[�������}�n��lTP1�7�y�xʾ��x⏲;$���J�jJ?��>�PrZ��^H��g����ھH�ߏF�C��K�7w��^U#ۓ�s�-3Aa���ϥ�L��ZO�B��J$�"���:rZ�'Na���$��q���[j�1@	:
I���i���k��f�� ��'��@ZE�ƶ%�^�a�N��F��I,B�^�w@��"�����I��K��$-��*c�)�t�����:jW����-m�36�~��E�����kң�CP#AƗ�Fj�l9ۏs)�m��s�$Ûv��d**!�)�Qݼ9�KK���W���v��?��®P��md+�!O�Y���C���/�n�2��D�/g�6ҡ�{Q�Ѓ�r�4�:6o�����U��5#i~��w��RͿ^R�!dg$vǑ(\14�7S�+��ySə�JdPFm��f�~��2��G�H��ۨ�?��c�5�ۼ����:1�`?A(�A��F����>��e'���o}Lm�ɞ�)	ESS��e���=�����/uyl���B�:/��l߼�͝ۑb�:g{��0�k�'|]�����i��� ���~V�P˪�q�d������k"=ɼG��QJ?{�����_����|�z}��@����.a�h��;B��TR����hN��I�0��N';u1-�n�^��Dͽ�!1FHӀ�5��;���ڨ?>A�q�:��1;o�VvJ��B�^u�Q幧�^V(c��(���R��]1�S��ԥe����j�L�1�)����l����ߗv����Ic4Q,������N����8�$�s����Ar��h�U�=E�gl�v}%J�\�..�65�S]^�A��z��y[F֥WR�}��������¶�>��r��N�b�4���*�wH��ȓl&����ٜ?,X���mA�>�#��8�/�;�J9PI:���,x3i3gvR��O�o�S�3ɾo7�wl%}f�ϺXR�͋�����ciYMϤ�_<��[��$8u�i�����VB:$=���H�I���ݕ��\���4w�(򚌫t6��~��mt6��(uW�sr���{e��u�aå%�:e*��I�����^2Q�mwс��ဳ�{� ���0�G�����[���SkI�v��l?�2���&�Q%��H��9����1��Y�X�Z�M*��:m��4WkLf�Q<jZ�>%O�"��][#�B~Ya�f�8~5���e56�=ȧ��Z�% 8$6�@���n���ͻi��Ұ�ג_�-�{S <4`�d� � jH�Ϳ�0�����_{;9��&�Q��2���'Ǿ=lЍ����v��bu�"��#Ss���W]�.w�nt-��/�?VY
l���Q�N���T|��)y�)�@=ضmfƏ��RCv.�)�均�(u�Lu�*�d\���/:�ԟ��Eq4
�Գ�^�^��LO]bln_P��md���z-el�I|������ꅧ)}��ᤢ����lfUU-ލ���2/�T������#(C-�qp��TO]տ�5~���1�hT���$��S͙�aS�~��Z���+���)����F�aې�m����E��=�8�Q�\��ӏ�������Um��P9���\�=��\�>���u���j$��5��/K:I�d_��"I1Ί԰1GVw��@׉�!f�Ŷ���n�^KU��;�N����$����h�=?����D��J�tH��Z7ү�Jby����}��E͟.R.☢*u�S����w����:DΊ�1��:��
=Z��Cbt��||�؉#��l/�8
����먍@ �+7J�7����U������5��l�Y���x}������U��V�E/=�J,g���)A4y���g��{��tdRwSǫ�p{��zIos>��b��h��k6��k2�Ќ=b�bR�l�~�0��O:Y�¾{b~2+�!OS#i���L'�#��͔���.�;8"���۳�fڤ�
���<�:�#���Q{N:��(����f��u/3�A���F&��G?�a��Id�:���d�|
U��7���G"��z���C(@s��l#np8�q ���|fӃ�$�Ҭ���Mi�^(���Q�`��HY������J$�}��^)�_t�'�{�Nኡ�G���k�>	^�"-��Dp/_G�	�2P[X��%Ҕj�&�~��)�����h��H��ۋ�]��~�����_o]��NM��1%�����91bנÑ�:��������]0O�K� WEi,I) _+�鯤F�ط+1��R��]ĩ<o*����ǔ.e��4��w��g2\�����ed�@�F�زA�m��GvD몥�;m�٤MJ���g����B�SN']f&տ�)	���$K��L�ܺW���&��[;��7<�Z��6R���#V{����?��uN�\;��/ī�Ŀ��~BBG'U��N�](Z�V "1�6G���b;"��Cs8܀�B8&:���E���vQ����wC%��:I{�J��,�}��>16��%I.&V��Q��L
T��Уi���䶚U�eK )/I<�s��x�Ib94����C�� R`B:
���N�,:�TX�(�g��^q�B�e������|t�&I����QkN���9�ݮ�Pa� )�COkKw e�&Pw>/�%��K
����Rj���`'�3�N��n�|^�s�5iȈp�7<7�5�w+P�GR.}#}��(@�ʻ�&��_W ��9/����
�[��e�wU=�u�А�+��rE7K�3�@����ʵH�@�`�<�"�:�ϴ�qG���|ڮ�s��K���5���Hy'�uR�
��XH�w�.�3�2	�x���%i~�7�ar���Kڠ��ר�W<�e~�*�N9M&��V��/<{�{�����xgx]z���̍;I���R˘�V�5���g�Ď��F/��݀�͑@ʚ�@�2��_��ѮN,��3�G��Ɖ�W_ �9I�ƢJ�9����'�k�K"UY�=��k�7�ңq������|�M�J؃0 ei�F������8z�ۿX#X-#xX:[*�JT�!;Gf�*�����T�B�(U���[���ZLWz�L��z�л��|�5!�Q�"�>)�Y%� =)�jرm3�^}����\�-jx����X�����T��Ӳ�F?�7J>�$���3�$��~���\�EʫU^�o�i�� l	��z�C�����JM�_��n�ݳ���{� ��)�*�zDj�� �D]��E��
վ�O�1q#
λ��m��j���M)�+\�Դ�#*����p0w�faD���ɼ*X�����5M��Z��['���^x���)�P�zW eYM��krㄠ^]�ʨ�gI��$*�x�U>��h���\�~�ujg��֩�˄�v}:����L�{�e�����x���5��+�3Z��֢v�k4�R�"�Z��6򶷩�W�S K*�i��OX �JU�YsC�Z�{"^� R>E�w���s=x�(=m����@ʃER�P���v�D�-�<H$�������]�$���B<Z_�ؒpF�"��,N�mN )$��g�Ry�Tj�0\ʃ�n�M ���)k���N�' eEMtR5[k�z�����*��:�kN?��;�$Z�w?���|W�_���_��"lh�Q��C��0*�r��;���@�m=)Ϥ��΋
�ܴd���]s����y2$�B	���>���Tw��m��S��a\�VV�#H���~_����'�iaAPry����>�!���U��z RNY7�͏�_�B���]��>T 嫩�q�+�r����Y��j����P��������A|��ko��8
�i��-5ұi=���Mu�w��L�Fd{���v� �d�o��򋧯Ӻ<Ot�߂��E��=)OGc�����@�$@ʣȶk;�wmզ�����%~��8��ق�Z���H��.*���A�=�����Л �U�6^�I��sP�䱪�&�!|c�C�ŀ)���`\94�N��vP`^q�Mw���0<6�P�~D�����Z/�+���NeGi�ߠǧQ���C�m<0��-2P����|MH��H��S�����I��M��*5���Y@0ڶ}+���d3N2��h<���i���@��A� x����xL��Q��'���kS�Ԥ����d�=d ]>��g ��DuR�B]���^�Λq�V�]��J)��X��.Q�j�0%��!u��!<;t�i%Ji�O�􎭬����5A�0�Ct�@ʋzRƇ�m�$�)%��a��0�Xl@*��&s��=RkG��g����A�3���v"�,��09T�55�Rђ���Pp8�@��ߞ�a���:���°xоnu�q��F�,���HYÙ��N6�4
_C��9 �'I��;��>�J�rֶv����+_��r�d�{����r�R$\I��C��C
H9V	|ue��m�h�W���lo|)�*ag �^{�DY�,P5��zY��e%G@��3��FNVT@1����Q�h:q�wrp�-;�-�7�1X��̠o"e�N�a���Ϟ%RoY���͍�8�s:�����`�5�Z70]��*�AD���& ���H���H���xe�Οd�<��I��<�=x_��J��@��h���){9/a m`�����7^�iH�c&8<&�d���ԱUzs�u��2�i�BI��y;��
<�&j��lZ9���8j7�]�)���m��Z���=d �=)C��H�|^ʹ�[�p�g�P.Hd(N,����H����o�o������I��[Ը�hg5�k��9�C��8n	�U/���{� SU���+ҥ�s�5�� 4�!GJ������gI�������S�	'I���dpa���6-�5;o��N���]�E��'H�铙u`��@�k�!H���P��&�
�!f>��C%�,4X�����{~��\w3U��I���w��2��3�A��n����W�|��e���?�"�0�!��Q���� ��,5����H���oJ��ѡZPLpRP�Z,�ɆCc�+������*`�H�?�>�WH.°��s[G[϶�C^�ilC.EMA8x�j(m?)�4�F�Y@C��E5]��9��c�����|(6�\:Jp�CYr�
<�`{����ى��C/�N��(���RVCȫ�BXtΊ2r��B�N
Q5�����KQ��!��W~��k�z��{_��}d��?r�w ���W5q^�'%�ޤ�Vh/�
�,m�AAS�޹x�lo)�[<e�L��<������^㲏�g���t�paOڈz.g8�����������q���!#a�ң�L ��O�����#�5z��>0@��	���Q[C���������"�D.ַE��.������C��)k@@���'���Ǯ����R���2��.jxX�0A�8 ��G��G�	J����3 ����$��� ��u��p-K�]&3�2Z(��
��x�߲���r_���wʠg���R���P%8*���۫��vZ��
tT�<�0xG89j�����|M�$��&��F����|��H��̓o*  
���@ʈR�IV���hq⦖�^�M���i���+@�.��C`;��6��Hdg�]�z�̏�8S��)7�ڐ�;ev+�>{�vҹ�с�sVm��b@7��w@�8�3��$�i��0��P!d{3.�M)��N��WJ�2 0��:�l9j)�������F�o��ᜧe���@�g1S�g�i�0�g���тڊ
�,�cf��B�[ e�� ��v�9*��EHqv&d�S�D5�+��]���<G�����U$��xa�Xd�%R�<{�����q��@��
o�SEnBA����oIF;��ߕ渲�>���O1�ȠK���c����#o��} wR���Ԗ�%�Ih�֦zZbԏHy؏�S6qn�;oPΕ�Ȫ���z�Ob�@��N������~ZP���65����
f#��+9�1��ܖ�k.�י'i,�eM�@�{���i�HxQ�|;����֟���M��q��$����[���w�M���y�l�y��8�#���������j�\�]�"����e���H�	�D�	�|)��;�𝤎�m��p^�A�k/��F�W�B�C���F��^�s������*� ee�U])4x$%xJ�p�%�3��I�����FB�O�QI��N�wN )��*4����]���C=T�%���@�1D_.�r�KС|�wԗ���LZu~Dwc�%r�6�H ��r@�R;������ )Sg ��+%e�#���*P��s�q�!C�ڰ��\�:�D|6���9`D�1SH�oI�u`.�@�vDRN����D-KS�H�PK."L�z� c��H��s�^t�ݤ���[���O��ѣ )7�)�_ eS e����P ��y+ �<U@е�s8(���RX����J��)A��_:�r[+��u�$}��#�+�#�>6�7�򯻙F1���i�#os����.-���~��>��ɇ��Q=C�j�v�Ka���D(3 ,����>5]����ץgJ�%�F�%)��ޢ�b+\���^�~Wd>�!�n�&�N:S�P� vI�IShă�r.ZMC���R.� Rf��B#�>�3�&��_+� {�j�`v�S_�	���R�х�@�x I�#,�t�C��M��-ư.! �"��ݱ�UV<r�rrHg��+��)�Y��B
	"DGi �) e?���^za\7[{��G�K��+@��>�?[N6~q�� �L_)���C�w�L}]K	 �X��R�k��Q��գ°(@�D�?4���/���?@�.w���t���.��[{R��A��Y*����Z��f�/��E�S��/hH�Y���{h�����.�v�h�H� e�#__Dk�`�Z8>�/H��k��?��[����H��,G!�8Ԣu$�Ɵ =�]]%}i�w�����܃>ߺ��&@Q��'��S�l������s{R�� )��>l1���%8�����m�
��C)�M`�/�s���ZRF��M�t
e;��KI&�k��)�y���R���r2�
��U#~Æ�	��P��h��)��!��}{X-�u�S�,��
J��GJt ee���?)_�){�[�y�BJ9}���A�bj�HˊOy�<%6�\:B=$�����;�G穫~p��[C@�g����&��4���z#ıKj�h����: ��XVߘ�q�R_�}i@���c�����b����r�'{�r2_��*�`�*{���C�+h7cHF|h�!���i��)��ǲ0��x^���.@�MQrZ!�,��r�QH9�(�C� R�!�
����^���� ��W\x_.��O�7O9m��[�-!wc}\���������˱���.���\D�p�zj�_q �E�M2T�w�@��i�ѽRf��y�(�o]�\Э�8��r�4��uU"�%����F�+�R�E��e�i)m\�@j\&箷oX��& Z#��!�x�@ʂZ��H�
;�\2B�rWe��F�B�"â�I���O��I��N�c@ }���l9�s���5����':���C~�K��37��1�xoy����A�(H�e}�2A:�x�!RL&�GB��!����?팙rh$N��x�aI��vn#�I'�njX0O�J�HŞ��]����~M��Sd�`z�z�l��.XW��fJ���ѫ�Rv��ɗ��q�CAGc9�
�=��p�B�6�+��� ���lK˾+fQryM] Rnj_�mm e�𞁔��H٘�O��g�i�M�C�B�  yܳ�P������M� �U:BE�`�d_�-��5�IuQ��G[��p,T�:8@�8^z�*��k��l/v�x��t���K�R��oP��P�Y�J//� � ��RWv�GR�}p�����;gq\��*h��OɂC��c7�v�?�94?����
������K� �d����r�T� �2	p��O��P�w����^b��kd�]M�:��Y���kC���,��W���vd�g�Fʑ �3���PXr����2G��j�Ws�
�04AhXRSS�10_��q���n�HYgs���l��{@���EKP������ Ԍ��U{yCH��^^);H�H���w�C�p�J�r�W �l1��3nRG #H�fڤ�
����<�R��?��SO?����'��?��#�7.A�Y4�#'g߹�ܵ5�4�Dr�'�	F�kڤd�[����y��%��>�Ȭ%Q��)7��!�g2Ύ��Q����l?Y�p�H��!'�R�8�:6���&9�
,����R�D�?GƷ��y4�'�����̿��Qx돩��gx=T��#�C�4z�s�2t������\R��3;��W�)�D���� );������N��,>5�	����g���=<��F�z�زQfӑN	�& �R���G�<�G��DC
){yᆀ�5��Z��yأ)�N���ER�N�W_R֐!��|�G���)�I�8
5qKl#х�ij�g_�m�.�ïd���Ւ�`p!,^�H@��ZD})�v��"��wuR+�sAd�#)��iM߱��с�7��d���Z|�J�|�IyS�Q �3���vl��s��L�JYU�)}��;Ae���/&CV�v���;��*����5T e�.¸����H�Uj"��ysԢU�,��r0S��.v�|��%���I1�#&��s��
t�#-O,4�������6����\��@g��o�)GxS�	Qbh]�Tv��O�z���?G��ؼ^j��C�#��1B�LL"���Q(|o��ǡ[P�)1�� ey�(x�K��/,��=�<M�O[�  �uk��7�<P��p
Y�RvH8]�q7� �4��@�1F	 ���R=V��R�@���f�սRnm�C��!�8R�.a����)oL�}���%2�4����]��� ��؀ )�����.�#���|Uf�C.b�zGQ��=�"��eoji��M�H�g8�2��8�	өH� ǃ:Iۺ�	�#ERVT eT4N�0��@�&�$�@8,�¯ӡg� %�3ER>c��%�ɏ��R��]�
H���W�'Ǿݔy�7�m�* LP�zOс�W�Q��=�aM;�J���ۣ)����b{���O�$\�c�~RvVVH�.�t���At끦~R����py�F���$q�4@�	:p �8�r���H9A���r�Q�@���݀ )+������kQw܁!2 �(��hM�/����N�o�� �#Я�����@/��@�Nw������y�`?27�NkY|t ��I��0���o�	읧���B��O�^(�!��X,�{�դ5��x%��(Õ8�k�T��v��K=}5.|O�]���e��~�^^`�{F}P�Ї��`!d\p���\5����H�-@��F�����26���:�������Z���@U�=I��|��f_.c�J|v;Y�M$�������w8�e� t��3�&�D9,�J���GX�'K;�����O�v&��@����I�'�!'WZA[W|J��c�a��_!��8{�����d5����:��3���q@ʾn@��H e^�TPрx%�sOPI�Ge��G�:�A`���i�,�O9�#������Z�2u����w���W���ƿ�c�����E�[�_���O�,ؤN�s��q�$E!���I����5x���x0�l�3�2V�)�hq��
��	���OA����k��2Yx�C�`��P7�����P��?� �h����������X͢�W����L�K� ƒ����YP�6�+RB�5կ@�@1�8�B�}�5J:q2�w���.�{b��qV?TO�9���ؼ�����`�-�u�1��dmqP��g!0vN�^�Nv]�YmZ� 5b_|jq���B�q���@���#�m!wU��/�w8��#	�[;��z�iվ�����XW`�����a>�:�1�Һb��� q��S�R�ME���������_۱ucx�a��^���;*^� ��H�}y!�9�{{�y�q}x�'`��]��\�&���ӎH탁P_ￍGbG��3��d]Î`�Im�1s���	�x��8�T�j�l�k"O�@�W e������*��*#��(����W�An��g�.���o���b�ٌ�u�O�aP��
�cH�0Ew��U�.j��a���}_2�)�،��.R|x׆0 ����9��qH��cHY�g�v��]�����b���pAЇ��̋/A�m�V�x�d}��U�c�X\*spc;6}��I1���:m�����4n�q�a�7/["�硧�XQ:Z���eL�����2j��Xaҫ浗B	a,�'�&�rp6u���p�����UY!v��>#C&����D���ʯu�/X�����k1Ҍq�XF��I e�+9f�v�[D�\��������F�*v���n,lI��+��$(�{�5A~+��N2�"\,��@�h��QHl��`��W��E<S����扎�@���m@^�G��}�w(������*�;�� }z��qa�;)۝?��d��}���@�3g�TQ�� ���_u|�B�20���R��)�n�/�z����P�ƃ� �Ð�}߮�5���f}�q�8�{���)3�LÆ�u�i�Ք���o��!���PS"���E!{+ �Rw�:���
 ?H� MT�2Ln����?�Ԏ�����`�%��%#�=`���;@�'�=)��HY��$�� ɓ���ZN�&`��@��'�D%?��d����g�~�{�LE�R3AT�<���*�*�%�F�4��Q٣�W��
��9�2�;�k���v��B�a�N�Q�� \g�#���36���J�>^HY�H9x�^b[�>:.�B���p�<����N��b��%�J��2��Q��
��d#F"��3��bA�`&�,)i�@��q�e��1�44����4��Hdj�!ȹ�Z���辳�@�& )_u�����ѵ��6�0
��Z*�(:Hٶm3�G��j��'_kK����%�4$�!!����xmJ��O�4!�W�k8޸D��PiO>D%?�������6}��Z>Q��?��ζp�=wҨ??M��XƎ- ̖�9/��w�`؞�@�N )7�/(��6�X'��|@R>�|������*#�� �����Ծ�s���m�(qv�Κ*���t�3t��\P/�z���`0C���M�m��m�v���)	; �G��	����x-$���<��R^-3��3�3��1z}'E
Dh����/� ����U�u��*�2�nGY6ﺛ��F)ZY,���*��M�� �B�X�y�ly?�����K\c7�]�(c��� �m��'�� u��;����������`xW���XW��O�9�����*����>xH��L�wl����_(��1��y�1��|�8�D�Ps������C�A�{�"�+ƀ�;�"�é�.p!{%l������Y��i�au�V5����!�,�]�_~h)+�@�1F	 ��~R�h���S�@�z��1fk�{��;4�!o۹�s��NQ��k�<����k$?�[ e��"ŝq�E�Ɔ����S�H��ST �U�d�\N���2����>H�s_��p+5/YH	:6�
��_nf�����)#Wd4I�:�V��)�����	HY+0M8 �T2BRP_҄mL�X�����R�jݼQ���	\j�k/���	�=�2��@ʬ�����m���T�NP�������W1i.oߨ@��~�=��Ӎh�NGR�����>|wOsׂ    IEND�B`�PK
     ��Z���  �  /   images/7260fbed-8271-43c5-b1e8-f8e9900a221b.png�PNG

   IHDR  �      ��֗   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD ���̿   tIME�6���_  �IDATx��ܱM�P E�g+�^ �3K�Q�53�`�`��HP�q�o���ra��FI�                                                                                       ��T&X�&g���gg,(�6?�^[S�_m�< y@����$H�< y@��A����$H�< y@������$H�< y@����$H$H�< y@����$H�< y@� y@����$H�< y@��Ƀ���$H�< y@����$�$H�< y@����$H�<H� y@����$H�< y@��Ƀ���$H�< y@����$�$H�< y@����$H�<H�< y@����$H�< y@��A����$H�< y@������$H�< y@����$H$H�< y@����$H�< y��	@����$H�< y@������$H�< y@����$H$H�< y@����$H�< y�< y@����$H�< y@��Ƀ���$H�< y@����$�$H�< y@����$H�<H�< y@����$H�< y@� y����$H�< y@����$�$H�< y@����$H�<H�< y@����$H�< y@� y@����$H�< y@������$H�< y@����$H$H�< y@����$H�< y�< y@����$H�< y@��A�& ��$H�< y@����$H$H�< y@����$H�< y�< y@����$H�< y@��A����$H�< y@��������k6���&�^�}gg����ߋ��[۴�Z�uϯ���a�˛ $H�< y@����$H�< y�< y@��i�>�.�i�pN2                                     ��*��s����%��Ȼ�'w��������H$H�< y@����$H�< y�< y@�䁉[�ԇ bv&                                       8����νzȋ�������=�`�	@����$H�< y@������$H�<0��[�0xC                                                                                                                                          ���+b��0   %tEXtdate:create 2023-04-18T17:15:54+00:00SMK�   %tEXtdate:modify 2023-04-18T17:15:54+00:00"�=    IEND�B`�PK
     ��Z�wp�&
  &
  /   images/e3aa425b-adcd-4ef1-9309-97e806748a2c.png�PNG

   IHDR  �      ��֗   gAMA  ���a   	pHYs  �  ��+   %tEXtdate:create 2023-04-18T17:15:54+00:00SMK�   %tEXtdate:modify 2023-04-18T17:15:54+00:00"�=  	fIDATx���!�Va���1�l�tW�&l&�f�=�Y��`uF NW܁#8�~��2s��<�N}�KߝB$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�/8�{����a�$_�~^t�a^;'yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yHYN����qr�݋y>���y��r9�WC�ݫa?+����C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C�r���-��.����`�<�!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�L��<�i���l�6�8�n������f��5IR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR����? bw.g�����9���<pM���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�H~���p���u��$���y:���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E��8�w�q·H~����-$yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)���C��!E�"yH�<�HR$)�#=Ng    IEND�B`�PK
     ��Zpg��>� >� /   images/1c06f444-5387-4cb2-91f2-17a999ad4bd8.png�PNG

   IHDR  �  �   ��ߊ   sRGB ���    IDATx^�}��U��s�v����d��@(��(]E��UAP�����]���޻�늲� HDB @�E���$��6�d�������{�o�fi��9Ǜ�s����s���W@?4��F@#���1?=�WF�VY����;4��F`�"�	}쮝�F@#���q��Bq@T.M�c|3��k4��F�Є���F@#��h���_a��y�r=�1�����eӃE4��"��ևM����{�����h^c����ږ[�[#��h�+c�����yi4��F�!�	���߭�h4��M���Ai4��F�!�	���߭�t8��@U_s�!�	}�-��Jg����'���O���iB�����h4B@����F�U#�5�W�~�!G@�!�\�P#��h4M�S}�q������"�)h&��'؂��j4���D@��\W=+��F@#��`hB�`����h4��Q'��7�}���gup�ߗ������D`�	}b®g��h4���&�W��V%^-R�}��F@#0
hB��-5	-O���sM4��&�����F@#�j�J�>#�	}���h4��Ⴠ&��g-�HF��q1�p��k4�M�p};��F@#p�Ц�C�����,�&��
�:��F@#�E4��"���/�����T��F@#0AЄ>A^O[#��h��K�Z_�I�F#��hF��%�Q����F@#p8"�e��qU���
����J�qj4��F�/ �	]o��F@#�8l�� �})4��;v����F@#�8lЄ~�,��F@#��h�M������F@#��h4�6Kq��#���N��F�P!�	�P!���h4����&����A@[��*���F@�>��&�} MD#��h*��*�����F@#�84hB?48�h4��F�"�	��«/>����q��zB��&��z��F@#0�Є>��_O^#��L4Ư�M�D��z���C@79`P� 4� �%4��F@#0�hB����h4��@@� Q_B#��h4���&��^}��F@#�� 4��#�:f���h4����&����F`�"0~3~���iM$4�O���s=0hR;08�h4M�N}1��F@#p���Aw�_Z��_C=��F@#��@����F`"!���q�ښ�����i4��DB@�DZm=W��F@#��hB�K�'��h4�
�Wp�hBW�='�zcq���5��M�ߚ�i4��F�5#�	�5C�?��h4�;���	�pߕz|��D`���X���b/!t�td|,���F@#��L,��>��[�V#��h�)������ii4���"06]���u���4��(#�]��� ���_��Ǧ�r�a����h�}�#p�cZC��ˮ'��h4�M��mE�|4��F`B"�	}B.���h#��������&��zF��F��B@K��d=4���M4�	��&�	�ԇ�D���}�-��F@#���?��?��4�-�뭠8lЄ~�,��F@#��h�M������F@#��h4�6K1��a��5
��}�en_y_iBe��;4��F@#p�#�	��_"=@��F@#���2����畑���h4��("0~	}Aշ�h4���F@��F\�O#��h4M�T}I��F@#��j&(�k���h�~��,��j���%��tz��F@#�F@����F@#pPЖ����^T���[�M#�x-hFx-h��Np4�O�����hZ ;`P�˅4��j�3c]�y�,��F@#��hB�O ��5��F@#p8 �	�pX=��D@[?���!�k4����Փ�h4����&���d�Z+'����x������A@���U_U#��h4�M��w3)��ƶm��=	�A�u~�. MA�R�m� ��D���/Z��P�#e��a}&�cp�ǜ9�0B����&2�݃�f- e(�0D�\� ��C�:	� ��ń%��)� ̥y��)S�{H �C׍~6�z�F�͖@6k�Yy�,��ay�Q�͒��,�A�/m��2�t�@:��NX.��� a�LӄQ�P ���Y5O1(�%�2̲IY�@�,*�g�R$$�t���	�8A*�EB�K��dRJ�2��0 H�����?���_�>�85T|~K� �0MA��mt�0dK�&@�bQY�
��SLX���K�������}�B�Ǳ����5�M��e%�<��w[t�݋����J�/E�����R��ZA���3<?�1`�i�2C)�v��>/L�&�!!/L���� xB��0�~���2LH�ЭԹe�9���0��D�ЀDH�0!`H#�!$Q���

i2�S��HL��m��2�öJ�.�� �	�D�O���iX~R��=�
�eE�Y^%��зׇx��RB���0߶���؞c�eXF 	;aKC؆�x�0-_X�A�Iv��)HB�ZA@�J�$�_��G�)�iӶ}a� �a)��-K��!�0�B"�E2�A��K���)La���P�
� ��@RTL�,Z��C�z�^(J	X�D`@�R
W	k2�!�N�R�f	B��0B�4BiX��O%��e�!���!m	�J��(��Mؖ�I�	� RJxp�ae�T�$tTH�04� �Ah�$�H�����AF���u�T�J)D9�ŕ�+��{�Ns�HT*�w�8}�ޭ��=r9��N����
La'�aقd%�5u�D9�-I4gClK8�����6hH�����cȰW��Ԕ�ԓK��/�`ME?4���po3B1�!̅�,�<Bb&L�"�M��<F`���rX���0M��	�R�[)��z@P�����C� ��. ���$��o�^z�����°`��M[�S���D �H}u�F�Z�e�lu/��B�џ�I���+��� $ B ���tUK<'�݋��4aZ�^�;ۈ8��E���?�dBs��O��< ���4iC�ώ��׍>�x�����C�5�}��j�у e�4{	���!���M�d `|���j$,��ş�)���"�^*0� v�@¦{�jl4����,��<I�!|}xn�o��,<~�|AXF(󀙇@	�_�K��D�2���!�t/�CJli"�&�xD°B~���!�"@�τ��O"��T{��L�� C!B�y��Cҳ�a��	a��$�Z���քiG���p��$�=c�>�4���&��E� ~���ӫf�Ϳ�һ �����+݊XÈd�������EHD6����Y��F�B�j�
�o���3&�����B�χ�"��ot`�y�A+"ҍ��%16�CHσG?�2HI&�2"�T�ϗ�C�?+rf�^��L��/C��%˄A<Dω԰���AS�- �2i i�P,^���u��[��0��D�Hѿ�+�{���$�:3V���WkB8�4h)�o�)㴖��T�D4�"$k~V<�>
2!����A��!� �<~ S�aY�a��0� �!%Ym��[̓+"$eۧ�"��d�`I$$Y �$#��$���A[2�T؆����3�l��BI�3C��B�wiH�IX�0
ad1#4�gqTJQ)U,!`		[J؆M)#)JBچM#��2�p-4�Pt}�� �
�,)��=�HY͵V����[�*��+䤩_�,<��!���g4��3t����6/���'{ׯ}��ߛ�=��� ����e�RtܦGD!�D��%����<DHtPyJ�Y��YJi�k�W�C���+�L$�G��X�����HS���)�_?V?��C���i2tO/��� �D�6Q)�JGg;>�+"X,(���FL�F�c<)�����$;7��L�D�d7LX��t:�D6�lM�R����>�����6Mئ�8(!�݄ �IAg�f��̖F�@㏯'�@��a7��CWU��XyF��}���b;f�rPa��lbK�}(����X'z/�S|_NbB'��$p�Q��kxi@��~���Jh��R��H-� �K��H����"�]���s@
<���XI�
eTQ�chDB'��p�y��ɫd��=or!���0J(��Ul���LYv�������>��αg�i��*z&���&��@�0��\}Âm�n���U������u}6,��"&d�e��l&� .�HBg�=&X"�����N�d���D�D�t𪃔^�Wm��C���_a:������1�(r�$cS=�|��I�]�Wc/]-:�I�VG�2�����eYC���� B�,x�l����b  ��Jں͍�* �u�q[61��܁".����D�#�"����r�E`FȂY(huX'~Wl�g�,�3$��e�f�8#п�tb�eو1R��у��da�L�q��#d��F�|"��ei�t	�R �V3b�0vD�
��-Jh�����D����zL���1��s��r�Ƽ�����=�{��b8�	�,��PL�d�G�v�k$X�"�Ȱ�7C8�M���X�s��>�Ü9�����8̎=�1��&�1�`c��k�����c���<)k�#0B
�&RP�B�Cg�H%7�:�F:�I��0��С�\D�)`]�F�NΘ�c��9���.6�2�d���N�%k�U;�	<Ҿ�9Y������\i\�}�ͩ��b��PB�!2��"Zz����L9]�#9R��tΏh̑FǶe�XRH9:�xM&8�Q����d�h���@��OL@�$q��E��?!E!���^�������ڇ�|���Y�"k �Pp4�B�A�^�{Ci�B	�"��#�0G{ ��c�OzH�pĂ�޿�|�B��;�� ��weh��=jq���+��9�o
k�a��i�l *�Y(% gJZ�;����L��%�Xxa���n9�o}͉��&��{�)��=t�Q[���;n]yL[� &��^�A��|ȇ��̙�I_�����$��(r*Ҕc,}�HGu+-F�(�:��(��2��A� �3��lz&Z��aKY���]�]�F�8�+���,r�2I�Vj��SՋb���O�`hף1�k����Gf\��bOz�Ͳ�BD�ba��PԅYCfD͍Ɍ�Ou][����)]�4B��Y�V�Yh�6	:�f �,�P���'�u�ˎ4-3Ҽ#���r�O.GY5T���8Pt9�ɴOZ�	V/���'�f�Q�l�����uCS�ZB�d2�&��[aS>�R�!V?^��_�^-��L�#��iL�QhB|���1�{�/���D�ݣ5M0C�Y��v0c:�-=rޒ�k�x��_n��u���A@��Ai���i�fѶn�d�n?ur� ���U<�"P�G&]:����g��^e���;>_z�*��i�4�$�Y���r��M+E�`i�*ZJ��="�H�e_������ql&J��׫�9F��}@�B>�H`p+*��dQ(K�nK~m
�I�11VQ�pYl����A�ie�\�4����w��8P�(m�#���b萢aG�c&�J��JwXk�y���>2QG�%y �&�S�u��a�{Dpѕ,$x_��E���,:��=�C i�4,R�%3=ŵEB�J�'�V�]��C�$�D���N%Ll"��ESM�,�������^�?�MC��H�!�u���>`A��z�^J(�pi`	�f �Z���N ��b���K.XrA��u5zj�a������cy�&j��7�xI��+Om��G#:W"�.�+�8Szd�M�*�+"���m-��ǚzd&�H(�bTX3%�DPV�A��b�fK@�{ �%m\��"?�ӣ�36�F�J��0�4�ؼL2	>��
���T �lx��`��fz�
��֬� �x���p#��p�V��%D�G�[�DIJPry��o�MN\Gc�)s�H��R<��h釃U<�ܨ��"�j�SAaJ !��A8ȌL��þ�a,����@��H ݐ|�#F�jȄN��(�D�|�Dɠ0t�tL�$���(��a�r��@�V|��H����-Up��5�9�+b��޾���{��
Tn%�?�e�~�o	����ux|�Ā�joD����F�����}A�>p��98�@K4���r�ń�
w�x�Ov��㔖�~ԅRe.���
��`%>��C��v3T��:a_�$�D�'����	�|'ϴag2�^.�" ��G*��HeJ�b"b���8�^��k�l�Lض��ɌN�l�6@d�uC�aJ���%"1�:d��40�t�NN�7��(补���n�&��3	(��!R� �d�vPI�^ցL;�SI&JT*%Xn�T ��-Ec G�H�f��	�Ķ��W��(6�H���rc� 0v'�~쪵�S�&٣y�(�:
��nr�T$iJLD�4T�B�J��0��D�F2aA>L
*.�
��(������o�k`E� XpP�����6���F�Y�.%ƒȣ\C>t"��D'����p��aMi@벣�m�ܲ��^Pw��:t��	|��n��&���<6������n��G�w�<e�� r��:GKC�gQ�5�)M�	��Q�rU�p��K��oI�#��)z�>�J�nh��҂|2���@�H�g5>DҢ�/�4��=���Tu��*�-�B!nv9���I�$헎b+���L�Қ+%� �Q)"�{��-�����`z!��5�(��5n+24��7� �欔�ᯘ�Ţ~gm�,��
�71l�De�Ơ)64�jm���7e�<(��0���2�b�`9��%��A�d�XHR@";����1q����A��hEK��:�����y�UGYoq�k���i�l�p�H��M�jmEʹ)������rمW(����� ��E"_��/���,�q+�h}X4P�r�Y��z<��%x�6 �JDJX��멚�i/�T�@�gJ2@�	�f6�������ֶ�[��������0�V��KЄ�7��^�w�o�y����� 72q�QAq���I�#ܢ2C��F�4���a���ī_�4^�2�
�<�5�͟����M�66!��!3�	�l~��$�%���B�QEW e9�-*�
����U@>j�`�����Npŵд1���X����ݍ���!S(�ȣ��� A��(Z3E[��=7Q��]F)Vʤ=��/2S[&ʤ�Q�WmܺzȖ�/8����Q�#�1P�}������ϣs�F����9�G��!S���#P�"k~D��${�&����Ji��c��h{�3
�����-i��B�&��d�ysмd	�σ3c��dr@2�F18 ��B���[�"�e+
/lF��m����)�QGV"*�C�NT1��:9���ڞcg	�}�Ui�@��j+ǒD�x\�&�Me%�P�#Y�B�c��\(��@��i�9hm����X|�5o8�~}i�M����8��\q�1�����Ε+O��?����Y�Tb�'���:���,����^��/}i/Z<��5w�0@��Ӧ�u�q��>��X�P�;%Ȧ����
����ډ��~8�ɤ�VJ(�\8&�L�L$&�TǲQ�؀dk+@DI>��zz�����o�}O=�\��c'좏t �"�r����"��9�ʑ�
�Eߴj]> ���!�P��`���E1���H->��r5��T`G�
((0�v#��z�x�	���|    IDAT���S6oC����<r5����?�����M����Uթ��v�����8-8ցR��9�Z:I�@M�̩p�Cݲ�h:�8`r;���h8*L%�)"��	����@WJ6��sxa�(l؈�|�e�|	� ʢ�i�j\<����Q����=R�F������R�/Iͫ��M��%Sp\D!i�a�L��φ__�����#�~��͚��ɑ:j�Є>j�>7�+}���^�����Z��ۇ:W�by�����C�W���ټ�_Gɿd�&G>S��J9�4գ����),>��8�w�M*�\ ���p�ytl݆��3�<�4֯]���Q��rU�"W^+q�S*�ᠺ��!]���%G�SNƜs��q���3>�gV݅���s��؁i0���E�H�D��IQ�M��Ū��U�T���Ճ�����A�Lb�t�6j������� �ZTy'�����P��S�S.N�t.���,��$�������W�ぇa�؅��X}�o�!�L>鈈h<AD�,�� ����x��dW88��0�I�/��ނ��Eo6�����-[�o{0w��F~έ�^��\B�/�����J8��K��e ���U���7���є/!����"�!����� Qu���l��$�!�����(]�1���\T�	���{[�t�=��X "-�����B 7g
���A����6��p��6����>���XD@�X\�<fy���+n����\vs� re
2�2���D��0�Nr*|���ԁ��!8�٩���B'{s��rBuE�p-�"��[���!��۶@,:
���1m���.�f��x����m�v�޹/�����x��D���g�Nf�$N�ȔZ*�8ݭBW��ٳgc��v����s�X��3ؾf-�e3XZ[����z>��7 [񹤩���E��!~1�Zܐ�N��L�����G�@�p0�c�(T�⠷���hmäe�ㄷ�X0H���ۃG�<�'֬Coo��(P�j�X* W�CsC=�?j)�\0��L�U�c�}���C��>d:��("�q��O�} ���44/����-e8�<�w����&P��{�:��0s�ؙJ�8k*���[0����)m@�A�PƋ[��\�mچ��.��"�R!�����4աeZ�,:G͟�TyO_{�����ص�
��Z�'గE�G��|ھT�\}/�z�A�!/�}.����R�@�3o�(�2��еb!���̨�TJ��A0��0�أ�I�TXfCqѱ5�������6�.�	}���^�+�e����Xw�5�6�D��#�U��4�(O(���\�m����[TU�}ɝ���1����Qkp*�9����x�T�ݝ=�}ڙH74��6`��mشi:wv�ܧ�j�$2�,ZZ'c��E8b�<4761��eaW�N���?b��gѱc�j�░˥���pu�ΎN$*���6�cy}-�yĶH��PQ��A,&�7*U��R���+��֮tqN�B����nG}e,'�߃�P�m594��v���&��/q�w������c��y�:u*��1yr�4G���vc��l޼;�u�2$�Ι���;
'Noǎի��-���oNg�B�5G20��A�m��E1{�m)RI�L�#��Q%4�JN�B���[&a�_����z3�֌�����3�?���6#�ʢ�e2����f`粐a ����]����X��y䅋���{�)8k�\�Z}��u껻���Fr�VYY�$�JD���r����3*CT����������JikAL�Q6W��v:�`F�����VkR=�]LnB��u����տ����8������q�Yy�m���~���~�Ά�L�Clw尩�6xL���)��T�L�3}����od�7��.��_�5���b�m��^@o:��b;{{���JE��YK$k�p��o�	ǟ��ӧa��9�k�WMV�򳤁ww����������O>�'��'$�Tt�G2�ww�lS-���aY&���k�N�ݐI�"���wK�S��ú�S�5�\dE��ӓ+Յ�B9e�A)�FW��������A`��|~#����r�*��p�;ޅ%G/Ŵi�P���&*��r�:��Q�_�P@Wg7z�>�}������\�G86���bj�Em� ���=$�����p�8D�P8V;R+�:�<�0�U�{�oP#t	���������w������c���u�x��GQ���򓖣}�4��7(a���)*���K��J���öΝxfó���Zl~�q̮����F�<�����R��.�ip(8��h5Cp�%�N�j�s�Z'�ޏ�9q}�/=���S1��g�~�k���^'B7��иt�ڀ�ں��ғ/���ik��L�ihB-����տ_P���o���ڷN�.��r�UxĠ�[�F�jQ��"eXCI�q��7hƟU�����M��%&��qGbs&�_>�g�yWR��+����"J�
�Ϝ�?�8���;k.�0� >z��&TXepp�d���D�^���;;p�e��+��_�&������aVB`YS=�� D��iW2��䈖�Ƨ4t2��=̩��;j��\�*�␖�I���N	6�>v���Om����������6n��#��C�G�[t$r�ZvP�Z2�s�4��'��`��䓏���^�'�غ��)�Ј)a�T_?D>�d(��u���܉,v2+�IL|��?.沇�%���{߰П�1�Ԉ�g������{6��<~p鯰n�z,;�D�}�YX��H���W\�\���9�1)U<"�t.�b����[��+q�M7�!����ƢlG�6�{�)az�6P�CL����lB��I�욪�|g�0P��0M5h>j0���ċ��'}h���z�at,行A4���E;�C�nk=�^���������	ݐ�i���e8���m�r�q�HB������ԃ�~Se4a�B�E߇5}K�`C���o[������@$�D>?��9��B�p���d2<��ȩ��T,����/O9	n�J�:Յ�l[�nŵW_�[n�	�E.%睷X6��86�2��H�JT&k�	�4t�-��j��w�_Z�����	�p���	�����O@Ξ���׮�}�2�����2u*ѡ T=.iS�TZ4E�S�O
�/�gz���!D��-����ꪫ`l������I�%��-�ȓ?](3t ؅Uf��b�3���3�7���|`�7�A��c0���'.C��ݸ�+���{��ރ7��fU{�p2)��W�#B'2'"�g*����P"�H"a�Ky<��}���s�ӘX��b�t�T��*�!��p�_\@G��}K��}'i���
|H7���U:_�(�:6�мd�o���ƲS>4��O�zC�o��,���怼��E�W_��w���ȕ�o�SIN",�����2*a:�@�*���>li�K[L��t蕄��L�rr=J3��B�}���bg/j��Z���o|��8n�2��/Uos�F�I�fn�*������1~���޾nP*ѣ�>��_�l���)�ꄝ/ai��Y-�0�RB��YO�'Q��G�S"B���m\i;q���K�^
>s��b:�M���o}��}.��^���Z�ya+���Ex�E1�q*X2�d*þ�D"����f�����IX�@*�B�r�e�z���U���Ka���,dSh�|$�h.i*��"<D���k�qM��|1����
����F������h|�۰��׬�7�|;�~�;�}��<_*��.ô9}0���z 	�a�	.�mp�5�\A�P�Z)ۂ!|������~lق��
^Wۆvj-۵���IC��{r�p�=�]�0�h�F4���p�Uk脦�5Q�y#5t�v��RZ�E��9�fL���&g��><�C���q��-�П}�7-�������?�~J>D2_�%l��ci�1�SL7Wu���#7�����4'��=;[)�4Y�]J+3)�'���Qt6����۰���� R��0�	�4���/�;��W(�>z�y�	�t�S�جI��o��\�#<&v�?��e��]��~�q<���x��'����0�Xlo�҂鞋dw/r�"t�H���\
���Q�����j��O>^'��d��mX~������o�;�K8��3��|3�8�{�*e�N�ǛMexN���\߅�,G�S5� ��۪"Y��M����-?��Y���z��ԺҤ�s�9r�PG�����=U�[��y�Bo��S'�ԋ?�|�$|�����{Ƽ9�����Z'a�X@Csjkk!=_[I%P(�9k@���j}l�q�^�~��ea���JX�s	��F�<��u�X�8h�F�\@�5�B:Q9V�"G��K�3PM���Q/�����,(D�#D�mO����!B�2hX0��fl��6[����٣nrW�)�1>�>J�>>�/_�����^����V�ў�`�aS[S*mɕ3B�P�UIZ���4����C!b#^�G���1Q��X�i��M�V���/���]`;Y�d�����|��@&�C�@?�t�LFԖ�HO��T)�5'_s�R��2���������}��^��@sm���,f�!��Ed���׫���Z��so��0"ǥ���Pq�ݩ���&L���+�_�+V݅I�g����<���������i"����t:��ю��!WfG]����\x�6P�[Ƕ0�/!e�x���֧��O=��M9,�4�T�H�.G�'�=�[����dȍƱ���F=�IC��6^pL;�MX��������u?�\�	���O���'報��R�D�'Pq]$��
�CT\n�A]Լ��S�|"}!Qѵm.����ܪ՘�8:���� �y�+)N+�dIn�K�bBjq�CE�������KTÿ��!΂�цu�/�'.�`��?~�x9S�<F�Q"�љ������z�Ϋ����;�<uRo5U��}�\�]�Щi��0U����U�BCe1��k�0�2���R�P�Ɩ\
w�ڍGJ�@&�|h���_����o?۷�D*�A��6"O����v�7��U2���0��6@z�3�L�����+.C����8!����Cc���5t
4�
`Q5w����i��P�p!�T~�������p���?Ľ����7���ů���^��I%���)�����q$�0�,w��tB��Ns0QqCX���!�ۉ���Ǹ���T��MMh/�Q;XB#
$� ��UDnV�U�cP��Tzc'L֦w�['5������:���ո��Է�+_�:&Mn�GA��H�6�Ї媘�{ݓ���Ʃ�4��OMw���y������q�5W����̜T_���A^�LY��Q#����	.�D)m�zDMh�-��/�}�8�j2��Z�r!�?����o�T��	��$΁=g
�[ڞ3��za�/|P�Q��A@���7N>K����W��s�]������C7"n"t���(REF(Bgm�J��e�ܼ�P���l
�vv�	x���x��_��_��܌�[:��fQ���;�v�!kelҍ��ߪ�����\��-����������_�
���Hul�1���Jh,���O��Ps"
&��O7G5����^r�-�ٳ������7}����?�ۿ�o?p>�4��|�$t��ɒ[ �K�Z,�8e!p2*�J�.M�2�B�n������ϡ�f^WW�����A4� θ�Y,�F#���k��P��yyA�N�D��x������&\���e��x�y���a��\����AMWxo�Z+>��w,�cC�&\j1�,�T0��.� �t��;p�%?A��k0�\�$ZU��t ��'#0���^#����������ցj�K���T�I4.�LoE���k"��~��qr��i����Gi���y����tߵzy�`�T^; m�|�D�q4;��IS���W�9����V�:\��#�������R�"��ۻ���T4$����M���ܔ6��T7� P�7�K%��,6��U�ƈ�H�O����N$�t쵗^�]O>����q�m��0�Io��8Ց&P�?�W(�R��ԩ�+u��b��9���ѿǕ�����<�~�����},=�D����Q�dNU�j�"H4~��� $,���zp�w��";\ >��[��]|1��6c8�����}����N�Qsd@����Y��jl������4�]�����8���vY�����>��糟Ǜ�x.Lj8�r�S��9_�֧B�4��t<�RB
� "u�KԆ��ɚBF�m��﮸��~2۶��L�yJ�H	r�*ƃ����+qL u����3v������A�
�,)Ä�e��_8�}���k���_��>���П����>���c�]����s����
�����˵��׬��p���
Ñ��56���&
R�Lݨd�RC^�&�r�n<��@������p���Q,�P����$�ԸX��Ը�yl^%�6*0çiD�L����(�e&���n�t��x��[��<���Ke4�+C:Y�kK�0 B���_�j���E���	���e8��On�w��I��_���1s�|���WN�%0Q�׸c��^�b����s(��[(����Զ��׋�~��X��_bz��)�͘�H�t����P�?L謡�]q0c�<�4���.�B���8��	k�v�W_�������p���Hfs�]�;��J���L}�AŦns&R���%���%B��"z�Ʒ����^ܵ�n�	���r��qf�Ĵbu����j�+����Jdu�����bB�6��-꽺v�޶9���X���ڗT������*ˑ��L���IL�ɓϸ��=iB���~!�	}����"��W]���{8e�LYu�"[!����,�����L�����y5ZqMp6��6
���C��,��m�xR� d'�K/�	�OT��-��ҙ$LǄiZ*](8�lH���c�zl�&_8����5������bť����"S}�r�������r�V$B��y
C���L�d�3�BÉ'b��މKn�n��ȵO��~r	�ϝ�l&�I�>�Q�Wj�¾� &��S^.�N��`�gr'��9���RH!8���0;p�/~�+��m4p\m-fT���ua�e��(�-Ƈ�CMG�X����ǩX��.�iȞv
�������M����@����_�/Z
3�F`Rq"�1� +�!���-m������z�9��@8�F*�d�w,���r+~��o���Z�����V�����$h�5)J[T�΂��Z��7"�߾��pd�H���W���Fs��\;D�.���$аhnL�k�O����'���#�	}��`�G@�������}��2y0`B�P):t�I��q�*�}CG����j�J�,���|��
�)l�$pGG֐ɝz�7����N�nd����Q(*��s�ef��D�^�U�jL���Z.�y��	��;���[oŵ��.���Ч�d}e��R�&9�e�Z e��B�um�:7"������ɡ������𳕷��5k1i�||�G�`����湮*�c�� w���9�z�s�3��%�e�R�� Gm`�z��@Pq������Z�.NikEk_/�-�0�&T
�cY��3FQ}~E�QeT&s�بC.��iL�-�)��ܼ�ݹ���/���;g!�<AmC�R%��ھa� �]�3(����b�		54�J���.a	
x(��؊;�ߟ�2
k���k2��yhLd\	&t�%W����4���� ����D��_���j��%�܈��HNrm�AqU&�5��\��7�	}�Oñ= M�c{�����s��+����}��8��!]�/��ۃ�cu&z~��W"t�e��Ǉ��oY(�.��	�I��<����Tc3>��/�M�8N"�r��4Y:�mǾXJU��������e�v�$��%=�}��J���,    IDAT��c%���w0��X��XC����x*(��퐆N��5U@"���4C57�^S���I����3p�}���-[�NƷ��c,9�X�>u�S�udF�1�@����gNU�l�#���@�R�]86�O�ł�З��ǟ��?�)]�h)�1y��[�.=���-���*������j�J,h��}b7}9v)N��|�ܴw>�]�_�f͚�]�|ҸmZ'�S �1�rD%�i�<t}�����h������U������w��������,U��1)���B$(�����A:ZC�lՑ���^�yGj�{�W��WC�H��6�U0�����ܾ�>�ԋZ�V��ȁ6�/�	}/~<uy�O�n���>��	�]��ˇ|�qs�y�Պ�� ��W�S�ب785h�>ѡ��yL��9��ׇǽ�A�I�_�����,pTt(�H�TQڔ�N�R���A=�+eJ�
�GM��\A�4_�d����ͮ��������8�6�i����Q�Tu����!堇�f?*��$�g�T�`��DA��i�����ô��W>��ى�P�k��1N=�LeM���P	[��-���(�:��C���4�O ���P>:5���%U��N�/�������g�����o����\K`
���U4=�E.���l��>�R�%��@��M�Mi���'<�ׅ۞~J��_���N��&1Q2�ǟ&�8�9Y�ɷ�R������#�l9����#��^�R�N<�b.�ܗ��NI�lIi���uHh�z�Qf�ae/����$����A�#6x�{b�J�*Ġ�:���=
���J[��k�n[Zo�t�������qT�q0=zhB=��;�~�x�/��i�������B}23۔�aE��Q�i@ �t*1y��͇ې�9�<�AMճ,~.�W��,t���P_�Oe�3���J����ɏ���DU����*�yC�Z2K���q8hΤr������Jo��LO�N&�|_/���Oq�UW�ڱ���Q�݋閉Z�j�ϔ�ÍR����~��&�ss�A�\��$����Wx�\ƕ|Ot�¿�+���?�)Z�������%�~*��KZ��hICw�����ũ}i�cu*K�I�tY���r]���������{W���Z�	���,&��F�$<(�A�N���{"^�.y,��:k�8����F +֯���;�����t�;9<�f�SR���-
r�ht��Sk��^��.d���5�QVJj�t����\�+��M����i	S�Y�A2`��z��ͦ�=�D�*��j�q�����tO�=g=���N�Q�]�r�<�MB��?��D�M`Ң��ښ������|�E����A%�����9hhB?hЎ���g����'����PC�Y2�rO騇v��Q��䂡��J��DJ>�8]�ηH���s�� �P�` ]��]55�����͚�JX�t)���`֬PV"B�ّ���]�L�DlD
� Sy�~��p�J�fk2}��/�������T�r0?�AC>�:?@�;�Ek�Sι�> �Q`��i��E�W$��8h?�u؞M��5���]]8�mo�������<~����[QX��Em8˄��B����b�0�l����=��&�"^on������1��3h+�X(���4&�}Ԙ�q�YT�(L,Lc�<:%���[�`؝��v�2T�۱!���g�䬳��2�u�f[����S��E>� ��P�N+A�\�,-&YA������,YF�0�{ݳ��G?��+���R'�6��I˄-%��P��i��t�f*���,�"t.�E��B�v���qG�YG��M%S{��F�Hp��0�Dˢ�Z��ܴ�9��5���3�p�+��R�q�ǸE@���y[.��G�V�zôJȄ�Q�����|��T�N�����_��b�n5T,66�*͆������ ��I��kj�C}�x!��7e*v�<tK��g��}�{P
J��A��L��X(U:Gzs��&��K���Y���|ֶc�R�����{_�:�X�00�I���XCOGy窎}LJT!l!�y��5�(�9��@R�>�w,����9��o�S}}p����|'/�����£\|�E:��떣�хT�4EّJB��s�z"B�d��XvlX���#<�r%r�=82��<i`z �Tr�$r1���)��2Vԇ��E	�D5��,ݶ1��%��T��'��'����O�_r�2�[��j����Bk�R�3
�t@&u��b­�p�)UhpO>�|�b�~�O�+��m4�>B0�S�C~��H���T:�ߕ�]�?Uǫ.h����`,�V�r���ɩ�14Y=؀��bB����-Y�bsz'5�M�r҇Z��t��q{���)˚~Lx�.����k�����q�V�Q��A���r�2�S�ё���V'�*�����{�G�YxU�&d��$�Y3��qwO��0u�QX�a#�9���Ũk�U~�"����u
�"B�*jTX���(ŋ���(��)�[U���2�
��N|���A�ڵ�� �e�.+.j��	=��T�U\zU�|=�"�iC�S	��4L�H��su����:����2�����O��?��<w
�}ܠ�Đ�˽*3k��O������{N*�R��mU-�D�11й7��WX񿿄ز���v���`���Ò>ʆ��lT̅ݘ�c�H��� ���w
6������G�a���O��c����G���������(��!i�,l�"+�[���O�\j��r�Y�$
��܅���p�׿��b��j(�ۆ>��u"k
:�-u��PM�����U��h�T�����?�_�;��o��ؔ_zɒ�Z�Z���Z����O\������&�	� ����q�i��_��v�oн�����HU"�"GѨ4�XCg�&R\�]�12H襄N�M���m�%�9����D_&��ң����>� �)Ӱ��c��Nlݴ������w�Õ⼢����p��)_4��1��@A��l��J�R�E���6q�������^܉�Xh̶h�|�>�	� +a(4Gj�fF���iҙi~!k��K�(�ݧr���T���]��
o�T<��oy�;p�EF�������}���2��G�㨀���e¨�|l��#�"ӼD&���W��
�Om���61�f@�MP�W�ӻ�?Q��\.�T<E�da�I7�Pak����X�\5i�20f�`B�aYx�pƻމ7��mhjm*Y[���ȳ`�kB:�SN\L�T8�\�Nz�o��Ͽ ��#�)�2ML}���T��z�Suxe-�"�)� �.ń������@���Q�{%�X�%oQ�����_��2d�ȥ�v�b����ҼA�~�W��EOb�Є>j�>7���r֦__���{�=�u��ZH�ÖJ�F>t�����AL/�Z+k�U�:����&|���	���Hc��9�ɐ�@��KZh;�T����k7݄�~��K��~R+�9��2���O��3τM�\E�}1Q'/���Lp�W����ńΦwӀ�lݸ���<rǝ�^��!0��fr����d�`i^*�9*/��%�h>L��L��O���Ʌs���|�A>���d���Q��C!�x�;�
��<�D
e2�g2��x�>+.5+aڷ`�	���Hf(?DǳO㻟�,���`a���P�51�r��<��ϑ�d� B����CB���&NAw�t&ʩ�<%�E}�M��a�ߴ�57�+�C����:ls�8�}�O;u��0-��0*RC�{�hZt_�%���Q��S���W��H�{������}y��岼�����I�!��*,3���&q���㩎l��Q�Z�R�ʶ�>���ntrƵ�_��^����<5"�K.����mkƎ�ڭ��K?2������9�H�"�����1��{������w�����J�J�\�>۪���6L�4
����J�Q.*�JĠL��T�
+x�@�
U�F&0ݎ��g���SO���Otuc��'c��%x졇�����Q|�_?�D2�|��]p�S��r�8u���ר@=��(E����v��UW\���۶�k�&Li��&�+�����?6��D��\���H_�X�@D$H%sÀ��a ��t!��L��v��XHd���D}�8��y���2s�u�\/�4�	���Dx\ߝ�M�J�H���Ѓ!�z~=~�ӟ�_]�fWb�e`��h$ZͶ��ܨ�*��UI���az$���b��*͝<�cӻ�i�.o���:�$� w��$���t	�;�L�1��& ���i�59V��/#BW�	�U/��C�9�4P�݁�n�?�җP�����<;�J�w�";i��(VZ�"t��6��9�Q�$�}
����7�
����P�]��&bW�s�=ae�L�y��d6��&lͥ��G-��#?��௶��C@�[�MW���.��{[V�8��`F.�N�80 �8HIu���9�d���젮j�2��ǁVQ�2�$�L�Q�L"a	�p�Ȅ+Lt
�Y�?��~=>}��g��<�8�5M�p��g���I}�2�E#-�
Ȕ]B�˽r7/�R��h�T]β�J|�+��
��fT��ѳ�E$h0װ1˲�"%�tU�S^����{�����C����C�qT�4����z<��	ltl
4L��iG.�_��`�2����ģ�)T�F�r���ي��p����?��ڲ�,�N���\��Rp�r��eI����n� =`K�4M���{���Ջ� �������`�m��dɲr��P%U|���'����sλ�J�)Y*���*���;q�}������V�>����V|���i%S�J5LP5I0�{(E!<�me=$=�- /+䵋�=tF�E�\���+q��6�2 �N�闱\���v�!�۶b�UW����ob��3���*5tJ�2z�F�*�	%���<Q$�KǹÇ���K|�cCg��8�s��:��F�l�'��G�z�h��V�\�q�[&����w-����w���LN��=��WB@��g��*(��J�i��/9_���M.y�������˃�h0'2@?��;E�M�����s�'�~�Ko��	)�U��6}z��C��)��e@�\��ލ�'�J��T��������3ž�e�\`�+�A������opǁpF&�xT����:<�+��o{��p����i�&y����V:o����R�4��Z�&n��6��?|w��ǲ�v��o/ʽH=t���H1`8�IQ?���?[ҥ��**���T�:�z��.�gTZs�p���(���8�+^�z����"κ���F�X��\/==z�6�.�ٓ��<��ַ��}~��n�qz��9 3I��ݥ)*&�m�gȽi9���MKS�q�a�Sz���"�b<t'Eh���{AUB�O�1n7�5��������x��*�Nߊ�\�[����0eAÀ�
�j���m~v��W��/��;��>�m� �]sI��N�a���=���+n5HKDF@W��,�z,��P����X��iC�4lÞ�.�
���a���k�����=;����]���w�q�{��YR���;Uo魯���4�ⅻ���>{��������_�����c�W�\ֳՅ���-_R����WtmQ��]n7��Ҋ3W���z.��_u4_ ��c;�f�������H�󑤮x�ʹ+M;�g�q�՗�5�zv���gףZ-Kʀ��\C�lH���y�q����o}?��N�ڽ[�u�����VPmw���n�����4E��8�(1�KE�ІX�d��li���I(T]��H�P�QYr�����B���T/�! ��6፿�+�׿�o0�~#Jr�9p�{��w"-��ۿ�o��������;�\�a&�"U��	Y�'L��;�R��H��� [Z�J*D/�wS����|����q�QO%�RD�v\v�}��qɵ�aj�F��
��
<2⤁N�4
�]Y�S;�������ޗ���>��$��26��t:���C���`�B����e����:��֣K(�P�kd�C�����f��2�_���5t����278�]-�Z	�:�e�F{z��6<X��7��ʠ���
�g ���O�.�/|jǽ���͍�n{�i!�Ʌ8&⩨���j�Ҿ�(:��lh]�n�Wnf� ����d��=��m�Pu=�]�����8����@�^��"����m�z��`btc�c������8f��051.ـ��:�&���{��ȑ#�?g�����I��֑b�c<���q�)(c<�	�������f�k�6ϰ�=z��GOP�z�v�[�4X�T
��˞V��N�`Ùgb�i�cn�l\�	CCC�2��&v�ك�~ ����z�-W0㺨�z�%0U*��v�S��x�G�@�tO ��LH��,�]��J��@�x��7��a�2S_���>V<���n��z=�C�L�׭���9��`t��oނ��I���==���xr�.,�ۏ�S.-`<��|�%��]�-X�����Խ������.Lu�P91���r���9��{�Lm�G�d*w��X���� ��YI yv��=�Ts�Q���9��mڌ�֭w�\�;�o��;O�<��%?@�O ������G?qk��?�vKc��Q#���+:�)�ǆ�UT�\���g�W�Z0��f�	"�ʎaq�nʐ4��A�Ž�vpˆ�e���K�E�l�������mw�xO��k
���ʐK�<`�z �J%�*���HU�Mޥ[�- ��F��̖}1+�gC<�Ch��Ba!���98
�h�ƿ_���m�H}=Ǎ��^7�-L��{���+��0��Q�N��>C�>|�i�E�u�HQ�t�����)�2��k�9���;�ݖ�n�0�R~N���x>�P��RF�Ršv�XfQ>��/ҮC�:��2�Nq�)�3AS^��R	�����xPB�MvC����:	�`FF<sa�S����3���LJ�zږ/�%��ȱ���Ra���v]ǋF� �ډԬ䧼��U=Lo���@c�ƻ�^��K�������� �DF��7��Ϝsχ?vk��;���1�����6�]�:��F$܆�r�w�Óם+�k���Q�D9J�J	[�0���n�<Hw��c�T7���Ĥ�����;�cM2��d�3�����5ϐ�U���L��=_r�%��4Y�	�R"ETO]ъ�i�&�䤔͜O���C6�I��rI�n!���>V®���h p�x=Fդ�a����F�d2�4�Q&�蚓G �ڮ���C@'ӝ$9F��LHed�K)��[��;��G(@#Br�zo��wE((r<tQ����XJ���H�~��%��'ngxz�/���b�Th�t[�,3��E�sQ1�u
{�0�y���0�����N�ܬ���K� E�y�{�g�Ş���̢'�k��}襻��A�9�����J�=��$�lފ#���L����6��_�O=E���6��B��It���>�O|ꖥ�~����G�j��<��O.��0\\�BD�3WȔ��R]B�2�4/^Cφ)͈~�MZ�	CꞃE��SIWX�tHy ��(�FQz�n��(��I���RЅa�qA�~�v$�1��=�=�0�����C��Q�P�#6w�X ��(��
�,����M�0�S���N*���i�X�HX�,�3	}g6"鲜����4+	k,S�87ewC��Uj�E�%oL��¶��ui8HRWec	0����Y�E���	U~.y�D�xDA��>JŒ��ƀS��5@f=wTF���*5����X����e��'1\�s��p)��HC��P2V�}��N�w�f}�æ{ιhL6�MI�� p!]$ M��l�Wz_����O��]��V�$Fs���2�W�K�ݾ麍��$    IDAT�x�R~t�կ~�����o�D���R^�#0 ��C{�/9����{�㟽u�߿f[�֍�4lnC��t���i�ve5�&)`i��)�3�E�F�NY����%�n��:k̻��צ�NA.�C�\�^��0%�����Ǎc�'^[�O��#<G��=E�eh�
�UK=�Ҝ��	_[O^�"�Cy[gf���a��-�E��!����)9cY��n&���N��t�hi�ݎ[��,���&M��=.�
�ٙTEE ��z�ڱ��Ic��9�|��*�=�Ͼz�ŁhܱtL˵$�.���/��H\A�"�)�sY��iQ�>�8�#���[�;ڱޜDL����4�� �Uy�^�<g鍞J�M���T�0/Y�@o���_hF8n2~J����~�B��4�N����X���v�ޑ�}�9��?}���n����������w������-���ug�̫�eZ�خ��Eh6�H���6��x��y�9K���)u�R���Z�y�]&�>����(A.�%j�;:I�yZ�D�#�^Īf�}D,�6�7�ASg�5�w	�R��(�W�M Ƞ֐:o�8Ӳp�Thb��H��˛o��5,�[�j�'@PױUr��:pcӲ� ����u��<������e�(ֻ4*r4a�[)_CsX6�c9@�qPv�k]m�I�Ј�5KT����3 ɳ�/iϴ��4<(W�zZ��NwHPvU�W��EZ�Fc¤�E�]C`��=Mw�V;(�s�){	b`����
ࣧ���+�<�L�͐�ro����r5pm�uc7��Q�W�?�n�H�b��jIr���,�x�ޡ�{�@��'8@?�<vO������-�.����7w#��:�q`Mm��}��))�[r��9-�gr��E��ַ/�Ye֕�4�2!|]��%Diޙe^�g/tɢa`��%U��r9	�6g9{-��0�-��Ex��fr�"Pbj�m	�CKL��9i���u�۴�d�W�eSf�0S��&(mD���n�������\e�ִR5ear붳W�H�����,I���&�r�:�'oY�ֳ��|6��R�n��L/x��a��˳N2�w�@�/�3M���0��QS�Y�׬L4�lݿH��f��U����x��3#�0N�~�ΡR���+�SZب�q[IG>B��M?uɊ��2:�A"R��It���V��0�C�����ڷB��j���� �_�����]0�Y�u�����[W~p�[���Ek�V��3DH�0����	Ӄ*x�Z��YgY���U���Y��2���M$c�@GƦ.����6�g�����%�ܮzMVԆ?XC�$�b-r��VL�Mʢ�_�:O�=�8Ôp�#."04�"wK� E�-G��]�[� ��2^����!�7�X��@+|����:3�qv5ZlEGC��;���'�'Z�|���s�TNU��������D�մCCψаь�7+\��4�`n��S��<=[U`Ku~���9�z���wցs��"��wb���3��v����cQ��(yP��0�n�v��5d>ңV(��dƞ�a�Q��:f�;��Yyp���޸�߾���+;�l0k�� ���~nǏo����w]�%L1�ѐ���E Fs��dV/�KW�k�Iq�gV�2�u9S7�6H�gT��ؽM��x�lb�l���mk���J���7�kkL�na<��Zb
j�'���CՒ4g�q�e��)+��l�n��,1���	j��&�u�pNc!�1��E_��Ld�`^���R��B��<��m_k��E@����(ٶ��aT�����b���U�E�V��`�V'h�Ĉ�X�s���!|�S�;�)9M��!뜠џ���&���HW5�b�،w��Nu����u��z�ROZ��ħS�sK�ؿ��<��s~���9�э�����*_����Unbs���LM:�ӓ�L]{�M��z���h0'2@?��;E�M��Ϝsǟ|����w]���J��D�<I�Nf;�>	�;D��p+j�n��M�����:�7Wh�!$��{�E�k,9i�� o�G���_hb�X�8�.g�ϊ���<?1�<?۹�2��]u��B��W.}�c	+K��up��c2�Sɡ�Yh�Wy�_�~@�A7PcC���������^u{l�<�����c�^�:k��w�?kY����$�%?�tk��>u~&`�;��BR���r���z���t��m�R�p��q��c���M��7��v��O	���_���� P@'?�����o�^ͳ�sYk��w=�R�P#`j�/<˓h�����կ�q���|�)��n����@2���>����?��U�л���� K|���;��TE6�fz�?�����w�E`�ɇ�U��f��7n���G�z�v��AЅV�����z����
���r�1�x��ε���SnB�����D�j%��%�x��$��$t^�4)�^�6�x�0f�F������Cׂ��	�{
z�WOSF�ٺ]<Q)3���Ce9��W5צmV�~4�B���@n��F87�V��)��d�yp�v\�a��Ҭ�Xn9���>���'�Zb����2-B~�tyO�ɏ���顳�,_4|�A�,Q��Q�����1�^�ÆK.�nk��sw�\}͍�?�?�eN���Ex-@>�����C��n��u�]��ڋ1����j���$Y�s�E;���;"ۜ��x|$�"k���|���s�-��3��g7.���?s�R�K��tAUu��HV������~Ɠ�P܀�*�s�z���@���nS�i;S��Ҩ֭׺w��#jh�81!�TY�&�Jb�>Ѭ\J��(���b�s�2Oݸ��P(z��S7��A4�F�N���_/ӕ*�\ą��qM�h�eH��J�oV���6k4B�����@s��:q��
��/�5�4ڣz���*�ky��

�����hE��[������|L��^�ѕhF�q��F(M�a���55����kW\r����?�����^Z#�L���5/ѻM��g���[nY�����%gk[�c �5��)�(z"�\�خ� ���4�j] Ĭ��K�Y�Mxިx��d_E�n˗�e�X@7uƺtkW������v��<^���j����A_�L�����d�h��W��-�"��.�j~�$d�n��F���y�#!W-U�Z���е4>{Y�>���.%�q�?�j�%�a�365���EJڴ����y�ݞGs�6�m/���2?��W˾ȷ�GSCB�3S�B���yf�����eA��q����Xb�T��%߳��%�d<�X��I@��B��R�Cyr.� �	<��;�_�����˼D������\���8�����?p�G�w��NLRԨ� ��������`4tY����U�1Q��BO��B�[��V�K]�D*_�j!�@(�t��&{��@��Dīb^V��"B��[�g
A_��5�#K�
��K��|?�u�t�#�W���%4�],./��
�)]5���i�AǪx���	��Z����ۭu��X<���nCҙ�c"&��r�
����D,#4�����+S
��c8������ǒ�,��>w�JC ٸ��λ/��:�}�R~W�K�ë%|�J�0Qs��g�UMPk�Y��(P����W�ӓwET�5������a�У�9<����.8�ݯ��~ ,�����t#0 ��n�����4e�������@�>y��>LR�=���1QX���j�|��w�2���i�N��;�:K��F��yu�)��l�.��g] -��Z�X� ��n�)z@T�3*j�G^+���/�w�Aa�������1:����4,��dCa2��?�D��My�=o��!�!�0�ȅgX2X1T.�dC�f���b���=�cK��c�~��p��	��)���@w|;5HXާ�Z��]a��S'�z�y�ߵ&n�)�;��+�ךװF��~�Hj��ԥ��1�w�p�>��G�^C��Q��@��=z���v��%�X}J�R��b�A�{",���p�U�ah������{J^x�5���}�YiF`�x��]|O����?����������Ma��XC���&�hp7뗊`R�����_V�ؘ:鱔{q�ϥ�t���qhπ+�=�;��s�ZC�&�-��YW7��={7��,�^@9�	
^�\0�G��a&�v=A]���ӳ�f�w
����I��t(�so�
�����V ��<"`r�k �)hxҡ-��V;Ť�r��eV�����u��F/�%o ��Ĥ���53�l��Q��H�������T-�8�*��^�B����5(��e{"^c��tFZ�/��chb\��--���!���2%��/�%�+TkA:�ԍF=��l�N#���76�ӯ|9��i�Jҝ��^~������g�s���3/:@�<���Nӿ���w|����m?�!�1%ei$�qU���&��C�:�Ũ��}.D1W�c"cV�@3�x>�b+�y�d���4� R�V
QJ��̹l��ּ��8Vx���Kͱ��ZO9�����v�ϙ���j��fk��id�-�Ef�Qc;F�o`�-�v�9�M��� K�a��кޑ9������bE���0W̈́��U8d�E"�k1$e����\lh��J�k�D�m��o,Y�?wn{��M�ס���X!�Q�ȉ0F����Dh�=tY�F�� @�GsM���	�|X6Mq�8A�hơ4g	Ƈ���<<��#C;�.�����{���}�g:G` ��S�)�,�����7?���y��0��ٱ��0�L�^��r���S����'��	ú2fV7Fg��\�XƱ������/`�ń�����U�dJ���Te�⭗������eR��V��9�쳪1��<QL����ym���ZR��z!�ڗ��kȓ���O�[�1�:��4!h{Ӓ���B5�<siEbX�@3�>�xmʦ�A�B�R���I򭭰����ge��H�tT��0~}Wr<N�%^Zc��k��)�ӗ�J��n�A7R��n�H�6��%��hd���=݆:7EˉQ����y�љ���j������w�����_���X5@L��g����?��c_��7�Lqab]��)��#��Ԏ�`N���T�sa^6D�5֡����h� �-����0����l��Y7�PE���#�h���V�o/�����x��_�L|�^�-B�_����jC�(l#Q��Ι���𮀈u)��ټ�=��g�ݿ� �a�l�.��������d���[^���q-�"Yj�𙆾��yzi+�g�%�o7�B~D����g��ȁ�c����ϽYr(���Υ!s�/9��T,���$��C~^�{޾5Kgpv���v������A }d�&���t�F�=�����s��[����z|B#�, �~�N�<��O�H��O�}�/�����o��'�'�;�������]�<O�+Ӕ�Y	��U�q�N/D��E+� �@�k�k�RA�y��y��J�t��6C�I�tj���h�n1|���B��s���jo,��>��E�����Ӓl�ɡ+y/_�mH^���7���:��%Į�ߔ%m��Ⱦ���O���rf�������'s�Ű|�A��C��|�'�q��()��*b��qQ�3{,�=B���̊�|+9�ce빵\���h�ZV���-g�ˌ)M��M")�l�]�1�������RwNR`���:�Dx�����T��8�׎x�$�9c��چ��33��.������w����N&b�I�<�T��, ��:�`��t?���v���~`�?|�U��c�,"���@<uъc�v����0ʕa8��n��f���F�^O�2��{�k2��6u��K��.9G2����O~cU�Z	I����nZo^�EOR�L�� N#��02��څ[~7�i�HU��x�&�7i�j��J���<�{,H�,-�s���\C���YU��b*##��V���\F"+��m�_����ϧߨ��8�F+ƀ�� 6��w�9�A
+"Dr�6��|� ���:����g�D�
�����f���X)�����r+F�-� �	Y�R�g
E���R����6��7`��lT�d9���A�n�`���П����{�^t����;_�����O� �I�0^�K���G����/ݼ��|}$J�F�~�N��w����VZ�J��,�]J�:̙S�4B��*�Er��!�%��ʐ枪�]��l��XЊBP2�2I�Գ0�ED9VHXz']���0�M��Ez���x���e�KFTH�*�ݒ�,H
>��b�����/����c<�5 ]�� ��實�QO>kN�u�Z�-�Ҩ^�!k�G.λ��$�b���7�'��5�rf:� �l�j���R:?,iO�Fd�H��6�Qc0{�biqo�=b��X+j��썡��Q	�+'����MwXl^�XXFɒz~�y^h�*�^���;���]�|g^r� �C�&s�_|�;/�������{j�� �O��xBw�~�S;��������_=��b�TH�B�'�j�sQ�W���CD�+��t��HTD�Ò�zc* "��"Q��NH���r��V!�+�dæf����lӪަz��ؖ�5$���R,[��s߬���t�ܧ�ߩG(��jQ.���P6��L��<P��}�5:����..?���9���?�n��J��V�QS��,nq�4�`��<��L�W&̣���Hd��s�����A�~0σ!y��43�˜�Q�8!�R��e_zVK�Nj�t�J�~R�gd{�K]|>��|2��3�Y��R/�����Q�͎��55c_�G�p���C�PQ�KR�ٴ'��J��o��m�1~�8X���=#_�?���|���ȃ�_�#0 ��� ҿ�����>��?���ڑ��"��+9f�$��nkd���r{�G$¥
�h�u.�yn�?BlKU��[e [�`.�� ]�]��v�."�s�@^C���<ˠ�^�z�yW2�Y.������J�`un|��+����gX��~� |U=[^��C���.��W���-I���ѫ�n�弾Z��nGc�e�4�4bR <�N=9��?�[��sBf�j-��+"�b�Ȇ�9�Z)bFJt�d�{&ԭ�tyǸ�yM���y`����3����Fs,��H �g�'�v�##c�(q#��>�TtR̝��;�ƣ��+�v�^y��r����<X�#p"#0 ��Sd�Ο���?�����wo��&�"$"�R�Ii�j���M�,*�1��A_�̹�tujr�M=�z\�x��n�C�����*p싣
�Zp/ԢK��8Z�0*��x\[�e�as�T$0a��h~(Ы�NO]�����_N.Yc B?��5Za�/p�̣�:޶����:��^S��&�ҳ��F@l�Y�L� ��N'�X����5���g߹��үn��v�䋑���w�V�?'�茔d�B���/
�y�F�-���`��|�WUc���W`�s��RCL73�M��$�e��� �8��ksgn�����b��}��_w�������)���P�1 �j�O��6>�'���?>�ҏ�vCKȝ�C-c�5�y�}���I� nC�\��гr(�PtUMKk��{�0����ST¡��-+�����s��pixh�W��"��[o�� j���m��9�Z;�eޢ	�Z{��5��c+���IJd�`h�1�h����$b]�����[�"�0� �6�c�C�� ���}�虮�j�H��<�8&B� W��_�߶�n�#B63���iL���b��<GіJ�����\1ΎG�2��r��L�*X4<��������"�CS5�����Ўct}`��8k�+hL����7��w�{�[�?������G` �/�\_r������|��������a�����    IDATChg���4�0�Y�7�:#����x�>\C��+�W��&�auۼ� ]!����l^���bk����ƅ:#L�CU�0��T�.ԼNV�.�y�[�4{L=5˔��ZG�/K��ר��yl�9���g�m3��9�(�e�n[���>M�}22�ݿ��f���|�/j����1Є�P�%�odZ�=*��q�9������}yə���s1b;�\�R�u��U�nB;�yE�7`���2����H�c��8��سjx֫�Ǘq+x�E]Cwg�"~9(0í�e������u:����[��3_��wO���<�����^Z#0 ����^�n{����o~��[���jC���C�^Ք~��p������#-Um(^kz�nê����zh��-J�� ��b���p[nU�-e d�q�$�ꐻ-�"�!���(�O�X��j���,�"|��%�#1����-�k�X�O�A��e0�z����kV`g�ae�;�T.�y�:{a��w��# �8���8&��y�3C��3޹�7Jz��(Wt�x��p2��c_^� �J�H��>@����2��:����J""��ܒ2��m5�-9�����%Æ��^�X��;���:U9Y�Qй�*	6v�2��f&��sМ��~ۦ���M[�`5>� �	�ɶ{h��\_����O�����R�$�Y���T�{��3��g��a+HY�]�MxU|��HY�7gY���4����f��a�������}��f���j�z�Í>�0l1W���a.�l ,t�ay[��@v��+Y�¹��zn�^��Oخ%١*��>B��_u�����r�ș;��o��7\o1 LZ���P��$�b<�)7S0u}c X�|Q!��F�
����`˛�h�Z�f�S������D�z���U�%��?�Uϖ�eQ��y,�,q�~�)��q���1�zI���	���r_�c�5�������=���:�f0��g9�x*� =����}�bףWIȝ�=k�]j�3�vzR�-�*W��;��V��v�|������M��L`���4�-!�9�,u��y�����4����@��x�*l��#zܦ�.�fk��k"�_ý�C7�hi
"��9.ah����ZG�HϮ]��f�VlԒ�v�\�̙-b̮=>��9�t4�yy��"�G_�p�t1�l���|���߬�0ϡK 1��Ͱd�,�ʂ6�!�sQ�+��v;^���m)�1Ux 	Û;�v��7SL���-�l��Iyd�n�qf��<�B+Z��N�s�}���X��0�+��F�j�ptt����^���~e ��:�|�� П�Q>�����.��n����ѫ6�	jQ,�S��S֛syO�����i�'`�������d?I��`+��Lm����i1~�j����Hv��ܞזM��550�x ybz-*��D-�F�mQi�a�)�4v�����+�J��/�MpL0���&�+�)B1��г�R!�Wo�.�Q�d*d��,��*��5��o�#[�M��tB�A$�0~�ٟ��:������,��z`/�BOz��Vv��ٶ��r���*4��Ֆ�g�U��(��4�,3�~��9�lVP�+���N��O����7Y����Á �>f���K��ahn
׼���������6\��w���_��$_*�w��� �O��|\^�S�\��?��-ޞǯ\%��FIL�R�XB�$DI>Ԅ�#�V(	�K��+� ׿6Z��5�,ڮ�KՓ�f&�k�&&��*&������������'�:�~`�˓s��/��?�����/R�ٌާ��5�m�s�'Jv�����>�q���eYRn�֟"���hK��5���1�H}��KP>OFK��C���edjjVz��A��v
��ں���<ݡw����b��=�!�R˫�Ҫ�:t�g�O6�k<��XZ�e���0��#&$C�����H������:XNz��L�oy�t;hNN~wӵ7�{��_ܤ��6��Z?�9���?��
z������n�v?v���	���J�,w���
J[\�l�vA75�V��*��L�Ze1lo�Y�5�y8�.�&�.ch�ic�T�Ҫ���}2Ϯ�$�k.6�_�[��L�-�#Q��	�x�Db�ql�ގ����=�=$]R)Ǻ��HU;��\�Ջ��vR_&���M�ت���#�4��8���;���1���g`D!���M䁥}�#aǔ^�z���3��*��&3�
�Z�1gfq�
��yY��������N�Ǥ<��'_� ����9�Mh�\�l��
��0[�	Y4��tR,�!*����oV�u��x������_x�_������ss���|���nv=v���q�˓���?�ELqv��x�+�]�WO�J�j�ՆX�[ߌ���m@W�X�V,#���l������H�$��Ƴ!g�RkeIcyG�~C�D���2�$lU(��濄�ϥ�=�fQ����)�h��i$ja�r�,�֣�W/���,C���V�[�.�� ���R��[��4&R8q���%�C@�c$Q��wn����>�V�/�= w������$=b\d*��֩��o�
�jd𺊤�c����.#�{��И4@JҠ�jPr7�N�&D1����<�Ⳳeg�g&B����lE�����檰���6�������h'�&�8A�����b��n�x�����y��6|�W��̷�ʠ��Y�^�G �K���7���͗~����O\�%u1��W����$��(�]��ԫ�c~�~YN�SH�r%>f�~ư-��WB���4�0+w�ۂl�Q�튬f݅��%א��g%ǐ|�jNqa�kΛMg����x�Ҡ�8����y��O�8h�)�H��S$�
J#FG�c��TB�����e�*eT�v4�m��H��i*#�uV�1�0B��Q��^���Ӄ� ��Z��p�s�a�8���-�]e/@�g�\�]1Ϫ�
�8i_���T�����뚌SAIM8���P#(��.��y&5����}̥���!�bZ���4����q� ,�;Wd������Cρ�t�;�ubk{]��?4�!��A7��u<��)V��3��߂�Agb����^������,G�8� ����)�o��7����������_�)F#� �wY�CP�L���4�S
��yi%TT���0�g�-��\;s���f����ѻ�WK�Q��D����z�*��i��q���1^���,i��I�]T��|�q�I��	'XQլVC0<���8�s3�ز3[7���j%�8���V=|�����qA�ꦓ��̓�]�����[���.5 ��;=>x ���Cgq��"������!��a?@��Br
���a���;O#j���qc-{�T�Ҿ��-��~F!Uu3���g�pչV#�Q"�KAq��'�L|b���;�%mZ��J|yDFH^��Ց�����H�����]��P��1)v�c*��E'�����h�+�/9	js���ބ}a���{��y���w��O�%ep/� ����+v�����v=�ʍa$�S��Kd�	�
hkh݂2˥�D�$/��p��-E������m����(d����VmkJr!��G�����l�GbC��^Ⱥ�����3`�0��s}t�:�F=������m^���B�C+M�a�VTGG125L��a� >��՞v�! ��)���H�V1\S,�����TP*#>MD�S膇�|��#y� I�fI�����������p���H�VP��{!�0D�y�(��B�qQNS�Q�2\	ߧ1����B���q���9h��j�;[/� �@-��D��\, +����A �"�Y�V��d����X`���vȋ����~��ٗ]��sD�@o��s;Iс�%7�#;�q�[ބy���+����>����O���'Ӻ0��� ���̞�+^��.��}��=�_�)ƒ�W!���E�,y&w(���B��=VL�0�U�мƥ{*Ú�3��ϼ���i��v52�x�z��B�2���{eJ�>��-y�,�l�х��Æ4@�:��>zC#ټ��9S;���� (���o��|�T�$���4�Q�'��L'
�\��3
�_⫚�5+��놫B�O7�%t�s��U�n�+�ؕr �׼:�v�tVZ������$�8��)��.t�.�{�(ʽ�58�ЃOc�lP�F�#B�r:��`f߭]�Q}FE�����g�T�����l��+���8FFV	���'G�>��̞�L���\�����j���g6�e�T�	�� 9��6X��`�IQ_?�k��8w>�p�����-�������|I�� �_R�{�]��{����ny�оC����>5F�sGʆ������~������K;�0U����=ۅ�J�Z�LQ���}�#+L#���vWzSR�-��R7Al4��ԗ���M#$̅{."�]8h�.��^����,fN?������06���P��C����z
������I����n�%Q)ic9X6փ�zw!�y�-;�:tC�SO���RU~�T*XYY��9��@ch��^��g#y����xe���1 ��%c�� Ir���~,>�>�����}�Eէ���;(�@9�м�ϱ
B��K�3K�&lh У%��q �pi;��>1�6�&r���7�<}�7^��~�E\�<��k�����1��DQO�F��z�$F#M� Зt=5����Ft�;~h��������{�,G/�(�m��; �s1�/�cPX�����GK��b�t[�P1%L�%��@k�4_`��֋uԫJ�L�i��s����{Ӏ���ʮ����t&j�]�1
l�7�B�2����a�WK%x�o��	� �r�F�����
���5T7l��s���]l�
��@J!v-�#X$�-�)�ͦzudg�_<=䐥c)���[�I� (��^)0ME<4�˨�k��pJ%��y�N��N����Q%&�\�cyT*d:�g��J���r��N�#��W�^Wmv�xB��~~P6�rP�V��zJ��9����X|b/�>���ޅ��#(�	j!Q�S7��aψ���M�����Zw�9�"�SЊ��x�|F
�L���R����@Z�����A9�����<��.�υt΄��
˽Չ1\������/�g����������3}���Ӎ� �������/�������4��P�C��\�8H�&#�@P^c����@����� K�����f� ,|���2ყ*���zqOr���*t|��,#�𦍘=�LLlۊ���s��P'!q�c��G�Ѱ7#�v[<b��V���X���E���x���j������a��N�&!�F�!@?53�v�)ǦA�\���IP�+��P�T��pp}+͖ {m��\�Z�����%T����>22�RF��x��x�R��<=K��>ڽ.*A��Zρ�3:��CG�yj�v>�'��}O���`�Z�Q~���jq��y����0"c�E�\F��QR����[�U3GluEQ�eUT�8�c�\˳.��"��8W���~C@E�L�_�6��A�CO��CwR���LT�Fq���a�VŽ++�nx�+~�5��_�,G�8� ����)�o�����-�C�.>�P�t�3*��ڔQ�\��~J@�!*����Tpǵβ���tl�x۶i��wM�^����%�b�4��K^	���8h ��v�#��Yg�����w�Ś/�4��W��n!L�5�H�1z+�|'� ���l,#�E(�.�A	N�m4�f��y'�MNbˆ�ܻ߇V������b�ڵ�]�Z����G�j�P��P�V���$�W�U�*e�a��=�u��!���lu��t�'�g�ķ{ϣh�:8��3$�h��g�əi��D@�u}LN��1�� ���tՑ:qO"%_ep˞�z��R�1� �8p��;o�!�~�F��za��$ߞ�4�8�>�8EG�]k��KkTC��T�4Ri�"!�Γ� �z��W�{���ɯ�Ͻӄ����k��(�8'�J�`9M�r��렙�����W\��j��wo� ��yb�m��������gnn���K���0�w������ �U��x�Z�K�
3�H���l+�ׅ!�$,��Z�'�S8�:�,'�4E;I�(�X-c���rF֯Cuvʳ뀉)�V��p'I��Ń�w�ҭ���0A)-������ʰ&��}������7�D�y���"@����Q��[��W�)���$6n�(a�V���{�b�֭N�u�8t���2fgg�`8z�D<����Ҟzj��&�ݠ��V�$�����#���0f7lP1�8��Ç0:5���a<u� ��.f���%��2���?\CZ�����_s�0%���@&��yz��k7?��'���#���nc(�0��(��U�J�CH���	��F�"9kB��V��ny���v5��B�������ݵ����[?�7�+I� -��O�9cs���0_.�V��Ӯ���7���H��s�V�p/� �K�a�V�����}�3���ΗoIa�W}H�ˮkR���Ӵ�H^�0��"�NH�>3^y���]���	y��z��d7CsW9N�%��9Z/@�+	)i��c�#��a��af�Y��Ӂ�zL�Ü�V��aH�b,!z�6R�����z!:�:�&�F�^n����
��݋m�6���{c�Caۖ-��M,>���Gp�Ygadl��|�VG ����c��,--in<�25���н�9�$������"LCU��V�G�����8j�#�&&p��Z/U0:5����E;l�<T��;�i�<u�*##R7��k���(��4TUQ!�	�G9`��A�Z<�Rc�:\�,Jth��Fؽ~�{�s��(5��Jⵗ����L�x��g���U"ԉvL�rS����>�Ĕp�qѵ�k�ɭ��6d;�ٮj�Co$)4
HZ��$�X��;^���0�t��r���s����������L�%gi�Hox�����O}���w����1P��P�wNQYt�@_��1����e��R
����&���X�E�4���!�Ů��� X���q=6]t>�.>�<�uv������	M�l�!�bQ[#P{q*%}I����2ʮ#��2T��j��a<�����1Z��^�`�}�a�\��ґ�X�?���֣6<���
���8c�YB�{��������D{fyqI }||\�����9��M��-����0��!�MNblj�Mt�U~6=����Xh,��nb��0:=-т]�?���*c�H*e,���u8�@J� �||@�Ro��ЉŰ}{��JPB-���L�dq��#����w��KM�(E=�d�x_"K/�)s�ϰ��"s��*��e��Z����!��c���[4V9���n��ٮ�!wz��I���Hؽ�yh�1�mތɳ�Dst�t;?�r�7��{�C?4��L��`�N���7~����?��_�#o�S�Y*a��C��Q�u�^��.�����4U��k֥���<�tx[��(ͳ�yK�S�\D��=��hs1u��s�|��X���i[�za��R�%�3��iD�P��R���Z�����F	F�u�Y��i���'�n|T�Fy�r�b��۰��]�,!l��yn���X^8*��Z�,�k1F�P<p�f *�J^�f�!���vi��Μ{v���k!�5:mɇ���M"�~�R�
�hk[2�	��'�u�C����[���ppqN�Ԫ�GF����&�$���)IK�h�P񈋴D�|Y�6�a	��.�ת�|-��_���o����5,�yca��$E-��0�0<����.
���d8��ټq)c��z��'��U3��M�Z�������4��F�4(r|�\��h��x��|�z��0u�8��x�۽k۫����� ��������g���/~p��;>��`���ڟ|��۷cb��q�5yꡕ�ؔ    IDAT[@��%�j��e����-�S\�]����X0/vҲ��=G,#�u�~Y����͘�mV�q��������������K��}602�K�:i �j��O���Pz�ђ�	��|�)�և112
7���|rdL���؃J������y�M)W�k�p��SB�c]:��O�����P2	X�$���נ�����U�|�U�A#+ f¾�&9eU�����F�����}�f�� <������Ә�F+���n��p��!�f��F���Y��K}�4Aml��
� �W�y��z���v�x�A�h7�=���bi�.�&�&�R�P7� eY ���.�4�b�&���
�L��ZӲ�e��s6��g�?]=���`n(�T8�Dh;�t[������k�ƞNO �k�5��x�{�3��k�`�cG` �Y�C��W���v����s�VZY��mC�t�8��s	�
8�ۗ�km�z6��M� ��hңP���8Xd?�qL���瞃���g �p.Z�����t;t��8����Bݫ�q�����e�և���]¦�A�頹����0FGG�ߏ��{�ĞG%�P���1F�e�LilR);�TE�PǪ��Q�3�n�K�
��]G�!^s�1���2�lfCӺ5s�,S�s�W�N`]��������*c����_�blvS�6�������%�^ jhCc��+���F�f�2 �<�%6��4�*B!��u�]x�����{B���,|��.���!�5������̐���u�3EF�l���F>__��t$��-Qk�.�m�@gĨ>>����GJe�s��׾����{����������4u]q��i?��7|�?��ѽ�ϵ{1j�A��(�� �H�R�4��r��K�16��B�_?�A�a�Jc%,�,yܹ9l{�5�x�+�v�VB�hDm������V S=
�tC<�ȣ8��>�s�Y��/<�ɱQ��Cu��=��"n7�!<z��&V���Yi�D�6�����TM��iS�,�oj�	��N� ��~�q#0�C��h�\GK���@�-#����E���d��W��E'�D��a��̓�G�Z �2���Laj�z�������b��P����86�K��F��KP�xPD��Ntl���m ��}w��7�޵ӑ�z7F-JP7Ϟ���ة��{��Q� d��̏G�\K\&c�Ks�\��:�)�"RD@Ob��?'��IQ���_��Z���۶���7��K�����������O�q>�o������߼�Oo�>�ԅ�{1�Y+�*��l��&�$��u�Yk���>@�wiC�JzӗNTO�{~e7+�ڽ�/�����R�.��/��E3Ӣ�~h�(Z�R6B�PT�������,���8�O>���n���(�N���vanz
ӳ3@����܏]��/d[�Dj�݈c���8�*i�^��UK\C�
�
���qC�,��d���eQ[�gI��`�x髻���UOH�������/��yr(�ʖ���	��'�0Y��Loڄ��$J�ѭ�G�QER�	�i���F��=l���^�[���M�&�c��8�(�1�� ���N<�����~l�˘��(u:h$�P,��q���I������Ǜ�k��e>�i�g}�2�t���!�y*:��{��C�8�ҋ�X�aqt�g��ڛ.��_{�D�J�}#0 �������u߹��=y�|:����_�yK!���O#������#VR��e7=�-���8{oS[�9�4��;-�������l~ͫ�-[��|~eq��V l,#\Y�vu�h�, n5�=4������3���؄��!�FRS�\\V�\beqQ��]��=��遳�Vկ�NiW��%Man�9p�iD;�Z���/��(��_�}�*��PL_n������-�JTr��x�� �79���N��w��#˽�9X�v�&Г����q�Mϡ29����6l�Z��KK�Gw�e�G�P���(���U{)����/��JU����ؽ��N����1�K1S^ ��@��DQG������<�gtg3�kt�럿����{���3w~D����Ն���̭áj�������+����?�1���F` ������w_��[?�����mYN���0 �]������!w���IM����P�p1�\G\`�E��e����)��,�X����0ő=��i��~b��`��'1;2�Z�b������@5����,<��ţb���.OP-(�}G�v�@�K֊���Y�G��&tI��L�V~�����,џ]jU��t��B�9�[@/N�lc0Q�"}�}���$�G� �k�i�.O�޿�
'�]%M��p�K�V�gǹ�iT''P����P�I�}�"Bytq�GˉD��21���z�:	k�=��j��b$���Ů�܆���T�1#a�JK3�(	1Bސ��y��Hq�a�p��t��H��8V�{��0ϮkF��$9T��x��(m=G��?���7^��q�`9����� �Od�N�}������o���?;��cc�@���o=�5 ����A;r��^�xM�Y�L5Io��� %���LN`��k1}��(m;M���G]!L��|����"�?��^�3�6����'Bʤ�9�L�۹i���}����i�,a�D"dSӳ&�V=�3b��dV�r3^�pJ�1!�m��o�kg)��U�E�Lv|S:��楿�P��+7��,� �Lg��<�����2A�pEֶT1x�4a��<>���Mc��8C��y*e�/uY-��Z_;N023���[�Q�TB����W�+l 45���
���(�)��K)U��%<�oc�]p��{��:!j,�k�1lJݎ��$+8mJ�֚��Jq�ۦ��3}�y�z�v\ϙ�{h�Ê��w�R����G27���џ�^x�M�{�*�^����� ���#w
��~�_��G�;qh~�F����p;���X[������7m{_��hf�*�B?f�,��𱅽.�3�Ԭz�ۉ��e���:�6�8��������N[���ԡg���%!�~l�h���6ҥ�ye��ae~�x �}z+�ػs'�z�<�(�����ԃ�E&bఎ����Ą�/�<GۜJ���9ii{j�$Sֳ�gY/pM5�>�:�`��y������A=����^�<�I f�U�\��h��QeH�B�&p$������1���X_BӅԩKj�uЦ�ņ4�CR�^GT��:=����N��Xn��HCTf'043������������$�.��h{Ý_�{��L�.F�c��r�d����X?���	��~-R\�1�A�?8@>=&���Dǽ%!�Pj�I��z.��0�^|�(��ׇ�9����_~��ShY��0@�d:%�
������|��>px�t/�hT\�]e�8C�[|īLU
�7``�Y�Vզ�^���}-W�9Q2�W��Ҁ$�u��q�o٭����31�͗^�s��x���B�K�%#��.���%<~�CI]��a������1��jc��!!��ԈS���0�G��(�n}j�>��_n��!_�89^��F�du+��W���C�}�������C�\��Lm�`��)�k��~>�����P��Iz����M�D��`|��86��l�&���ia�����c��mpF��M��C���:�rI��+~��jXi���Qt�<����5,?�(N��1��b�dC���Z)a�A����0�,3JM�}jF������x�8;f�[�:��`�|9���8XHUϽi���(x��!��Fsb�-W]{�eo{��'��p�ky�9�⸇S�*�~j>�g}W����{ H��w?�����?{.�1L��Jh��^���6�A��f�6�BW�;Zvk���o�9�0��W�����5��Q��qp	�3S���B�����<C�+��U'��G��[XA{~��%l���O"]^�\���'G����R���,5�n�>���+޶� y_�Lx����|��O�}�M
�k:AY<{1>�m�	Эa��7��<��e�tݯ e��-���f��/	���|;R̜~f�lA0<���,F1��I�S�:�t��p��6�UJ�g�y9�QjwQnw0׽�����]wc+�����<D=}������El�F-��+*rm�շx<#�nU4�8�V���Yу�旊B�|��-�U�jۯ���4Y?���/ſ��ַ�|�_���'����� �O�i�\Y��/x������c���ť3�%
�AꈗZ��HT���s-��K�A�NE�\?W@�bJ0�襗}����<���n����w`��1t�y*�B��3w�����	��r~���>��7l�\����v�#���B�n���(�XY�4`�wf���Y'���ъ��О���0�3z ����H�5��t���D���t�.�Ր�
�-��GU�˯���eNM|�Y�I��F�����%�nފ�Mp��¢��45����@�z�cc�y.�S���򴥲+��U��6:X��=��+���w�s����Z7��K�D�f����J�z
�J�4����g�G�Lύ�QT6��n?��~ V��U���Up��W�;5��l�7����m��v?/_��IN� �)�h�ݍ��>p�����ozq�HQ異tF@$�+��� �~�;�Y6砧b$K��Ee�c�g�����D(���ֻ���F�b9vЭc悋��W���|`��n�����0������[�N/��hԛUl5W��lcp ,�0�Ɣb�y��%�f6	�PB CH_JB1�{�l#aɖ%��h�̝�O������{�ѹS$c�ҽ~�f�����~���S���Sxs�cS���46	s"��=�ػq���}�%F�QG�ꦁ�WZ���핓��tH�nm�k�P�L�ҭ�s��?�C�⩊s2�,��="�
��r��A�u�Ի��g�<�^'B�f�=I`��,G����(R) ��Eb�;6��"�x������-�$\$::QRD�[�4%aE9 �0X�)�
:���c���잽H�KXoB����y���t�k� �#R4�4��âO!���e��4� �g6_����� ]�t��C,ISȝv�Ep���CG��s~���7���͛�>�e��U���Y>5(�>����Ƈ����'3�z\&�f�T�D�Kb}�� ��r�B��2�й����K
��abd��G���MW }�@*��Q�i�-��I�#GZ�ӄ��a��زb%��cp�^���1D,��m�S��2�u�Ǧ/�����G�r��X�+>���XŃ�^��5�s&���`-@�^���%O�nQK�k���]=E�B��Cg�����o	@'����	Y
�b1��a�F���-T�`��[Lj���#�ݍļ.�5�KÈŠǣ�ڛ!�4M	8�����F��"I)����s�C8���&r�Sbh�>��ķI_��2�ޣ�gJF����&�4�3�(�1�{��G�iL(BA,w�i	H�rT�&��G�cQ�c~��iL�wεo���믯�Y������TG��?���o|��������׭ʡOrg�̗r�o:�E�iJ�#��jg:-���vak*K�-u�*,����]��@W$�M
��!&x��fv6�D��>��R,aaG;��E�1��о}�c��U�F�/�؛�����.gk3�	�s9DV��j:��+���ӡ���ƹ z�*�ȡ�j����t��߮������KidHQ��k\��;&�u�ѐ�M �B:���؄��+��ѐ�@� #�ӘDCgg�{�Zb��MGp������pG����<�bQ�#O�^<�3�y��̓<t��n���&�o`Du�kG�>�:���I�EF&�Wj�h��_v)��xnx��W]u�5𩺰�|==ݗ_���~�'�B�ï�xãw~��c�{�[�D\���^�RCm�d=@��L� �s�y�����R���S���@	���Ж.��7_�����r���BV� �u(E��P��Jc��`�Ә:v��a�����)�c^�I������2y���N����W�텍��
^ٗ��$w�Ha!ioǙ�U3=���^U�x)ᡋ��#�y���U���"��Ϗ�R�ʙ�W���:����-D8�I@�yL�dR�z�DW�߉,&���;���Ձ���aa�c��R\E˂>D�P	��#^vќL ��ݯ��O��S������ge���P|��j�3��ܧt�)���C���!�\�]�1�9�S�֐Ĺ�_������{�%~�g?[/[�酨?� }.PP�3a�GQ�?���O����mc�����4���eDB�����`Y���"�uEs<@粮�C�N%OvDÄ�`TUкn-�y�ۀ����ym�eC.��'���<�%�V3Q�T�@os#��܅������ ���FYA\���)��v��S�!�"B�X�Pt�/�x��*�1����1���\��=���)A���}!v�;KdPD���/<�.�����k׫���01�7�S���:"�S����eU�IZ���:G�s�E�r̊�1����[�w�:H,X�Dg��67A�f/���8\�D�R�80:����þ�C,=��$�6)R���)�y�		|1>b��u����i���eXȝ�Tt���^ȝ�;���3�^)�~3o�[����~&�)��=ԡ褆�԰�9;�>���}�[�o��,o/�h��|x)oJ�![�ek�a���˗p
-y�'a�ș��H*ݘ�"�k������ף��-@c��g�r0��6,�Y8#Yt+Mh*I?؏��W`�'Q�:�|1�FL�����GV�=�jϺ��p�53#9R�\{������C�	��qx��Yf�aa|)]�W���V�Ә��9�]tA��5��}a^�8o�T:��.��ԐA!�,b�i�3�B�>�0�C�H��BO$`$��,�t+&��0n��"�z�AK5��d�qDR1d�SHj*:�Q���zrv��4��|������6"$z�:��Pd��ͳ`��Gk��41�l8���2>��\�M!�B�Щ�	"̨�	JQͼ�b�UW�jkÞL�77�zӟ��g��zZ���z�չ�#
�O�{�_��W���+�K:U@�$���duf@��E0K"�iC��*��\4Y��jH�2�m�܊y[7!�q�D�"���J�(Ԟ�c��z�@c΅������df!T�F��U
�����P�7ŅP�x��k��)�����&Hq3z�>�������5�	z�U�聧 m�ޑê�WL�N��B�ǥZn��Ȁ�y���!ϟ��C��.q~f8]]���Ƅ�j�	�
����Bijƒ�>�Ձ��7�J��cDۛH+vDb�t�Pm�8pt{�{��	m��<u
�s��2�1�C��A���c��~�;��s���FQ�1��E��ҭ����7J/vn�|K��vշ>q�8@�?乍��c�6��}W�����]jxty�A�� զP�\���eu3"��k2'��ia>!��zHC�©��K�ސ�6J($�ټ��~-�U�F��I��y�P�4���աg�l�OB��+�C���ǎ��B��Y$!J5Iq(�@N�1WʋȨ`\vj����`J�����碏���A43��E���J��@,N$B�<�@ej�{�r�^�� �k&@#�Ia4<xO�i�n�{�>�y�p���q�AnQq����N�7��;.r�Ĵ�K�(���pś wv���(yt�\�x{+U��� 3"�h�0��ͮ���p��gp�m��ba�1��)�q+¶�r�]��3�����p��a�-8.y�l�H9t��v�)�K��_H��D    IDAT[{��|�f�.���ݵ����O�t���������:���3���/��wn{��_��_v�
�{,I�K�$�H��B����X�>@�E�}K�Sz��zV�����'�Y&�D&�5�,a�嗡ㆷ��0�230��~��l�D� TK�[2!K�d���:sxq���+��$����,�T=U3��1���� ��-��+C`ƚ�W���z@@N� ���^�'@�� $�*p���e�r'��Zh?4O�<_:�@�n6�CQ�����E�J���UT��`�>�2r���%��p�zȝ�8�g�lіVDZ��lA)JanjDCJ��L�������ϠM7�!ɈQ	#��y=��r�c浢%@/�,�Y#ĝ���
@��{.����[6+[3T�˖�w�3M���7]��:����p�u@��9��a��O� >��K7���_�|g.���q�0x�nR�ʀ��4��:yf���2 /�ʼ��y�Bɖ�hi ���\,������� ֬���!���i�!�:r��f�4�f���e�%��8҇�b��AH�,:#$��4]�N�K�a:�x��1I�n8��,��^f���t5 ���gi��AL{t���,
1C�B��@�<~8�sdlN�p�r�����+.�bljY����cx]˨ɉ�h7�]X}�pۛ1��Ѻ��=ГI��l��&-�����?�Wx��|ɩ<:eI�fM]�����ȂWw�̶��]�gM^���E��y	�  W����d`�9�ѹb9�:$�Hq���/��:��Y{�:������8z~��w��_ߙ^:�#�i��X�q���e�~�fK����6�!��ޠ�@��$�D(�jĐea�1�ŗnE�E�{������Jp��SL"f�h�"�&s���I��B��1�SS��Z�T����" ��B���x�|�{�e6�4o����zd.�O���&D ��O�	������
g9x�>�.��0V<	v{��5
�j���k��� �[w�8��E?X���ɧM�&���48'���I"�q�;�v��#tjo�F�� 	��浣a�t�X���47#����F*'���u,4������_އ��MY˓I$t2��9����B�A�\�l�+w�3F<Rܔkc�2��IO�U�,_��V�D��!U�ٵq�-������O=���S��:������'@�_��g���G�� @o���Y�S��s�X�r�u�|�f^:�7��S!��Đ�-�9�b4lZ����F`�Z�YX��l.G���� y*GK#^����12��� }� ���UA��A��FU��~�xR�gY]�K� !�Y���ג��y %���.[�L硟������W�N_l#
Ђv�>6�_��)n:F;��˅(�+�8��B�ſK[x|ѕ��(�� ��h��
���QUeeo9׆-��S��Z/BӒ�p�Z��F u�Aio������T^KDSgƟq���?���k,"�����&<�^�u����G0��+�7g�Y�]ڱ���q�ۚ"�P5,[�֭Ł|�d��s7�r�w�:����	�*�\'C�a���2�޸9��'���^�����WGƖu{JqԼ�D6#��6�U��$3I�]� �כ��E�+kV�ʬWv)�pDA�uX�;���"���SN��C��:2�C��l��$�ۣ#�<ԏ��:Z)ʃR�:�k���X}�D�E<��@�k�ʼs�=��T�aR��㑺<�샀νUO�&P�V�<��&���������/�D�_Z�����zu��ek��p�d&&�`�s�w�Y�Uo`��%��,�Sg�t(�Û��A�3��ݰQTH榉lX��)IAÒEXy��H�E&��y�
�M)�Q6uk�)$c�i��?���L>�K�Q�m�Is#O��V���%���g���WE:�"|V�S�s���L�}�x#�]tUŒ5������������6�v��?~z������W>c��g�T���F~��u���G�r痕Cǖ���_4�����w�2�7�E��[%oī9�4��,
�FQ�U*��������n4n�#�`�X ,	v����0���P�9:�VȈ����~X�@!��"#Aet&��]��L2
B�G�����0�g�B�7��p@��pu�Xb�B��j�?��P�=�HW>W����sظ�\p�يߊ��ſki�����.�H�/b����W�郆�	� �R���J����riUb��Sd�-[���>��5%�����+�������y�ӖP|� v����؉YF3\�Io�h$��1�e1�Iuy�~�L���|��Ԥ��ڞ{�@I��s)��0�1ܩWu�k��`�x�d���|b�������C�3/Y�-��:���Ӄy���^����5���e�����	Щ��2�
F�t��y�Nu�m�����3g��sECZ�`<G��`��^�\TAN!�(��i8�&�ǆ���0�sd����!�f��9h���d�d�1��r�V9ᚹ_oq��w��`}���C��,���Մ�.���_�u�>Cf���Z��S���|�p�����i��{����^�A)�@Q�����1�¼�Kз�\�P�ZS
����[�dNL��P���t]4;

�ދ]w݇��=h3m���{��� ���9�	�%D5����~E�� �S
�K���;�P�0A5�v�����Xy��ȧ��3=�|d媏���/օeNeB�������9�IqG�>��o|�=ppz#,�Q�w��N� t�PYj�S�Ӧ�;����T��~�]y1�b1
z	9S�m�@ހ>��؁#Ќ�j&ÈoSAG�uШj��2bC�E�������������̞� �`�
P��ȕ,�H���a,�<5�f��q�����2��Gj�����)�^�h	��j�@D�����溦!mеږ/AlQ��������0�*j�
�)H%`��g��{?���jM��8I��n�#:�sZ������ftF�1�Z�Rؽ� ]`�E`D���̒+����n�螚c��o�f�ԷyuF��<���zuF�up��Gb���]z���u����n�X�.����r��j] :�9y1�u��MSd8����b4�!�~5���>`�|�$Mc`>|t IWA4o";0���y�c(=���1����S��ڹ�f7e�IJ��!���^�7ez�l��]�g��M��ܸF�{��}��:����;�˱W?��Y�ܭ֑*�P�O�V�!���D�t
	ţ)P�"hY���AO&Xw3���ݰ�`���7EA��"��q��G������O���0�L��WU	i�SU�#Ae%zd�IpdO?�k�J~=c�{!w�g%��B���K�6wvbɦ8b[�������S=_���G���Y7�����Y7�g��O��~��_��W#��/�Q%4���ƞ
��_�U�yh�y1��,�`r6k@�4��D�.Y����-��	�f���,h��Ɂ!(�"��"�|R���� ���� eh�%��]�������Ty��O��C뵞����3�e%�.�2�P�t9rqn���
�/q-o��w\���7�_��=@�S����Iz��X����bQL�@˲�h[�Z{����#�x>J�(��G�!�.Zdz	~��ɽH�Lb�CʶY9�Gx�tHl�E�<@gO�ۄ��8S��. ��k',�Sw˝��-MXx�:Z��lC�����{>��w�ۧ�u�շ��:����B�c�^~�_����t+@�c#A�-m*_�$'��&�A�-���pbSh�-��˰��+���"�1���u�>2	'S@ap����d��rã���ˠ�v�$Iz�P��GN��@�����^k@FD�^�t1���."�,���Eޚ_��'�L��@�Y�@[U��]T5���'�ث��o+<�*=zaY�12̘��b�x-K1y6�b�u_���Vcr"��P��-�@���w�G}�6� !b�Hh2S�]=�ޜ5��tx��
��(y�yȘ"b����*�t���F,�p.���Rԧz�^��+n�������#�T�U���7'���n�}Egr������O��������^��LI	�x��\D�X���N>2o�A�N��J�Eɕ1Lݲ浢�����֫�6a�6Q,�:��4JC��>�NIe,�c/����G`e�H9.�-�aCs�܈���.�"-�eH'E��A2&f�0�zśO��tܹ���s|&���0�����Hx~���7����Z�M�k]lJ: �H9��5�U2cQ��Z��ի1QPlN]�L^kjf%pK��<��R(�t �<��'�#�ɢÖ���)�:ĕ/���Ih��|��s���	@�p�'��X�Dͺ.M��[�vw;���+����O��O)�L^uf3C��mN�(�-z}B�����]��Ƿ��/}�:&s=ݪ���#E�G�/:�u���C��\�'ɚ
��?\iH�lmD��-X�֫!�Z��bˁ[4�L�P�Dz�G�X��nY8�krc�,Ğ�%D-�XH���ڬ,��O��@.)�^��Ӕ���M���x�����9Y@���� ӼbhԞ}~�>��O�	Ԯ֯U�&�^�����WX�؞g.껽qF2�>�穑�Sg�#�@�9�гe�e`�uмx	��G�5��4X�,��Z���������X`�h��LU���������x/�r ��NQ+��FekE%�QC�8գSZ@S��l(��V.C�ڕ��]��~ߟ~��7Q�������{��+����4�?q���������.�Eʱ�]4(�+����G'R� &�X��(r�������B�ۯ��a�5�[.̢�����qL�8�@_C3��������s��bp� ���W:��e���y�mw7�<-S;X�\��/B�b�rUT�]AX���T��ǟ�fjdA��t����q{����3��k��|�3�#���\fzO<����#x����.zB����nm%UFNS����}�:�߸�L:6�����D��!8q"rФ�����CO����=S::t�.I����XTX Nju�W�]�$�I�A�N�G�ٞuL�e!��ĉqT�ni
�l<�nk���M��v�׻��4���O?u@?�g��#?i}���������l;z�m!b;H���z�3�8���e^�o�0iY��pW,Ĺ��h� #9(�wd�a���3:��_B��c��U�<���ێ�^����㔓��.t.�pD�puZ|��)-�����h5��@V�"�\.g�s�*�	c���ܹ��?<bP9RX?m�]ؔ��g�G䰃u�'s�Z�Q1\*7:#`�W-8����t�ζ��i�<(�b�w�j�Mh��h_�����;;`���Ԙ@co7Ł��PU1�Dt<�}�>��?�������<�Da}���J
L�;)ݱ�b�}*��r�i���c3� �"n,����c�>��Ϸl�rۍ��/��S�w���3=���������Y��+q�I�+>v˶o��g:3�V�i��-�5�`u��V���	jL+��zH
bZ�JE�,D�[ބ��.e�˱,5�T��6�B	���Q_��QL�rK��Q�Ⱦ��^Ee��M��t6j�b�%5Ot���<�0P:1<�s�ܧ��_"F��#X��cP��읪r������k�f����\r�Fn�b4T%>��>����m=y�=�:QI��ގε�иzr�q��Rh^��*(b\�'Qص�}�N4M`����!�y��	Ts$�6��r�:�� �͔�dIa`>� ]FVrQ Q��� =�d�Uu{��o��#��Ӳ�Ozƌ@�ϘGyr7��H��������o6/Wj�$4:6���X��4�Uؒ'�r�6�f�$��"g������k����@okƄiA1�4��Ґsy��݇X.��8����J��h�f8�X�nJt�������/��\�IO��j{�e�+�*K"�L�NZ+�/[�:�+{�8#�_Y-���5�� 0��>�R��x�n�C'ź�e��t���e�]ފ1E'ńa�(khX��kV"�l!�E�`��pdjc�`"� AOsd�x��}��l)E�l�L5��dqB�8׀�<:}�T`I�N�2i�~��5IBNv�wX����#�b�����ο����}�ɽ����#����8�G���~t���_t���.�A�� �8�;'1J��2dVx�l�U�m�a�Z,��7#�q=�F[F��"?0��}��r9$�%8�cH�,���v&��a��d�N[�����ނ5LҳB��:rU>@��y������+E
4O�9�jàVź_�տGY�&�W;X+��ݟL�6�vaV�Q|��.��}g[x0]I���� �"4LK�k̪��o!�|z�J�Q�F!�t�炍hܰ�*�&S@c#̸�!S�')؜�]?�9�>�Z�:�5	2,���(��:J\}���	�����s��%,:�\$/�������.��>P�C?���S����~�C��>�����/��g�v�}��h�:\�:-^�I��Y�j�z�Q	�Ú��G$������چ����]�u�2G2���yn��Q,kk�5<��}���@��f����3�`��vӛ�����$˭z�pl�d��ա�Z�c0d\Ԣ���� t?����eb��u�Gc7���">o��C�3y�s	{�	8�c�E�{CN�G��8�0��9�՛G�)���,iQ�EF��hݰ��&(��a� �5��j�j#&�h�5�_��w�3���豁NEeM��X3M����� ���QI�����&mcL�]B^�9tKU�x�y���?��y[�~t�;o��{9=�W_���N��;i��߽c�?|�SJv��1��4x䴈��(
���r��I@��Bl|����6dsE��p�=6�x��̞������Q: �d0@�a .ɈxR�j�B�,tI@I!w�/�N�3�i���s�3}��ʢi��MWV[S��w H�.�9���W��A@�!A����]��l��Z�^��{��=x�aFK-�W���+EnH���=V�'�U�1��8r%Y�a�2RO���"~�Ƚ�@C��
%�`R�	�EC����>���Fb`�\�7-"��cC&@�\����8�8G�N!�,���6+[�����C�/Z�����/�����`=�>Ӌ�Z?�@�k}U5�7���us���-����/�=������}��]d!Ju፶�8�yYkT�=ʒ�D]�k��H�5�xc���/Xp���*2�L��%L<yx͙��d`mP%��(5~q	�]H��<"���{��+Қ�x�'/�☇&jҧ�0 b�dߛ�Q�% =��۶U�w.NO &T�����0������B�a�.�Aָ8�}���v}a��A���L����C�2�E*�B��_x���IS��qg�v�mAڤ�pm�B�e���u�h
�dE���e4�
��_��g���"��oЖ+�)ݖU�E�������{ٔ�9t"��E��.kE�ڧ���I�&/A�����.���[?��dƪ��k~�6B��Xs�U�Z��?���G���w�˛���`���DT��Gw�1g8
C�b�ԑk�c�5�����z��+�:��	%�G��C�G��;6��� �l�� .ˈP(ݱY����=���x����	�Y�7
����Ef��C=�t���?����Y�5����hyu���E�ƫF@-�}���k*^|�~����k�u��Mʙ��3M� q�ML��D�Hq��9�����l�!�,�6Q"^���ԐĢ+��H2�����z�3>���0�TT��>r|�QڳK����$�È���N"�
�!���C݂�IrL�x���Ĩ@��%,�`��1��w���]z�'�>ӄ�?���,� �S�u�?p���-�� ���]Eq�*k�    IDAT%b���Al�4d]V��m�.݌�o{�r�l%Ä���� c���i�~�װF�Q�a�p	IB���5��׭�������`&@z���g��R� in:�����t� y:�yv���}O<��t1/�WtY�+oIѴ��,����֧^)"�W�{>�6��|_'�yh�'CT�r�l��������BoV�<Ȑ�E$�0��e(\9�դSG��cp0��{i$K���ś6 ѷ �xrG����]Z��gz���0u@?˧���#�>t߇��?|�k"�\䂅�U��X=85�P���l�DTL�5࢛oB�MQ�&2�҇�C?:��q�J*���;>
'�AB���(���I�G9$�L�l<\A����Z�Jn:v�ߩ�h��q��g���L���J���g賽�ZӜX�A�<�2���'��avL��AȰ|�8�4�U?�AX�?�ྲྀ�,��$�EAZ�����Q��D���笆�J!��۵��lQd؇�������_D{�DD���B�vN?���l6��1��$�aMY�N��;�a�y�!��`"�|���o���O��9˗����r�>ˁ:S7�︷{��'n~����L��d�B -.��Q�	��z��1d�������=���B�0��6�����$�)`d�;~�����qh�,SGB�#��(L#����}D�����jy�%�)�O�t5��c��+� 'vC�^fx�@��)!!�jO�Dն��U?�����_}�3/����.�-]��Sz�����7g�J���Ty��I�x��dX�bl�nZ�|{3
���ϟ��� �-;�4�������)��GѭE�	�a��Kڎ��C�M�*�]��t�� �݇*�i�bɦ��;:0�����o�����)����4,9c%����<���d�?y���_}�/�өc#���Vb������H�R�c<��]�k��V�睃�c�P(Bqd��G���@/u�zi�^�-=�Fx�1���?h&&��;@�Gtx<�C��i瓡V�xp���Z��a�k��1Ss����ܦtŜ�GJ�<��s;'�z6�{X��xF<�N?�z9�P�@@���wq�D�˻r�:7�G��U8B�]hZ��6��eZ�\m"��?�����ǒ��h��T�I!����%ˬa����p��!��Xu�E�;[1��j=�mo����'3��}�# F��g�\(<�����/�����ßGm�ql43���HqD(&d�Q��D���k�2t�J�����1���ci"���^z�Q�׬H�Gj�Pi	��ʚ��׃�'�e���A��{����v'�3M�0Fw�߂�'�I z�<��yŵ�s3��<Z/�m���j��l y������L���h<7�o��y�LO�Y���-z4�|2�W^�o>ҩ8"}�@k3MI��,$�������F���
��Yo[,u#�f��T�.aJ�X:	��ݲV֦��X}�%ȷ�0�i�;7_x륟��W3ͷ����&�L�:���Ov��E���}�����o��{����2�(�<����E1 �����O|X�S���cA.�0v�0rC��T4X��GG���a��hXJ"�Q'u!�&�ܳ�ʂ���RH�p����ߎ���|�l�2�b��L�*����`�3�]� 	����
eK}6E�l��{�a�Y�&��\��A�C��	��W̑����c�ST��,�.���\��z	�֭A��ȷ�@Y�FSf<
DUȒ���"^Ա�'?�޻�GA�i!I�/5#:WΔ%�v����J2��lb��p<��뒋o����u�l�Z}����:���s� ]{��}����?7��O��:t���,j �jz�؊o+�y�������ߏ�;wa}O�\��W�ٲ���$�/?�����+�8�E�R��f ��>�	�g��I���w��{�ж���Ô��^� t��ާ���c��.�k����	{E�
�aƀ�y�zg"�9�	��P�(���2�%��
����q0��cSg6((�㈭Xe�"�֮�D��q8���4�Tҡ��p�_~���(4&b���k)L3��!�y�$���>��a�y�om�XC|/������Sg�rT��S�:��� ��ww�eo�׻?�ӿ���HMN��-ͮ���]U#��̂l��fȫ�"�j���\�i`蕽�9�.EE|*�ܾ���w
���+$��1|ɏ�d&>�x���Vj�p���8����w+r�\N�$��g���B�����A<x~��K��Q���g�O?G���@ݹ ��}��2��F@���Z��zB�����>�l~����S �Z���.0�߃U׾R�|�m�pۛPT��ѮF���;?��_>�5�$Z�%$lqI��ڈj*���:0)I�s��E<@_tw��Rqjݚ������o���~��w�~z�����x�O���W������h�T62ϱ�!Ɉ�64"�Y.ҍ�}�5�y��0Z0Q4����J�#0F�a����4P�?�l�(9	Q�����7�1#������>@�k?�k!@���0��3[����B*�
��HL-@��d����Y��Ǭ���o̳��ʖArb��0��a��r!4v�Dds5�]�F6��֊��΃�݁�͛�v�c\1aG$4(*Z	O?��w��}X���tU$%	�m0�<tKS���1��0y�2�qH�0��-�`����6��V�כ?���v����G l�~���mO����6�����<UJ�zҖ����Ə}X��EVס�LGQ8
y*��1ĳy��a�M�Id�O� �<t�am-���<(ߊ����T��YYӉ��L䲰:�0௺_	��N��rc��9�H}s9����/y�G`|*���Ze}���b�Ey�V�a��?�#�G yp\�dp�#@7e���
�BA�0ֻ��N]�p��CY؋�(�6���&Z4ё4^��~>�(Z&�h+:h���Ng����j��R\^��[.�Ă�j8�����H�at��O|�o�<�������-Gub��F�����=������?n׺�d��2�hq��*���a����ъq��2�t��2�f���;w��<>��i��4�������vO���% �Jju��o�k�)�?�����{��!�6G���2l�2�2��0{�s����TT ��tL�����;�����>W�"�x��̅� @�=���_��y��I�QU`X6L-��,c,�!�l)�^q"�!�����������{��O�F��m�耂��-����P�%�:�] �����[6�hn�Y�����O�e�Է������7
���V��Mܧ~�p򹝷��ů|�y4���Z\	�$#�*��8���@�5�!�G�Ը,���^܋�T=��#��@�@?�"܈�.+Qc,\�(pl���B��Ljt~@/{�^�<���l ]xoe/ЫO�k<�O?~�j�z���� �V��l��傞��Чؙ ��1�	
���f2T�{DB��i�s�������)�0l�u��%�0�����в�\���%�{`��X]�k�#ak��3�����8�(Q�(Qh�/�2������9�p1���I˝�ٲ��u�a�bG���.����>����E�~S�������]f�D��(=x������]_��';����mĨ5��aL�0�ӎ�?v�sV �((
��`4�¡c0A��`�a�յѨ(�l޴�L~s9�sV��jq��D.��_xx����d]��������9��4����AZ�����c2�����=t��O�v|;�����P���n������~Rap~x�pU��7���i01*es�AK2��΍Ѷe3�С�\��NL�mY������!<���c$�^D��m���:�*e@?΀�k7��W�]�
х}(u�=z��o��˯��o�=����:��Ϲ�]��k��m���_��3W�|�:�Y�J@�%��k.ź߽��L�&����I((#0�~�(���ٲ�&KH)
��j̩N�`[f�N���?�r���?�~���r$�;s�.eAP��ڙ�k�{#�*����Ӆ����0���jq� ���A��
' ]�OO��[kM�0�W�����0ÄW;T?�`b�8U,}���V��ե6�.L�e�o
�G/B��-on@��a57BWI# �Cb�2��0~�ӻ1���h��R��g���p� &Q��q�Щ��I�p�"c�����w!����e���]qË���6��5u@?����ϗ����z�[����\	�Tb&�����$6�G^�0�/A��?:gp��(���8��yC#��#�� ;��0=2:!':}�@�w�i. ]!�m��@/��k|%��j�*L�.��t�����)�B��O��O(�y唷 o��Ѓ ?W@���ӗ����т��tb�[e�Z">b�DH�Ol<a.м*7��+g&C��-WU�m�|�i�p�*&mFS������ǲ����c�%AK�Vf���g����!���L�]#0w,(�����:����:M7EƲ͛мz9�d�v,�z�G����������ToK֩�����y�'~��ȃ��C_����
&�!�h��+��bl|�M@O�
%؆	kl�����0�D|`��`f�H��+2ׂ
	�m3,�+�V��
�UB�U�h��T��O�)���'LC�zOH���4��@\>���_�~{�4+ �_�`�u�Ϧ�m69f����d)E�}��T-��-t��0���d��g2���#"��/o�g���\<z�Կ=W�f�T�w�~|ؽ��®�E��v��N�"HԷ�Xڄ�ᆬ ��s��-���W�ZЍlstM�*kШ�e!�-�ɯ}ٝ��ihW5���r`@�$���<#I(I.��W-G��������ѕ+���/��c�絢~m�������V���v��c=�'}囷��Jht\`b�)���z�]s5�)L�pK:��qV���� r|�v��m��?4��R�
�xE��K��$_�G��p\�D�U��P��/��=��3�}y�� <^<\r�|���{"7~�����Õ�uu��*Op�O�
��_*ҥ� t&�b]��cL��_���W�g�8���3@�����7]C-@�&�k���ZĿ`�q9x����G_������a�H��!+)��a��W�8�����IHr0m4�
:���wq���A͍z""tϦ�"@�SK֐���YQ,��FӚU�>8�rr��?���~��S�R���빉�)��Y�s�Ϣ���l���#����W��xK&�8�ɩ!��%���@[�i�F�d�����ab�4er��"�s7�l��x�z���v�d09�HL�2k|���gY�kӽf+���W��[dV��\��k�Z�ȫ=I���Eĵ��g�"$-������<|���Y���`��!�s���l<t~Ue��Y����`��*��9� `�xE<�Z�?fNC~�_�"�����l��I(:��%%-�l*�o���^X���6�����ͦ�C�?�'��;�W��#ry�dKL�n�ڧ*�$׆�`�y��r�*<s��ˍk6��ǿ��u���|=>�ۯ����|�ү~���C���Ǿ�7�d����(ι�-X���Í�1iX��u����aL��2�cCp�6<��m!"�,�.;6j�JݧHP�C�
��R�C(���Xt�eM<<̻�	@g��ˈ C!�uWc�q
������l�<7Nd����.�ţ�|�����*u0���S���.a�=]�?�.B� <5@��@'�q���d �mx�����O�R�4,������dh&�3�#W�!��KOG5,��J�l^�bo'J����@L�Р����S��{0_��MA#i/X.tGB�u1���3�Ę�r\��-�ѱf��ͼ.�Ȼ��g�y�/'��?�#P��� N���ܽ�����g����i��jW����1e��n���(�s�2E`p8v��/c�嗑*�(IPI>�Tx:
ʅ�����䑘�J�j@zVe0�P� �̎WU�sڢо#����T+OM9<����%j��c�lQg5�'z{�{�� ��g�Q
�Bl���u�b����j)��:>�3�>̐�MȪ��x~@g��u��*�,"����?��7a�ߏ�DD������^��"����$��B��T4�Ě�X��k�%}Ȥ�(P%�D�b���L�|{~���,��"���+a�61�:���224_�*6��R$,ľ|n���r�e7x��^��c�@����>��������>��Ｃ%o@r-4�Z�7�٧`��H۔�� 74i"ix��Ln���h�4�D��='�K�mǮl)�J�T<A��{v��. ����ۚ�)꣥j\0Ĳ��Z���(o�LC�R$�:�0b]�eЃ�^Aᓹ�teSt,?�@O����g��E.���E��X��4���dC�'�t?a9�WЅ�W�Ѕ��:'Kz
�>@�	2tHK22͍Xq�5h�h3JM�D4�h��.���vہ���|럡AT$ey�F�41
 9H��{L�E׾�y�8l�;V]s퇶��z��\_���U#P��|B��ź=���_������B�``�e[��7cR%�
�=7��@����_�ml�p�Ty>��(�ډ�F�8�3��S :��`�'I	�'���7y�~�/�rM	���"�#=8���h����0E�(?�։Ů����w駚�=�)Q+W�w��p�+,wo܂fX�8�6g�o�8�΂!�Zە�����j�t�aV�wtʣ���.?]���	� g㡫>2%��"I�K'��QMEb�J�}���=���U��&Ⲅ�^BS��ǿ�/�ܱݎ�F%��mc�61! ]&@���p���?_x�s˅�\���=�ټ|�mj�@����1����?��_������R���&6�x���:L�U�L�%Aϡ��՞m�k���.���źI�q�[�� ��u?��9���;����>4�x���@� M!��c+��U��5��|�&����"nf:�FU1�#��贿E�U��F�`��w�&=��}�#
��Ix}��)$D�v����;���$,d��.Xہ�v����Hi�B�ec!Ȝ�z�تX3:�6W1
���*z���5��@�K0�A-bo i�:4_��: ������#��)\p��AZއ�TF*� =��4�u;��C~�	�7U4kQ�lS����)긦PԀ+n�m���P��B���n��#��ס���1�!�\���s�3l{}��v���m��w�o������[ރ��_��IҀ�i4yp��q��m���åv��J$6m���{��40�	Q�>�O��s3p�Յ),4�� }^+z�РF0q|YJ	�dhȐM1"�1���-f^-�d$���A�L�Q�� �Ǩ��l�@J������b�h��y��Q!��@ꂮݯdJt���W_)D�@<�R�L�K�C��+cq" s���PD�"2���n�w��|4��)1`�X2��o��_�LSS	v�j:l$�.���`�w�^SA�e�5�z�נ�����T��p=ܦ&�
;�6]p��'��4^����x�����g���oi#@���?��s���k�\��\���#z�*�]��dJP'���ŗq�ɧё�1_�@5m�L��7�^@/������)$s�H�Sa@Nb!�6	`�8�q��e��q�p�"�s�0Z*�#tV�]��
��k��_0��ˀJa�>3�D��p�����z�}.���qg���E��
_6_=���L3�ܒ:����T��1MC|����Z�z�o�A��p[���    IDAT%��ݛ��/���H��C������3�E�������\t�5H�̧p����|p�{o~a�n}���0u@?�'�����/�}�����_m����K����A�MC6��<"Y����	��܅�O>�.�e�rQ�r�$)[�=6�7�~��r��v'�uޕ�X�$O���򘙢�B�q	�I
ǆF�.G ��m�@��Ӟ��������jm�%��`-��ƀ'��;x�g���;�t9|�M�[�A �����N��e��2��#�^|^�t���<�8��W�N�:RKU�Ƙ�`��	���.�6�G:AQS`����X��撅���O��G�
QIA�4���)8Ⱥ`��X�_��K0��8o�7o���g\Ƚ.Vs*o����������}���^y��/=��߻��>��������1j�Q�l8�9h�<�c���Nar���t:6b���!=�0S}�T}Wy��:n�-m��ĕaftb�IO1N�TF�sm�1(�����iI���^��-4d��Iia�<F��u�lpBr�\x���Sje�<C�G���L���ٲ�gzY��[p��}��RQz�9���X�t�+���G�@z
T~I�)�,��)����el~��z�V�)�TE�L�A�f1?و��w��b�%�m!m�,l�o�ID�n�EH.��!��ݱ��]�wl��~���G`�xu�U���k3��~z���?����e=���?yi/FK�0��,�(����^ڋ��{ѥ(��6��IH��zE�S�Lk�E�yP�����4�-��7.���TYeǷ\����yP>U�5�y���t���ޭ�p�E���02������GޟVGx�̸��A����ؘxu�3=��S��E"�?'��~C�����	���.�
H�W���(���㲂%W_��s=Ҋ���d�M��T4``���0�r?����q1�,����J"s&���YЍWJ�=�n�����';����#�֗�0��#���.9�܎/�����M�o�U�{7�0b�aY�t���}�0�kJ�aA��m���E~�J�E�x�e.?��0x<�J�(שh\�C�j�S�0�r��8�x���+��۵���C��?�!�*�^��	L{���A���0��үA����
@��ɽG'���|¸���5St�����Wa`�����k�"EL�F%�U+q��n��ӆt���&3EDŰ�u4m<��⥇�@��0�}�2��n�6&SX{��,�� ��l����a�On���F�$_����)#���Ǘ�������MW��l��j���lV����������up�bI�f4��ڀ�
�XG+q��=�������ԅFy�� ��^]31��^��0M�¨/�*Oo�J��#Ȳf9n_�S���z�YE�'t��`=~���w0���k."�HT��O�a�r��)��a�~ ����"
N���6��'��&�U�c]�|���V��uM�4�Cj�䝓����ԉ�[^�`\�`�9�-�{/��aX5P�i�U*�,�h(Z������ߍNGE\�1a()@FJВHb͖�.�ư�����n���u@?S��tu@?M�z8�뺲��]W�|��/>��#믻�F���Bd�
v	v�gp��#(�f/�>��:�4��X��F`�256V_U����iA���+��Y���>�)�4��o�����M�<x~T�1�!!������xb�{�!�]Rr�V�"M,v~-"ZQ'o?!�"�-���'�\��A�C�� 7V��$ĵ�q7(a+�����b3DA�i��u�u�_�@PeV�E"�M3�ƃSa���w����hnг����7���>�Ewͧ���(���,�$ !�!6���<���l��Nke��?�V�r�Kr;ɺy�{�In<`l0�1l��X�4vK-�[=�>��﫪�Ӎ�� �����}N��_U��7�o�x�->tz�}����P_�2t��4*�k�I
�Eg~�sh��|L(�T�ɝh^ �P���^�s�<�Ӂ.�(�.��+"`x@sC#6l=~G3�`��[o����ק¾0�9����S��>� ����;]���×�y�o?��s���f,^�
U�(VK@�
ul
��#p��'��MG�r��4�x�h�<g��Y��=�/�[��_?w��_��!�x�F	�B��<�D�����4.B���o"��5'�p@]_��;���$��y��R__$������9Q Mۅ��:Xr��L[�ٵ�t�Y�nN�;neP�B�%��F�A�����Q/��U�o<9�,��*i�����@�<̮�Q�$��w��M�P���p���j�D>������׆c�3Oě���w��;nR�>�T��9��m|�s/��#:
��'1���J�'�)�T��	�|#R��M��K�G�����@WЈd�B�'`�cO���R��Ūc��%��B�Yg\t*��a}�g�uӟ��j��;m"o�`W`N�� �����?=x��m�>��~��W6}�[Ѱd��F�Z�X)C<>
��18���sh�/@V� z.V]��p���Cv��u��<�\~��p}�xs&�"@'H�����.fю��rp�t�]��YG�M�����7�Y=�8�� =~=i����
,�9A�=��(�����_�qӧ���dDcw���)�!�V��l��?�a�#&"ҿ�j"`dNB�ʞ����VoeK/��C �𹒼
��*g��>���ឫ6!���N�1����2�Y���Y��>����2���:�9)p����b�!�/�'����)	f��� lo'������1NĢEQ�8���c����GH�>���\*�n�ؔ��K.��L�`�pT\��?��w���|CX8��
ԏ. ��t���=�sO������������o�i.��j5����A����x�&�؋��Y� )�-Kߩf�|�>@�H��&X��f��̸�4�,^G�8�6ɧk��Q�����zs����&V�T�lbDG�5�Z��B &%��(���f��M Fb�MGY:g�Q�<�������W�YO6�9�<<T͋Aߡ��j�q�,����Ř)����%�~ץ��Hd�1�+53���C����l�S�q#
kB|%���+�ʫ��B�Ϛ�|�j��a��֧3� 4��C���B�@�#)��F}���,�/������B�$(~���|` ?����J��8�=b�0��&�[׬���G͎�?��_��GO��h�\>|+� �q����
�W*��W���762��˷��كذjUSH'`����K��?<�f�Ȓ.en�x��3�U�j��AeVZl�2+��zǜ�F����y�B�g�M:N}̰P��]�гA=��� `�ed�J`@���V$+:�{���8�L����ʇ��a69s�a�<[���%H��Y|����ܢRv�1l�WA N�a�<�H����!apY�>���Ѝ��lf*��`*��v�87��q�VB8��|l�e���]_v�{:m�^s�u0C�'���g7Wz�W���[辅�����F���EǂGU1�=V�������n�,ׁ�yh4��2~��{q��_Cs=���EB����26����c�u��=w}�O�����7}���P ���f���<��<X�����k�4W_{Í�.φ]����:4���=�<��1t(Ҵ�Z&4Δ�/�����������1 D ��沙c��O�0����&Ck��1g2���l#��Rw=�OW��x#�ۀ;Ǒ�KhK�@�raa��m�!�,��4)O�����hf֖�*�E}���jCmz2�{}T`b�	Jn0�
��^"t��E���O��C܋��%����Nd�:���)���NaM�樃t�p�%{��N����$t�HYp:��^@�� �Æ9A`���f�Qŀ��p��|^��U6Z9����B�����xI��q� *h4<���Ul������HI"D/�(��8Mº��m�Z��aq�;���?{���>��Ѻ������҉_JW��z��UI]���m�:,ˀW��Aph �����	{h-��FY�oY,kI�o�5s���n�'7߈�]/*��3�X�6bf(����sZ!q.����<&Mg�y.�0c6ut�$B���sc�[\��O�BY(��B���d�i��C`�J��k�D�cvAt�H��߾f�li��@x!���淂����\b��ܹUU�P�W��|������=�,t��D>�?oz~��S$'�����k����Z�ga(~;��0C���(f����z\E	�/0�߱��ǟ�pEQİg#u�i�t�($i�*11N�<���8~�/���ǑC��Le{ׁ�+Xs�f�8g+^�G��;n�������x��+0�`G������ ���ON����Z�x�bT��j~����]{Qڹ��P�E4"R��u�ֹ�ͷ�o�1�ֿ�~�8��������\��|C�%�zP��F�R0_�)�9��c����B��ʹt�ˠ���Ds�\��H#V��(��:��?O?��9%�W�bC��|b�n9���GYo�r!�^<M�����:{|x!�=�����̙&/�<;��hL.^c^��t|�"蜦G�J �����L�1�u�?f����W?Bᗹ`>�^TϹ�nD�8�Emx��I�5���d�?��X�Ɣ$����vl��׭@N	��
�@�F�
 ��x�߾�}��FF 4jm���L*Xq�F�g���Ƚ˿�G��/����FW�n��B��n���}�Y����Tr?&V>i�r�ؚj\�'u����.�j��������ES��..����i�������K��[�>����|��i����}2m�q�;,�ϔv�%��N��Ik`p��g�.́GY�,Bb->R��>k�l�2</�\n ��nq���t�
�7�X,&>��s�^�㽈z.��sv���"����=h\ގN�A5rZ�r\���Ku��0@�b�������ǣh���V _#]G��y����ֻ3���t��Z�+���foas��~bv}}��ȖqxEG�q�!�>ϯ��i@�	�,bܵ1�ֱ���a�g�BQpPU���G3T8cSx�cǓ/�A��YQs\�%�������3�+�~������޹�ү�g x��x��'�Z�;M��ri۶��j�}�1��s(�����f߇��Q�2&7���ÿ�|Yc���:W4�d�顇?�%^R77��1�Q��y�ٓ"K��F���DT
G��J�m��Ye.!�!�I`y.$M��%�t�@ZQa�60�4M�$�ϑ�Ta�9��G�\�:"�D�o{�����ɀ��$��H�Db`�%�:]S�yQE�~D��zUQ�}�2��%Tm�$!`��p֝�?�ӿe2�	��t�G�h��]>7�"�siR��ˌz�)%�q�x���8���6p�$��H�4�,H���p"w<U�a�&mLQXF�fQ�f�x��$��g���h�^� D���axVS�U9T8�VG�P�ð�_����U	�`�S$���`��5<y����g�T�u,ׅ) [?q:O_��w�8ܼ�컿�?�鱏���p��
,d��~x��קa�Е�Q�vs*�L���6!�(�=���O���t�Z!,��t��d�<7���]�qY��V� ��2�(��vVH�1m�4?m�a'}v�W@��<[���W��� �Y<g.�!����B!I�"gyqQ\����d.�̇4���׍zݴ�,5@�<�Ӵ9b�&i��z�
:����Sr9P�\��4�˜ђ9�J#f��:��"��xHH!��R0Ad����kg�:�(��-��A�`z2$��a�B�L`F4����(3'�>>1
Lh	�	�E	Ԩt,��HI*WG���f��'��<]'W"�>zН��^��Ϟ���)7����D4�F����Y�$�� ���x:.��Vm�� �{ۃ�x��^��x�G�tnUѽriM4�]�I(���}�Z6������X�o�!,��-W`�?��\<r�[.~�A՗�+�\Ȏ�XBm?=����'���� "gQ�8�<OP}�|nO<��|'o�q	{�T�O:-/*WG����%�dmYj�ms&I�yE� x$�2P	�c�ά�� �5�m���4C���̲��I���(Y&�  �l3�-�a];�+���\�Y�*4߇&����}g�z��YV���.<�b�5��NUt�DUӡFmx�T���4��Dlmj(��re�r��mq0#**|�0��,$���D�yo�9���K�5��	�E�d2�<�3yI�[�T᪇
K�1�0t�'$�FF���E(����|���`���i*A�Ak��,����~y�)MX�	K�Y�rK&�3K�\ՉL������� <X����o�	����S`�.4Ӄf9x��G��� C�L���x�ۮ����+��vn�z�����S?���q���n��oq�Si�� ]�^���I��RxrX���"��Gp৏��{K}	�  �,ՃOL�,�|¬�o��u��ہ�;���F@����}@W58��*ɰ&<k_r��j�5��!�0\��B��I��0|�kA�e�d��C1�Py�JӢ��"�$�(P�M����H��4���y�˷86��붃FȊHj}(�eՊ]���p�<�U���2�����ԭ%u��@����j	H��R̀%��p�އ����%��肄͚WM讏FY�>�o�<�'��P2��J	VB��N"�Yj&�$	)R�skH�2�����I�6�Ēn4w�a� ^���@���hI�p�3�i����3]�hF��J���?��T����Ia�#�������c}WJ�wH��l��۴[�~��S���X����Ix�������Y Z�I�õ����'�5d1!���{�W���z��J^��oZ�@�?�C?Z�ʷ*�Ψ�2��|x�2��	X�1�����cY ���6~b�#���y�yֱ>s�I[�&�S��6yG�9���l�
U{ɤ���IF�2���z[��F��$rNU���E=�jkG��(���i���]˗"ӐfW-Ѳ1t�}Ͼ�Ŧ��/@ѓ(r�RהF��Ӱj˙@K�̹M��]߃���^����A��c������jB��I�c�j>���$d�@��!+Ш�1��o��T2onA��t��a����h�DȆ��ABŤm"��ɕ�H-�DcgM�MeuYF2�CU��`�N�؎�(>�6IE��B�]j�c>
���-�г~-&��`ߋ/A�*�3�As�wA�"BF^�1��иa=V_p.�n�<�v?�,j6�� )�e��S z�D��Q�<R�㬺��g��`�C��g3��Ix4�N�vt�a� �b�`�
�z�"0D�n���`I+�5�R@�j�"���Al�����@sJ�kX܆��	\p���%4��+�κ�n��}��h��߅X ����.1�߅{�"رC9�箄Y�NJ�z��NT*�\D���x~�sx�c)D4p���^����z�ц}Ϲ��v�y�i͝A�βXl$,��X�Dls6@a�5����t�S	�/؊�K/�@&�![6JŔ +@���P�^O ����L��������'Qx�Udl����y�ۛ����uѹ���@@�{�3%~�4[��a0t��c/�0^B���
2�_r!z���MX#���cl�kp���&�HR_��J4yE���r�_�	�=^ω1<��"�� ����UE�^\r��5+��,�k!r1�����ȡ1    IDATWKEy���g?v?��͐�8�E�4Q�fp�'/E��[�%]@.������O ]2�H��[.��V^�e�l�3��>�Z������=��O?�Vb���$�C!@�h�[Rؤ�\γ��Տ�������+���Åu��ըt��ć�T%����+p�m� XցQ��Q� A1}4
*~��Wx�_�7t'@k2�48���)���R)�ө:��v��_�����~�>�+� �����O�'^�Y�NB��S	X<��
�B��0v��}��`)$dI�;2��Yvߊ�Xo�I�)���"���2�:o�Qٝ6hG"u/`D�����k��gFJ*2��Ry@Y1������̪#6����U�
F���Xs��a�~��8��(&�{�`���벋��*E�-�{�Ě��"T*�2���F���c8��9��yH%�(B[ك�o�X�<&j6�?��?y ��|���VY�躰E���T[o�2�+/�2ρ@����q�_a�3�3}��MX���]���|�i�vd���B75�`���i���;��O<���o@,Uay>ο��?EG#�J���c�=�cj�Nt�@� �
�%��#
�����O�*�҉4�w/����K$Y�㠅�lX�.�aa�(����H���:	���͓���tR��C3�1�P(@�ҼO:٠��)��Ÿ�ί��bRP��	"A�\4I
�^~?����f�-��g�p�G�԰��AnoG5�ya��o?�/. ��x?~7.}�ߍU��#��K��Jv��$euy�;<i��&� �`�=�?0�%��e���3�z�����|KP_�|����|*�m��p,�3�z
�Fޢ.�~�g�-��i���&-NZ�%�m	I�.���G*A{���)+tlh.�H���xv�v������
���te���T��DZ��
k"�@��@K�81���>�W�x��Fl��J�����Ċ�֐�]>�8v��,6�b��������Պ����Mk1�ָ'.����<z�O��vՍ�C;m�I�Z�ôض˙� ��Y��RUYW���i�_���O����r�\��/��@F�Dq
���v1�̋x�������#+�,��a���O�B�ӑ��G/A�*2ql������EK�B� 44q@�����X�4������ȃ~�*e�T�|�')����a��D�~�R����@���ȝ)	��$L67��o�q�j�UUQ�M�G�B��c|?���߁7UB3������ٗ_���D��sϽ�n;�!�JN�Y�@?En��N㽮����W���uM]!����4 �M�����ϑ+��X%�M+��IsѤ�2����Q����f������7��'[�1��7:٘����զ�U�1�6 Q5L�y/���O]	��nk3,���dx��jJ�%�!���˺�Lbm([�,gZTM�B�ܶ���8lǄ�܈��7p�|�j�� �>t��r��&(�l]��		E����l�\��q�ΥK�wv _�3�ڶjh�=T���?�1�1,�Ed	xE��wI7�����^�l�B�x� (U`RP�ʠ���[�Z	�[���l� �̰'�J���qY@"�1��5	s|{v�Foo/ږ��i�<�e{t�6���ځC̍�y�H
TÁ�)<��p����
 �u�Y.2���~}�OP�u �T�~��K}�p>������S{����������${������ٲ�o����D���H^�kj���_����b*���DP~�@��Q��������c�hR��� �c ݜF��k�l�f������n��m�z�ގN�S;����B�/�����-�����~�%�ص�mH���'�Gr�qdŝ{p觏 3^@���-*�У������^���x�?z�q����W��'SZ+��I�!I���4�^�pښQ�%�I�ؐ�ӒR
dI��s�xq=Ȯ s� w� �Zc&7��GeS1@sS�+{i�e�c�L�^������;�*j���-�����P����E�+*�����X�\��� wtb��l���=��_>�Ş��w4_�#��e���� V-C�@V�o���
��P4��Q�r�|��Z��b�s���	HJ	,I���S�KS"���!�ˡ���R1�;<ǇD�^�
�� ^��A�G��,�!��,�g#X���5���>�����ZՀ82����
/��E>��W����e9�H���"�۹Oy,;[@��҆��=��{����6��y|�����d
g|�z4��E�%�($u�J	�Cyh?��a���R.`�5dZ�Xq�&t�[�!�ߙݸ��O~��]��N�pV�x_ �~1���y4���_<��1��1��%@w�OL�>:����q�އ��,���f�P r�"
�]�fo��8��M���N�������deIFA����!vw�QA�������!���2��B�K�bA�X0����ރhl̢�����h_܍���Q8�2�����P� ��*����,AkiBbQ��Ȫ
��|6�ф�/6cE�.�|x����e�|�O<�Ʋ�,���b��u�b�s��W-E���I���6�&IH��d՚	�r ��(r��M�5�C�:Rj�{�r2Q� &�0�}t55��d��̤`�};���
ġ��!8�nH�m�"�h`C=m��y����$@�}�"��	L�|Gm5]�����p��m ��\b�����7�FNp� ��.��DZ�1�%�����oD�U� ��0��^���/�xt����c�o��1�aXh+�:���`JQw��q�W/���9uv��3�0�����E���3+�M�F�j�N��HT�wLhF��8����� ret��le*�ŀζ%u��o�u����:ˬNo�a��l��xdM��5� Xt�&4�Z��(bԬAhh��քĊn�m�.>�Lm���*��w�_{�d
��_�20V���ڌ��7����<7ϥ��6&�8�k��4��#p��#�cə�u�B��<.8/����Ks�΁��(�K�j�8�ĳHC08�FY�ypt�l��`E�� C 74��,h*�Q�>$�TQ�Gul�D)�Pe�Ka���_�uBR��i�=O�R��uj��D6��aBp}�4W_���N���g������N�8
�3��ۿ�ta�*���J�y�<0<��(���Z��tg:��Q�u�=�������܀r���w��D�x����XO
�ߨ"��&K����v�GF��*%�X��nk��=0��wv�{�W���m%���f�>]�)���{�P�~�x�X���5�W�r��@���(r�y}?�9��U�X�l�xr��=��&Bs{��]I}f�VW�V�N���}Z�sЉ�Db)� @���4���y�r�Ǩ��ф�+���_U�$5*�6-(n�ʱ�#y�c9�GF�����u�TVI%���-�3:jP��yV�2���q���/�4r>>�ǔi`�E�y�r� ��0�r "��{�L�{�X�7p-$]�}}z�Edsp��	3Y�ҵ�~6}�f8K:QD�a�VXu��!�Z(IK";�	?_���>8�9�����ЄJ��J�%�@����' �S�Bfa4hhX�ʭ
ۡ
���x�/�+��������9��(�~��c��������_�3����P�^�w|ޑA��At8:!0�ˑ�{�C��?;s�Mz,�;-<�N�=����8C�R��Q��(
�]�i���e��F�5h�����'��x���H8Z%��e�I��υ�؂r:��k빷��կ���{��yow����]�S�n�{��C��i���>���(��A*W��}��8��h-�So7f�f1�(�i�g�� z���\q�i��yz��Μ��>Μ�F:���I����4�N�dKO;^6�1�C�IGv�*4�[W�XI�#xہP�Q=>�d��L�ő�{�!8U�[��Y���+Q�T(�iT���	���	XC�r4��X��|�́Ś����M(fTe2űC�tEbgKa/��xvY�(�*�<r/����!��C�l.������/�hˢ
U��=��K�	TBW4�]׈@૔jp�&��^��@��FER
$��T
��Vt�ry($�NCjj@zY�fnB�GNb��B��d��?{o<����`>��l��X}ť�e����	i�SU�P�w|������O����~3��YxS� z}p?��=tt��	�^y���ET�**�0G�*�J^��G�}{"��:4~�BoJ��.��މ� ;�7o��ү����{��}䏾 ��[<������^���TB�H���G�{	���J��J�(��E"1��+�]��͸O���}}=�ǀ�L�
�)�&-�t�ԢS#�2;y%t-�74@h��-ȧT4l\���6�ḭ
�|ǅl{0GP;x���GO�E�P-�q�R��o@�E[��]T)��m�4/W0u��=�\���GQ�](MMh[���0���@����=�.��l�Du��UD�<ԑIT���뽰�C�mnTm�mAﭟG�Q�������4�R���CMp[!�E$<��$��
��t�(t��11z��{���ۋt�2�F'�/�P#=��ft��
bG#l]f=w_�x�M�,����(�_�$mOpKU���&�ڶ��L���dۅT�@<1�U�?�6�Bg @w(,���� �dx}�f��o�9���zR\�#M�j|o�4��	ЩC@3� ��߂ӿ�eTS(� �Z6�|�U����?x�J)��oh/������j��o=��o.H�~`��G�V� ����0)������ߥ�D/YW����F_�5���΀�HP��;�~��dF�>���qx}��y.ʞBG��l;����_����<tm�ԇ�V�cS���ܲ(�F����'P�$�}��Xy��:P�s�.mʥ2e�=��{�� ���@���?6�x-J���k��J �/��w���@˗P:|N�OԀLhk�ew�
w���p]��i�F��m�p��Q����@m�AtO�ٹ)��Ieu��_���
CQ`�yJ���|2|!�62�Q�U�by�F�0��=8��a���j��Y<�F����.�߲�G�
Uy�C�ф�3�#��Ì������Lh0j4�Z�D�ö���H�k�=�Fɱ��x"=sDӂP(A�Be��?�$��Ut�3�N��_��<�R=ɯ��X��/���k�z��.� � �2�1I���tl��WPjL�@�,	��Tr���q����UI eyܒQ3
�m;eM��t�+K.��M�}q�?�m�C}����}���S�X��=����t�(�\�M���I���<��M�Ǉ�D���)[
=�	H�!���It�˿Ʋ�4{����1����ai��B@��%�V������1߉�/(\�}f �ȩ�5Kp�-7������k*!�ۼ�I��cط�)��G�8�.�����\�_�S��:��E�D�P@��a��x��P�&�U�i��;p��lX�Q��
n4�E�$�ȢYC%��g@�>�^݅�����P=ti%��٨H
�^~1�����:,U�ᇊ�1��X�D=����L�D'^܁���m��&ID�Hh�Ś�$��mnA������$��l=K�݊��@��wI5�y�L~|)IDJӠI2�G�r &�(l�Rw���r����p|�}r
�EI2ɡ��m�{zo�xb��P��E�?�[��W%�{��Þ|��F����$/L�^I}PF�[����c�*��/�LA�w��������v9���zs�7o��ց���{��xˆnz�{�����Sm �T�#���0).w�ӮQ���tz)�d�4�b� �L����������# ���x� �6M�8랤���/��A-�0��N�r�d��[���n�!��M:��X���>�լ� 9IB�r	���e��𮬲u���0������ǡ����lK:	ko�V^�)T� 5ʖ	�L�Bc���#O<	m<�lAj2&}�G�.��w�z1�����TI�M�L�S�cD��F����ӯ�96�%iY5UG����}��(�UؚWa��\�tB�r'w��LN�0��u�z����9P*�;$IA�DqDZ	5?@Y&� �]�	l��u�%uTABc+V*���:e��ź TȊJPQN��=$�)�=��5R��� *oD��_��:}0)N�k�"M��;=�1�GD��gj^N�o�<�����;e�ò��W\�e_�S2P%�\
x)�#���1<��ѷ����6��YK7�eq�!J�;��/��_<�>��/|�Gp �#xS��%)n��j�2�팮��	e��
����y��j6�a�i�$����w:~6W�#.���;���i�'�����ķ�K�j����^���V� �ǯL�\'��}�KlVB%k�X�&ن��$����Ǡ���F����Q�ƪ�>��WՔ�gd��y���>�v�� �� ���� �D������o�{18���e��@�u6��03ulB��%��qT^y��!$�}������_�,�-YX�ģe��Φ+�VB$�{�D�#Ӕ��N<�v���=M���|Z�^ WV�)�V��b�6�s��8��FE�P�m.�����iá)��C�b׋�-��9x=��+R��˜V5�=���^GߣOb	D$S���_���n�=3s'/N�[@�nMd�Z��)���'�I���Uh��3ȋ>�dDm)
�*5����đ��Ь(hU�լ�e�N�����w��\|�]��������V�d+� ����Y^q�p���蚲��'(4��Gr~�%����}	i�<ؑk��M�G����1э����Cr�L6�� y�mx�R{�Z���̔ܧ��ĸ~`}��&���̹������/AڸՆ4,�2k�U4�=8�����:)��.V]{�|�
XI%%dr+��L���O>�Ï>��E�C�"LI�8��.��Ew�	�_�1�fc�PR�g�.MT��
k��5R_:8��WQ�׏�\�{�"E����I����.��/_�Jk�3E��!�W���u�&�4�.r0��.Z�&��?�C�>�&�Dk࡝�sU	~��π����*܄�)�����Æ;nA9�@٨A&����3,T�r(N�8S�d2\y��ek6���%��T	��B��+�*0<
��a�{�14�X,+a�N#���q8G�����{��K�'�O56`ݍ�A��b��T� A˄W,�6<����'8z` ��&�c��f4,�|:��W�@���q�9߸�O��ɏ�v�p���
, �����Cp�<�i�1�6�*���ǁb� O�ĳ/���G�@�3x��J�ă�r��g���|kL%���t\b���9i�S�L�й�?MfÞ5���G���]=k#*YX�{MYV��F5��v?���h%r����u�%Xsõ0�:��*�' ���zG}������!J���h�\����Y�q�`�t2� �*( on]%��Q3*h�TL8Ȁ��a��]HzMFEP�����s�ULΪ�>�v�E\N�����B.T�����TǞ~����-'hu=!��!@�UL�6L��e	�׬E�\���LY,�`.��;QL�(�d�o7,U�����)�5LL��2i,?m=��,UF����0YaN��s��x�Q�rytݱ��2a���c����Uf�ꟛ���9,��]�f���E�Nүl����x�I��H�T9�-x�"��~�?��G���4M䤂�7�k���OXt�E�]������^�pާ�
, ��q>��H�Gw^����S���u,��jG�0�̋x�Y�Nd�P�5,��g�q�_�t�{V�3�i���b9���#L    IDATV��m}N$n�3�.��k�=3���rTQ&�<��@��[o��YQHꨑ���B�Tፎ����Avx
�
*�S �ܺg�&8�M�����0��KU}�������L*�S.e��u�p�� ��a�3C�3�{�k�
��"���PKe؇�b��w��$J\ I���|
�����*$�����{k�sŝihČ$U]m0�s7�����M@^1ќH�hZ�Si$���jiDǊ(U�8�߇�'��}�*\~��0u���. f��pL��N�t�F>��|ɵ�&Tt��eG9!����2�y�R�?4�,�?��%w��y�rF0b>2��U~�Vu�y�s�}��Hz+@���p&��q+��Ę,��y��I�b�|t?��{0rl��Z�$�,�D,?c#֜>�k�>Ɋۮ����d#X�Џ�
, ���VNg���E�H���^���Li�%D�"@'sʔr����?�N�F7�ܹ;�cp�3�7m����)y�o(�9S��������^]��7�ý]��.��g�Vb>�+	��jW'��~�3�@��_�)S�_*��w��>�(G�fr�>.؊M7�����r�^�]�Z>�{�-U��tBøicB�=s.��&�D�㒻�sa�c� A������0F&�r�=�x�ߋ���h�E��;���_��O^�BCU���>g��Ӗh$�diU"� ������?}�h=P@zR�P�]��:V\r:��tv0����ӿ�%�����W�f(�Wl2X1<c8#S��oҼ��:�Z��@k�"�C@Huϰ�Tkp��@q�~����v}�ӹ��h\��1���%rg������M�U����" �ފ���Ƶ�$R�#)��F�d@Ϗ�Ь�!�����8s#V�w,��������Ͽz�w�M^x�{�����^���s��v�>/8��9:�;U�?z����j�*��R�m�����p���BN*�4���ǀ^��6�#@��r�#�K��P���:g�Q�N�i�{���&-�'�gϣ:��@�ne(�	0����$��َm��
q��	����~4��7t8:�}�lGz8�V2��ϥ����x�K1x�s  �'�����Ο=u2��GC*��m��аx�Y��/�jJ��Kni������6���ƴ1�w]�<j���oǞ_=��eC�%d:�q�M7"�e�����y��Qi��Fi>ZU (Ta��v@����=�8�_{5˚Z��5�ށC����+.��f�d��~���h]ԎM�WWPp�ϓ�*&��O��w]r
v���mrcfJC���PZ�`(;±~�Y�\�AG����Уh��袱u7�ç*{��M��Tk��<�s�h�c����q�����!�g�$ck�A �Ť,�^�g�~3��0F�9׶��.䪉��}������Z�$tr�!1�������~�V�/.^��[��?���m��Z�@��V��\�Z߱�$���TM�!�&��Z3��Mb��x����F��MN\���:�N�8��A����f���!���$�F��X�e3	������R���I�Y�c��e��\?�9�ʣZh\%��2B�f%I`@/��ಯ�	�����%��vLR~
��(��GGb��V"�9>�k�c�u�����t
'����hM$!K(��ԑ$H�NVP�|Լ KO?]�֠�P,x��~�R�D�Lg�"B�T�z��2������;���8��zׯC��RW�P&Id�y�4x�4]�c���"q�;��@1x�۽� �s\l��Bx�$�=]@cj�����*�J��%&I����lVـdXFs8��\�Ш#��ъ���^S�d5�8ص2�j�R	����ᇶ�!_Bw s#�sF�})>��<����fg=k̥�ið�@�����C���2��1ْ�(�>���5��#�8A�	E���[�vW#r�_������l	{��?��s,�r�#�d߁��p��Ȭ\�����.�r�����@�{��ŏ�_����Щ�q��}��W<�/�D��#�T�2<���~��?�9����e�$q�#mpQ�C�<OQ=~Κ�t����<s�%�G�hl��siiZ���8J��ۈ�Onf��śxݢ��+ZS��;�Įk���Z{;.��m��5(>,Uf�T{dޱc�a�/�>YE�JD-��Y���o��03I�5�� ��P<��-@��-�B�i$���
�n	�c@0=Ԋ=UM���;�.M%��"|��Nm���#�&X$�E�ӛ�a�X�y�RA@e|ÄY������ MdÚl6�j H��:1��}>��wζs�lk��J�����R��Z��L2�3�7&آ5�T��}HU��&v���'�X���g�َ���ukQ"Ec!�ٸ���T��~�����5,��u@ +�o����!l�D�ܠ�����d�N�=Ǌ:5U(k'@'��z@��@��"�<m%��������|��J������c��a��߅3^@�"#��'�`�%@�Y���ʮ5]~��w~s穴?,�ˇo ��w�޵3&@/�?|��Z�L&�H���P,3)n���p�_��@nk(3北fmC@w�򢯘�Vw�1��z PٞJ��^��0S�2dp�PU���2�bu8��w���%��̽�?^XH����9w��_�i�K���PJeT�6<����e���T�����	���r����1��Ybc���!A6����n�t�:DY���(� ��l�*�c8Ї��6�X���r/!�ʀ�H�B�"�y2��a;����<ͯ���B���c(�O"�����-�C$w7I���`+!^�\�e!I2`� ��)��=X�Ƕ�2�8Y�Q��1������(����� �*��#;^E���p�^�8�9�Oa�UW�QT��p�<� �e�9�G��G?C����ć�<t좢x}��d����L��A@��ӴA4u��	Rf��|�������Ms(C7� Ê m�l��&X�inu؁%���+P,'�p�d	���W���z�ւZ*��i�_qǪ������r/�c��+�I�bp�E�92y���i�R�?�W�Iq�/���0�K&�d��ن��(���E�^�	�o�'c�z=)�z�蜡GO&U���"0P�a��A@�/��G�H|N�a��e@�nv�b��7�6������j��>�&��'.O�8��\#Vz��"���uX�m+�E��u����	�T2\/�<�]d�B�wQA�K�-f��Z��r1:p�X��å�ds#Ԧ,
~�j�U�T؆	E�x������it�,ո��WL� !i���B�6��t��Q	,�'ѹd12z���]�iM&t���1Tb' % ���(�Q��Ѻ��"�O� 

Wo���|��򯿁�WwB*��T�	��z�=[����EY�#S�����ơ�Mb���N�C�����y"�����e�s_���� O�v��J��$��/<Z�:R�(J���	ID�5Wa�篅�QP�&őg�;Q�UF�p�w�?�y4Id'���x��Z��47������<�37��(�7��ޯ��
����,|�o�4���s��Y�(�R*��H�,��I�>�
^����Y��TT�p(Ks��s�%�Y��Y�y����ǎh��@d��P	؉LE:�t9���O��Iz��)�db)Ku�2�t�g�ܺ�����E.��q�Cǡ��8��SЋet�	(��-Tv72i,;o�ս�P�q,0U�@U!`�2��@�@�1�C�FC����X޹�)�'&��u.E��Y�DKjX��%�=�
p�,±�?p�K�Fϲ�jp
dE~�Dq"�Ʀ&Xİ�U�ۚaP�)QU�)	�0PSX�ݬ�$S��BbY��������TjC��V����(2Q�<:	�j"�ˣ��g�>���[��}���p�u��o�@����nVP9i2���k?~ �e��˾�A^Ȥ?n^�t~��.����~v�����)��< �v��@!M� ��#��?7�AY²>�E��4�I%9T�i�`��\Cub?���9����`�a�N`ӥ�om������r��ο�����f[x�V`�?��۔D��c;�Q<�ojb)�+#��{P�
�7x�{?B{�@��!�y�U"@w��J����N�5��yq���EO{i|)�wqY�1Y���v����@�n�P̦���K�ݶ��5�Ev���$��Q�?�<RU���}]1"����Cj�
�M�a�4T]�,"�Ͱ��Q�!�]4g!C�/a*M�|7�@4�=��vzoW�8	5���@2����JL��\Psm�m�4��ï�(��#�AWc�:�5e!�u�R ���I�[�t��p;����P�N�%8�*`Y�"���gq7ʦ��d�J�lpqd�?{�$�u��>�'�l�Xl�"�L0ILJT�"-K��O�-J���{�W���u��mYV�,��]�,۲iKV"�$��H����;;y:�zO�����]�+��ΰX f:�>}�7<��ƊE@��_?����LYO�����Ng���V�����ܽ��1D1:��1<��_���d��9({
A^���\�Ӹ́j��8�S��?���:s>V��LП�؇z���yE��~�y����i��DÆ�*@)8}�%��wM32��+�a5�{�~�YU{�{��[����#/G�{�͏@��c��=�<�N!��������h$�OJf���X"ĸ~������JWB�
M����\h1����!��T��=�=6;����N���3�D�k�x�k����D�"�HE��ر]�v��a,������ڠ���i�z�I�8,q�+���(���uE��f�z{a��ԋ(:z�WBSTL�O�|voW7#�e39d�9�65�L�YǱ�+`zt1�Z���6#OL����O40@�4R�.N6��P��r��	�DV2��{��f��=���$���]?��Y�KcJ޼i1���e#�36I R�G�%u�b���.� ��ĺ�kX�V�@�B�!]/��d��$��N?�8RG��WVqE�6����D�|-"����5L�s���՜@�L~�������us@�]�8�/���{�CFC�1��N��xgгܺ7Gɐ"����₪`ӭ�BǍ�#%۬2�!�.�tJ��g~� ��}��&�C��������{7�َ	Az�wϞ?���O>��{�oW�j#P�e</��~�w	�����@DQYN\44��|�<��?�=~�E]D�2�lqe9l��g>���t�Y���y��f���i��N��@���Ԏs1�μ������� 1����еm��Vd,����nhD�61s�Nx]��0I��K��M��"1�흐�;ѹn�hČ��������051���Q��CS4���,F&�14�� }�����䡋T�]@k�
D;;бv���Ίf��,jA��|.%�"�h@&�����J4�UR��8�z��NL���E�^���Í�,:Q4,L%gY[S��m]ЩS��Z�AO�a
X�����䩣�e	�mmhk'O݀A�2��ƨ���(ZMG�5"�t"�Զ@.Ҫ��]�!vv!�;�t狅,��ۨ�۹s8��#��:+��(���	����m.͘J�>�Jc� ��:s���g�}�jX	��{�N�VA1��Q����!q��0s({ݴ���;���L�������bX��2KK�X1o����}�v^\���[w~𖺇���㥸�:�/�(^�� -�ӓ'ߓ��ʮ���N�aO͠)��џ���{��Vǁ�j�=�9���C�B�|:[�} g�A�ā�Ҷ\ ��)�^_l�a5���cu�s�3��<��|5��}�:؉;�03�����)>3�Ybk�h�D��my�4)�j�
l5
����}�tv�m�c,�d޳���ڊǎB%$��Y�Ξ�[4�ZkP������brDC�@��F�V� ��]Ӑ�,��J��Zr2V�`�WZ�c
w+1}�4�O�Ffz�L
��V�F�@/�׬F2K@��:�{NV��Sӳ̫n"��b3."����lŁ瞁a�Ʊ~�fF˘y��^#��ؑ#�x�0�^�%���eaV ��ֵ� uu�y�J�{�8�|N:7�B��y(�<�E��w��>t��;t}�µ�_0BS9W����8/��=�x�aerT~��������5�p����ׯŴ`��K�6���tq������܏� Dd�K��&lQ�|�7����q�iÖ[�}�,�շ��@���2����������_mZ�v���	,DT���@5����ёqt��y+��6���V��j����9���ʂ����:Wzc=�7գ��I^�`��ʓ��X�w�("C^Z,�����Bi�`�m"�)�	}r�y���h�s�g|�^:���)�	\���4�#�م��I� ET�����n��(z�;�Mf`gs�֓)�f�gҌ��(*�h���X3�Ěa �aj6�$���2Z[�k6�+d�:6�ښ���(N�@�呿0��W^�D��$�H%�2��݉�W���45blf��<Q��� ��2�PMj�jM#55��(&�G1;3�\����>�Z����JN�v-�F��F�E�$\��=A�Q���,!�щ��A�R[R��Y~9=6���g�OO�2�"
n��6��˟{8���dB޹'K�	�ЇRৢ͋'@�2b	�d�PtɆ1؏k>w;��ȒQ���3a��,�L��� ^|�I�EQ5V�M@Q��Mנ}�z��6n�t��|��W�����@١��Ų��O�;��G����s�+��o؀t1�V0+�E$�E��8����y�8z �UVX�gZ�(dY+?]�`;kotڒ{G^IR���& �:��+տ*�	�;���`lq��SYkY9 ���VL�̲�2"�gf�d3���*P��r�)y�,h�`A��qE�z�16���@����T
�x�y�D@t�|��$��$�:�Q��ڜ��u[��xg:׬B�������n_�B��\J?�p�cv��."3rb:Î���t��͘�t=$�c$�����R,��n �h��7�}��<̙₈�sg�d3(�Y��I����݃}pE�Sc0�y�����8��Dk4ߘ"�*����vȝݐ�H�L��rr|��q����h�n0/����&�y�m.#J%�;�a��2����z'R�҇
!��F�k`���yE�bDz�t56��-�4�Q$��@!�e���,"9���8w�Dۂ�)L��`ِ�*z7l@��hX��`���u@�Ŀ�����Mel�<���v��	ǟz������ʝWo��J�9�"��YD�9$Fgp���Fn���4��$����J�b����_w����t����(�����燕�v��ЫIQ�S��0 D58t�M��L������D<��{�����e���u�.����b�����(UC!_@�2ID!P��\v�����E�Ү�ʸ6���
Si�R"�1}�ƮNH�t�R*��� 
h�l
F6cfى)$H���n�x6��k���r�y)'A[O���1�I#��"�D���=���#��D���i��LJ�rV����Z��L'9����72jj��(Dk$���4�1��L�8N��ƀ�ܨ4Ma)�r�8���k!vΝ�e8��݋�{�d�9��-���"aLfZ����B�u�#-��0W(�*��y8��hue������^H��FΤ�Fj�kVy�><�B�����u���.��@З��8}���xd�]���_Z=�z芫�d5�Y�ϝ˲N\��$^��/0z���,�dD]�-��Jq��d�Z��E�{�v���Z�qX������ee`TCL�w@�]Ȋ�l(�푧l(L�0U]    IDAT��$V,��j=�X�,��X�"lR?#�c��B�J�����	ޱ�晩ߑ޺ y0"%Rn�<HYf9�ez-QU�,�����T�L��:L#��;NJp����uY��ȅ\;��=�3b�g�y�Ѧ&��y��5As�N�@jv��̣Y��@V�$-�a�Y0u(��Z�J
Dꩮ(p*�I��ݗc���4�M�	��]+yͱ��$�uj�C�����L�+3��IR��Ci�9�	5�	�w��Iƚ)E¨8kV���
�Fr�΄xT�ȍM�8?��h�����G���8E��'�Q����hܸf[���[w�v�'�h��▩��e�UoV�W=t���T��:���<�W��mCW\s-�x�F�|�1�;R���?��߃~HX�D �la'��1��jD�j8��D���*����v7y��N؁5x�!d�(,�j��	���Ɣ��m"�{�z"�_&;ѓ"����0t��mCt��mC@��>�7�z~��+�㫬a��x0E���|�!�]
��2����r�$Cr���3��4r����V%@�eOޕ�G�*����[���=r�ɋ�Zk�`�޳�:t�T�T�]̳C4�2BǁQ`)���4Qa�""(윬��iܹ,�Pj�#R4Cf=T�F
����^e�'��u���%���R�a�O�7��F0$Oc�}<���������:"�hH*.(@�5�����'�H��fuPo�Թ��3�T<���q��#L����I�.����W�Ct����];w~��?������|]��B������4#@���wz�ѿ�)сko���2��[EDu+�6N��>�����V�����$(�(_�"�3/�������.&�.��|�=�U����k;��([ңwH�X��;�;��0>��L�@� �W�L��D�#����0���$C�)���`1�W�~>�7�J��4-#ky�?ʻL�I `�H݌�R��6�@gY�3�ZYd��t|&�#y�[(jN�%�XQ���:���ԧ�cF�I�*$�c���m������^�5ԑ�����4�+��җ���j)�Cw϶��Te�w�1|)_����N��H	��ǧ�ĒN�����Z��}ɰ)MV>����?�(zBbѓ�AJ�Y���"�&`�ކ����W2pYn�H!�L��i$�6�T����B��3�T���z�o��J���H5��o���n��٥y��GY�#P����i�:qB?��m/<���C7��m�b&23^{͢�C�؃O��܉�d]���k#"��M�����9��x����.��%�� ro�����QD�7���4� :�/���I��<5�!�+%�����j!!&���!dt��<,y��
�B�'�(i{
j�>�TG�2�J�#���|�{��N���m��'o��g�����>dD�ƽM�UE
�SV���(gZ�^�6��b,2\���X�"3@�MR��m�3�!SU�q���P�ix�\��F۱��tq�W@ HƖE)_����:�4c�+"L�a!|�Ż�w���U���ąH��n���ά/�O2��� ���s}����e6l���C��`�I ICƶ�R\�����B��71o;E`튌���Y�Eb(��=?�X�,���z�&39��(6�ۋ��R<кq�mW~��:����vsu@�M��ߐ����d~����?���lz;7]�h{#���\!�u������7��S貀�£�GX�=uB�����恭�+�$�����&� (yP��)�{�-��i�Z�}Gyɒg*Wc�f���&C�=��4��P�3\���ׯ�Z���m�C����}����l�ؽ�G2"�������7.��S~�\�����xAT���7��`�2�X��KIpa���{<|^�d�y3�'\��F��<	�d��j/���ldꃾ`QМ������:��J���ywH#�J���"oژ&cdh�>�(��bڦ2@v�:����ˣWS�����7������(��ӱU	��섲�BO�3��\}����{�[�G`��}�
��i�~��3������6^}�u���fr���by������S���!��!����0����#���',��g���GL�"�N:�|�� �{ ,��5͜��GF^s6k<� �{��Ç?�K!�@)�3�)��^�W��q�|�j��j5��K�@Lp g�g?�_J�v�
{�����7xB�J8�\�<����W���B���v5�i�W,́��mU�#���*��<��|k��g�}�����lF^�r4"8R��Ӯ{�ۿ�)`�JL�:�Q�seL;���sh��(���G�S��;���(1�z7&c���h߰�k�>��[�'[���C�x9����@З`/�C�����{����}���r�o�C�F�zk�F��b������D�D=�������(���� t
�za�rY��^�Hb���H�{�A�{��Sb1��e�0N�
��Z��򺾗Xн��@�!�ۧ�'�� ��^��6(@T	�6�U"�A@������}��`� <�t�9���-Ы]%+=�S>�γ��+c5���q<q�K�)����j�T8k������]ټ�� �-$O���L���/���s�9I�� �q桻�6�ۋ�{� :8��3���u7���/n:ַ�1u@_�S�ĉ������ξ������_�����ѣ�-�P��$�oC��t�"����=|� �=C>�#�eE�������6����^���B�{����s�� �T[�Qx+J��~h;��'p��Ϲ�20������x� ��%n���9���D&�. ��"���ju�<�Aǟ�Ҁ�]������+'�X�%�e1LLc�m��^JQ	��r�	�)eB��+`R��y����#�gt�)�.����i�uc/��O=Y��6Ht�d�]9�J�T��b7��N�--Ϸ���'7����_�0�w��@iꀾ�'��'��j�^�������_=���a���0�}R� ]�a�"E�1�G�xÐ�T����N�]��� ���y
\<��ղ?0y�}�C���=@�$�7���a@�-Z� �	�x`䉁�� a������祹7�N���C�(C�U��-��U�+���׺�T����׹��/A���V@w���7ea� �Vܛ�&������i!�Ӂ��|MW�¬*"]�BvEYJƄ0�D��9����^aM|ÂN:$&1��"����;��ix-I��غ}����۞X��Q�֗`ꀾ�x�����1��7?����ϭ,���'>��o�YM@VX-u����Ň���/:.:&�����P�ܷ����D��i>@�!�0)�Ȱ2%���3P�-��t�2Y��=� ����>^o�J�n�17���J	�&X3�^vW�u;�<�)=����{X3�j��c8X��s��z��ʽ�Wr���WsO����:&�:e��1'(� �����?�}�]m�4�ЍD݂1�g|����ԩW��/�J����ۆ����u�K�_q1�}Z��A�|Y^5��n����u-�_��h��	D���;z��ӎ�'����w=����+G�ZA�Jo~�۰�#�GF��E�l�E$R�GO���S�q��J�(�NzM@/����zЃ9]�8�<Zs�Q����K�)/�]�� M�S�x���R߯�+xL��WΛs����áv�3�� ��x�;Ѐ��7�t��R���Jx�3�k��ݻ�ꆚw�*�x���>�^��˒�,��� "��� a��	�?�Q4��:貄�B�	�8���)�3���4�����fSL��0L�l  bϫ.��mÊ��!��<����M��̃��u�~�����}v���	�[�������׏<q�7�E���+p�'oA�A�,	��Ģ�hHf�����/`��#7)c1�q�d��s���A�[��E���y�����`����B����}���� I8DO�-���^���+�=L�z�ۗ�����H�a@�����Jq��Z�^�(�A�t=�:;~�`X=��8��_�z-�|�j�X�*��9�sJ� <���ч�rݑ\9A¬�"�ۉ=�`�*��"U,��ga�����ӈ$ӈd�8p��9h���� c��i?tS�vlE���HE�/E7n���?���;����G���}ϋ���]g�x�W���W�y�?�j�����a�%0��0f��FhN�q၇��O~�A�E�a�NZ�/��HJs<M4�u�:�r`�QE���ja�px�DH�i|/��V���bTq���\��@�T܊�q�ewabmW���%�aC�J��	�T��8�:�<��i���s�lf�C��|7}�f��Ǜ������I���7�̬�tX�sb��擄g���
FHc~�fl�ܧ`t�b�v��C^z&��+!Ϥ�nژ=v^zn.U��\�:@�r貈Y�D^ �wl��+ߌ֍��W}q�[n�7gY���R��%�NKq��1^/#0y��D����r���������7��z:q��?
a� f�#*�ADw�TБ=�"���;�<>����fIdaJ�b�u�� �T��#�`�}�&���U���C�p�q���d��{A��%{�lS������$�|����G6�������T�
0+q<�W2���/��R��r�(��sr��Zs��g�=�j$�j�s~�0���X���q�ISA���\�&�?)�i���0t�M���ۑ��(��auL�9����T#�?���Geb|"�i�E2��Yǁ.kvo���=����u������_z����<G`y z�8py>������5�gϽ�����7�y��ّ�EUl��Z���Z�+:0#�pT�i#�[P�_�3?�wϽ�n�E35�& zg�8�0~�Hi�yKp�r�j�-2�=��<� ����U.��k�îθ�4@����Y�����U^��� ����Ѓ��j� ��z��+���yԽ��� Y`Z���R�ZޝI謐�i�{� ���k"ݐ��mCݰW|���0�a��B�e"q�L#�-���Ȝ~R6��&A��lS��$� �ڰ4`�ޝhZ����{����o{ׁ���G�9o@\X�^��UG� ]������[c�>:�I�MMC}�~��ߺ��
�!�$N�|->�ı_܃�}�D-����5� �ϓ{���2�6�3O24#t���r�����`�w���������*��9g~���<�x%�+x�Zh�^j���^C���TKxc��DZ�~kY��Wq�ٵ��U�_�����+����������/
�B��(�2D�g�"���� aD���o���47`<�c�s�L�� ��BN�a_š_݃X!�V�3t�fF����gvDĆ}{лm;��%iժ?�����RU��2u@-�w��K�.]���w|k��'VG`��k�}�=X��+�N4��B�#�-��R/�C��Ι�u\4:"�?R�t��z�2�<0��m*+q��Κ�0�:��p)Į�l��Ij?�0�kn�~~@�k�˿�o�
�^�9� ���W���:��'�b �>֠�N��[� �F��`ʤk>�mW{
A���i�s��'b\P����
��3	��(�-��3���y�����C�X��T����Ifq����f�(��}`}�]`��tL���\M��+vbh�^�D#���U_��n��2_R��;�:����o���1������3/^���~��<�zmC`1��~����CojDJQa++��
Ħg�����_ư-��t���Y�I� P�s��C/{��nȫ��W�jcV"��%`��6z��͂�x�*�Х��|B�U���r/qjs��;�`;�d�x���$��K��{�FY"�?�� ����E����)�v���95�A�N�_��Yg�v��,�q�1Ѹg;�}�6Xm	�L&u��Ч����aONC��A����g���� A\�@!v��Ӯ	[�����[���X�|�-�������lu@����}��Ӈ�}������CO��ע�`"%�hۻ{?�>�-m�i5��oj��&���Gá;�]cIt�"+�a��lb��/vjS���Lp�ߠ��H[�G���'�B��R�?2��y� �/���Q/Й�`�W�Щ[X���J@���=l0(��s����s�Dt?� H�HL�k����B^zУo��QV+�>�'��5j����[BR�1�IX���1��w �Q�l�Ev&}|��4Z,�x�/����/�	.�o�s.0k�0�	�d\��`���ڰNw����?�����]��.��u)�]V��}Y=�ʛ%@�_~�O��O�}���JQ��ȉ6������A��G1фb<G���6Ze	�T~��!<w����$A�-HD b��=�D���,y�O��I@8$ئ3H +�J+EP(���� sR\��q3,}���g]q<MP�#�J}� ߀UxWV������*�_KX����2i�S-<S��޸��_���1#�,<fy�M5�{�w�������>��j�9��R�F���R�撄�+bJ�Ѱs6�=��!����/��`��S��sh��⹋8�yX.���Ý�9� ]�(�M���(#G9t���lG��Ո�zIY����yc�2^jk�^���P��N�|�����#7>��ou������bPl��p�uh۽zO'�1�!Wס&����?�S��KhcS�E��E&q\�LR��vX^�Gv�j֙���Tͻ��U������X�+�y8wJ���.�R�f>�9��?�0|/��^����Qq�̯���~�ߗC�g�cBp�d(��cu	����BD�S�)�G5sf�HG��mJ�?�$�U����,9ޓ���(�fX?�M��ӫ��",ۻy��ܶ��z6�t\î?�0ڮ�
��`��C6�YL���UP�H�>~�;>�x.�VY�h�p%yQ�`�5�&]��&\U`�Yz�lA˦��;����|�_h��������{#�X����|��i��m��?Ó����~d堠 b���ʪC}X{�[�m\�dk#�D�n@��H2�3#����A���E���4�l�b,�9��ːDd�r蔏g�S��Kt��h���3��,��{�
{�^���	nO�m�G�
����j =�� ��-<7nx��"	�<�^����~�e�.	+؅K�eOǢ�
�J�>��%x�NF$ݓj�"#oZd� "��U%4�؈]��n{+U�Db�Ffj��$Z ��0r� ��+tH�E	�a_4�Dc�6�8F\i���.kMl)�ƽ�ѹy䁾�޾/\��O?�и����|#P�e<?R��h���3�������C��ti�"b�ށ�7]���F���卪��i�9xw����	�bH��hQd8��<`�)� ��U�0�"<�;��H+�c�B�s���s�A-��|�_����x�:��A1�Ɂ+8d��L��F�,��H�� tvDr^+��ᩁ�rᵆ�v��6�y����esA@g�>��G^:�t��d���t�6$4�n�@awY��$�Z�}?�}�`��t&�X�Y�iع�\�����N��{�F���յ�� �7hs��i��t-�CO���G6\��6@\����?���?�'uR�2^����뀾�x��B������������_�6G����-UBR��0��� �� ��3��H�ZN�hU���$������`P��nXh&0�b��g20%` �\\�	M��|qf�#�o^@���|�+�`YV���e/�/t̓�
�{$���܃߇Ǣ�Ӿ���Qh2�贁BI�    IDATm0�Ήu��:�A�S+���n�֮a@g�#TfW��������`H���c��"��U�|�>�n c�녂W7��Dab�i!�[���"u�8�<�.ME�("F�ˁ)HH9.� &� iA@�N��ظo/V�BÆuϨk6|~��?�̥�]}���G���xN$��9qa�����L��hߺhZ1GqpHiAD��X���"�ނBS#�
�1��c �jh(��<pO�󏠝��jIE3��f��X�T��P��u����@9u�JV�ȓ�����dF����d-�n�TV�g|�2��.�/�^�ti�î5]��!���s	m�t��b��3�|�.��=ؐ'�,��ΟOh�������?L��O0o�86�	T#.`F���iŮ[?lـ��"�:0�yHE�x3g�!��'���8���0&&�Q�-�T�A<IEҲ=@w��E"
�AS��ʽP��иq�3�;w�>����_��Q�֗`~�����-/��^��z����~�[_���ѡAQF�k"B'�H���_{�5C��.��8��tE���H8"��,���_0���X	]��MD�瓭d?4Lwt�ʦ:y�a����o�bN=<�Zn��r.8�
\�/�a@���|���ڊj���d����sUˡ�<j^�^��gW��àl�2ߤ��`)��g|�\��j�k��\�Wk��<,�^�йqA��8� )��)8��u�l��G�� QAfl
��IDr:���Lm.P|��=�8D��h���?�� �D���q�b�~t:��0R���{�q���w��/���~������vL�ͅ���|q��{�����}���>W@��"B�e���*#�fZwnC�0����4�Lh0��w��=����?�0��E¶w� ��q�*���L9�y ����D���s@Q��~�Z��K�9�������.t���p���u�a/��C��ZFV�(�|��z���G_䤸rٞwd�[L�=(��{��SyW�`�)���:��Ŗ&$�iR��ر�h4$lJ6��Ә>|�l
�(dӀlڈ)��(�.S�K�&-)�Ќ���E���;�"���Rd������/<�l�Wy�u7p��[�r�*G����z��q��w���~9���\�ŶaRnQ�T���ft�݃�}{a�t"�E�%��mB��76A�J���!�O@�a�ʹ�Sm:�;���:��� �X�e�\/��z�9x3Ov�Od!�d^�<���i��\�� �"��A9���0����p�[��`�����[���kEXʿ�����M%��3����`��X���xlLDѓgU%�uLt\w���!�=�����p��9sq�F\/����a����[ ͚�4aQ���UMAҦ�s�5g����oQ���;^����3���o�ܟ>���Y߬>UG`��[}�ހ#@�S[��{�����$zjh���B\�r޺�T�&�P�����a������IǄ�i�l͆��^��_��#O`@�Ф�h�ؖ^ZtEa��"y�ˢ���Ԫ#�4��Ѓ��Z����B���u��Tv)��[�[X5�^��������J޹�Tlx̸��{�_|o�JBЫ濇�U�жИ���K�Q�=��8���J�x?�S��=����KIr���(
0,�_M�$X��%\,̶%���[�z�>$Y݆�s��6��r���ҳ��yȳi�<���I4@��$�+�t�@$8���gm�$�:�IC۷�^�ex�ptӖ/^y�m������������"~�w^�������N�z��{���������7������gZx���75�m����{e7
=-��1��
U!��ht%��:�g~t'b#�T�u��ˉ�W�f�.[leWbd4����|1���TV�r�z>@�ϐ�^��Z�e�[ܣ�	X�l7w�E�8���kЃl� -��X(����Kyxn��R�+y�K ��t���9ƌ5J�+� �#�iѓd��j�FM��F������&��ȸ̜�HRy�.�MB̦-�?s�WNANg���"4�K�dD �I� 0��M���LߖMp{���j?޼u�����߰�������k�:������'@��9t�cw�_f{n��e"
���&� "��eX��X}��!�D����nX��t�M�ab/��S���!PN��vq-(����0��ǥ���j\ʃ:_�֫7� �Z��?_�o�R�Coo�Z������]� Y��𺘕��+�RI��Dx��s��\�^y��d��1J��e��"|�=�,"���ت>���;��B:gg�5�K��oN�iq�,���� /k�R%�\���{+�n���EN�D<�`��Y��S2i4:������5>�f��]
9����r]�Ey	H�.f ��X���z7oDd�*L�#�Z����M^�ſ9�-��@З�>�Tc�+����~��ӿ~r�J�E�� .RN�eqC� �� I�.��r6�E����J����Z,
��@�
����?���� }��eBr,D���tlQ_+�Iq�Ϡ,2��։svw���Kto[O���.=�w���<2�{@~�RHb������[���RծL6z��������?�	k����o����T�+��1� ��#(�s����3�<�R�3
���鵓�!�8r1�PV`�'?lY���\wf:��%��0��CGХEaM�"f1u�$��	(�"�e*S?�4h���tF]}@w0c{�Nw�ЉU�b��׭�tS�D���z�����x9����@�k�9s�YK0�Kt�%�Q����u��_�y��}��Jqbp�Q�,�3Fn�%�hX3�{w���wE��NT	bDE��C�� !(��<��w�=_D��!j�P
�
<R����<�[��(qବ/o����z��>v/$Q�<�Λ���y�`n��3����'3�k݃�5���	j�����8�ev=�����ϥ�
��w������^�5����/�������T���8��"!�Ep¶��-7`�G��$0YH�%dǓ�
.�\���Sؾ����:}
�'����ФJ�LMfu��E�`��4��A�u�t�5�t[TX�]�3�wDX5��?�g�^��~�e:u@_��n� =~��M�{�y���WB���r�I	��~2�����֊޽� �Z	�����KO�:�ٶ�*ʐ/�����#���a@Qѩ�syV����)�2���m+Ҥ���*<��gV�Q�����2+\�Q+_�n=x�Z�o�ҹZ�N@\5���/EX��`Z�p夽px��*s����Lz�k����b �z�y��-n��TE�a;(8&���%9�Ą "ٻo��аu=t�ER/@$�i�=�fGD��(�bq��G0v� ���jH�u$×Fr'�tEȺ62� ���)�.	�E	}[��y�zD7�?d��nק>U�r_���R�zЗb/�c��'�?}�#����;4<$(�Ɋ�X�D���F^j.���\4��P?�wm�6< gE�����&�1�B��b��'��O~��E(2,b ;�+
��	I�f-�\2w4���>������ ���ǈ-����[�tϛ���j�g�E5�V=�|z��Մe(� �`N��s�XX��<g5@�S��*�Gx�י���K�	I�Y5j$F���&�B[+o�	��{'M@�,�hZ���8q��t��5ez�Ǡ�=�vM�S�20'�(#�U ����]�)�.zQ 0\��6�m�&�7o<�w�}aﭷ���/ӵ��r�u@�<���u���g���}��������T�����iᶨ�#��[��X�вs+f�(4%��6�P���d��\G-/����]`���Hs�"�����C���B�8<��zy��u��C| ��xS"C-Ċ���^�8���Ig��:�V�o9��@��� :�U�B�)!�a�Iq��Q����ơ�t��_L>����5l8���s�t�P��.���J��V�6��Cu6#y�@	��{�	y�H�E����J�.ds�[���ګ��{�Vt"��A�L���c��(
c�Xѐ@���8w'�B�Y��Aʌ���W
g����B�E�Ӗ��t"�m=��A\����N`h�/����?�,�S��F��o��y��rq��X�ţ7�����/��Lp!�ǅ⻆$�a�
��3����>��ڊ�n(���[H�]c���SGLׁ����;�	8r+�]�ѤF�/�YW7������ �k��ʰdV0��d2�����UZ�˜:����Ŕ{y���H؆��3\�`<,�9�Ӟ��=:t�"��{Z��^j�Tw���;^%���s�)Vv7{���n�z}�9��@]1��[�{_���|պj���Dظƹ\J(���G8J��F�c�w�f�C�Z���T\���ڎ��=`�)���`�(�dP�LBI�!gs(^��X� gb�S�@��X{`�uY�9����ǒ ���{A$q&����H��׿7�!�v5��M'�v���������W3���G��@З�\pO���O^��/��g���h�M$\�����IS&y9�ۜ<u�b]�����֭E��� u��h��(�pE	��:3��)<�/�	�daZ�@K$�Xd\w�9���_�d<��ե)pؐl�-Ԟg�[9�.�<t]o��4����AV|������"?�
��ƾ\��eR���ur��A�r�����b~3�*ۆ��b�l�6�K
�3�gmyY����"q���ƺ*�0d#�"`�v~�C��܊��C�0 Y"TKFn|��)h�"�<��Ù�59}r��Q!��^Q�F��ݿ0"�9�� �B��ST"� ]`�w*�l��C��5P�W��׮���/��}ͷ����oꀾ�燻�b�?����՗���кURM��F�F�����S�ȥ�;��lda#� �nzv��܄�� ���a�V�4���m���>��K�"��ez�uj���I�,u/$�Q�I*���&��pR-{��P��� �0P�Ie���A`� F�4aָw����: �J�Թ�N��T�ZmL��<N�:��e������1pB��F�J�?̠�%{��� ��`�h�aǇߏ�믆�ڈ�i!��A0(��8���8"�<�����H�r�՞GtQ���#w�(���]w�sp�}��@�k���޵u:wn9۵�W����ү�x=^�[�z�Q���b�_�� @���+���/�]�6
*���r�� �4�	�lb�z� �d��*#ݽhݰbo"k�`w�æ6��(��<A��lO��a䡧1�(hM�hav>�YkW�u�Yn��w�>�,�/� ��؉�F9���L��zE/��m�k�C�����׭W�L��G�� 8���7r��%�ɚ��y) =<���k>� ���U(zr�a�Vq�|Z0���f/���G��L�����L�!�,ǧ�N�b��!y��Ϝ:��G�$"�P:J�`{�%��Q�3��� `�qý�r�"th�C疍hڲ�50�ūn��=��u�~M�����yVK~����_�����o���	�D��� �<t����`��!�K"1(+��غ	vo��hY�
n<���ÕlD%-	��g����ǟ�@Q@���5��Eu
�z"3��E�����/�#�n	6�%���� �`Y�ЌgZ�>@�k��%YA�z~�Ҿ>9��úT@_��=l��+����W�V&C��C\��L�Z$:�`��R<����X>�"�qgD?�B�*?SL8&��a�;n��ahm¹�1� ZfGơ�M���I�kiE��Y�?x��83J�ٲ�Jd��a�'w�q� ���.x��<��7 +{����}��[?[�~]�d�oSs.	З�׺��
��cW��o��٧^������У�0=�<�()���A�K�ݲa66���0�V`T�бq��f�CTb��U�ABQ0���x�����*+q�k�E�-���yd�w�������)��?^X���l>!t�A���:��*(�tN����7|n��1� �~�oz-�f�{b=�*#��n�T��Ό�{�Vй����.l��R�8��*d�	����гoֽ�z(뇑l�	�L��BO�1s�<���0{�$�L�3�>{�y筊�'�&T"P2yW��.��I���&
H;��T/ Y�{у��4�F�����u7}v׭���,v"Է�:���1|c����K�ub��w�+�,�yÐ� f��6�N`N2`�%H�˴�mS���(�.Ihܱ	�[7a��Z�J�M@$
)�!X�b2�$�16�ӏ<��<���z��	.c�ɢԢw^�VG�w��M
\$�i��bZЃ ����������+�d�W�h�}�k�)�9ls�e@^��ϯ��B��]�kp��5#s��~5^nV�ؙ����۝e�2@���ٖ��&#%)��D֭ƞ���a8�Ȫ4R����<�cSЧ�!����ۏ��y��Ϟe��m�QU Q��v���s/J������a@'A��ಲ�� ��N@O����~4oX���X׾k>{ŭR�7��[��:��և��sBt��3����_��y��U�� ]sLD�;���K��;���%n�,!o�D���5Ћ�k���ى��)G�xZk3��܈�)���:����ơ_�
=�":]��!�;'+����l%�����--�h���'�{L�!��j�d��{5�;�t<k���e�U/g��B�
�Tk?Z!�*�*�T���2��KE5@�v$9	k�Ӷ<�1���8	6���a KâK��,aRQ���͟��e3c[��I�0�"�t�lN:�o#��`W_��<���W�''Ѧ�,oN+��j*h>�1+����WI���À�� `�t���nLQD��ܳ�`��ѵ�o���O?��Y�Wr9�@�/ǧ�D��>��\�=������o�}~�����z��:� �2�W�u�B�~�-:=U���c��}�Fh=}ȉ*2�okC��bB���,�p�4���'�y�Y+*ZE	Zр������z��A�(��V���h�/G@խ�L,�AN�$�1��"�γ{��w���$�@y/��Pm�L�Hq���ռ�j�=X����B)�����K����t�ϠX7`>U?nh��Y.$�~����T%8���$��|��5�ڱ��AǕW�����/�I"��d����pR�7�"u�H3�L�={�,���fQ��X��I���W2x#GY{� ~�T��sm�X�ݫIg�(�8h�Ǻ����Ǌ=}�^��[�үK��-���}�>y�����y��_��w�شJR�&�,���Q�]"b�?K��&��bU*��53���4tmڌ����V��Ed#�W����Wl����:�/��߇�S��R\���ZP�3�i��'D���[@y��ڻT��@9�|!��Ml�W��Am��WK�W~ �O1�RN��z��CN�0�s@]H.�
����vK�|����B�E��a��LDF���{3�������	3[�[( 7>I7 ���&�����g1}�(rg� Z, Q��@��ʍj�{����=uC�nB �Sբ9
�S�	%+6n@߾�L)�����[?\�~]�����«ؒ��~����tD�t 	�ͻ�����7��|��m�B�)��Jֈ�F�L���ō+���9��9���i ��::Ѻz-�V]���H��8��(���1���!��a��]�:|}Z��대$"L8>�]��5Y��@�[@˒�����R�8��j��w-�|�,�(Ɨ�FD����}f9];�W
�S)`��7��M �O8��� ?$8    IDAT��g4���r�a@R�Ѓ�GIhUQe�DQ��ȸ�g1&���*l��G��.��:�sEOA.��5�An�ڟХ�aNM��u�<}
�WNAG� Dm�&E�k(B� �_Ά�k�{ �r9]X���( e{��l������ݻкm-����������z��.p���^����C_��f�/�+�����=���WAAh!3��a!wj%͘�>n(~}8�Ԡ%M�I���%R���޼v�wlŤ"ݝ��dĺڠ$b�,"fِ&R���= u�z\���0��f�ߙO}gM0��-�0rp��QA`�x�,�V�;<�a�{�g�/ �aw�N���Ы�������e>=�E��ń�����2�?�o
�k=^J)B�-H(R�YĤ�"�n��w3��[P���7l��������Y�]���P4��8H��Å#/#^�!eӈ�.e����[�H�t)���ѵ��B�9�A^��ld�D*9�E�ڋ��[0۔8a�IЗf][�G��2~��늅����_�;�N?v`�*WF�D-��Cg^���ӚN��B|C����G�|�敠vv":8 ��R�
dc��=PZp4�$B�D4D��|z?���Oa�r}��v�1/z�^���A�@��79�8�z�U������!����.bU}�R��/�
z�����������_kM�0)�V(=x���V#�TM)�Bx��W��oX�Ô���l\�9Cg��~�@/Q0[�#g�ЋE�`�09��%@)Z��9/"n��x�$�O���m	ɗ=�DR4ʣdzQ"�����)�=� H��vYD�rX*ix�Nt�ތ�X�i���^u���2�x=^�[��R��ez�u���~pՃ���wҏ<�u� �qu�C�<s��E�x�C��D<l���Cr�.y�^H�R5��͈�@���lLC��AH���[�F��(�)Ri\|�)���{�?���vQ�jyfb��*�
�`�..�a@{�a����i8L\�3�8f н�ޛ�H]�[��yz�5)#l;�t��r+�g�{a��������R ��H�}� �o���#iL�hC����W셩�,�I#�JB�����l)����$:�b��q$G�A,�1-�H�U�a�V)�A�v���>۝ƚ�ד�˳��cQ�Hp�~;�C�u�^��ׅ� ��7#�~��g�M�%;��s���ۗY�`f0� ��2 
�(ˑdR�U�+���#.��R�$�R�TR�(n�,ɥR�%)���K��U"	�W� 	� �Y0��{��M���ow��`���m����}�w��Ϸ��|Xm�N׎�ٷ������t+)O�ub��_'7�Z��D��|�7���[2K���)Ud�C7��^�--6h;��8&[�($�0g:.��`v�������k�th�תH�3�����翄'?�Wȟ;���B�z��\�������@f���Q�Ji�Tg)~���k����j ��"�-��;
���9���H�,)��YHWs�0>o�{����Ž�u�N�r&�з���I<c�w��@wi���a�4�뇒bgj=m�wڨ�<��z!�ב-�bO�ř�{��
&,BTM�00ƙ0�i�� ��F�'гT�M:4ؒ��, 6���~��l�ic�C�߱k��3�;�~�C?��|�Z��g�8(�ƹ���J���Ὗ������Ï޳�@R��򊖻^)[ ]�� �T䵈�9�,q�#�Z�sj뾃�÷�?]��k�=;��Z�fݓ�\/%˽��8�����������Q�x2�R��(�Y���>�B!�94�̘fW����Z���]�Z?)mZ��̱���+��Q�g�#F�����E����Mt<�Ќ��R)�����K&�%m��4�a����b꽀�.� Y�~��E�hgiǱpٶ��\�����}�B�Hst�[H6��_ �̀�`r���&|:���v��A��
3	%2'	���9<
��ī��>(%f��qU�qG�ָΤ�n1[����5(��� wl��~S�܎�F�t��;���O���^�&V���Ai����g�ӝ���G����Wz�!����m*����2� ᠕MotT���9�vQt3l������A�V�λ��k��KX��#k����Lx�f�~�s_�:�������؝ۘ�bL�6�<F�G0\!�>R�,a0KԨ���p�A�3�����z
�d=�u�`w%-�W�,���e�0-��R�%[�c����p�M����wa�-���B8$[;g��9��2;��שi�t���̄�Q��B"�d�g򚂄��u�����L,�<�yǂ}����~��['���16W֑u�ϝǔ��H�ds�s�ѰLL�V�}��<�	�L�E�Hg�-rĊP9L�ܼ��{-�P�`}�)�\��B �D�N�?��g�����м� ^0�S�{��3�_��O��uV����r,��Mm��/���|�?���7��t1��s:Ǟ�d��x�&���L����KEQ��ﬧ+�,Nisе,��:��h>����38�'��<IѴT���gp��/���'��9�بS!1r�":*�CEJ�zX��mn:�/@}��ǔ�^�����x�h������_�@S�]�8"��}k��:F��Zz��)� ����}3C������r:	�1�^�5�� U.��e�C�d�_���p�;�To�p<t77��7;謮#a�y��J�	��fkh]:�����1oP�plʷj�5�Ռ�-cQ) �b�R0T�qXd΁��H]:���A��1��.�n��ۖ�11qһ��|����������&:f	�7����R�O��]����;�G�V�@���8�3j�>�1@	��Ls�Y!>c �\t9עREǶ��������]�!ڳ��$̉������f�D��5<��O��_�����G-Ie���)�''I�w-Jr���$�p��r%V#�5[��lǌ-��ht�U�&ؖ�?6�}�v5ڢxﶀ�9���X��_�������r���s�	�$��<�Q>��8�%��cR��T��A�yX��V�î�������L���:��]�Y7���F	��uiO��-�z.ܠ�3O?���2&^��:�t������Bߠp�j(��#���0�k���9:i> sF�l]c}��w�v�-Hv�8�[n}������Xk�1��xu���ͳ+��i��������O���h���x�8�� �n����$��R��%�Ղ/:�>%���E�5��^�!v\t�s֫@���ÇP9x ��,����
⊃�4Ps<xi�
_�2֞9�o}�s�x�D��q�f���hJ�[)0g�S�eh����K?ҷ>��R����k�������h*��X&ۥ̋����ǯith�-�cj'M#��U�Bu*y��(˪ pk7���i=ճ�>z�a<I����g8HL=���<�F�Ǿ��w��v/���"�� A����α��>ҵ�?��N���B�����K0�Ӟ;I���K~��[d
�:!��ch�v���	�ʢ���K�I�ѥRIqz:A=��r�n4�<�h��g��{�����/�k�<��k��o�{/W~�?���>�ۣ�ޠ;��q-Q�^)N��A����ze��I�;Ҫ����[ǎ#�^K{ѫ70q���f�47�H\��JӷmL�+0���8�������0N_ƒ�Ĩ��N:A`�*-mwŹ�{M`H�����v�>��FIeߩ�p�V���p�t�#�t�`��R��a�_U|]}�9:
��� sr$	Y�C���:z��>LD���$A˵�/���}Gq��ux?V//�<� ���Z^��X���;g�a���Xp9t(���ѿ���e�bYȢH8"�(Q���U�]~/$^u����HɆ·t):i�FƧ"�!,�F. �@ާ����>���h�Μ�w/������QN[����W{�%��Z^��?�w~�}�h��?����ng��KPt����ʏ�ph�L��T�o�e�$&7:vQ���;![�A2?caqŃ�0+��Ի�[6p�"��38��G�Xkc&KP���i�4r��>�W�^����I1�}��
	٭����w��<^��\_j�|'���oi��ɿ�㎷����K��+��=�#o��L������sĸ���7���R�c:h���M�;q��;���`1�8�)Z�W� �}�.��6���:��?���s��N!�wP�_� �0(�{�MS�}\!#�@^��3��R�f��[��
@���a��	��+���eښ��Gc��C��Ϝ�w����������vR��5�@	���\ˏ��>��w~�������{`)1��NR���i�m ]����yHդG���"H�M�+rU�ͱR�?7ka�U��4*{v"�=��=v��7Q�mԙ�����/=���X�/����@�傌�V��:?��b�ݬk��uN�rd�V��Ѵ� ���r�8�"g��~$U��ʆ�JR�v)u���H��7�>8��}o��]�ɭ���+U���
�
��HQ�(2:��{�*(�3�����7d���t�����C�1}�Q,��s��<��t:�[]�(V7aF1̠��s�,�K�8�8��S�q�&]V��)�A�r�.�+E��Fm�{(·v�{!��b���;����c�qm��npF;�)�vKR��`��;`��w�7?���ܿ.�Я�x|�M�_BõXO������>������co\JMQ�k�$��Mo 2P��؇���eT �!Ӄ��2��&���$��[��oa������g7.��Jӷ,!���=����8����bt��(>���j��j/�D�a:5Q�Ɯ%�q,�s������Qg;������KE�ڭٖ\���.,'������F�e�
Gct>�v��������آ3�J5����g@���LM�~<̄�:��%��v�8�y��N��ozXc�Ďy���B��J��1��76t����g/��M��F�/��"/p��'�����d?��A��u�D�pݥ����g�3P8L�Lv.sQI����1,dpir:��ٌS�1�g9�F�X��e	Sw݊���;�ј~��˔���o�ϼ	��{�����w~���h�o<��,ti[�S�K�N8J|r��Q;�j��l�aħS�#���`��U♜H�eʲل=3���Nр�fekϵ�����z���Ѭ#��P%�)����'p�k���W��F?��G3NQ�)�c�E��*[�	��e�{^��Uva��r5�Ѩ�Ji�tG�Q��� �:�t�Է�?ǗjK�R��E���� ��LE��P�1�<w%��o���x��iw��led�񰚄�t,�kUTnY?��w��2�l��A��o���uTrI����Ac6ν cs��L���O!\[��D�DSA�'�� ]Jc�Orf�04b�Q[�9�CM��_a��fz�Dz��`�:�er �L�����=Gc��m؜�<���g����o>�|��C��(�&�����/���?���N��o��c�RCף#@���R�R:�H���	�/�!�2��I��H*՛�����l��Z��-̠>?o���0�gga�	�^��8����W����e��&F��R�9�k�eH�{")w�{X�'Á�ۦ��"��:��J)��G�y)md��K��t����UJL��3��l/�*�6N� ��^������p�w��뼆��T9n�q�ܮJ���,�F�����޷�����6�H:��܀�dX;{g�9�}3shZ�v�'OK/��c�ҳǥ5��r	fЃ�ƲX:��!]�ʕ����Z��+�y����a�i+�6g�.)w]����d��JP&�-t�\��F�=w�����<�����%����kp�%��F��A���(,��7�p�p1��>�� ���D裀��U�."�+��j�e���4���Uo�Eu�.$S��>�����X�e�v#��0�U�f�I���g�B�����g��S_y�^�E��I��|#�`�Ԩ�Ly1�]�yQtT����4|4
]W�
7eo�o�dl�R�R���j�ۭ�����U��-�C����?�i�cW<�0�����.��Zc�*��*f��Gn�������J H�4f�;E��[Y�Dh]X�b}Y��jj���S�;���o#�|	N�fR3'�;�.�I�#��l�Pp�ne���
���F&k�RQ~`�b�n'��lK�q�,Yؽ��қ��Id'*wyϛ�>w=�%�_{��~���5=�����(S��/~��_@�F8��Dݴ�zU�̀� 9�6�$)G�GZ���f�i
��Y&������c3��91�v�ˏ?�=b�]��5���P��8�4C�r`{�Ϟ��?�9�~�8����Y�AӢ^|;�aID6ܦGS�Ҳ4:�K��۱�_.%^��-������$���Z��* ��:ߠ?|�*����.{���65����P���V�ScD�%w�j�62ۖȔ !C�vqִp�C����u	�-t�k��q��!nwd���S�q�ݰ���5_;�j4,���#m������<AͶ`�����	C: �(]�Z�~Tm|��8�9
�K����j�CBs�G��w-ʿ�9b�¾��b���XnT����[�{���G^�N��(-pe\ݷ�uj�����o�N�d��,�Mp d	��M�h����\��e}������ӆ�@Lj�)�jM��f�/���Fufg�]Bef�ܠ�'0}�-@���wḜ��\Oz�پ�p��=�gy�ً�7Z�w<L�6L��NxI]#�X�cы<ڳ=l���܅є�(3����_.B�M@چ�~5�U80Wz� B�t��Z];g� m´�jg#�[�-[����2<�\lD!2ǁ������`��#����w;�E1�8���&�N+/\�ޅ9k��<�k�h�p�fF����9�=�,6/]DӴѰl�I��QFu=Jvj,���p9T�ಶ�9���{�F����� �EPFd_9�0�m-�]�?v*wc�Q{j�[��w��_��KWs��ה`����=���-�����~�/}�IqE�nf� :7�� ��ڪ�<he�a �#\���t���c�Un��i��T����--pff�NN���7 ��у�K��f��yv�`�����=��e�[�uaQ�����8����G����y��>�C�P"Ks�ul���i�A$|��� ���&�z��p�f;Z}Ng��4R�j�/�b��J5��ϧ��GO@/"sUy��E��h�Z�z�b��\i��[�w��� �\�n[&�A ҭ50b����8u�8�t�0�}��_6[��lSLq���V��c4,GM�#Dg��dCS������A�i�u'��}=���g�(hKt�#�УLɾ��N`'�����:X:v/��:�3����Co}�=�xW�wsoǯ����U_}y ��w~����0Bdo��\��'n�Z>DC��i�V&��_dWB��T[����,�]a='�
������F7�Yo����F�`9�`�Lb���W��:�3H]N���q-4��˫X���x�3c���1��U� �8#)��հA�|�.�E�ҕHi����pF��WKnȡ�ɑ~'KZ �ez��Iq[2��"�2�N�s1�,Q`�J=����`��a,�uj{v�3��$:�.R�A����(�q���	a����N������+k�$	j�	����g� ��=�p*p(7�E��8�EHj�"�N��;g��!�;��W+�X��]Ƈ�U�����vYܪ�D@�d�#�NpO��~�Q��{�\�������������ܿ�W�6o���^^���en��k*��?��S���ﵿ�����T�B�u�r�Ӗ�O�G�V%��b���97��Us�Jm�bC,n	�\��MU{U�h�i��UC]�
ï�S\    IDAT`���gp����kj��#�W�T\X��ԝ�/D-n�3SS@���/~O}�a�����	PO2LX���4e¢�{���mҏ�P\�����_Kڴ��k$�` :2�D�ũ[]�Ђ��ߪ�@�G�Q�r\�>e�y�|�c�Z;��@8zԂ; `i���ɇ;�:��M�F>7�[�����!`q`69Z�^�}��]�b�z�_�D8���/���������#��D��%��k�⮌�eх���k�z��?��e �r�y��0Kt F��܋����q�j��ϛ��^���Y�K��]����瞻P�}?Zӓ'&�=��{��{~�[W>_Z�,������jE��������wï}���4A�B�_WA�0O��e�)Z�c��� ք��YшԬq>��@bp=r�``�"�إ>�Ӫ,�C.1,tȂ�L�y4�fa��H-KX���:�i��}~v���Ѩ��|0�l �.�K�蜿�K�<����d���4�1&-���KS�
��c���ܣ\��#JS��bU��� �M��m(&��+p)�Jz��+Dt�O�T��킅GG�6���`p|��Öc��`J�*',U�1��?9��R��mq��3�5�����3c`�Tخ�^�!q}l&VL3w®7�/����(7��>�D��D~�f�T;��'O�%���MM����@��J�"�XG�n#j���70a�$���t��9T.$}օ������#G�'GK�&�s�I�S>;8t���V��4�@�����K��O�w���c?������~�/�;���9���]�@�gx����~��-�$A%�tM��&S�:��͝�R�R�4)����0)�PU�e�`%u��[�=�"�)�l&�I�R���im	�Q�S�v�D�ٔ�z��i�v�B��+ˀ;5�����0mnŅ���=2�]�J����|I���s�9��4Ǵ�	�'���OZ���
P;�ئ�2�̒� ӼU��tE�;�̨���l@����c�"�y�ã�/����}45<�-�g���0�8dl��_"IQB�Y>%��%�!�厅�NS놉�8A�h ����o���~LP���	��5�͵uu�0��[�"�,G�讬��2�jN�s�2����/b�6��1�ϞA}F�5�ˬ��|4��p,�Y���M�4�Z�����#t�ڨޣ��QE�bz1K��a�r�B���ѷ)E,���}�wo�많��{����U/}X�z��(k#��t�_|�W7��7�(@�Dݐ�jܴ�ś!'�Izq팩%����b����B�S�S3�qS��Z�$t�ـI�@h�ߗ�a�La���&"��T��ML­5�{U�	Tv, �h�[��k]�c�9?��TA��LML����֦J�3Z<~g�&��	tϝCöд-��PҸ~�a"I�$�g#�؀�0SI�
9L��u�����eBG�N��"%�a�..�{Tz�Ǥ�E{�#n���}�E�0sq �����6+�Rl�ѹ�%h&b�#l1�۴�~Di�,�&:6A�A����I��>��(*��wQ��nW�n�eK���2��T,�8[-x�#�~�<vMN�����E��9xq��Ewey�+��o�J�Pg=
}����*~����^�P8�|t)}0����nbh	(4cr�����>����	����������o���]�+�kt��Ǿ����?��~���Ǿy筶�F�[>L��};@W�Z�G%1 ���A�i��ҫ4�J��ȷ�|G��o�� �ˆ]� HSl�{0mͩY,�݇�^��VEu�"���*.Zf��mbb�̚������mQabbBΡR���'*&�.��翀o}��˨Qd��nO&�5L�.Ud+""��Cฑ3{!�
��R�.�!���Z��� �Y��|{@�5lm7F�R��?@����k���*���GP_F�K=Q��3�5��N��#lK�鴓XZ�b�A7�a� �:��i,�~�]���^�}� 07���֤N�J�s�YóLl���^m�7��,N��9�p��'�^v�G��'�Cu�(���[2�fN��
.���AB|�׼�yMg@�}��D��j#t�ץ��i!`�={�{�;��m�bs�q�r�џ9������^�@	�7��~���������>���'n?�8h��[���/�E?zPҾ�#A�3��XR�#K-Ka&l˔����,GL��P��<A�8��I����v��вQ�����C����wm�َn�Q�<����P�h��0r��,O��]n��6�ԗ�^]����3g��M�N�B���y�E�-q��mdp֊p7`��O0�E����X�+��"3�ǈr��`���N�C�Gs�� ���0抐%��r��Nrߋ;��)ا�]CM��
n��1�-��0D�4Ѳ2���m!oVp�ؽ8��7s��¢��1�@���!�NN�#��Z�[�r_ܵ�4O$�������e��8�cVϞB��E��ҍM�V/ˀ7UJ�(�N�Z����#���Mn�^���/���R: Eʝ�AE�\�*!�����\ ��e�-r���{�;���[q�������7�����7�vT^���@	�Ҁ����?�����}�#�cO<h;h&��h��M,#Ì��Xʝ�c�m@�)��XC����qdŨ�!��	Vd'3*g?���6��0cFs��sJ�%�ޣ�GV����O���[@m����A^��Ϡ����C2�c3aW��&�p�8�
l�FQQh4�U���T����8�ه��_}Ʌ4�\��T-��g U�; �0��1��)Ep��h�Ɵ��h!Qi�:!����Զ��Qv�S;@�!P�Pj� S�^ K(|:�B�����6ݤ����iw�@:��$�03���.��S� �礤�!�(F��H8*��C�飒�0�!��6\��a����طo/��ƥ�+L�54\�g_�v�u:�\���ŋp�n���ڰ�Vµ��:C"�{G�s^g�������Е�3\iW��-�����v�u�'�Y�f�@ER/g=E��xtv@a �l��(v=x?N��i���y�{���~�o����K@��7�Z~|��&�����'����N�����$�bT���4%"�n*����8-tl�zcc�J��[f����U�Xm�ܔ���s��1��bqUu�|�����mN}s����aT��/.`bi/�G�()IPm4���Hޟ��Ѩ��%h���̤��Y�g����eA�^�tN�D��%Dkk�n g���лtY���*0�NNqH�Nk�P�TH\Z����A��j��"��$���b|M��]/I�"�̵���2&����)�e]�ړ��Xb/�Z1%W|,:�����;�+�	T|�s���f1:�6\�A�Z=t�7����6d^y�� �X����hTX;�_[:j����b��9l^>/ҭIkq��<�����9
bӐuP���H��	خ�_�cmzW���~n腛�l�R�t2��L�D!$�9"��=vs�s8�q�=|��o|�/�Z��g_�(������
��;7}����>�[���������hG�/��p�c�׭�t&ƥ6�(YVQnj�˸q1��Q��65�\E���P�-Hl*�̄3�]� V�u�F��l�*nd���!�I��0]����ar�nX�M,�݇nc��A;1����X#<��I�؉ٝ0m?ۯ	�^��]G��ޝ�0}��vK%�N��O����4�<ӵ(������$���v��E���K��1��AV1�k[��G{����"K�z��Y�f灀Ɉ����fH����Ad����5�����?=�.I	�w.b��-��u?0?ˉ*�9L���a� �Bq�N�F��C֋ē^��j]t��N�������q���C{ys�L�w��XYFocy�#��JS��*B���r.:�M�p��Y�#d�� ]�݂��� j-i�kh�mm�Ѹ���藭pNy��{X�uꔻ�ۍAn �XCg[��mcױ#Xx�^�w�ӕ;�~�=���O��/s�����yq�=J@����U_Q�����Ͻ�S��o8O�ر��h�	<b����;���Q�Z43z �R�KU��Z"�����Ԏ���2�W"�"���Zo[Kr�z�p�JqAܐ��H��� ��AN2���ڈ*R����p�5���\^���^�,�)n�z�8���N6����NL��ժ��=��y�+��Ȼ���x����Y�]^��fR��m��r��vG$K�[��	Z�:���2A�b���N��/#w��RO�/$�1'"i�i�$K%ca9>r���$!�.��M-S�G@msW�S��r$�6�8�o����M�������C
?�8���꠱0����^����BrcZ�uau�ž��v{�Da�}����SO���vӖ���G��B�oa��E�7��9�&[� &L�C7:�T��U���W�⸌m�[6���|@��{-��/⮎��=*
&t:��`I�ĐLu����C ���!�����\����ԏ���o��_.S�W�{�/��%����"��j�ԣ?������S'��9��	�K��lb/�$o[j�pn\���Q�n�G@4�e��U��ǐ �~�>;�k�5�--�#����5�-�iH
yfq���p��BV�ab�nLݲ7װ�� 0���&�f�;]ؾ�ɹ9��9Ӿ5N͇�YH�P"D��f�S�M6S�D�88���(~}��&<BL�����8�}�	�1��� >������Z6��|���\'H��UX�N93뮃�NW�vf��FF��$���쎝�ME��5T)�뺨0�혨����ͺ���&1bF���C��z�}Ĭ�w{��I�k��E�\Z�ыp��}���d��I|�������-�a�ԌȻ�=�z�Uqʌ�o[p�S8«�	
�_1�M�����:˼ ��6�b����_��z���b} t.X�8��T�r$����G�����[���^�q�*w��7��>~oG奿(�50��zz�����'?��[O_�`����#�Hj�@����Z��e���r�oJF���9Y*Qjb��V��� 	�M���#t�A�z����[��\�ؘy�l��;��Fj!�3���-7���,�$}�'0����`�ӁU����}O�rJ�ږ `7�`86�Sd6ێRT�x�@�D�a�^��Z�*��Û&<ד���M0fM=N�������a%9��˧N�K�^��A0�mol"�C��d�0BF�6�MR%h#��'�6=-�u�s38�����J�ݢ^z�� ��<F�4�mˏ(Q���'�v>:y�I�M�ʳ,��=��]�66���i���8���l�wvLي��z�&]W���#�z�,�E�p��Y�_� �	�!Z���5ׂ�<�Q�;��~���Ma�ȅ�����ATm���J�g��η�h�ш\�F�s�_��|��\b�]	���cR?A�ϑ���5Jߝ�N2����m�q�Q;��~�Jqe�z�L_'�]���F\��ȟ}��׾�O��}�a~��.F�
�i�[�k�R���]w�Sۛ���0Wj��.��(��M�LRX��D���!�Z������H6ۑ4,���-�U�9#�� ���$��:hE	R�GuzS;v	v�>��YR �į�ܜ��?w�4,����]��ֺ�N�19لc0m��I��0���!�y���M�ı ��K+mZ�]8~E���S@��Ћ�dv��p��
�N�©�G�q:@4��ܿ+�}�q�j�V:Z�'	B���#���$臁�A��y�6�A���C#���NM��"�v��lazr
�n�jS3:	:�m$�.vNN`��I����f�>��+ZkȣI�CgsQ���nۨ"��{FI�8�H�u3�P�F\��h��Q@GF�m��j�Ep��w�>�F�E&h�Vx5$9� �Pz�S�I��ҙA�i��gy/͍Hs��w���7ރ��؜�>U��Ȼ�.�_��6xC}f	�7����.&�1�|��~���������F>��s�z����� ;�4�ZZ����k*�5����l����
ZkkB�㴳"�*�{m�
���l�A$/N�p �
� p+g<���K8��B@��RCc�n��&����Nmss��^k������-{�9ւ.܆/ ��&]���$��~U�CP���eY�I$�&Ή^�1-x#Q�ͥ�m�������<G���F߭$r	^R�t��E0���!�R�o����G����E�dA�8�t>E���3B'ؓ��H��j#���{n5����
.�;�{F��������&�k3��?{�fj�6j9$B߼x�˗�][FE�`H������ER9(2���H��2�$��y(;ʑ��*Wn��ng���k��^�K�]z��5�5�t�,$��xiQc��K�(�c�Cb�	��n4ｓ�~Һ���x�?�7��7�|ui�1g�4��k��s����yۧ����r�~n7S�L�3X�!�DF��Z��)�"RR�̭q�� ӗ�Dǁ��0=�%��ı��}Q�H�oQ���z�������F�Tu~��$�/Ln�>U?��_�MU+�_� �RtY�6\l�1����ۋ���Z�F���$�K�h,�ʈք��5�~W��>=���0���"q�R�
�9�]z�3���*�:eN��ՠ�5��	X��*���=5��)�(�θ�},��I"}�l�2M[&��{�#��{����e'�.8����H�˵\y}E���^u<�_���'O���ݨW�hQ���ìW���Ο9��d��.�<�SO��,��Fh���2��-�G��ڹRx}R���{�(oR���tu�l��ʋa7c_��X/���n�-G��G��~u��H@W�8�������V�yL~�t�=�@���7ae��}�л��w?r��F啿(#����1�Gu�'��������̉��:@�٢=��n*��(����A�-&��ʍ�H���a�*o|-#U����0��b֌�v^���cL�oe1�x�*t���l�T$B@�V��zp���!�o¶=�� �c#pm��L�.`rjv��N����Fڨ#kT`�kh�a����Z�0yS^�˩Dff��Tx�c��*A��*��S{�yN���
���e�?��T��n�D}�_��z��<���{����X2L[KdF�(�0[�L ���3C@_�U3�)��L�Ã�N�-�~�dQ(��v�%}��ϟYܸݖ>�hcI��If!H �2I�gI"�	:/�N-$96�h�N�E�(��âʖ�2j���Ì����o;v����hk�k[�ЅǠ]Y�3�0t4xm�i��fB`Lr]�lS }���p�Vy޿��w��?S�O�N����i���z���<؇}�o�3���Yy��ܞܐ�,f���It�:'��hU#�/��	'j�J<j@�=C���q�EW���5�#���F��|#M:�2����xTLs�>>S����Q I�iN����-��2h�6r�%A_t�St�~��������v���DR�`69�H�T�V8ąKJP����)���>��k��m��3�A`�iG�	r��2��eP#fa��J�uSm�� g�Ū�LMh�S���R����8���T�@�߇�yℐ�F �si��<��f�$N���@����C\����������
�7/H�p,�q���cݷL�Q��1�(&�<R�x-�L���RJ�&�[����{knH��u��U�n��_I�ҡ���s�#�b��HGD�!��8�(�����ǫh-����\�q����q|�ǐ���z���7������\�m����W��o��-/e�H��<����ڿ�<=�]E5�Y̭��G`����#rnbE�FR���y�ܛ,u��;�?&C@�b'�1���E�\-�q;�=�  DIDAT3�A��8H��4��_�liʠJ4,�}���֮�A�ff�
w܀���0�ua%ۓM��݃��4�Z��i��Y&D� �$�N�&��IFc��-`�߬kp�lA;T���9���r��,[�{qH�X��5��]�E����xYN���CDV��a&�Q1%Y#����S$
ڎ�<	qԡչ �oڨy�H�������~�2�/\@{u��5�c�|Yƚ�1��)�#�?'�䕤�f�kq��繱�?�ZW]_�9抓����QsQo�g�ɮk�h�
'�(�hQ�A9g �c�Ie	��<G��8���W/\��5G[�ξR��GA*�	�2�F��,)�l��_u���;`�ߍ���y�#�|�=��W�UZ��X��Wc�����?��o�������~�VӇ����J��)�u���7a��
�yZL�CTR]=K��y��.�aɦ�{v�����幅��t�nY�',Y�B�{�x���m>��6����/ף�WE`F��3t�.Vq�N3!�ٵ
j�S�߽��n��aT|���U�TQ��.�wU����h���� H �`0��3Dl�r�3�y�x��9�T��T�]e9ؔhe�]�����fk��X��eM��戓P�è\&P�Te�
ǘVY�"����U<ӕ�Ehon���S8��X;Fȑ��H0�p�X�>�C(�y �j��6�:t��FF�J��5Cu7�&��й,"d>/�څ�8�Y��l�3PkJ�+8l#���Y���ס���1t0e�X^(���n���oےjo�"����cG�Ҭ]�mw��=���,���=�Z�~	���\����'���|��~+��s���(��sbI@�<*�^Uyh�+M�+�=T�Qm�[����Jn\�oj����j�Fn�*�?�`��X�J�S��*٩ ^��jGB4YF�A�Iv<�"���e�0Rg���(�5vүq�5�`[�M$����,v�ރ��y�&�^7]O�t����� ��6ef�\I>#0;�D�l���Q}�(R��!�[R��H�4�n�+���g䞨7f��1��gdϿ��P@����ܓO�uiEZ��ϳl@r\ �u�0{����-[�o����:atN�(�i��"â$h�wu0�� =MNdW���5!��K���D̢E;R�.�����O~N^�����x��P,����L!����q�$��9�E���ވ��G�����N��,�!��O�
I��C�`���p�w/d����{�Y)�z���K@�!n�+����/V�ط���~���o��*�d6
%����&Kimvʻr����L�p]#?Ւ���a�s�m���!���c0~U�a�/����#�9��Ԫ��� �Y�ju����;2�}����\-�I"�L	�P�%L3t¾jw\�2ڕ2Ｂ��
SޭVPk�a��M �=��Ήn�]�O��~��Fs6��]��:\��$K�1\~&{������FN����w'��.��X���,/���4��z��A�����2�nN�����_��e�*K0�m��95�N���è;e'�eI%׫�I�[���e/b��cF�R"w=u�%��j`<���lW/R��X�B�uJG�?�7Q ]���r)%�h5I|�-� �M!��tU�њ�ZmQ�Y����F���N2��o����x��/V�>�GJ@eY���J@��C�엛8�ԏ}�#��凿6�3���	��ɜd�My�Sf4GD�jiS��jOS��h�;��īӜ��Fj�^�1�[��h�(�!s����"+0�뚒�ի|(e[|�������)�f�n������<��%������/��t\aG��-��&��Y�(�:|u�3��m°.�5&������Gc��v���P����e�h6��
°�o?�������bsu��;���5x������rw؏+�]��u5��Y��&|�a�*���չ�,�t%09�A$Z	���W\�R�H}d�ْ�m8-���@�r�T����6\�w�0*WN�$D�F�
8 h�
��e�S�&^ ����x�?Ce|T6�p#G���H�L�Jֈ��������7��C�T�#	���Iz���܆�U�����/��w����x?~-.�����1�g�������?�O�r毾T�/������)gtn�5�JזSKzJB[��iy�85��l��t��*�p��"����]߰�+�p�����yut%$�� �8� #���	�(��
�d��DU*��ד�O f�\�d��&�=�>W�W��,���3$l����cR�ڶ+$6��S�Q�8E��(�3�v�Q%&�;���L�3��Q�UP�*2�t}cC�U�@�u�ř����n�S�(���{�l�G96��U�kɣ�yi'��n<;�t}^�W�������L��%�U�o*�R�J3@���[&%�{i�[ֆS�Խ��n_T�m�|Gժ�U�/������%�"E,^��[���(��xnt���Ћ��W�����<f�RX�#1�P1.@��G����ߋ�������ΥyGI��N����i���z���<z�}uOe�����ڗb�+O =yhpNu�S�84VJg��2�6Q��	�LV����I�\E,J�F�T���E�� �����>�"E�C��2y}أM��C�п��,c����:d�6�L��?Sךq'�H�7���'�v��-�bE6��3U�ۮ$�ͥm��Ϸ��+#q��dq�S������](^�37�<0K:�է>�Q�B4���`M��g��-dlUc����ԐcEa�"oaӫ��8��!�Jڊ�1��9-kJ0�*-#��s�Ե�xEJ��iz!�鶳�!)��߂�.wTj��`��S�)K���x1[ ��b1,e�'ϟ�K���"5�LDѱQ�#�Y2潜�^�Ez�R�v9с�����o���yӨBH��=�C�0��}�,�\�}�������O�G�|�xE(����xS��#����}g����2���p���t�2��i/B��Z�H,�����IW�� ����R�M����G&�qD��Y�G1�Mj�|WA ��j財�X	��i'B����@f���- ���ޛ+�U�X}(�@�^�E�M��)��4=?��`��B|/S�"�"�%i�6Rϓ����
mJ͍5m���$ئ��������H�{�I�����	l�=����JVS'���2���4�����2t��GRi\=�� ����8J��11 �8��O�D<�L�S�Xl/�ի��O�7��EC�Ӵ�����#�����h�c�W����dd��rr���@��ʺ2�6��(���MRV�h�;�X��Y�L��vK�h/�sP-�:sA[k'����m�UМ�Aui�;!ٹ�����޹��}�dՍ��W�]�@	��u�>? �s������o�����K���K�H/���S��>�v^f�J�4�$� R�lk�F��E]X���(�˩e!y��`�����yh6�0G��Z+��s�)L!�1ꥬ*����mʟ�Y���5�)�U�vkC��x.�jg���aa��\%�mnn"�By�ȤF1�V_��~H$�x����ךA_"i���Ps��mV��ttx���2Z���"�dK���5�����I�%Y90F��I��~�ة�����!0|Po�����N��^�+�tmի.cM-M�x��C�@�JJ��.CZ8/�mv�@���r*�W|��_уOD���`+V�E*G�6漾��Y�$x����dl�7��t�62ރnO�S: t�����"%�Q���Wd9������s�K���-�=)��̋�(,4:��V*y\˒2� ��Z}��C�{k5e�4Fo�%���09�8��m�*^����xY��z��%�}�A�������������/�>w�����^������ޝ'���_xۥ��x��;A�dy���p�LX̌>L�cY/�uO�c�V��^�¶\A�0��9
�J�(��-ѱ0��)�T57I�L�\�܍ @��Tڵ
�SQO�\��ϊ_��(|��F '�P���HM�h�֐6/���f�aï����������Q�,������d#�9�I$;Ǣ�U'A"N�h�K[9ea�-�P�/ѭ#���ܐv1��8"��q��X۔��!�� <�G�^���i��]I��u3�����rE���Hz��k���ʲ�q6[ey��,�y�{�eX��܈�Ԉ�����Q�Np*��a���j�L�4��0O��a�8A���a�h�N�c��m��OLLd����m�y��ٮ]��z�aEq��6[l���,�{�~����o����$�r�a���\�6|�j�c= oKjԖb�6�w����<M�,M�ܴ�s}�B%;�jx�H�4�+���h�GYy�d�XH�Ȉ��G���ǰݴ,��h�e�i
/�6u+��l�ˌ���:�ͬ���ϛz8(�� 	�Z��{����*���Vb�6���~�a��t*k+�������|�����v����x�����x����h��Wp�G�'�ep�����|��8Y�7ͬ$�̸XvfYndF�Դl��cY��1M�,�����9#:���z���ڔH��-KEO�0��^a�����fa�'���yF��¢41���/�8nnC���41$���<�'Fr(	?��=��ۮc������i�΃��3�f�EI�D!�(5,�H�0D��.��S���4�T*���9ACν��J��2%L��9�.���Ϋ%M3n<I�)#o�1<�'�f�~?��a��y�O�ܰ�GDr���Y��j!^�0�U�
��I�Q�f=�[q�f�m�j5' %I�f4��s�y��r�r˰�x�!�wdF�N��)309��u��1�����R��i9�N�:=)�;���Id�if��c�yb'Ql&q�������/D�<�(�����v�kڦi��m��='#'�cG�y�I\�
m��,��\�����.#�"�=,��M��&�y��YӾ����;Y�R�l�����ce��D�����432>��F��&	�ku��<�l3w[��ȟH�,��,1-+�\75m��]��]3�"�33�����4O#r\;wk��V�U�^qèw����7W:����������?u����w��^�Ʒ@	�7�=��>�쳞���lo�ҮN��`E������gN��57[��]We��L";�2rFVAh�Q`x��Z61=�-ˉˍ��za����K�qν��ߣ�YE�C�f�[v�ǱА-���,3�$��^���{nǺU�d��I�o�c۹e����\�Ź�c����$Fj�Qn՚5�s�$�M�ô���%������5�$5�]���;inA�,�M;M�*.�wtkr2��45�0��8�#�x3�l7��q�4�,K8�$��԰�JY���v�؂e�F�����-��Y^�qf�F��f��>O�c���2L'��ض�$gt�ش;�y�����5����eFB� ��\�G(�U�#B�U��2��b�S�Jy�����	����W|Q�ct���i���gq�Q�5<x�������Æ�EIbĩ:f�jQTN��]�ʍ��h �&F'�f��]ͳ4�k���t��{ >r�|]P�?1x���Yb��5u|�)Ni���l6n\��^��$�_���=�v�9�G_n�;$QRA�tr>�����j��K�<s��j�"J|ݴ��xQl���h_>���
�Yͮ�Ks�;����;uoI奿J���*x��=�?g��zxn�Dm�B�.E� ���!m��`�5G�&Q�.��$��ɜ����usӰ��*^�gi���ѱ���2,���e�M�S6p�/��E�Uן!v6
�le���H#����[nC�nO�VMs>�β��P�!��=`yVϳj�00O� ˓�<�M���� ��#'I8`�ٶgX�\#]`�9�ʷ>7�7�v��$ٝ���p���0~|��s�)�s?l������Wq��%�J\��� �檪�\W{�S/-PZ������K z	�ں�J�(-PZ�����7]��=��u�1��v]ܦ�$K�(-pU(���T���@i���J��-P�����gWZ��@i�����%�_����(-PZ��@i�׷J@}ߟ��J�(-PZ���UY���2S����J�(-���� z�v~}ߤ��J�(-PZ�UX�&�2Bk�|ki��� ����w#Y� �M�*�H������J\����Y� �_?_�Ii���J��Q,P�6w��8o��]^Gi���n��~����J��.�us���f(�%/6}	��l9�\Z�����޽�F
Q ��ь4�%R&��]���u��ҡQ @`��@�g�x$����g�.	xc�S�z��Y<�t;� ���  ��Zx�ܺ����ک�* лv^� PJ@����9����+S�p�1�Z2aA}�! @��n����*�L��X?�t�Z�� |H�]����N{U�=[# �G@��q7+�* Чr� ��{��J��� ��w���ys��nu%H- �S���	 @��G@��	^����%�|M����v(  �4Q	�U�?K~%�~�@��A�'@� ��� @���O�5��
h. Лo � @�@�^���h+��Nm[�p��-A� 
�MT�� <��s�T�>��` @`��@��nV 0U@�O�4�# ����� ^8��8�㗟�������3d�muG�� 0C@��P4�, �77�� @`��@��h�}�Y�73�z�vX�bn��5T9�z��X�( �/B�8̇�1u~c~�&@ �@�@�w�η�\�j	 �] i�wo��	('ி\KW$�W���@*)��]�Z@��n��	 @���@��Iu @�@k�޺��'@� �*�J'�A� �z��+� ��*�T��/�=%'�K��Y.0�ܜE� ��=bW�� ��7�V���*i� @���@��GU @�@s��|(� j�}T|���R�/�跽⚊ �J�y��qg�*� 
�
��S2�+*�}¶+	 @��3�P���g @� }����-�&%@�@a���.oO� @��U���~�R� @� ���ps�F� }z�^�� 
��͍T�Wǻ��"�F PY@�W�����ͱ4)���Z�}c�Ol�'j�!@���@�y��~{�v�$� �Z p��v�x �T�V���t� ��
�8�VB� �
���&#@ເW�	s�G� @ ����0�X�����d @�����Q	 @��R����d @�����Q	 @��R��@���҆�� �$��IUg��^�B%	H�!>'胀N'@� z�.X胀N'@� z�.X
t_��w:�$0��` @`P@�:� D�t�ÈWXR�/{�l�E5��޾d�[�  � �ۍ��*�    IEND�B`�PK
     ��Z�V]{[� [� /   images/995ec925-f4ba-4c8d-81fb-fe52a7fea57f.png�PNG

   IHDR  �  �   ��ߊ   	pHYs  �  ��+  ��IDATx����%�u&���|{��+���wq)P�P%��hfB�FҌ=�1a����#��v��8��Xֈ���"A� H�+�X�k�km�ޖ��9�ޛ/��	�� ���|`�U��/�ޛ��;�I�P(
�⪇�� C?
�B�X�PB��d�P(W$������J�
�B�P\&�Vd�PBW(
�b@	�e��g���@��)%���n(�	J��ҿw�׆B��\儮��b�����r��B��x\儮{�B�P(����
�B�P0��
�B�XPBW(��P\2���.gT�B�O�k���E(��3(�+
%�kJ�
�B񊡚��ʅ�B�P�b(�+�\(�+��a
��j��Bq(�+��J�
�B�P�(�+
�B�p�	}��M��U�x��/
�k��N�f��M���(�d����e'���J(
��
��+���B񪠲�B��@	]�P�R�d�xY��wi�맄�P(��%�K�_?%t���j�:�BqC	]��P2W�;�)��å�2%t�B�X�P2��p)�L	]q�A�
�B��h(�+�<(�+
�E���jb
�B�P�&����d�P(*P_�x�P��B��b�d�P�z(�+
�⊁փx�PBW(
�%�W%t�B�P(���
�B�XPB����
�B����~B�\�P(���W<Ԣ�P(/%�W%����
�B��PBP�Q(
ŕ%t�B�P(�������[
�
%t��b�d�P(�P(�+
����5�)�+
ū�6��~o��B�P�J(�+�$(�+
�B����P(
�:��B�P(� J��P(�+	J�J�k�7�G��ꡄ�P\,�eR�V�P\PBW(.Jj�˅kY�T�,��
��j����%���P(�T�_�PBW(�k	J��J�
�B�P�(�+
�Bq5�e�%J��u�)
�+��l�J��%s�B�x-���P(�u�k�����P(W�V:�r�}e����y��MG
��r�j݂��q��G�J�
�B�P\}P��B�P(�p�.J�
�Bq�B]��,\�K�2�~uJ)
�B�>��{������!t}V
���A�`�+���
�B�XPBW(.ԙ�P(^k(�+�J�k
*��.PBW(��J^�C��u��@��t+�k��).^Bק[�X�Py]��b�&w�B��d�P\1PBW(
�b@	]�:B�
ŵ���߻��}y(�+^G�E����k��]��塄�P(
�:��%t��*
����%t%s�B�P\CX���P(
�5%t�B�P(��QBW���>�
�b-�QB׭PquC�`�B��(�+
���$��PBW(W.��j�{}���P(�\(#\]P�B	]��������/�B	]���d�P(�(�+�W�~(W��
ū���BqeA	]qUA�����
ū��⪂n��z��W%t�K����^j8r$����\#AE��L���n����%�l�}9�F�^�</,�(l�e�l��ay9�޽9U�K�x���N���'�`q��P����:-��dV�����X 2˽Fb�Al���l�3t�!�oװ�ǌ�X�z�8d�|b01Q[H�q�%Q�&Ѱ��Qd�4F��4BڎP��Aױ�Zn�I�n$#d�4W�qD?1�>ͅNݦu*&�<Ͳ��kIb��Lб����8��ai��Ȥ�����V3/z�����f����*�N�̑�2dt~�n _��o�40F�in�����'�-g����S��ҟ�i��1�5Yv�rh{���%�,�.��Q��{_�$�P\~(�+J������������̚M�O�l���ͭ(�X��O�i�;͊�I��3��s�
�f9���Yk�Ȗ�K�<�����>Ki�+�Il��O.��ʭɣv�gF'G��4�0�M�=";O\�y
>EL,م��8:{~�.��
���8""�3��P��8���.,3/E��3��&�m:"�Nj�4|<l�X�k���F�%9�	i2�5Y-eH�gy����5�2}��Ւ�ׯ��zR �r:w��Q���[��(N2�D�$y��FEnx���5����FEV$�d��&���HY��B|=�RfLy��W�s�|��vk���#Z!C�llN�Q$,sE'�d��|��O��Ɔ�YQ���x����� ����^B�O�#��<�0�G�<��YKk����k��Ț��O��l	�{�=>&k5�E����	]���#'X�Ԭ,�`SKl�K���4�4��e�c��'-IGy3���C�Cc�׉���dvf�U`�/0�,������FBө��ȶ[�ӧ��4}�	��w�ar�`�T�������5L��̜|o�b&�t���Hh;����v#��?ԁ��)�t�Vp�NMM�͎_�C�x���c{<K��m���뉖o'�����Mf�Mn�zYg#�i�(�w��l�ĘuYC�?xc�u'��{y�ؔ��^l�d����[Yޠ�bQ�yO�ì�}���^�%�w�]�,���)���)� ����A�ID Zk�5�V�eÆ����\J_,�(��x^�x�7�^��ȍy���sJIV��yș�!�ŉ��m��e��X��uIGn2�����s��]��x��{<<b;y)�y�����.��q���ؠX��aQ��`4�¿��x�����t�B�T���#G[y,�w�M�E)XL���'B�O��|k��_c���ΓN���&"���pH��u6�,�u�\����Z:�|a��X]:M�$�>}��E��]�ű���4�����kS����Z�\֫`���&a�l!��D�,||�D�˸��,d5�YsS^ԑ���{f,	 Ku:w�Ғ�_�g�d�o~&���L�����g1��z�2���4��ɸ�*�u3Xʟ����4��k��P\"�Я0\�� ���n���c���m̷��9EZ�#b�оe�d�ĕ�"!<c=������?���ܑV�ɐ�d�
YŤ�N
A���M���=x�g�a2�E��y�9Eai��|ޢp\	1��4m��"�YQ��`h,Q���`
�$gQ�-�/��f�7]#a�DDD1�k�56��8x�5s�C?m�I�= a�G?����Xs�s���R����H�w�J0��`*�����������㈄�1<v���d�1�����`فm#EX^?�����2�]GNK�������~b��Gf��� G�.�b�:�lg|�؀ӏ�"p�e���as6ː$IG�z$iM���-���ԥ��@�)	'��I�/�6��tҬ�Hr:Ao��Ӊ���#:��Sd��0�a&t�]�FjuL��~!l-��Ȳ��L���]�	4?:�����D���Z4�l����l�Nfo��M[���Y����ڹ��ǡP\�Я0\2_��?ܲ����v��S-�wj�5��B�Q��l�l�drVt�l�q���@�Vޜ�m̯%!�F��i�f-������^�dӗ��;-��W�>I�Y�^�?�X��D蚤xY��=��9��>�uy��^f��k�����Xl0�y��<�б��@���_?>"vb�B[��%be��k$L��%���6mLLM���byi��
�9��~=�I��u��u7��(���"M�};�#lB�Mk�
4k��u��>�Z�E��ƌ�-�ױ�0� :���Wc�d��C2+��Y����[E�u�Bg��,p�{^�w����<EX���	N�4b%r�'��'�V#��xW*�,��5g>rK �+�_�(Ș��B���,P��s/�ƅ���W��(�H�`�	e|ܐ��sj�&n�}����mp�
ū����~t䩧~���Ξ��x>�%�9C�WGșX���8�	��	��%tѸ=���W��eN���l���u+�X#5��\�)���$�1������[�IS��o�lەx5@�T�M�w���5!M;h��@D��Q�5��.
m�,��͉5u77����n�h�YR�B�֦V��;�D�t�c�#����r��A� x<��g��n�mG�|O��z�['&vF"��{���*E1����1�9�>[�i�1�;	�/�����>�_[x2����3|nF"���k�^���r�8��/"��^}rG�2�S%Y���P�3�#Dh��l�����P�v>�X+�
���ԻM�Y@>���Z���P\"���d�x�7Y_X��� 8k�O�m�Lǲኆ-�M��F*�s�Zh�J���FY��@L �ԅ��h[	b�Ѹ�6�:��9�+h��?7��r�R@Hr�Q�ǁt���۹"�X����&�p�k�l:6X1X��ՙ���
�u�ν�f��O��b O�i��]��1Ss�u�oR�k�׭���5��y]�@@Dz	4~��@T�b�S6�D:�;w��������k����G+<����B_��c*kh�~8N��%�q�<r��G8a��e���g��h��d� s7�����Cl����ք0�p�؂O�[ny�{/������Nw|1��Yx�B~�Y��C�CT4h�i޵���2�[��~
�%B	�������Mf�~1��&��ah2�ɧ���s2"OY��jQ��C���t�v��~#���0#������{Vb��m�kbzf�p�Zt���ySb�X�����e�D��ǒ��N�4s�^�[�C�q0�(ʑM�M�r>��e�9��w�b��
�� #��X�4hc�Ӳm 98��!���2���'q&>FB��8f/Rʝ�#� ��P8a�����ܤ��Ow�@F<~#��sl�~��o_Dr��i���'	��[	�����H2[&��3,��#1
.	��o6�"|��eS~QDb2/"��CP��\��@ƨwx��0���8��\�J2_l+���g?������?rB]p��"�^wW�b�A	]a1�R�ەDL���Aa�ռ45����${цB������kǞ,�|+���-i�c�26��n׌jpi�tq�p1���N_��qs�h�L�6�a�L�N���y�fM�c��!����Y!Bް�u6�;��hz�<���g���=G�`�Zc��n��_1S��%���G��/�4gqH����.��i�����V��|O_���=�H������7�˫)M�n<��Rk6�����x2+��)D�E^ ��9�=g"����bH`1�Y��y�s�g#��u����2	��4H0��Ʊ|�|0���3*|0�{��#⋂}	�7������\�U�y�Gd�Zy�Xf qg�=�R�FJ�K���x�%�k��L�i�i�Mr��;--��a��tH�Gg��f�Y�W�Ȝ�Q:��i`�7m��H���.8�7r�oD=ƀ3����S�P�᳾2��E��B���u�E�7��Q�k�a�f�
L�}T��o36��a&�u�I�;�I.�uX�UEa��T���ڱ@�Cfm�O��x�����3�G2g[�%��	���x�	8p�����<\�a!�u����ג��/!9a�p�:
lD�q~�~ܶz��`"�������L�u��+v��S��G�4F��̙}to�l(V�Ȱ�<M�.�u�I���YNq�A�c"`�2%/
֠"Ü���p��ݜ��Wo����g͂)��1b�c�Y�����ljP(.�L%tH]����R B�p�U�}Zgˍ���W
O�Uͥj���U5��{��#�͓��䬥O4К�DVoK�V�ӑ�t�#"�k�h��VG̮U_	bbb����E֘t�ܛ{�<kĈ+CgFgM�]�P��He������99
4^p1^��ķo�S��.`�7�����c�÷����رA�6kX���u�v�VS�؜���J�(G�m�\��GBͷN�٠��i]xMz�!��O����s��ڊ;��\
�?7����ŕ���}t��D7���lג��hry���ROP��4b�$��F�F"q 1��p$�{<ǔ��F���p�d��R!�ob���1�^�������^��������`x���?�E!���XV��y�aH�LI�L�x}�Z�]WPB���O���E\�~sI;�nc�g�|�ba,�Z)b���$*i>6U�l�a�BB����4�U`���v����m�Ы5�7Z��9m��p�k�9���l�B�l�Dˍ� F�\�{$���k�	MB���a�x4졝�� �ؐԐ�w�t����i�d����r3��vW�k���L�B欠��:��&t=&�aDDN�]��!ٺ	��0j%E���Ľ�D�[z-Q�t�X�.�Ed>E�ӊj�� "�u逎d*��0��=�1V��F�5>�-�Yo�^NM�	��O0j7�%�нN�h>[1�s;:�6���	.����
��.��%��Ѡ�Ի=$K]�+�s\ݟ��˼b�q f���Q�b`W�n��Cf���T�i�$I
�s\���s��w�/�1=u�j��)�3�Яqp޻��A]x���H�F
�8~r�ml�v��6YN]��!ʕ�f�$��8SsAZ�Ԯ=���6ĭ&7lD>9����LL ��Q�'I�	���d�D���/y���41�g¯�h�m�nK�G���jD�q����Y�������i�˨e�Hm�)>:���v�(e^�eB�&�@�BF�	(9|M�`43�d���v3�n���af&�Ob�,,bx��|��� ܊11�@�2��r��!WW��q�̹N�2�.��A/�տÈ����]3"g�!"ܠ�Y�б}"�s�&oًMw݅�[oA}�n`�&�Cs"�J���>����X<|�������i��~��op�������S��*��+�N���1�S���j�YS�B) k�Y������Y\7h��0t�]�}��Evq��Bq(�+�Ffr.�ũO����~c�k��4y�e���YFI����gF�|yی�5l�M/%m�G�^����,��w 7܀�[� n�]�W`��$�D;C���N��]��!&�Ѱ�>i�\8��l#&�W�0i����$mL��r��ϝ�P@��Bdx��'0K�1�廂h�کc��6��U�&k���z�y��t�����a8��҆�����.��|�o����M��^Pi���F�g�4�{�Q��cX|�:&E�n��0r�a�1�������{?� ���p!�C�^Z�] z�}�\��н�5��TŞ�|�-�y�=���7ۮ'���ܐ0_
�K����{��o�����q�����x��q�~_�0K�iv#�h�y��#����^�k�B�2����X�]~aН[=ʷ*��1���$v�f, 6�>goؑe��Bq�PBWH"nۂͿbiDmBAW<]Ҿ�8��zSyt���:WY�T����pdt�v��!]���q���I���oy@Z���,..b���㇏��GƓ?�z9�t{Bߓ�k}IujMt\P|{zw�u7���_���nBc�.~�'�����6v�	��Y�hd3��>�YW��>!���#�RW�ãh�g��Y?C�e0���'gq���;��������-��|��s+X<s�Ů�h�l8[ ړml���Ļ߃���ܼ���}8����c'Q[XBF?t�:0 ����?!�c�3)M�ុ���"�F[��A�6�z�$t���a��|�o}�i7��:�sH�b@�_"t��V0H�bj5ꘝ!�톽h���o���]x�s_Dw�"����{.;a\�nL�~\!���<�u�W_׼W���?��� ���U��_J���T��`��2�Ӊ	"t�/޿�⢡�� �M�m��`"�2�T�H��VW&K��2ƙ�5ڌ��ֲ��Wn/�R5�zh��>�=�)?���b�?����8��œ����~G^<��'N��^ĩ�g$�A�8�]׸�j��WGB��9��~�/�n��>�C��7��]��ǖ��58��8��S��H���)�C��a���xy�u��d�؄`� vP�rə��#�r�b9�+�`ȚZ�Q����)#���ַ����0pۭ ��N�ŏ�܇G�|��X&2�/u��G��W093�Ms�x����$�ܸ}����1�y��gi�:$��K='t��CW7�G2|��!�݅�+fg����;>�+�
���N4���;����ۉȉ��D^/��_�r�#8w����}���s�s?�q[��{�wߺ���o&����s8�i��A��=@\h��~�ev��]5.[�	3�i\k!�a�㲮��R��U��ņ,�q6C�C�BRp��g�gF.��������B��[���$P�2݊�}��.X��>0���O�r��x�t�f[� �Ւq�Ir�+~)8-'���j)����~���Ꮉi��>��/���`߳q����{�N�?x��ZML�&�e�6�~����[��4z&vQN?��y���}8~온u��=�c��G{�#�秎�Bc��iN'h�]�qu�ԗ�ul��8\.�W�s+%G�>2\h�~O��Jݥ��82�A����:m�wZ��k���� ۶ �����}���7���3�{�-�A��]w݅]�vb�4_&����8v�8��y|�k�ė�~nڻx��x����x��������`��s.���ڴ�zՈ�H���ؗ�n��S/(t��C�-��l���-�~���6�G�}��?��<����z�}�n�6l�n#�$4�&IC�D��=yO=s��������c��~�W߉�t6�~'^<q��0C+��Y��p���߁���*˕"���N}�����|.Z���~EeM��U�M��!�#W�'��/�3��Ñ1�tMy��⡄��M&ᜣ���򤹾�����~kW:cmP�Z�%�T�Ċ�q��� Mfvv85��z�zD���4I��aff�4�!��f�������cǮ��q�^̐�*MV�yY�����3�����>���x��aH�럛G�4�t��ÅkH��dI{c2�&�0�»!�p[�m	o�ʲJ���w�����2�wjg1n��{��c�K�wN:������������F������7ރ�;wbfrJ���Ͳ���k,|����̩��������~�����;H���$׹E��Ĕ�`��ɚ�gVpx��J��|P1SW"�B����4I�oL�q�&�M4qۇޏ����Ñ�����.~�`�3�w��]�������8[��7o���Z���M8r��8���?�����oNM�M�6`��I�D���բ�\�IGh��s��x���T�A���b���"��g�e��,T�o+p\��ypyy9)�K�W(���`�y��uN��.d�h]����j+$J�VԶ�u��Ff�K��آp�Y�R�W�t:BFBkn����f'&Npn~��܈?�o����w�nreX�H�/['���m"�m;vb����ַ�'H���������"�9&�5���˽��!"ϰ�]�b���C.���\	ې3�>�LҘ�V���X�zT�^G�I��l��[���>
L���Ï����_�C���[�g���[�xi���*�V�{�s�G��͆���y7ܴw�s'���O�o�#8|wҜ����H�j6��mh{�3��)�W�ޔ�{�K%(�9W�kX$�w�q;��v�~���-xn�~�_�����V�>���λހ�A���h*u"��369���	q��܁[����n����X>~��s0��Gt�M�:-.�;Y������4�x��;�0V��]�{��``⬯�⒡�� W���5��<B�i�+�TM���Z����J���]X�ɍ��K�k.�椁p��qI�靝�i4�@k��|�;�_���m�y/�Dl��F\E�/:���HjΟ͟���u�w�ٍ?��?A��ė��I3�!�[��T�������`�r�Ǝkл(oS�Ab\z�.;�yJH�֙)��Q��v���[?�!�/}����׿��� oy绉��{lٱC��tC��k�i�k�ʑ�����H]����;����a��,����}G����z[ZML��ù�4��O\�B���{u�aI��f�*"�#�8�G�Ӎ�h�r��v�=;p�ȋ��)��G��?����?,��O���{���6W�c�ɜ�Ⱥ�}�9w�X�q�k��o��v���7�S���xa�$��s@s��kq�}�4�,� �I��c����?.���!!8� R+��s��29�_�)@��@	]!M��Q*����.r	�*_c���YaVk�k����V�eK+,�N�����i�n���1�fץ%�x������o~�[%Z|��s��k5$D"�x���z[��Uo��������z�6��]��c�=�C�!g��I_��e��%�}3�D�-P�ش[���Q]���,���p�$��I0�q��{��.����_�"��ӧ�䳇�G��O����w?��f�#�}�S�*����ӡ�dl��qyq	-���܁�&�j_���O�#��@�E]uX����J�����	�����r���%��`��`%&!ez;�ؽ�=�O��m|��o᣿�1��?�C!�n��ٙIѮD�͉)�� a@�p�w�f���~�5�jM��~3§��_`���젏tͩ��|�u
	Γ9!�k�G���J"-}節�_�F|�I���k���M����%�u��kښ�5���5#f�M�쟕�~s\�k�K��>Y{�f���^�Ӗ���7ő����_����N�<	�s;ySӳB>۶����o�G��mo��2�#��Fd53=')j�����้U�;s���_BZ+�Hgr����S��<���3ô({�K�:=��nq6G��q�P���>���`���m+n�������}?N������5���>F�&���8k4�,	�;�X�U'i�����He�$�q�NWÎ�o����?Ewy_�����.f�5Lq�(A�k»��֣.��9��^��#2�Z��(x�}���':�La�]w��[��������n��v|������9zn�LNOæ1��Vz�ι�<[iz�b�c��@��?㬅<��s�w�#x����>�g�܏mɊ
s�:R���Q4n�j�������4�p����� �Y�7�xq:=��uQ$u�E�E���,���������e"���x�D��Cq,)iy�S�aB�uu3Z��o톹f{*�_5��L���>��4�0�.-��
�H�emƦw�}��k���ˤ�����iӸ�ę�8�-���q�>�RG��#���w�ox�]8x�i�����S�<�]F<�L$ąn�J�V���ȷ�����e��	sJ#2�ҧ���������ןÑ3�ؼm~��~7�|VFd��6ZM�+h�'$ ��KZ���7u"1��L\"��p�_������{n½�}<����cO�4��V�~k<o^Xd�@;�R8��}_�>�cÉX$*�-���8�;1�c�7I��w�3�D��������]��Dd;�e�6m�9��~�"q��N����(<w9i蹔 nuZ��m��"�}�wp�駱��)�9m"��i�,�������)U����\���&�Zy͆!A�
�ѯ�=y}��2��X�u�b�i��ä��oG�0�h&jgT�֭h7f�K���ƚ�m%z��|"aͭˍH��XJi��m�3�������D�=z�f�H����\��c����(ؿ̛y�M�i�Q��x�ے���ؽ7ތ7���x�}h��˒���PV
�F&��g�uq L�.(k<��.Zu,���16�r�++x�H��x��x�[���h,���s��lDڛ�|O��͝��j �I�H��>/��z0�h=ZH�)v�~;��[���r���e�ڸ�����}4#�1���Y�o��%nC�v��Q�O�f.l��;c���v�+���2�?��;��mo{��mO	�3��i�t6JڠX.z�+o�5�NB? ���1��y/Q��^�%l�tz�����y쌚�L��܇ ��ڈ���<6kI���}U��Q	J����&�X<Pq��]Q,�Ƒ{���A�YB7���A�쌠P\"����-=��a�aO+�}�e11��gF�rm���Mhw����Ľ��+Q��CNi�n8����7o~e��M��{�����A��"�͓��\�̻g�ؽ���h�V��E�����5�|��k�ꢻ^6� 9�z�KU�A��|��6��i{�y,-��;��Wބ�ԤktB��f�n\d�O����u����	വț���O�kp�.W��f�p�܃M{vc�Ƀ8;as���4㌈�AZ�H����8�Z�6������g��3A���	�}��0O��ɳ�$8�C�y��~�̝+�%B�C���ȝe�<q$i��P���HZ��U~���I���'�}�\w��Z���sgq@�(�u�2�g���?��ၫ�K}����z�{� �?B�99??���gs�[�����`���T�Ƀ5	Vx��m��_��l?Z}��w1�^T�5�i�ؠV���{ވ�sb߰aff�\7�ܑ���n\L|��:��o�����d6"�n���w�^����.�8}Z�!��X> ��1	��r!�Y��W>��픎_!�"�:x�G�_H~���.�p�֘��8�#�;��V�.�y �g��`Fk�_鑆���N#��'-��6l�a/!B?��ō[�����_X������ZH�r���q���D��w�}����s������8s�Xv�فz�.�r������{��x��Jr>�o���e�%��M�uW
8)"9��.�Zؽ������}�8V��0���uV�T�8ܻ`KW.���g~�p�r�������{e��W;�����"�"���o�Q�h���\�&8�{��������Bt����n�:ز�:�ƛ��dGJ|�&vJ�g/J�]��f�VX�v�;A`���[���#�Y�ʙ�]r�KLh0c|e{&��T�%!f�J�)b���j�wf~A��ݙ+s�9J�}�V5�.\���nA����:#@xYAe;���9lݵq���a���&��-�$>A�����~�*�ɔ���c]:���͛�(�,�4	B�I�q�Fq	�"\�Ć�~�ӧ�ٚ�ֱܿ�МI�D:J�>߫�ߏ\���Q+ƍu�ߵ�v[�tP���� ��A�!xϥ��Z���9� �^ ��g����0(#�#�
(�|��*�6�Lz��Ҡ�~�b�z�B�\@3�HOqo#����	�
_݇eI�m&S��F\��pf�ܧX����甶N1ks�����.��ݔ�.�IYL�I��]D�k��LLL9�P z��:��X��>&L|���ged8#�������o�ؤ��""��0Ɂj���W��tw�	�k���L�l����O����{A�-q�D�^C1�#�d�������ƽ���![^�JRC�}�l�'-�7,�/dmB��)�fgMI�����fn3&��OsZ���&�����(�&p"w�.FCcN����)K��w%��\A�� U7l��e=�~5:����5L9�ͦ�	�z���ɘ0����c�vR{%�E�^֏��zpՔ����ͬl�R�
5�+.J��,V�h6/u4���=��r�8�M۬É��6��m�$D���]ָr�|N����а�{�e�`1&��i�<�p��Ӫ"i�Q���}�]���"���׆}]_�;� k�\����\�[����D��ڵW�"�$2n���w1���n�u%����l��qYo�w�ϼՋߜC𸽙�?��rGe���[���2�I\!/jwh�Hh�n+��y�K��h��Mׁl�6{���h� ���J������$]�OCnHW5He;+�3�D8j^��3����	�HA�w`B�sq5:N]c�}��N�����M�����(ōZ�ӌy�R���5D�_�3���� ��fr�z�U�+Q)�P�Z(�+d3!�6f�6��X_Hi(����ꙝY4Ц������ވ�Z]L���>�:��7t>r�^:�=����c��4�#�fg���v���q	N�c6i�,,Hnpå���>�M�u�*�,2߉,
�~܋KK�1��IK�,���N�"+CDd[d�X��Zg!($ 0E�;w^9�,�/.�d)i�L�V��:�}��arz���F4Μ�4�I.FC�):Q0�{WB�<�>��}v�(y�LQj��Ҳ[��=�L"itn�ʟ� m��r^�>�Ǿ����E�͍�!s�߃B���B���'i��-h�Ə�{�
�V26���+�j��U�R�/_Q7�{��t۪#T(^���H-H;4]lM���:�J���Y�p!�Ț�6˿�)|�������f֩Δl�Y����\�#��*%~�:��;��ƦX1�F���d.�������L�\�� ��J��B��9=�/��!s��$"y7�-�|yτɚ���,&�S�N-�ù�sDR� ��&�K���\������ن]�eA��X�N\I�8����ZSR�$�|����O�O>�)��#ܔ�y��E�WRm0�>�i�AV)|
�ˀ(p��1dKK��Iw��XXX����D���.���B<9Jˀ�;�(5��# H���ƕ������u�Qg��
�~�܏�?Q�uc���"mq~���Ǽ��Z�C�|�E���$���"w?\�8�����+�aU\�PBWptTJZp�EM%�'�!H�Q��΍7�V��¤�R�DE%��j�g��Lx�Dd���H��Z���ۢ���]�؉Ӥ�:���7�z�����T�,O�2�K�Y��DB��헣�SO�5IW����,c��O��ѣ��ӄ��{�e�;[�4m;��QH����G�o��Kg���`�֩�p���(N�[�ǣ���쩓8t�)��{�-U8[,�����Y!���m�R�
�g"N���Ftψ3�-���K`�0��z�<�CģЭ�ts��-o���q��x�#��iĥ��[6������zG_�<MZ���<�;�;��珻�)/kX0I5<�JF� s�k�&��(/�,��R���S���Ν�p� vT4$�����ݴld��a2���v0q�>���5!�o�s�Ve�j���{��R��%#yn˪{|9�)�[@���6�_WF�|�C	]�A�S.n���H���9�c����h8��#-B���[>�zm0bga��Z��2f6o��R?y�8r�0n�a7Ws��Z\s��"/�ްٞ��(�l4DbSy�e7�R>�+�=��><���x����A�]�vq��
z���Y;��� ʵ��5��7�g~��6�9->��DS�����)�?�����hN��FCY6�[��^�����uZWƕ�2��ZZZ�D�%sO�	 L}����鏰��A\GK<�4��G��thS�٦\!�M�	D~>!�z$��/�{���qæ�x��9<���xׯ�:�~lU`A$����dKK���K=\Y]α�JB�$����-�������ҧh	��'�]����"�K��t�%['T����ţ�h�{��JT!� DH\�3�\)r��Y8������N��n@���8*�Z��c�&��ݰ�#��R^��V٢�Ҽ��l}dwH�>&���n�3jaC��t��Y�p���~��Op�-�1�`(�h[���"�A��kt����l�s�#���qC�����a�^��
Bf]�ɵ�<r6ݺ��f��	b�ױ�F_d&���08��a�=;��VÖV�z߇��ڄ�2	��B��l���t������ױkc�eJ�Vb�VҒ�t�vԸ�}i�c�_ĳ���#/br����&��:L��:,�%ć�s,@�Pދ
k�h�!�=J�z��$��+������O��sϊZ��r�8���*���H����	|mW)[[�-~H�]^Fzf�?��+)fh]�\��X_ltf<��
�¸��~���@�Ղ3������_W�$0���Ŗ1њ��[\� ��04\�/Γ8�=VqI�g�e	]��@-��Z2� H��������r�F,k�a�Ӕ�9�l�������b��4�9w�z�w�ʛ���C��O~���{1�aZL��0�f��g5B�F*�FBx�D��~<V��X�m�md� D�R����׉܆���r�b�%]ۄ�X�b�T�_�c
���#�򤋧N�6=��Dn�'&px0������m;��[�2� ������M">r���Ԟ�v�K�s�-�lMr�[� �Y�fK���;�}?���aH��R�1G�1I$>A�jsĸu%w���۹f�s��g�;J�:�����ӹ��V����O;w������S_GV�õ�� ���H/Yx�G���Ha�z����?�{��p�@����X�&�N�ʸC��>�u;ܪ��>>/�l�ow�g��lU�E���*�Q�*�~��䮐�"E6��kj!ow-��g.��K#D�yO�w�n׍��3+E]&''�g����㢥MOM`����Ծ'�/��;�Jqi�%c�?v��zm}JW:�����E�K0�t��Ǳ�8�<u�($X��@`�P����k�������Q'�Ԭ�sl ܠ%�s�V0<y
��6G1fw���}O�+��{�џ�+tff�92'p�s��#_��]���!�IK]�x����~��?��>�_0�n�	m%����̍�G'i������`4Of��.��T�gH�s�I�V�m?#<��9�ͻw��ݾa#�{�Q|�s�ǽ��[ظ�:����@"X���
�a]|p��AGЌ��-,���~��}K��i� ��J���LV+������ێ]�E
�����r�����\q �\�Y��%�4SFW\2���p\ �0\i�}�m�[닌B�IS%t��$ג��]ɂiݕ�������$X8m]���:سg:DLϟ>��H;�ݼUJ����W�Hd�������h��[�P�Bz��أ�%����d�" Μ�pv��Ç��c�����	^
�G!�p�j]eBN�k\2g�D�ߜy]��Z�?6�rZ[��=�x�F�� ����ۊ��Clٲ���a$�o(��bF6NX�M���9\ޭ%�?=�4�-���'ǧ���q򱃸���]O��Xm�>�"�?�&5n�R �Q�qeQ#���Q�~U¤��&!�?H��+H��B���$�c����կ`jvoϻ13�A��$���Ʊ{.V�:��<#Nxr��E�m��6��'�O�N:��$�mm511������Ǿ�kM�է�T:/�����y/��E����L�K��G��U`��*�_�nk�4of�n
�%B	]A;kJ�a� e6�s
T��(�j�-|��8�w�W�,KB_���_S��̜[$�~N���u�6lڰGϜE�����w������b�����q�N��$�K�� ��8���D��+���IѲ����p��I|���}��
s����Tv�����	�K�}��_���_h�*y�$$ő�Ɲ�tdJBɀ5�Q��G��[И�Ñ�����زg7&f6�����H����I�H#�8�����Τ���p�����?x���.:�"�M������]� ��&���Jx�k�pf����P���'��N15Q���
� ��Ͽ��7ޅ���?�1n��6Lu&\���S
�/X[M����WƢN�K��0�����/|���cji	�zV9�^]���K?���H��un�-�[/�G��g���3~A����8.d|}!��=�_o�?���֥�he�Q
�%B	]�%���1��Z��5��II#��X!W�}�6
��M��~�p�����q\eT�-1�}��8��Ν9��G��O�y�'D�����3x�;�J�z.iil&�G���N�/�kl�&�#�����},9|�ӟ�}�݇��"Α���crQ�2�c㰷�y9_��֓]�m�L5�"�Ikl$+�M��b	������Obn�.��0�|���[��XW A����bWi-&"�%K�|�|铟�W��?bO=��Z��m���%r����6ՠ1�iLΩ0.xb0�j�ʤޝ�{�3G�v�{��@�)iӳ�iG��x衇иq7�=�Ѣ1rPaNBL���cׅN4a�
�o�9뎜s�N�}��>�����Y\OkwCkS�!Z��ہ���pw�Qi����o����κ{?�ŭv�[�� b}��iu����ٲo���R��ЦG,����K��B��ǉ{8(���Qw$)�+mQ�B���2�AK7�clŤ��$�U������y"!r!
"��{gO�������Bq�Yz)�I����Ol����q�m7cǎ�wnR廪���>b��%�����s����}��x�˰��'_�!�H��F*��úL�@vNX)J�E��5x��A��d�'mJy��4C�^{4�f/C�����O���Y� �2���7�	��)�'Y\0[D�	 d��Ź�x���[<��w��>�5��^g��:	E����3�g�z�Y1�C_fO3?���U;��8]�u&9�܋���� �������X�/cff
������@ϩv��X�4���n��њ7����"�<�o~���/|��c��Y�N�l�inh����H8�~B�8㟻����P
6h��s��0�Y��!%-�%fK{�)��Wr�Z�L)����Ѩ�i���2
�k%t�^͠?H\��X"�E�͝���>.#W65k��2	I�ecM�:��ĸ���sX|�i����7�YN{�$��ę%|��_�Ï�o�[q�����wݎm[���j�ˀ	�_��.F+=̟=��~�S|�H�����yF��'>�E�m!7���h-1���%a�6X$
1��&�q�{m\}w�F�汫3����iZ�cGN���k|�[��o������'�u�vԛm�R\u.Il=I���|��Ƀ��W���|�����n�h�d�i1g2
$��`F��Y)�j��+�lX�d&Vomṧ��P��,��^��y�	"Y6�o��洆�?_���ġ��{?�O���wnG�h��j���\��ɝց�������<�����SO�@rg���IS����d+K��9`L�6�B�h�4�P ��DT����5�h�k��0fORx�<6�ϫ�,?ϡ����A��x�$@��)4��Q�9��:����%t0L��JWT!u��
W�J��^/�^��VGE{!���C:�-�	�5j���v��1x���WP�#GC	������ҕ�={�;����f6�`��-ذq[6m�ƹYɀZYZ$|E���}V�v�]�Ȥ�����$�1V���}�v�H�x�5�.�b.����	��&�M��倰
^��xm�}����Q��z[�����q������x���{n���c�����4���
�<^ؿ'<�����p�d�i�:�!Z�)@$�$Y�uf0���#�w�9@l\�5��܎�w| �`���E&�:�6A��L��4#^����<�o�3�ؼ�۶b��]t�6H���(��/9���H�q#��::ז��E�����D2�������$~��W�sO��~��_T�=�Of�|�����<����Pm�/VHŌ*Aw.ޤ�8�,%BOs��:Z��`bjRM�K���C�M:��H���w��ft��1RSČ��E��G~c�+��:�^�[��c���>H�����&}�����p�iH��zS�s���4-ds/�����ɳX�3n��Ӥy0	��#�pDZ]&D�$�K��������?Xnr�W�%K͘��*h�i܁��s!*5s�q6I7�C[��T�����#ҦI��	^Oǜ[X����>�'�i����x��z"ΰ�M�ۈ�gDxt�ɔ�G7��ĒJ�,�nT���Q��gm=����^3c�;��},ح�F������ɽ��v:��$h��IX�:�ƨ�©�N��Q<O�d�J�$0q��A�ՠ�H���&=�[kllNbk��v:B���8o��-
�-aV�Wzx�}�|�[�]2!ZΘ�����9��W�wT��2a��V��u���7r�	�g9��(kIS�X�%C	]!�si
�>�(Sk��V�q�4��;�NWg�!e����[��7Zn�BG���1Y��rh�B?l�dr�q�.k�U��E���.Bc�(���e����Y��ȉbt=3K��AW|n�f�BI�Z*�s��n�����N3f�<��a��nW�t�M���5�X����u�Y-��pH�ݣ���|˲I&%uj�"�k�#҂�yD��A�M��}S�5�<D8ӯufvI��ll�GO�R�"�*>t㄂.W<�c��H4�	�s|�6=[�#��� c0��0 �r�?�W�+C�n���ɤ�=�-����g84|U<nȓ f�?W�q=���ڑ�s��qEI��RTy�C�w��[������x����ĻYlI��w�~}����.Z魴��CW\2���{EI�+&S�	�93_��!u+�TѪ����vT*ڸ#�_䢧�5�t��<"g��Z1�u�bqg���U���YÎl�53�:�i�J͚�i�Q�y�Ќ�N�8+Z����i�\?�E�9A�M�y�T��[� �-&
���GR�5�:��[���Ÿ,)4#[��e>w���BA���.gJZxRCA�0j�0 ��&�~��T�Í�I0
� ����	w�s&_F�5[a-����k��w`K�8 7�:㱡j������6���1����*t�ȉ����gےb��Z��ǄO�uGn<���}�Q6r��<�B��ei�7w1�+7�a�n\�m,\KQQ��цV�e�ښ(O��^��U)m���~?�"��|��û_��o�>�L�����=sV���%ta$,
]p>6���!~y��7����v�`���LZ��*� V�Mx�peB��w�[}��Τ�S���DH�Y����L��qښ�s'61+G��+Osi�)s4�
�#]z��#G��ŋ��mѹ���`2�/)�¹��#�2�@����jf�Zn�0{30�h���oE�s�:ǌ�EH�P4`&vQH��&k��b��@|�܎U
�aLLB����(�U�\�~�o�L�>�½Jq���䇏�V��O��G��+[x�;^���h�9��C��KK�<i�EĹ䉌��(j��<��YH��:n��J�_Cz�GR���'ޖr�J+��h7�ˍ+��K��$\F�W�?�~Ǐ�ج>N�[]d�V�`�?��ܽ4瑧�t�WTCW\:��\̓�k�~I�9� �C�WZ;b�|(6�`Bw��6����d�@��#���%�ϵ�G9&k	z�=W:�6���'����W"��1�6�L3����.�:!�>i�p>zُI��Iٴ�mK-��&gH_xY�\��l�:;�cR��Ȇ9�s&�q�sͅa�w��>V���G<��J��f�t*��� �mC6 ��
n3K��cNŋ��{�qt���P�Sd] ������<̋�͖�~T�"�N��\3�B!E{����_�H��ȵ�\�'c�h�I�(�s:�A�>b�Ѻ���q�"��g�I7Ԏ��;yWM�eTT8����®�s��rU�SY�ݯ՘�ٻ�`�(�����Q^J�Uw�;�-ppI����S��e�K�����j�͞C҂�f\\�wAW�R��p�^e=lS�y�ϧ!*󳋊fΐ�׮n���r��>ܳ��b��2������K�e����$/0�jw(����#���[���Ә���5R�L���Ӻf%A�e�0�9�:��:��)2G�R�,��k��u�m�:�"���2w�,����-J2t����_DAy}���0�����ɑ��5��G"9�~^��y��J�i{l�����`�b�"_Rp
�/�c�1��oږ�A��c�(/\%����G�/��B�������1r��ӈ��n�C_y�\n�{����Π2��AX�@��L�Y{<�'���J��W�����%�f
'�qYe�疅ѢF����D:��P(.J���{/�<��qZ��<���8������c_��3r O�˺6�-��^�bQ�wD"�s�62Y$A���w5�Wg��2��,t#��K���L��;����d��-�Ƌ�k����R��}����焃P=�o�ӷ�,?��vh�|d����4�� V�0
"�����8���F�!����	5����	 ��8΂�����'p�������]!@S	�<�5~!h1X:�q��qH��&_9.�V-˭F��L�{�_#�q�R�:A;��7�T,*�T��nX���4�)�Ū���xsT[�˾V�_5ۃK�Ƶ:�F�~�z��ik�K��:�+&s9��� �����Mڔ�b�L�N�A^(V��뎃�$-xk����<�a=�F�,zR:�M�g��<�P}�J�A�x�Kӧ/�G
��8��\R�a%��,�p>qf��I�8m7h�L2{�R�xm��q5�co�5��
c�{EQ��O����m����� h�� ���HC��w��-�V)�����S���/��_��s���9C���L�K˺�>�2��V��;���
�/�� �*�~�*�o�0��ft�*��tR��[�Y�YZN�+з�r��v�8�@�ϧXb�u%<�!�q���u
-u���1����5�4jFjuW\2���a��vUδ�!�Ϛp���t���r�̑�V�������=DG�pP��ys}��F8�hw���ο돏ÆX�:VW��ر`�os�\ ��T~�
���Gʷ�����q�ǟ������h<).�R���:ӿ_�H���TL����B��Uq���f�L��NE��Q��� ��D��5�Ҙ������m�,l��f;�r�����gռ���)�	���w� 96��W_4'��mT��`|�l̈́�-D�;K�9�ဿ�%*�
�=���X�3n�N�p���:]�9/H�� �,Cn�����7ݒ��?�-�\++kGv IIq)����E3g��3�c�����;�9����hF�%�[RS�H�؁�+��=|������EddV�NTdF�jni�]��e]�i�#I��J�P��������bY�U)s`K��Z���J�ٲ��uu���ɭ3�y��R\�	�����eW��<6T^��8�t��\�[y�௮��~W���uӇu���%:�U��GQHƾ;'$�^	���?]5m�_�X�>l���Ӊ�?ّ�T��������^%�	m��E�ǃ����2		�]�e-_m�p������	�B�R��'ں���W-��{V���e�[��ʧ�o�8��sV��.Q͹�E��u��
�%���<c�O_V�3��g�a�� ��|��gN�D!��I���1�Y#��C@o��B\��1�³tMҗX]����K��ƉMʔ^���5o�v��v�r��ֵ!�=��p�+P:��]H�2#���[Hue�S��D]��\�ե���~P[N���0&�eu�-���ט�,x����)o������Ț;�c�NβЗ}W���RX���݌gú�=0��(���P%�Ƽ@Hp|uA�6H}n��5�5��\Na�ֻ�@�������8�Lho$���妊g��u����r�l(&�^�%�*�.�8�OY��
]'�E,0�h����Zy���w��,R��f-n䉥�D�����G�v��`&�,�b)��
�rf�E	�'� +��=?�+b1$�.�f�--���'1j�-@.����*@g3>���vh����L�:�nk��,�I� �K{}�	��ܳ��mLK��h �'9%����T:׉w#�9��}Y����]�|�\KO<���{Nۤ��+a��e>ؓ�u��˼�J�`�i�㙰�K�s-Ok���]��h��N�;ps`�e6X��1�����]-4���'e2������pJ�6��9)�O 4���V(`�T�{���t�3W��sx|��w��h��'���`/סk���gh��e��	��;N�e�U�F�$)�$$�g�$z��L<���f�:Z��X���EUV�k@�w���s�!6����[��K}��� J;K2�+��>���_g���ZΗ�=���zzo�-q��&3��S�*�ي�����n-�*�M-"�I���?M�8���ey�᫏WV��w��iI��ԡ�E��ʆ+d ��]�R<t���>N���aq����z���i������@O��e�=��l�,l�
����]�utO�V-y̒��ƣv�K�>����'�0�L�l4n�eybi �.�V�Y�2��Y������f5,h:�+�L��V2�Y!\�-8�,���.1��*�Ȁ���w�(�n�9��\<TK������+o�*k���tE����P��Ifra�UΕ[9DP��8��t6C�^�ͪd�����i,c��Ym�f�[�Wgw��;d�~-bdՈ�J���x���j�Uìk�}D��_�<�F-�xb"[�/�2���2�_{P��מI~��-~8B�?�J\�����S˞��e{0s�o�Z��k��M�oG��a�.�n��5�a������)�������r-yQ
��\����q��.n!x�H�I�$�5�����6ɧS~c����b�*κ��@�u1-䙀�$����-�<�:Q"	V��1�2����&��m�\�.��E맺+{���Պ��3u�n{�����h�sƠs	�}\ҙ0�����y���Ғ�s����x��PZ��,��-�G���Ek�Xk{Q���c�� ��{���?Ln���� s�Y_%�j�j`��{��n�}.|��{:e�W@���}`�2����*��RuuC��)��dKe�!Uy�����M�����P���GϦd�l �g�?es��p�xy�"g=;t�V�0����v�����l��5��O�7�W"E+�ˁuY
���:/1W��$�i��n::��\�?K����\����S1�Y`�F���Jz�˞7D!�͛w�w�k�=W��~?i���:@�W�ׅCy�g{0C�b������W�j�U;���L☳�]����r�,���Ƿ�Oes|k�W�0��g�	+�Fu?�9�P�?K�Wֽ���,p`����*OI���)�3�ЧK�1sЧ����p�l!�ynP�R#�1><���(j��g�02U/Y�i.ge��(���)��Œ�����^���;��w�tm���B�5���*�:@o�W qĭ��fZ�)KS6%ۜ�^�ŦM�Eo����>�{�>�ŭ+\s��oV� ��"����:i���F6���w�8N���������-�a\���W�Q7ǚ�����%��������5�j��}fU(e���ҕ]~���%�W�gKL7�AN?�}��c��>�����p
Hu���=s7s���**X���0��]�rQv�#a��Ks�ӽN�s%��ڨ����e$��Y6�,-l6`,�&��Y��M(ׅІ�,˽(=R��U����NLH�^Oz���V��tug?�F9�4���Z�-�H/\��dD�����.saA+��p�)�B`��˒$���)Y0��Z�0.Ik�K�s��� ֫n�F��*�Oz�'� ޻("�.�d)��	�����U[^�wͮ}ފE���Xj��k�~�W�Z�&��l��@e��6l���Q[����F}��O�mi�������Cy߹�?��ځ:�Z��sy���v\*���c������AC_k�s�j�%�q?����-��(����ƃ+:�Í��dh� ���� 7¡����n[w�ܗ?�v�r�8�.G���b�+�7�v;W�j��yb9�7�ϼ�ipP�Z-�.�*kT�(7�h���Y`�H��7/�(2L	�y��%�����OK��2�a��pV6C��I�zr(S�V�%j����N�)��om����+�ű��v�0�ZmC!k�q��DT�p�/���	V!��`R���ĭ{�s'�m�3U�cA�zz/H�\"�����&��j��ޮ�X8%��t�ū���;��Q
�z�L�Ч���l�)�q��=��|�K�_ߑ�s��1�Y�T���Qf?���Æxf?H�I!O�쾁w.aTu�@<�pǳ�	���h<�ZY)Z���9�oTb�gD���x�%�	�B��ػ��X�0���ܢ�ͱ���Zw����#���&)�l�Y�4�b��UlS)�t�f�+S׽�iZY���c�L[Vg�˒\5{�]��ro�7� �媴IY>���(ZՌc�|F�v��U.��	V|W�ρm��z�������D5g�B+���®��b̢E�]��,|τ��Xq�>�Q͎�6��S/������hfϥ*�5]���A�ዃm��v���
���Z��u7����rh7s`���s�*'��R(�����zwм�1�W�`���ڔ;�O7�ٻ��ŋ�A�1oZ�N-��H��4.�F$X�)i|kI�H���T�(�dN���CZ�F��q����b��T8����@�X���\�w�+�KiKP�<UW�;0Q0G6�l���-�}�,���Ѫ���*�R.�W����/�ߢו��Gwʋ�0]�q��,q�V��d���q&�>��W�á�X�SHB:*�8|ֺe���I��^��j�M�_�18]Gyʃ�6���2�P+�T���ּ�`Dv�H��%��EjӰ��pD)��j����K�L�;���(�4�h��20U����z�T�,^�\��w��5�;7י��P�tqs2��[����]4��J� i�J�<!�A�ʺ0qg%S�
Z�B�Hs6�a͠��--zW���lV�1��%P�V�F��)�޳r��f�ó4����j��Y��9#1Q$��Ҳ�6$4����� K/�7�ر�ۆ��պv��X�e�z�v�4����Nc���ks)6aj��|����w�)���*�M�\3H�m�b��e��p�~�]����rJ�n2��;��H�-^3I���.��$�Ҽĵ#5X�޸�M^���/U��g_�5���SP��i�u�xw_f>�
��T�~�������2����X���=�L�Ֆ���Q8�?�ByaX9��l��&t+�Ç�����+h��'�����f�:/4�>k[cn���f��Ģe�2���7QLk�̥S\�p�aio����
p�
l\�̓��e®��vsV���M;L���+lÐ�Lo{q�g6!����Y�e#GVX��� �۷��kE�P_�a�2�\��s?����sW�ce���c���@Ģ�_YkJp��{�KKk�+&7�����su�uI�!�	�SXv2�|6A�\/s�0�t����2v�
�Q��sF�e��?�%E�jO��K��Ii�2���d�����K�M1
ga5���EΉq�����4�� z#\W�O�Si慈����)3r`�(a]���{�|~����ªP�_�u�m���tr��=|�P�O�s+�25�|��]�wHW���44�6Yj~s��[�����=u�-8ϣ ')ء&���6�T��9?D�^ 0w�f�����<S\����h�KA&���eUۭ+*\�AoAAq1dwޒ˲roݵ*;��%.��*�m����%���U�ﹽg�W�<5ɪ�~2�\��{.jN�p�k�˅V��Sƫ$��zn��s�en6䰕T��&��l��Q�{k��KW���F�P@oy:nOG��8�=�sX~�P����^�[y���Kw�V�����$�{�-��U��\��ϒ�*�ت��,o�j�<y�1
U[���n��5A�K��jWn6_��u͉U�|�&������w�k�2�E��\ټE�ҫ��A�椳��O%������}��Pg�;	�g�������%��.g�4�-44?�k��A���c5����*�!���V2�''�qp��Ͱ��W�x�B5#��b�m'���-�B�u�d�O��^����+��h��'����E��t*F���:QɁ���UM��y����_��Y�Ɲ︵Q�C�ʁ���_&'�B�;9jU�uPѼ��|/���hq�ۙ�\�,���]	��o��(C�˃Ȗn�$��ST>�E~t�<*\L����9�@�ǂG�S�*K�T�C��H�V�N���*w�^�������D��^_Q����5���hs��Eq���&�g��T	���u����"A�s�(�6��t~1)��aB4�z�\-ϝ1��}��Pa���.�(:�Bi�� z#H�yV.˻n��*��5p��;����-{�?W3P� ��� ��=�����|�]4�M�2r�J��P��'�A�Ö!�5���WJ���v�~�����U�zz?,`��m�8Ʒ��9�y��X
��u��zhW���m���c({C��7{lTWf\y��Y���P,J��2��>��)�<���݃͌_.���b��<��*�0��$We�۠�b�_�-�c�sa��/:`:�)3g���a�I�a#��#R�T<���o��F�)��d޵{>�[��Y��;Lq���*
U�8���:�+@�=�`�2���];X+�E�E^߇i�遜%�q������XRl)�J����*Z�#iu=�P�Zicak��e������]��-��d��<�X�=@mx>�ie�\��(Jb���6c?�aUY'p��F pʅIӶ�ٵ��Y⢖XE�e�WϠ���J�����J�*��Q��u.y�k��^>'85#\a����޸�ʲFu>}F\G�r��CW��Ǒ� �ý&krUi���u�660$@��2�G!i�	��Ϙ|�]6�A�g�B���ƈ=��<��Hr�F[��w�yU,w��fIa�A���E]��%z���m��eq�$��߿i2#pfc�N�pn��^a)�e�:���Ե�2�֖����c���(lx�0�p������e���W�^�i���SxJ{���m�*�w����[��(U%xV�1�v�\.A靓kbǥ�����ߋ�;��'�W|n��g������J��KH4��|�Mƺ�c�\�,�kZ�[�J]�����{���(�9r��g�3-��m(�b(�Pf3�(�څؙ�Ya,��j#�<�4�ވ��ʸ�x�+���8�!��im,^�R��r����#��Rw�ʏ��	إ�Z���:�j.I�vZ��U�1�9�~��݂\Ope{�����}D�~�-q�8��n,�B��8w�IF����d9FZ88-uU�����+�$�&��\��
j��`3�8��*H�v݌�;xE(�zk�|�6��,~6����s�0<7��Y�!������0�i�fDK��yF&�Oi�HX����V7)U�<]RQ\��dWb_8%�n�_[fP��K<��n��s0gt�^'W��}���q�+U[�����%"�<�
��^���%d��eU��1¤E ���Ӣ�4rni �^i=*�V���.~�5�9���pg���	?����̌�Y	�I�ε�Њ[��|��]8W���<o�,��Xo�ŧ�[�\STYT�v���^��
�XE]���]oA0Q��	���"��&;Z�N[�R��Ј�h�#���+���y��ᨕ��z�}Kǌ츸�����`!fu��5j�QX���O5Z�ij�]�Ȕ��"�����b����&k�c���[�rU�n-�B���꾫) ����Ugٻ�vc�]�Zp��I�q�}�̓�7[�hq�����F
�f���~#$AҚ�3�!s&g�9�8>���p��� z#����#nibݜ(UY���uV1TE#em֚�2�Qo7_�^K���Vg���ܘ>�;��ߺ(�[`KY͆�}=��Rsq}wL�|K����u����=EZ+ �� ��"7g2�l�|{a����+ n�S��W�.n���m���ҋT��ʗ���%ٯLD��"�t��o�MrY�M�17>US�y�s�պ���$)�C����vi����'�͏����l��Coc��>����L��Χԉ�4��}�O�o��6�<Z��ާ��0��� 3��]:���b*e9oY�u�O�4`��K� +
E�sR�4�큎�:�X�U�Yf]�.'��E��H�K��v�^�^�����&�����j�=��y�\��~/���������\��>9�];�Y�t����{�;�	�<�+'�ck��ä���#zM�]�U�Vb�z��˞��e9ӵ���2�E1(�<�����+�@�ʄ�gڡ}����vI�Y!�v��"��ЄL����:āq��y&�D�o&d��f-2��^�&�P/([�JH^���oS�m�ŃaS2����uQ���f�nu������\{۸k\T�<qU��@Yͮ����IJ�2�*;�����$J�
��P��;�`*wf�#E,Ȧ��]s�F>~i �.�V:��>������p���/��L�VN��-�J��BYLg�����r%��&S>��߼���N����3��+@)m�8�@ P�H0p7w`�-.rN�kE-$�X�W�(8�>7��<���2�F�c2��^Ʌ5t�אr�;I�/6��V�V����3�x65� ���Ɓ�wQ�,7x��d1�W�x�t4F9M��N�C�!  ����y.=��p��G
B���^�g��i�"��2ҡ�It�0q겦�H{�i][��{64�^WA�?7$W#�K%��"�⠪}@	�K��V�|�[����`��^���+�����`��w7{C��+����Kj�(�'�t����s��M�xZ�`2i��F�X�I���0
s����V2�m��I���U�]�Am�֋mז�m�a-u�<���䧹�9x`�o�JG@���WE�s�������j
̕��/�3Uh��L⟅6҃"�4x�|N�q�x��"��k�VuLs��xu�[��v�.ܺ�KO?E?��X~dM��d��gmb�Pe2�JT���(���n:fdmg��-����C���������B�pg��>Vt�U��g� ��;$=$��X7��sQ�lB��w�C�|
U�Y`wO+r�i�����>+�*�Қ˦]��������lއ����̶�(�������ݻ^����"�|�����\9��xF!��n	��xrt:=��4��'M�Z#O,�7��`��2�[���&r��6�w�6�UV�׼+'s�֥�̴��v�>��û���\ly�K�x*{�y1k���҄&0��)3+���W3�MbR&�)` ����q�d��)22�V._��ͫhmn #Ӷ�o=���:�.n������l�+5`e�hŬ�g�+#P�e5��lU��Պ�R%��
}�s�vb]�t�r*/dp�(��诌F('c�	������a��;88 !e "K?�2:�BL7ަ��@��x�.%�=��bf0���&�#��,eAśo�3�[�ʾ��+�+`��#޾W
��d�r/\���H��v|m���測�҆w�����UKUU�%mR��_�˅gD��-{��h��)�J�q~t���F�P@oe��Y�pF7�t%#� �����~�� ����.fY��X�Y-$���М�d���p�����x����Mk�N�/a,|���h�hrʙ�����Τ���B_�b��x��Wq�����6v�2iだ��bg��r2"+2�d1�Cܰ�m+/lN�\�-]7<��`4�7����H\��d�^��(�fte�v+F����b�_~�i\��������Sz$���8xpo��'��� �4%+>@���6�[Bs�;��:7ey�&�9�k��m��]��I��7����@���U<��k3/��e��8n{����޺�K�:��#�1۹
�4��I�Ae�%���3�N5��>�Mw�΢7�Qʘ�'�X��=4��J�@��;�J�T�W��</�sW��,�/���^�bw;�8N�����XRa	/���s����!�(\���j�����]���6�Hd��9r�#��/	h��N���q���0�W���A��e\z�Y\~�Y�/_6VѺ�A�wX]��?+u��܀#��L�p��h,.}��9W~F@�$��k��g���.Q΀�F�6�NB@M?��mG�x�!2��1Z�lhn2K���1�O	��<��陯t{W{�:m�Ą8H�H����/�{p��m<z�-�%K�`� +4�a6C'*Ѧ{h
-�E~��9�������a(fCq�s��\|:Y`,p1ȅ�@���c���/�9�P(�Ws�j�jBc>���j.�C/l�0����HYP}n����Y���Sڎ��ʸ
��2��*'���fә^�&����?&i �2([�(��s�2��E�9�݊T����咍�ߔ���0۳z�B�]�g:��������d��ifv�$	)���&��cd�	��t�Yb�n�^�����_ų��<�4x&����������؜�.j4�k�D(v���������d�1w�%�,���!m&���Æ�>Y�]z��$����2��Mv������q�����ػ���'m�����G���٣�gp�ә$��~Q\���.)0%����/`�z}�5<���8�}��ƃw�����x	R�J@�J��J[�_���@��-a���`�"�3�������ǋE�VmYg`�y�7�qz'眝~M������}���J�t�����EQ6�!��PF�i� 
&h��'#��4��Yk�v^��D�p�Ui�{��#Yq���LG��B|W���9;L��g�v�q��[h�s��p� ���Mڴ��苔@2'@��.d�o�0�wgF�L���S���x��;�t��+��2A	���ٞ�B�""��;Y���D,e�p���yʮ�G��I`���"%��s����<�@��p(��KWN�O��B��ұ�t�Hb�}���� .\@A��`4k��Bw+!�x�������}V�I�`�@�n!eD%�%�Zb5O�^�;�I�b��Hዱ�m�}y��Wq�/�2)_�9���!v�z��sܹ{]�|��e���Ȱ��PL������Y^�s�:�x���|ݜ����lźꊹ6�6&�hA��監N�e�/֟�m�}��~���r�Բ��B3N�v�V��T���F�P@o���N�1 �����Z�mL?�&yV�0���N�+����Y}��n�����XF��L�!WE�)Y�)�T&d����A���\R6�DE�[�~�y���� |��&N`(�p�c2`@@���гL	@���@6�$�|�(��Ӝv!�8N��M2�;����;H��p����{�)�{�X�rt���C�?|��U\�v����x����m���{����b|���]Izc�N�S���V��/��a��]��)�y�y� �F<|���K�H�R@������18,��]YBJ�ZSR~�#�Ȑq�}o��du�g_ƭ�}��`��?�[��op��7��r����֒P�
�L#QZ��نq<�X"!�¦N��{�	�����\��(L�bN��eE�`|ϑ���917u��m!�KR���aK�#�2�D|�Y��͐�IZ��Ր���.��Y@�[�n�϶����E�_��R��lܽ�)��qۜ��c�\���ӎ���0	p����3�q��3X�v��WѢ.\�mh�9��G�T��9�n��J�y�����p��.���O߸.u�}:�*����,���L���6p���;��r��R���;��:'����
\nuq1��,;M��8�hFf���=m�1P)�o�v������W�`g[t����^�£������`B���2d�@V���V�dE�P��굡ڑ���cj(e� �)z�
��ma��/c��;�}�m����Λo�x2�
�jb(g��\�k:��)IP=�W�4�q�x�]����p~�zn,��?��g?���`�H���"��dB"�-i�Lx��WY*(�� sX��ϑ4��tϢ�IA��c%�*e�@vߋM/>��Ou��[�s@��bu�x]�nI7����ڶj�Q�VzAV^@�h�>}}��c��o]!K�5\z�E��g1���I�B���ө��ȒJ�3h�/���I\��#L	􆻻H��%P�Vd}��2N�e�;-��w�./�s�uҶ��� �/����uɪ���_`B�>���do����
��ci���RY���Ȱ{|H�"�k�1�K�I	�������;���L�C��Ə%��~qj��;�}\%�\���C���A{mM��^�J������I�p�]̂��s"��w��Cp�:z׮��կC:�;��������$4N�Ia��4))�L0�<UQ��%�&��'��,�E[֯ �2���@�*�T'?���e����C�ly'������*LT�b�!(�z�7`��G�_)��4�O��y�}AMR'i��u�9��'��8�9v`�m���� c��),qV�^�B`���;�����WzHn\Í׾�+_�2p��P��S�$'t����(s�k�*	0'���y��WNf���hI"X$�OD�{����<�G� r�Ӧ÷�gf�{�p���CD��{�{4�<:Y��و,��p||L�O	�7��O�2�onnʽ�
�v�-c˱����*שּׁb�[A�����G�#L�}F7��������n>�ַ�%{F�ԥy�nw�2OpH�d�)Y�\zr��Ւ�P&%ڛگ��,��d����6����{�t/����η��_��3��XK�Ҙ�X�Ҧ	���T��
��v��{§L��R_jm��_��,S���?����QZ�Q�t��9#J��JS�gM�F9��J�S�mO&����?��������߿�'�IRg�L`�stןy֐��QǺ�x��y�>i5���f�[����1�-��&�@�k�/o�o�6�}뷁gn���8&ˑ�8k��#'˛���T��f�r@֩"Pd��Y���-�;wn������ʥƕg��*�lo�'cܼr+����E��@��{I�ﾅ}�B%1�	����=�sv�w]9�ò��>�W��BF�X8����G@;d�]�����2�Y�	�k@�`�K'��q��Y��>]wJ׸}�:.0�g�3���:.��f�1)49Y�LX�BN��:^���S�3�[Pt��ư���ԉ���lm`���W��E����O�������a����K۲b�n�6+x�Q�uV�����~by�����B��=���?}O��M·�$���v�Z띯'�網����UL�S �I�Fybi\�sY}�"�,��]Q�j�`l���jw���<�/+!Z&�F�Cy�Q��l���/�
O��g@	k[�3��۴=Y��^~	O�uD/���H-w��Pү�d!G�a��Y�`̆�`��wȲ^��\�r��������+g� ����/��{�4c�����}���{���(��|v%R"�ک��@Y����=����t6�V�������0�I΁i���rT?��:C��Ʒ�`x�2B��8���˸��<�<&eᐔ��O���}4��(����h�x�h�8髻�!�)���A?-1�st��� l}����/��/�����0z�q�B�p�'f��\�-yf| b�0�$��fT:��g���ϧ�Vym���[�A0���(�;���s(��
����p��BJ���,��]p#��!���k���g;����F1A�	��%Ԛ'-ǳ�q�j��<���oB�YVv&(�ie�0+G����,�>']��/=����*Z�?\�D���ƴ=�^��l*�gC�z3�Yޣ�=t��HQX_�F�{E�Y�%Y��,lj��5�J�O���,��ޞ�'e��5� $B�R�K�s,
[��-p�\�`�k�1M[{O>*�r��Y�i�e��:���i�5�e`@,J0c+|2��;�R!"���G{�q�?)G�/���&T�ǘF�O�������. ���>X1\�rY��sN$�sB?��3��m���,n<�4i	{����я���~��p��~[g7�
�?S�d�����\��!R���Ԥ�!�>��ɖ����͆�8��b!�}�6@
ɔ��p8�ĵ��ru{�@#�<���:�����W|�<�J��R��T8���1K������:�r�D�ǘ��6V��HaH֧n���%\���~�{��;�5���%iÜ�2���x���W9������x���v����=�Tk3Z���χ�1><@A�ا�H�d���.piZ��%q��Pz�8S��Z&1��q�ڱ��G=.{���b��H�6!���(��v�bn�%����N2��Dr�Lv��P�Cd�#�qD�OW�n�`c;�.��Sװ~�nuV�{4$e'�Fg��64Y�ň"e�\�s�8u-u��߱������_�k/�����&~����o���.��cڶD��$JES�9�#Ρ��e�{�?��K�o�/�����r/��g'b��x�L� ��I���}�a�Nz�7�������e6���0+;�8Z��9�V)_�_���,�9K�?b�O��t��d����_|H�_m��k���7��� ���;}�����2�c�EJ�>�`w�� -:�:愛�����%��`gWz�oxa�Λ�⽟�#ے����JC���v۝L��B���U�������biY��+�q�Z��������wT��0deFi0=��y�w�.Ц�N�	qh���$���e
����P��dGC<�sｍ�BosIgM�c��=�4~[�.F��w�H�w}U��Y�q���̧�����K��.6/l��=��?�{��?ƣ�:)A�BB�l�JL�7.�/���4;�\������y�����m3�?�jL�j�������)�t6-�/�Y�yb���F~�R�F^`�~hqo��,J�e���^K�)�F�f|s��s�K�mI�m2�QDܖ4DN�#�	�ݼ�_�-������v���=�7��@g�!� ����!�x�`�߿�/>�2:���ܹXG}��>������}����[tE��mFC\��$���^�,�'����������n3n,�L�J��@�KWMj���U �8���2�I�l��*+����w]��i�7�}�	Y���[8�o������+hom�u�
֯?�.Ǌi�����h�%C9�ot����n��{��������-��X�Ƌ/����{����Ɛ�+K[m�㑀d;����Ώ�p.K�;�t���n8ϨE_f�s,}�
d�F7�U�s��F�P@o�k�[d=(n�I����K�4YLr]�����8IK:���1��{�6���e|��B��KR&5H�8NK�LgK�{��P�1�]����1����.�^�4��5:Vge��>�wq�������Q��]b=��e����:�Ɯ����h��00�6en �,+��5	~֞�t��
h���Ԣ��*c������XZ~iC�|.;�vгt�*����v`��0g;�٤t���#�9|1چ��!^�K���ǣ	�'(��C�B�/�����4�0��?��F��������W���г����9��XM�\k499߁)v�ט���u�>.ľ�@�������7J�)��H��yϊ����o��9ZDs&��y���'��A���B&1aq����>c1�0��Y�0iY1��dr�"-��<�i��[���~�_�2���r�=�gRr&�X����$%KT�h�sć3wq��0�t���{RV��@M'h ]K��f���M�ƭ�M]�i&��m�i�AZ�����M���߈�V#�3��[�Nd�$>�j/@՜F�1�!w�-��n�Yʸ:�����$%_!�af��g��	їRV�r�!�������1Y����� f��t	����p}]�������YAv���)9z��dLG9�e�n+��͛x�_�Cw�8z�mvp�����\�1��k7�s�Ϋǔ��!%3~�ލ�b���j��sJZ������@G�P�Z�x64��ybi ��L��6��Ѹ�%:0nbٲ�,���/��\�:E)�f��)\�U���6.�����d��f)��7_y�|�k���l��N0b�Z #���-��F�}��o�M�f������Z�5���_`�t%{����ѿ�LyJ���D,%:�,�M�T�[��\����?�9�K�ɥg�OGկ��q/���M721�%�`�=VlD�0lyUF�|ރ{7�������]�/Y>gb�],%i}0�t���@�yv9�1Up�3M�?.W���`6B���dsY�	���o�_���i�h��?�ڗ/`�Җ0�)��М2.G�!lEx��5��ﾏ��?�/���]�)
-�ا�&�|}M|O��!�y�9w����Rp�/&�tB�<	i�-��q�̶#!��;�M�4J�ӏ%����[@��W����C�I"�l������e��`�&�`����( j!���ws���(�@}9���i�Q�lak��C�6��+R��o�q�k_Í�>���	�ǘdm��% �mxO�r�G��=$�/�Kׯ�`���h�g� c��wv���;�<%��6x��^�L���W�p��-c�s1cqɂRo��0����:庝�����2���6�D;0����*T��������ק��K�Z�U�T`;����������]�zJs�|�k�ز���P�|.�v�����!��'+����=��>n|�%l�3T�1v���lw���Z_Axaӌ���Ì{�3�]���Mi��
���_}?��?ã7��3��H9�]?���'"v1(f�+E��ƨ쌫�W�V��j��),�����U��� ���B��]�&=��3�g�$������՛S|jdy��O^@�����*bs/^�5���+f���v�n�w�3��?I� �����R̋��|2������'��}0#+��W���_{�^V6���iQ��L"�L�������q����|��bw�����Y����� �d�s�3���bm�K<����e���ٟ��N��������8҆�xU���� �#����xYeY�q�k���ث�s>}ދ��?D��D�	.ߺE ��+4�G�8~K!"о�Y��*�PGm.��矦���[7�y�"�D��֏���P�M��{ �� ���$��R��k9؆�5����#B��5;:�[R�����IE��ni��������J�O�4`~�|��N�wy����&Y���(U[k��m}仅]�F��p�͊#A�o�����
mޒߴ4Q���Z�'�=$��_�s��m�|�K� �N5��2�����cq�N	Ĺ�Y4I�O��Ŵ���5<�����>��"�c����n�?�eсMBXQ���Z���y�3O��~��lЋ�z�?���9)O�����e���[���� p�uE��Mc��q7��w?�ѽ�|�il=u9)pGw@3e�������At�u+zZբ�C:6W���m$�+�ǰ�{?�R.��3~�)i�\�`6�N�9���a��>o��y8l긼�v��nCH�;�K�-a�ܸ0ٺ�ٴP���'��4��3Y�.�b�)�[��y���VT�������b���u�]�ԭd%O����oG�u�Ϧ��Vq�^í�~��_�:��3����uM�=N1�;&�{���!��#�t��6Y?��u��p ��%Y�\��Y�=+���e�.�X�ҟ��⺨r
������<��y|���p���å��e_���9�فz�Wa��Pי�\7�R R�:I#R��G#���p��.N�c��dw#��;# '�s��9�2}?�9��S��zX}���JKn�o`t4Ƴ�u����F�ʶ�ja�	������WDs����+	j��Ri+��y�&˝��� ��T��?Y�U�2o���H#O*�����������CZB�n׆���↉U�qJ�_�I	�� /�dc��od�]��/���.p����Q:FV���bWjJ�9�f�)BZ���Y����x���ٛob��'IYm�Y�aqi3ѵ�B��$2�����e��2�T�w�}~�"���ܓ`�N�[��N=�u��Wy�γ�1��}5�����K?�ס��d2��=��ݹ���콎t�3K!�:�v[�Q���5��^F
G�Szp+I�W^����_�����?�;�y��Ͱ��֊��17�F>�\s�rL��yj�����q�iЕ%��*��x0�>I��Gu�vv�H#O*�7n~څ���*k����2+���F��HUI��^�"e�?'�el��l�s���+/��CĿEV��M�B�Q6Ä��L^�#��3t�%f�!����/"L:8|�]�i������� RS�1J��6���R#aw7X��%�nf�pMD|9�h����� cٹ��a쌻:�{�������̒Դ�aś�P�2�}�c0�h���!Y�3k�/na���4'�=�A:���riQ�-m^�S���ʋ����5\�ro�ُp���H�α���K�K��f�O�]��|L�+K���m�\��n��3��o��o9v:�w�t�{�)[k䉥�Ϡ|������@���&m��\�zy����m�p���v�B��B)��H�}FX8�=�ؠ���s��������`cCZ���10�!�̠��Gc�{�h�ڈ����e#/p��7i�!m?�

��9}��o��(f�����I�qcD�+oZ�g����9����`���<�I��p��0gV��{���̮�2�[�?TL~��)lV���W=M�[ij�9��Ǌ+)��b��!_�r���H�y��!�Uz椰]�^�ʭ���5�?�t<B+np��]q[O�sB��Wq��!.ݼ������_�v�����t�GK��iH#w������s�?.��6�b<�ek�>�(��1�q�Ƹ���FyBY ��� �	no������19;��_��(�J�'2�\��B���8�_���`���ǴH�}�����;�_����&�b'0�Ű�lo��Xk���w�����GG�{p��,�lg-�c��@�~�0��;g?k&F��9�Kٗ�)ɦ��,7�_,�w��<��m�����m�|U�q���������\!��)�U.ꋘ�����������9}�0u/7X�R����O�6�ΛXY[�ƅM\�ކ��1,C�'��5G�)�b�N����`$D@W��U�+x�������>�Jz��>���K�9�|��=�%��9Z��T��^�e��/L��	���6��?>&\W�F��Z(�H� ��~E���q��r<�Y��oG8��u:���~��8r$��J
�4����<�$��s�r��1-lǹ�~����U\���_z�(��)�&S������\ױ���?���m�rt���1�d���k��v�0eK�0�zkX�Ze�r<��ު���l�X�j���m���z�n�ڔ�pv�]fQ���Y_�f��[\�Kb�����K���ew<.n.��n5������0?<=�\^�F�yi�p��W"|2��[q������{�q��W��������!O$%{uy eZ��6�d��hoo���}tVz����q��a+�W_2=�fh�3!ⶱ��b��}��~�����ʐ�{.�s�A��~x�����LCnv�<��^-�[���x�@�G�Ϝ˽i��!ewW�W:�0�4[�� ���0�88�QuI���6O�,�*V�
�����YXI�������m\����|�U�n��i9�����*��Qr-2W�97>�A4$ОNq��=�n����8���I[+,�� Ԅ�5zh��N"U��6�d~��9���E_��g�l�-G��ۻ�}�q�Y���}N~���e��Z��"Hb�6��Z=�W�P5�a��m�����,���~������Kx��6NS��#J�N�đ�߶	����>���3���O��/��?%@���S��h�,�8�z���7ߟoY�o�����=�ph��j�w��D�,4��� �9@o��Cʳ������u)|K�KR��K(r�p,�:���f曐]���dnoZ��fc�{�����p�~��O�1����"���uUfc�yv	wK{t�.Fwo���h��-��|řաVs�� G[U����{�-���ՙöô	t��",��'�c���3��u�r��+,����F_�v^�8��rDt���ɢJ�N������ifL"�y��P8Zd�s����o��?��}���p�����]���}\}�y�lII$��6V0#q�O�o\��[��6��w��o�>�ŭ��t*�5�h�Րu�<L�'^�����_�
��w��@Ξ	n�*�|`}}]@]�C�f�j��3�|H��	&���l:�68�6.�k�a�Y9<�4;B��3,Y���ŋ};䖬��`ʸ��4è����|���� _xF�m��#�W�����;{H�*��t5�Ť�Ⰿ��>� �������3f�mi����Z����'P>&8� ��?S��9��������&�s�oOV��,9y�H�z���Z��y��-��%8������0��.s�6!�(�$��N��3����C�����[�}O]�(ԩ���Ш&K-JC'��������xau��w~�cܣ}��@z��g�����a1��l�̯;�L%�H��\O��읲
�����ZyV��F�� �o�|BY C��0�/6bJh�&;+�Y�KD���ZZ����]��X�L�Vӄ��<\�b�����������Y8�$��h��;F6I�h�� �`:CF������x�K��p��1#��u��L��f�%e�<�}������Ŕ(�����\(c�^s`�,�%��y�ܗ51���7�T%w-~�2��	�{hrT����Y֦9'0�H!l�1���x�;���.nHk��Go��37щb��q/�I�������/��?@Ҏ���1��.1Q�sh�������)1��{�?R�eۨ��ι��*����^�eг|�FyRi �7F>9%}um�����q� 4�3�)3E�g[��l�]�\�PU��9I�eJIB�lN`��3��.�}��70f9���Grd��?<D;�؈��CDd����~ӻw���!�t}\�W.���qCX�`�Î,��Q�������Gw?�n��̗a�Y5��mO���Zտ���6��\S}��o�$˲z�����R��F++_�$�)�+o�X�.w�$2҈�h����?�ʭ�p���i��68F�w�(�DI��!��w0���������"�D����OhN��Y�ь��s�c|�d!iΫ�;A�~7l�]s8˕t��Ǳ��#��V�I7ԯ�<�4���$�d���S�x����I\�e6�-�n�cG��-Lia�q�N���s��=�/�ɀ�E��p�2%�|0�]SeYPm�H�3�;��;o�,s��/G!6T�~T=�}��ʺ�UlV��]t���͗����V�ˊ=��f2�JL" 2�����w���xz�'ٌZf}�j����_�s,U<J�تʳP5���,��I��r�!�b��OJ�J�B����NF��Y�)"B��"���������3B03|�'� �Z䜷Q�b�`��p��E<�{����{8���`6A�0�}�j��\<ݟ�'A]͕9.��|���k^�^B%����v����z��w{�����O�I�qH�m��Ϲ<���(��4�ִf�%&K�%\���q�k�����Z��j� �t�)sxwB\~�Kx��W��0�Fqf�h&�1gJ��d�+����i��vp���޿�^�a��|��b2cY)ܦ͂�2��ʰsձ�z������Q�<��v/N}�ȧ��xv���pvܝ�/��~c�?	�΂?��������d.��M���S��`6�!�D��d�)I6�%�Ԟ'a�-��#���93,$~<��|�,�1��fXYYA�9�'3�@Nf���;����������
��˟"��:�s�뷹 ����"��Pf5_Z17[��A?���#+p\��gn��ԡ�;�Z��� ��O1~����(+��%�L�B�Q��UeA (�e��+�:KV����X3v��b%�_���f� �bg/i�Ԃ��S/]�s�!���g�&��1m��:'��A�,�����>��x�r�ѣ�8|�]�}�f3�r.�(�qGNڋd쪇�䥫�Y	] Ƶ��(@��2_wl��~΅�,���=���z�6Z����'%t'�u\]�S�
�*+�^��:k���nh�w����v�e���sq�c�Ր��0��dR'Vr�B�
y0m�KO�V`�9��z��> K|��M\����w]�����t�Q�#m�K�}�x��-~>�����H�ؠIۡc�tL&���V$\�D4o�M�ܛ���m�+�P��;���t���<`�Wid����.6���=���a�7�T>���L�Ϲ�Nي�Tr���<W�f)�,�/�=�d9�En���+�� G�`��[���ob�W1�Si�n����� #k|B�w�:y�������d�����b:N��D&��UAY -R� ���K�:]��K�;�n�(dK�l��R"N)[;�;~�ջ�%~V,{�k}Y{U5�χ��e߹�;��_�9Xrݾ�V�&?C��*.���٬�R��P�7�=�)4���:��)4w�1tD�=����ʋx����G�����B�#`�we��
�X��4�9k�P��8?��9����f�|�j�X�t1>�G>88O��F9S@���խ��C��)ui��,g��c~1VzJ`.�jdj�9�T-�%�;���o����	\�@�V���>�i�|8D��~:�F-�h������ǌ����d��bA��Yڷ�(OEΏ���q��)�ꉺs��c����+������1N?~�Su㫺��h|(Y֝�q���Z>~'JOh��1ͱ�
%��{����O����f�Cdy�Υ�Bc�rrd+� ���_�
^&��ۣ=����q�� �T�U����T�Q�d�2�I��I�))��oZ�����}�љ�Ƿ���G�fr}vd�MO�Ӏ��.:Jj����Sv�H�X16��A��E�O+�qa���p凿<}�������hg��:��ݢ��#dG��~=�Kg�>���((L��P�~ؔ��GN��-���~'�j��]��������{,,��k0��C>Of�����{���˲m�o���-����x���7�6M[^�C�6_	�BE+HC%��Hid�~��/ㅝ����q��v	`�2ς�Ļ���{�x�g� �U=���>%|!��EQe�sH+�$9�.����\�<|�/���ެ��89?�7��3%i^��"�^�ȵ��r��"x��?s�����a���.���v���O��{��K@;��Z�`$���E:�O zuh1V�F;�ݻ�b�-Ĥ�Kf�������o���$�hgI�B�����gk�<>���2�q
?n>./Ƣ��ϳ��:y��TAd�.���0�����n��.\�ƣ;�%�ގ������i�vg)6��~�wH-�O�����!ZQ[��n��=������9a@ʲzP|/���r����'��h8:�d4�F>}rƟV�r��KkW�t�,�����]��M��|���7i�B%��eN��"C��-<�{�C��/
%�p:��j3�q�����T���vw0|����{P�>V�mR*8۽%�R�o��@��W��'�\����<R������������.���s�g����_<�ies�'��:U+p�M��͋���d�����V���v�G�$���mR@{��.��CN�[��<�����_�%�ƅXМsލC����oA#�d��.OމN�6$%t�t}����Й�A���m}�ν�|,1��|��-��C>���z�Y�e�+Y$�����e.�J�� �!jn,8I�ۗ���:�!��׮�·���w���ŀ ~�eDc~M1�����#tU����������#�����g�R�s�)�r"�c�ٽL�ޯָ1��^��G=��{��X�>���ϒ�y#��,�|X��lz��|L�Z�֋̘|���Z#����{Q+���/c%	19�GJ ���)����x���kx���'�,���[��ئ�����bds�xU�y�z�]�u�+A\7� �kי1���!�����Q�GYu0��˓(e�B@����g�.N��4(�<.�22��ea��~w��{�Z4�NxB��}6������~����-�O�"�K�֣)��c��)b�i��G��<:�-v\�&�98�,�n�,ˈ,�l�J����e$*ENK�s�q��u�P������Q����?�K۲m�c��m�%�U��p����,���Nub��E��f8|�]�׾��ta�}��ng�������
�����Kx5�����>�c��f3��c�q�kU�w0w���%���� �IA�I�<g�(�+c:��,���ͫ�Y8��F�gz�i�y��W�̈́�4����Y�a`��!�������$�u&��NU��Z���!���0������pvf����ٙ���q�@.���G�� �Q==3-JW�~�=w���ʬ���̠��TWf��G���{���@�e�t��0��́pqϏ�'��R)n+�����}[�b''o�!{���>��F/<s����ޅ7���fv�(w�TŗM17�S��Jt���,�Wm�2��]�yL7��W_��aV&m�L�m	����r���N������F�ϭ�^9�lO�L��$Ӻs����{R��N_���/���Z�7���o���gJȋ���'@~��w��7��5Q�>F��Z.1x�s�"�	�����������!w�S��ϑ��3�Xz��4�<{LZL)H��Cj���At~��_�4"�I᪋�պ�k-g���~�����R9�]���ukC�-���񫳯�ut+HO,{+�M��[��o]E��Z7@�`>��G�wv�3|��Ͻ��Q��JYOR ����S�2K�S�۰$������٠�yr�x�s��j���sL�I�ɓ�lYd�^����矷̵&�t�w�y,�f�:��d�QH�QZ'.�]���ZK��7�~���}�Wc�޼&�ڸJ쐳'h�]���xuk�����f�8E3��9z�90Ŋ&J�lk���{����c�a�'��S����]��2[�~J�f������r�Ԁ~�e�~�
�/��e��eR	ơ.}ω��?�H����Z�}b��p�������1���7���^�6�1�I���u�?����#��F���UD;�gz�cfӜ'�R���F�g�ʠ�kR��bU�Q-aZۖ�5ǖ��g@>p�Z��gϵ�'�r��)O˚��,�/#R��;�-\4�sf'U����}��ݴ�e壽���������Vq#Ā�2��5	�o}��x����!p})�*��LJ�TS,�=jZ՛M_����&nb�����3�(:���ٖS��Ej@?ﲾ�%*�Yf��2ˀ���dt�޸�^��k_{��:�(�1�����;�|��4����I� �����.։�7�z!���*��'%Kml˔��>��J@ݔ�ԙ�jyV�5<�d�U�{��e����^{��e󺗉/X6�H��z2P�2/�}��2ĺ��=�5?\G�BA�z+��~����� 
֑t�� .4g��A��$�H/�;x��)�{�D��x!�,�AL�ya,8|�\���Qg��n�I/��j�<�'�=!�ш�fԩMYj@�:�[�:�6��W���l��0�w�h����w�C�󕗰��˴��ybM>1�x����?B��c#%fO�����P�!�<M��"'�M��'U�X
�"�6aΓe��Q����L���?x����֟}�\�Y&}Ԓ��L��I�k�o�����捥d�q���/MI�[Hw�sć������`�����zy��h� �=�� �m��7W:x�~)�׏��_!db�i�y<K��3Oi�]���,g�Ⱥ�:�� T�F��Z�,5��w�n���(�j`��tU�~f�6�a�ŴE������o�����g)���s��?�����m\��D6J���_"������Ɛ��J���z�dȱ���[�a�:��e^�E9��kS�|�L���kc�Z���K�eL+��Y�\�䔺et�e�u�M�5�pYv.5�Sc߱���0+A�	��j#������T�CF
�w�GF���XC���Bb��f�X��������i,�8���Z	v$E@��|+e�Kb�4*lW<w�C��9/��E�V˗^j@?�Fn�%M�|���nТ�I����"3ɩ-lG�" ����NID�mv	��n�$�44����E����{��vA��任e���;���my�ް�������,��N�Ek��i3�,@9'@�3GGX� �	��O��ٿOo��9�Y.�E�wg�g�L��q�>�\�.�%��Q�$��\gХ�� �lg����	r?���Csu�j��%�`K?@B����W��w���F�� �s=)o�q�(�Օ
�Vɿ�9�;.폓K�,�����>A��*�KOX�y�b�gy�ɉ���W:�0��t�ⶥ�>�垃, ��7�x��n)�Z�����C���A�Cl��������p���t��J���x<�t �	8�2aW����,y�|��X�[;�X���6-��C�J�S�b��2�q.Z3AgKE}�pJ`��2(p��ǝ���ySX�2�t'4���hD��W���A�-��6w�[���a�{��(@x�&�o�F� ����12���9�����a����F���4P�ps Qhl�(����ud�#�]���� L�!ɑ����������(���:B��j�j{u���)m8�$m6.��'f�x�mRPvhs�4q�{�Õ7�B �ϵ�i�+�)������>��6��zp�!����!G����&AF&<��<m�M.(S��Q۲ڹ�3?N,K�Bn�z�b�Y̢e^�}=�Ma�7m�76$Ўj��SA{Gn�:�S>�Ʋ�L�$mjΩ��y��X%xXϝ~V���v\!�eeʕ�L�Bu|��=�R@�e �Q7�l��Q�و+��Z�a|��v���ߣ���n�@gh������#�����?|���~�y��ІT%�d������ŤG�+n,�a$A�� ���E.���Q�\a���!�%���K���b�Wf�-�3�G{�ǉ�*\�
b/^Ľq��_��o�E��"	��\>�Ig���@�r��Ύ���Ĉ�,���AQH�y@`��<\&pt�L[-PsO�/���Ǫ�͚Q�)��$�$���,�6���k�!R���s�}������څ�h�,��Z��?����׿���-���U�b� �#�Ϗ�;Ѹ}/~����G��bzŅ3IC��f��/��\[�DU�i��tfk@����JU:��>�Z�.5��w	B׉���#�����9xC��+̢=b+E�c�H�]\�\]���w�Pl�L3���{RεMl��A���s���h\ �D�U�ѳ&�Ӕ�'˰�Ӕ6=k	�Es<i.˜?�\�I�}�Q�z�����s���W�l�<�R�us�O��ƌ�uŪ"E���������x���]�'�h��I�Yq�Dϼ�
�^�%���3��s0��(���)�t;i��h��)�+sp}��yZ 
�PI�C���R�9��;�祡�+�l�����r�ͦ��ɐF� ���^D��mڱ2��N�`��Cb�Do�����!�^A�H�9wsdsם�x��}x�owY9�s�2�� )l��v89wq@�l��"p��
��2�\gǙ=oYY�O�t�����UM�e�l�"&�RX\En��)W���+GF� �&���6.��&�>��捫�È�t��k-X_]�+����ާ���c\C�le2u�]3�I�EQs��G���'��He�<w\�j@?FT�En)��s�/�b��4�0�{*"Lǌ�Q<��v��/�����]��U����6F����{ȶ�p��v���t�Ѥͭ�jS�2��Ր�+�=%��N_��B�y��s:U�ZlIX�aW�4~�9��O��Hy��u�Rn潇I���ٿ�[�̌Š�F�4�������ll��A�(B���fsSZ��(@�{h?�,6_y������{�k�W�˩\Wb"P��w��]l���tA�4�b�{a|�ǉS��RR�� _���ıy����7���c�ml"��uxx��߁�����KO��aj0�'�mo�h�`���V<��+���f+�2*�7�|��.*]��̚��Na��ޫ��Ī�l�=���{�t���@u ��y�TN���E����Th<�3��V��1�w�i}��[o��W����8`��Z�I
8��1vrtV�x᷾�w��'��>�U?�({�ƐҰv�7����[�Y����v����T8�e�����,��]��Z��C�F������<���j1��q�ڕ��ܦU�c\dp���>���q�����~�	F[;�ct�5�6/tz�5�r.�t�P�r��p��m�"�I׷
�< >n����L�9�޼k.��D����20n١�V�I�ƢRf-�g8�(a��8�������>��yWZ�7N����fD�C�s@L���]�����;���Vxh���XhW���Gr�ͧ*��MG6��%���s�������sR��<R����Z9���I	й=$G�J=ufi�܉�O ~���6�(t-봐`��?�����qcu��ml��>�J|��ֹ����9o������}���Sց�4��;d�/z�>�q����ܾ�6�VA�8����>kYt���O)��X,e��(K��PR���|�"�l���H��{�����
�FE��na�&/��x��}�-/DDX,�n�a��N񴶔[����	[ T��^�	�5ij�剤�s.M�s��$z����������\�}����x��߂���.3��6��>�5�q��D���ఇ`8F	��k�<q*�|g�[Z�3u~�э{K�NӯM�YϰT.*2�ܪL�QSy��"�G�O�҇LX�m�:۳�:^a��k:����Jv�:p�_d�(��|?�觟����=C;���?{n��E���m�P�[�A���*1���BI��٢��;��%Ԡ�uRN�NG�Ԋ����:+Z�.�~���������6�B�R��Q��g�5��
{w�D)�Ƈ!�ݾw�ӏ����3J��\����;ܽ8�c/"��>?����9b�}b��j/��Mw�A�j &�V�.r���<�ݦ�*���ɧ�=|��Ɩv�� �7&��¼~��'a��L���/?9�iD�WYcu�?2?,'O:�y��L,�|��b�l���&�V������'}ʢ�w�Yͱ��.nlz��OD@�f3x���w?@����7�Ak�@7��:��8����*�>��~W�ћ����Oi���:�U^��\�ZW�XN�I|�I�6o��+���3J� VyK�����Hy>�}d91bH��:���:���8/���H�#��ȳ��z<�1:��FU�r�>PG3t�V�< �O�f��L� wN�ҏ?c�/��F���e� �����*8��锛��O��Kv�D�Ӭ��-�2��c��c(d�ʵc	���?���s7�lS|�J��d���~���\��k��HCuI��� �^y�����.F�=�³%$F_�	x.��r�Tj&�ȵ�;��8P��Q�~�b�Zj9����0ą�ey4�N�hwڻ~(6�J�v��(��G��u`s��G����ܦ[���8>t�}�n��m�m����
+����Ê�ƱMa݂>ϗ~���Q�z��Y�5�$�D�/RJ��8>���Uz�..�39w��}�sΟsܼ9��9;f�S�Ǚ� �E.q#�z�H����6Z��0\_�q��9�0��'��tp�՗���{���"�[{2�v�d�z�U\��;�.A�w't�苗(���Z�(g�%��lO[�4��&N��*
ɨ�	�s��b=�@�����-$��C����&8�#9<D���
ۤM��w�(�����̔��YJ<Ě�IA�d����~�	�;[���ۂ#��^-�:��?���+�E��e��~�4�Կ�H�Q��Aڙ�Wϳ�/�S��c��Le��r�I������o!Q꒑�I���A�x��;{�Z�4(��g������:�Z����D��,�`O.i,,�ظo
)�X<��p��1:�kh�����5C����ܿ4�vN%)���N���W'�͈�İ	�Sb&�/݅�4�ot��h���Ҏs�mZ���8E�6���In.KمM9���ؤ��l�j�{�"V}�X��=N@�z�S�E���e �)�ߖ�4���N`�s� f�	�W�7~�yVg��hN�+�)N+���a��V䜆�HW@n �p=�?���9/���������
���<>��O���c@ǴHAi!T[��G����\=�?ˌ�����:�_~=E-��Qj�y�,w��貗�iA��1�K�Z��o"|�FG�H��a^��7)b+[�>�`g�i����'�x8�(7&H�-+�|Qԫ[�0����G�[�^��.sM�N�3Y�
 �s��Y�4���L�zQV��j������ՉǠd��������$���y�ٻRw�����L|���Tge��� ��%���M��	Ź��0Q�%��g�|�������i���^�(3��5�k>xn �o�$nR�5����R�9���:q<��fSp�s'@�+�l�㹷~�tmvE�!�M-�wb��b���	�t?MЉ�L�i�Kdc].T�������1���-zn�Sg�S�lη�%h�?��s^p�S%�OĬ�c�{R�=��f�	ԜcNo�\���$|�1��g?U�g*C`�yW���t�xA��J4:r�8�a�!��{{x��;(n�@��3	��i7
�lu0���������3$�>���(��ܫ仫J`�y��Zg��77�w�z��o���j9�Ԁ~ޅ(��O���yB?\@�0�p���Ѽr��J����H�}��T#=�����hP�,�C�c�2���D�¦�"Sj҈�D��F\T���t9B�	ӵ����4�ш�3�LC�<�uZ?��Em$*��l�R%h;s��� 4��qVgj��1Ʃ* ��܃�P��{�ŋ{jk�E_� ���A6�o��]����Y`>!�܎e?Z�:^g���n����gN���~R���6@A	��\Lfv���D6B�@�X�4��"�.�C���۸�j�{���A��AL��`4�Ι�^~��?����x��~ �p�d��H-����).�Dף�k5ȳ�f��n����봵Z�,5��w���0��wN� =b'�Ѭ޾%�F\D�A��eK��=N��ߝ=8��η6R�]�)�ٚ]��$e7bAVc]:��5��2Ռ��^�|W�*
]N�3�[���Y��R�'>�9�1l�!�'1h��_���*3�����S�X�{�_'X5N��O:��XV���?i �yX���@Xo�c֭k��\�>��9�m�@��ރ�?D�
�"R�����c,��7�˛���~�-Yl�R�(UN�Y�'���
@��Rh0"�c�W�W^)N���ٗ]j@���q3����4'X\l\��;����I��u��QL�e�í-eG�����!�gT����3��K̩��,��vT��\��n���F�kq9Ov�º0Q�:�g7~5}�,����d_��Ȕ/�P��'��?�7u/o:?z�'��/_��a�'w���e��u��q�i���w�	\ޯ >�Wm>zH����O	��ocr�huz�x�&~��3$��_�>�\F93�U�8�iK��'�_�r���˜yޕ�Uj0��K��\b'u���Yۑv�hDx�o �{K���p���q�����O�u��Iϡ����M���6U�56��2ˬN�TƍcT	���:�te��;pfPg:pj��T]�9V��
��j^���|����:�/ �w��˓���cͿГԩxj�īXF���`�s�.Kk>����s>F���9)^.��s���c��M\�{�_|�a��7J�i�ܴؚ$�U� a�@��J/^^���k9�Ԁ~�%-�7Lӆ2!�)�f~���_{ v>�b.1��.�z���`���y� 4 0�����Om�h�q�0����Vm�t���}��y\:SN.�\&<��R��mN����j�Wb+��C���w�ʓwp[��V�������G�|��Y�}�'^�DL�_�Ǭ�{JY�3\���T��9��^�2�,��˳r��?}�t3�ȫ�����Wζ����«/�I��}��s)WcL�v�*��ƛx�㏅�7+��(�xW��'����>�4������_�q��Z�,5��w�
7��P�Mt%we�p��t�1o|�֓j���1Bb$��a�!��!G3s�=�]����2N��P-0U����jRF֎��n�U	T����S�r4	��4�l�t$�Q&Lz�3u-u����ed�/S��̎��4�<����X�d�S�6s�}VO�殌Quq<=v_���9��N�����'r�@v)����|��+��B�=�	�y��C�z�e��W?���-�ЊdEWj:(�Е4;<������AK3������SJ��\����Vsڀh�Y�z�|t���S!fN\$���{>x���mt��G�4��jޭ'���_eH}$�ַ��n���ݪ����/ۍ&>���-�����x�1���R˱�2gu���q����)K��#k���lpW��� ;��VZ�{.��"j����Ǵ�R�����/�yV��ߧ�60ǅ1�w�b���JWF�������;���k\۽�w�>b�io.�y��+�&��'@�w��6�g��mh��قĮ�F�f}������k��K��\�u܂�}6�3�p}�/]$ .��>��w�>m@	�s7Ip��!��t�|��ʎ��f6ŀ+NJL�����<Sq��V�!�w6o^��7�
\��ş��nチ4�	<SZ��4Hy�p��`��SV�*��5=Y�OE��?��r�WL?��=�������$�|R������6�q��ӥ^q��0�:h8�YU]��%&�p��@ro߃Oh��R{9�"p���y�c.���.n �ؕ�"��)i�J�k�@wU��s|��S�^|��t1��^D�\ھ�D�ɈQpg�Q�p��ƍ�+�c�4�C���s��s�"�����^�t	P�#���޼b&E�+>�Fׁ{�`�����?E����1��1BO��Q�����
P}�|��L��g��l��]�7s�S=^w��uև�	��b�Yv�\k�u����{�f�N��E�Ry�n���`R,e�����}�9U�3��g�5���?;~U,p�)�S�69'w��#�x������IzI5p���Ǹ��m�K-v'�1��F+�W��˗�E�G4J�c>HIN�N��q�'O�� ��{��C�1?%[O-_:yJ`�Rz-�S�ev�KFX�yYL�y��^�ӆF|��298Ĉ+d͐M̀���/�}:��@ok[�{�饡t���#�[<�
7�C� c�][$��m^%�㎛������ i�\�?5߅��qE����UY����2Oq��>oV�\L���^Y��Σ���5��霔Zv;I�����W^�ۊ$B=� 7Z���$�q�ٻ�@ߟ���v��\�R[�A����.KS����m���K����S����K�9N#}E�<pGx镗����)����xqJ��"` M��7C��>3+G�1�C�E��)ƿm��-��&����HG7n���a�t=���4ybj]F��k�Y�?N&�ݴ��^�H_�ר�_4'a��8��@Z����V����5��������s�g皅��=�.kHkw���������N��szg���{�y�n��޽�}Z�+�R�Ѕ������!�\M1]g�������j>_���K^�a#��(D���g�x���qz@�T!��kS���9�='�t�9Rn�jvUkj7C���
F��"K��y�7����@���|N���6��,�S���o���q���t�� �����.���ֵ�Ù�S�������?���S=��u�<�">Sc���b�1��s	��ɻ}ݡ�75"��oJ#"��>H�X_Y��	���1��6�Ħ��@ȱ�b=R�I	�ow�W^)�?_y���}�|>2�#o��[�q�՗���Ux�9p�0�X��{��0�ޅ�&�=��ZF}��8�.�0)����sOr̫2k?b7�]0�r�m�_��_�F2�Im�bL5mQ�] �kV�|'��-p�	V���t��T���s��-[��[UT���s�ӟ��P*;8���~:�]+���sphNH��wD�`k1�)��yP?���gn�s�
?��P*Av��V���F��7�s[Q��"����rvy��^/�/�dy��E䑏�/܁{��<��'�o!0�l�ˀ��O �~��ih>fώc��t�Y ���T}�/�����Ih�R��*y�0����dg��N���Y�B_1�S��N�M���=0y���T�����]
��<�,rW��>���V�W�ŕ��]e���d`:&���8�ݏ?���.:�7q�gpO���q���V�^�'o�C
�']��|>�y^��n��5Tk��Zj9��&�s.�����B�پ~�*S�ҡf�6�ԫ�Pt8�چOL�M�kL��J�k�iq��t�����M�d�f���s������L�*�M��Ѳ�� �ѹN+���\����l[W5��ټ|��������foh6��h*�:�T{�\g�1��-(��{����9,�&g}�G^��^^�^-6HZ���p|�e0��B��U�i���J���r�E�W�.�IM��3AL���k��Z��\d�('�X�ݯ��Z�$5��c��Ѝ���
�$�Z�ꊄP�\���ki3*R�tz}wwq��և1\�� �j�����u+5D~�����N�i���ʗm���oX�(�d3�s\U��MmqL���U�^1��k�׭8�l���l�8�(�����WEr��$�L���� ���3�+��P�4���fi��H���B�k��3w0�]�{�S�]��LN�LԦ�U�Y$�Z���:Ƥ�;lj7V���|�(��@P^O�Bx���&�97Fu��q�(��%��J�P=B<NK�?I���\ǽ��I��I6����k��_j@?��9n����.ljӠ�#K!kD�6�XD�}�Cb�Q��މjH3GI#�Y�$53�Jژ��f)s�- U��J3m���n;o������m+/�����`�Q�)��ʋ��u��9v�׮�I��i��8:��7�@|��d��Z�}��������Y�%��e^�g<��xmoya���W��d�(9�% �}X%@p��Moy�4PQ|R�L-�֊���h=$��U��T,���mT��p���m1��3�Q�Lؓ�׵UÙ9���D�L�ҢPT�q�6��Z���dbX/	��}�#>�'�A�?��/�}eS���Z�g2N�j!W�s��C�I`�X�\��n�g12��=Ā�}�p��/��`��-��s,���/�d�d/$6�^�H��4�IR�ib�l�>�$�����rc�>�RWM�����ɋ�_���jҞ���\5a��q�N�n(��ϲ����9���\�r�c��&��V�M{?r�S�Y�uմ;��8�:�m�p�}���Clq�r����X�z�3�k����n�ֲ�W��mrw�9�d��V!��f�Y��1��j�#��y�f���L��2��*��)Jw�=^�4���s�G�#9��wѺq}:�}�A�'-2��E�jc���;�uNU������F���� 8���ZN+BX&��5���s�i�B����8˜��@��)w�bG�w����:of� $V/ѹ*O5+:f�'o�G��SQ���T-c��@fZlX����]e;������N�)-��W��%$1��*�{1�W|�p&�^GO�s2��=ԕ�J 5�ݢ�|��^��6��v�t�\�K�ʜ�I��;�o�Y��cS��-�����(ݢ�D=�����IqG>͐uƁ�ߧ���o!LY��)�f�m����JV� �mn�<̶����I�x��Q������A���a��66^!�|�ں�x.6�^Fcu��eT��WIC��~�:���v+E-�<�TS��~n�|�w����;����q4[��8�Yw�"@��e�Q���-x����l�vG�Rϛ��u'�ӼR�\3��6�U�f�0��i^er�D9-��|T�������-3`.v㕼S�x�*G�9�8�-�[0Q����vXC������t�l�ݺ�<� �Qרv�J:���߶��'���d�e���q+��B��	8�	�:�y�*\zȍ���ư���"���0*��P}~
����p�y@n��z�*e>S�<>���'I��|)������cc���5C���S��Gؼvw^|���1�Lz�*�`���(Ot�c4��䨥�3ʗН�8�g#�.9���AB;rgc]�h�n���$�R�m�9��ڬ�/U��t�`��t"'d��~ֲ|K� ��A���2��x�-������%t��Xv
XV�K�d�%���)F? ǘ��y�/k�����[';�W�F^�#���,�����M�F��V%�/��aA�k�����M��)�ll�����yQ��6��#MfR>wǴĵL�\��Z���)u�\�蔮��p毯#���,�~��[�@?�����sKsć]�kcp�H!ֱKQ��j��_û?�)��=rz
��%6��r�4M�1RҠ]ύQK-g�/���������A�vi��'���y�ܭ*�1>��Ѥ�,a
���!J7�p���5�&�M�*+�a�8u��
�ٍ�S�h�5@jİ��ܭ��\eM�flG3�	3����QFLe�9+4U�6���X��c"�6k��n�{�@�����Q�)�_�Al+���ͽM�"gj�&`�̙�;.�?��Z�̺,+/�NK��_}b8��g��e�ŵ��~~Ŵ��`2�k�X�Jߔ��
������~D�[�m�T����d.ؘ����?K���nj�{ �O(�&��Ir�G���{��u4/\@o�~✘�
�\ϕPRtVVom)5i����|�k@?��5�����N��Fa�=�iF���H����\ua&�)8��κ�(h�efӭ�[M1?���ِo{���K�;�;G��^Q&<�H0+��}T��NY�T�S::����j��5��ة��V&�l��Ŭ�pL�Z���c�3l�0LZ�3�Axf��*�g%i�J;��ۢLG��J�����%F���[L��e�(��𹞙o�`��e5_�hK�V4����k�ⳉ�e:��0*Jմ^q�O�[�i0U.w�2S�*4�����P5�������s��}��K����o��&@��b	ц�B�:,\���v]m�����Ŭ�п�b)�Y�/.9��w�ն��^���S����`6En��z��r�����:X,Q�d�W�D0�Y�1=+�Q��}�չU��g�,O[1�{s����*�矞%&����ڹ�T�da4�	��g�[�@�9�fB���Ca�늬(�0HV��s-{�t�e:�}v���$0P�K�X%@M w��uW暜
WZ=��fL$n�i+o4�����p����e���2��U��^i�q�z6�R�/�r�#�x���x櫯���(������VZH����)k$���,ϸ���^K-KJ�_FyZƹK�\���a��"�3�/�mJ�~?���mP\L���e�׹�2�9��)+��l��ͯ�v���J�Θ苩k�3��n��<洲�X"7�`{�K43N�2�T�b�s `�I@S:Ne�Ϛs�#�s�A����E2� H������_6u+s�|pf����'�GJ��2��ț͙�r������Y	N3��(U��w�e��%t1�Ba�I.=�U�A�3���B�%�A���:���ؔ�фb�!��t�=W��Mdl��f��pJP���5�� ��\��Y����C�~9s��� (Qlx�N� ���hW��PL���C�J:]5�P��B��&�͜�����]�>��������L�p��^�HY9��⡎y^��y��Bc�i] ��߳�hTD����Z�(5��cy/"8R\�B�m\�˛�#�+G�sެ�$p	���0��ћn�ێ	Z�)�V��T�2�G�a[(-G��_�8��yg����@`��;��fb��Df3��t������̥�+��,.LC� 5E��I�y]Gs\����y
>=sNa
����������d�t��R.r�jF�|d�b��HQ�>C<2G7�a��|��@=���h��Ichx���p���J�.��p[�B����I��uVv8�a��J���g��t�r�!f��!�Ea�
�MW+:<n���q��<��G?���B1�'*)#�����/G����>�JiB�Xr�o���<s�HDላB�q{M��Ǚ \�59�CP-�^?�Ex�+��r�E%�\
�\D.B���h4f�N�u�o-g��Ϲ���d���4lF��"3�5M (@.�n}�j!(��*�VOq�Ӕ�m��������������@4�c4�b��~��ߓ��
b��L+ �4��C'��n�F\��B;4rN��.��1+�p��xLǲ�ðtf��q�&������*��@@4�v���`ł��+L�FR %��G��	�(l��L0|�h��ڷ����X��@�t꙰�E�-�<�9�)	b��}a��i�MH)(�	���i�Ǥ�1C�-'t�&1�眥��t�����͊����~#	���J��$c�<Rz���
�s3& o���k�%P��0��~�_|z���]u���/�Jz�d<[��b�/��ϒ�[ox����4���5�~s
#=KyF\����cPtN;�	)���͍K����3J蟳|�r�=/P�v]�2���p�Z*�r�f�BqC�-�.*@]F���a��;?���5Q��Y�`�����^���%@VQ�����ML�������a�m�VA�E����(fB MЈv��0	���I��&|~>)=ǘ6�.��a w���&S��l¶&sf�1��J4�dsm:�!@U g��d���#4�a7	�����@���e�`	=���KϚ#�tL�$U���
�ݠ9�ҽ��lGt����s�*��2�J7)�Z\��I ���Y�hҳY'���I�!e�Ɉ�s���ul����8�h��c\�k��٥�a��<O�p?���=6�_�ƕK�~�Cl�b��
���$Na�*��</�m���f}�� ��`#D&�Y�Na|���p}a�:W��A!E�I����JmG�kR]���w,&�PWW;���j��R��,_$0>�ս8�M\�'+&�XI~l��˜���O���Jpج<-�>N�,.i[^q��j����@�X=&0ۧv܊�ߺ��M�m��% �M�p��޸q�.]���Gx�go�`<ƕ�W�ܳ�`e�#&v���'�x����"gX)��5��ѳ�%�]��ʛ��o}���~�bKg39��G��h��������^V�F@ ���T?`V���^���O��x�x�u:n��{���]����#R(z5}�26^x�f ��ѻ���O�b�E
H� p�VW�7������}�*֯^�C�L�8-�E����G;��~�_��.�B��j#H�b���`}w���z�e�������C\%@�ح��z�x����O
�n;�������6�k�����'��ȇ	�:)��u\_��Z�G���<�v���m���Ɍ��i��̦[�3a��؏dֱ�d�HUE.��e^�9^�cZ��=Se��������p9.l$^tL;�ZjYRj@��ń��O�cEO�:R��b�,$�Y��;n��"w�x\k���g|3km^/��m �e�\�K�wE��jDL���y�~�; g
h��Mi���ކع�Op�_;n����
��3�H�[7n�G��o�1��Y��ص�xỿ�k��6@�J��wo�-���4;(lHdX����0"E���1����bԔ�CZ��~���G?�5���6�	���?a���D�q�{��w>hVا�{��_��?�y_^�����c����ࣟ���(��b�������?/=lб� ���'I����X����sw��9���~BJQ���Uҳ�r���..�-��5\���x���_���Qw�Me�z'���1)7;t��+/�������rR>��tHyJ��_�%)5�]���q���X�V�x���o��̗�v�����ZŤ�L5�ޮWm��FO�R1g|�sbˊ4��B=�.�K�K���O��R�3�~��t��O߱��L��ZW˙��Y9/`������Iϗ�f��k�X1��&mǆtM*}I��ϫ
��DLUo��O:eټ�s�]bR���wo��[_�x��"��'������[�ѺW�������x(l.D��<�7���/�(���g�~�ظ{�|�wp���\Z�Aw��� �)����BR2�����W�ӿǽ�����5�	3��;�p���<sC����s��m�x��'X-\���	�LEKI�Xa�~�.��־sq���ox���3����D�?���«�O
͋w�/I����m<%���zJ7��iF��o�MR���
>�����z��T���;\��\YG�߇�n~���}� {���J\���^���K��o�|�%�@��wѹu������>�~�.:�|F�[�m_Q�R���=Ipc'�3�%`[{%_��&.�As�e*ިʺ�?�)����5�^vY��
!-suuU���-2C��r��]�B��W���rV��\��U��R���*���(mF,K�
��Tn�2���Eik��醘(��/��C� �u�^��$o~��k���J �v�wBd+!fH��@?�	{dt�2I!�p�~���q��靝O9������o|h7q��G`����$(�u��ǅjh�����`��;��?v�S���-�~��sw�7|"�C�1����;��4�~R���j�9+m4�\�I&x�w >qo���M<�{��/�I�����E�� ? �cL�s�d�
�B:�8�Q��G�d�.�_}o��<<b�?����_"��Iyh�I�M���>6.��ʫ/���g�S5?��Dz��r{��*)*=��d��@oo+׮��o��}���8�t��<ǁ��n��5��K����y5����JU����n�鍅I��O*��t0��N�s�vC�t���X__��棄.ާ$(�]Ɖ7��I����c��/�|�f�Y�T��F!�v�:��Ǩ{�ڨ�$�NC[�#�]��O�4��b��[���^{u%�ߺ��~O��Wrۧ��'o���eIMc�b%A�p���z�F��!#��xDl9
�:9�p0Gx'�S�AL�p�b:Ra�#�ؗ�ҍ|��w�7�q��7�W�7�{#�v��
�&�^W�r�� j���in4��^Q#����ߠML���g�f�%�e�O���6o_�su{>F�Y!B5�!�|� 0�p��P�4RT�Z�����	�6���WH�𱿻MJ̀�$���[�aL�`�n�~$6�w$��]=�������(Hq�{�.pu��fi����s$�7$�`ej}M�\H^z�g�5��eT�<��%��?[�I��|��~�l�ˇ��3�Q/S�E��t��WS�yR�i�P�O}�M��'ō0x��#�D��̀
Σ/��:���ZF�����Jpf�}4����?Ĉ�kr\ �ӡϻ{���;Ϡ��� ���E��^'�����~2���_�*'�H�7q03�`�˻*�}���|Y���f0ڧe�SI���L�7��  �IDATI00><DJ��Z�ڴ��� s��ځ|!t/vG
�0�1?<@Al�#��rzt���x�.W�!FNt�#� �&7C��9U+��w�lH�[�`$������Y��7WWp��M]���c�����li�&X�v	7_|�?�fvI�ҕ���b=������ �#4/�Ï"��w4 N��~E?&`'v�� ��yQ,4�1+�c�)��Wp�����+��O
���$N�;ӹ�)O����H��{�H�鸘MD���X��W���e9���;n��Ҕ�R�lι���c��+|��3歮���V�˫0]锵Hf!&w���8�k���d�υ-<gkHq�E��4�ɕ�RwQ�H-KH�/Z>@�>�ܿ@�\��Knބd�L]P�V��'e;m�o�J�����˞��lI�-8�|��~Wr�G�>�����P����˝�<awR����b|&6~��a}}��\�g���" W4��p�4
��V<�\�l���?�����>��E�иqn�)AQ�lF���tQ	�b �Jv�>
��3$��f�y/�5��=�yK~ER��ph:�;�G�
XF4�Q��(�:6�{���!���RX�	��G�Ꙧr�C�!Dt�	z�Z+m�Ʊ|���K�7٬�h��x	�OB�I��1����l���8T����\�����i�Ő�l���ę����N|��#͈�;��K��z˳����h��W�3%�=G�NOI��~e}��p�(�Z�.��ɽ�/�H�8�^993s6/�+�gvŢ(�  �J�C���f��g_[V�F��V��⭹#��.m��G۸�B�L��h8D�����U���Y����[1��Q�a��e$P��>v�t�_G�b	`�͌�#0����G�R��&�ۤ͛s�{4��a��{w�@���6�3��Ϡ]���l�n8?�����VV֐<�b8e$7RaPgǷ4UQ�HL�!�1���h)�B����@u����G!:�B�K��w:-�4������}*�zJ�Z�}�Rx��|��ɿO�~QHIU��p�:�� ZYG�tg5On��4;m�9���r��(�G�s���g��ig݌��T:-Q�V��|g��n���*O�}��Ⓘ<F��3و�ρ��rF�B��k6��
�@�m<�7�w.�^�v��f�썣��d���(ʶ��3�v^Ĩf7���Ie�x�)KX	��&h�GO9��#a��=׍�уGt�1�Kg����O��E�Qѹlr��p�?|��ǟJw�MR ���� j�f>����_Y�����a}����l���A�~Ï�_p�Wڪq�xn���EJ
�8M't��s�I�#��L$���%�8X9`�-�/ɒ�� 4�3�hs���X:Wd���>:���.��ѧy��}��+�7����b�n��Ln�v�p��1tw1VRRt��j� ��.�J�@H
Ԙ&����b{�1�A_zd��
��J=.���ʘ�K7�q�P��م��%:�9
�-�$��ح1������~7Qt�96"�o��}UZHwmk4���*��1��gǯ@�S��y�/4��`��kۅ��"w
Gw��H]O~�VS�s�	S�~�)1�*����u[�+�u&S����9Sb`�6������hy��N��s����Xf>�;3@�4,! b�u�.������1"%@��{+�.I��<_�H`��9��M����*���� }�]��/��o.�B9W�0�K3�6`�-�7��hh��c\������>�!P� �D,��������e��dӮK�p:�ޥ 
 V������ �Whx�!:P�a���ڗ/�"����=�� ~��օ5tV׈��4>�9��W����Z���������$w=�������Kh]��a�n���f��X�3)��7���O��ʵ�$(9�l����OؿV|s�{=\&���_j����2:8�M|l���Ӭ̫��w��:��2����(�z����/4���Y��	;�$�x�Aٴ B�'J�b�uM�Y�?��O�K�&�͂6����ټ��0��h0��;��C)��I�s0�)@ø"�a6�P�Iy�=�xk�N","�w?|_�s�+�H���P
�y:�c�;�"����ޣml}�C���l��]\~��ՋR��V��Y�;������:1V���T�$�d����b?�̸���K�a�A�$aJ��H�B*�i�@1���x��=�:���k���"ͫs��^�ݾ�B���54ׄ'%Hz���"�{�Zw��mN�S�$w��@,
�����o���u����s���������溫�������v���]�'~�c�m��wV����2�r���A���h�[s��L[X��/7f���6�E�6��2�R���UԀ~�����{/O�	�nV�>m�R�sx�)LS��)7���f�S���I.��cܚ�;�K�a��"F�"��?$�I <�?@w����MD܈������)|��@�'��������;��Iw{���8����	�8�� P��#xi���"����G(�C�H����{�6�� `E#K�{fP�=6�Hi�*��-W9����-��zg}��w%�k�+��@")y�ZJbᕬ����|v�����������������DL���c�1^���I�x0�gA@ۤ��}�R���*wM��!���n}����k�3���>b�]z6C~N�j��v��g+�����l�S{��Ա�us�QW�8�]��?��Y�H3q�3K3Q�ز¥�8�}eeE�G�(Q�
>=�G@�v��HQ�ٸ�Z~���s��ϳ4N1.\�X��4�k���ɓ7!����#\S�R�rt쮼���t�M�z�YV%Ù��-�V��4+/;\��>\`®,S��e��ɛ|e�:�R F�h�i�6�/��K�K�����g�k���y���c�;M|��G��% N%��(�q�_�]�\�����Jln<�������6�=�Z�he��J[*�[��W8��%�ʡ׹�ظբ�5q8ܕb@��0�2����5ϛٸ��l�^v#������ؾ�f�x���G�D(Ԣrov���yq�C��Ώ,�l]ۥ��q����פ(M�]�Z�\d���.���s���&*j�H������%���s��!��k�˨�aC�cBg�/ nK���}�ua��̚`1��ak"͕�q�PWF�[��r�rZ!�kg�s�Q�$�2�`���vL��:��%�|>�x�.�p����NQԅej9�Ԁ~΅�icq�����[�N��ҕ%k.,(EU�#\�j��Y`��=vѮ�I���<��t;�Jc��u����jf�L~�\
��^��Z�>P,~�{z	��W��@2W*�q��&�]��FL�w��8׌�`px����!���F�l�����`�vf��l���Pʘ�u>�/~�\���p������_܃�R��>G��M��V����	h��ؑ�:���6e����8�D����H		I9Yae��˦������9�`Hc�Ho�:������"�)���X�iD����?Ա�p��3��)z��<������M���C:g�� ҙ�ͮ#��gׂe�;f����R���ee���V�{!���GI삫�6� �ʚؙ���XQحHm'������Zj9�Ԁ~���"���f���F^�'d��S\u�#2crtb��c9�n�am��x��ި�����7o�v�����2{�����T���Un3aNEl�f�0o����R�l��L 6�2�Ǡ�)^>N;�<o6�����V����(����<](&�2����#>pSͺ=�+�<H�5]�;F��L8�Lr�C�J6Jc�9}�׵emM~[�O
�(=��s)�&�ͥ^RT<��p�U:7�syh�Ү݌}��Ȇh;!���	�v��!wd�0@��q���5얟K��F�K�+�kK�ׂ��}j����vlTZE&.5����Z�+kL���R�eǌ���3o�� t_�K�H}࢜��'�Qr�r�ک�=;Y���QK-g��Ϲ����aT���7R�%﹕m�XU�JG6-�r�GE�+&KkN��j���{���o�,&]�lzQ����$����Ӭ�pa�l44w/�1|�R섎���|Ó�-�rC�A�Y�9�g&����~7UR�Ey:�[��n�*�1�s@��՗T5q�˼Y��4�x��a�����+��/t4��Ag����8v�r	_%��I%=	��J���J��7_R�B:o%l�Id?����=`�2Ǧus����vixR���A n���p{W��̵ُ��ܲuu�n�F��s����Jk4ϐ����51c��=�|W5)utm����5��1�� =����Jg���k��R�θ~�\������}V�`X\�����Z�(5��g��KD�>�|�s�y6�����Q=%)�$�hB�m���(h�J���V5�n�����o�ws�mQn�q��}X30��y>�����L)\O"湁�o ��n�!An+@g��p^0��b)`�n��m��&J[����\j6
��X�';cČ�^"�f��,�9:R\����(�=0#f��'���'`$��nw<���b��i�qᐎ�y����o=�>�����%��m�K��P�j4����@
S�a�>���+}lt���t>���%�N[x����C�vM7�|l3���x�
P�)k����x�<_�s��A����U<����m��S���6�K�xNS�2����0k�W����3J��X��n�=
Rmte�{�*���Lg3�FuL�Qu���-+/�C�4z�� 2;��F7�Hd�;nY��g�T�:I+�a����8��S�rӆ�dN�m3Xq>�ϛ��~�^�P"�=����pS��@�+�5ڜ��-�y��Ս�;)!7�q'�rm��0��h>���(\���@2J�?}Gڗ����?�	�i�W�2��t��R���0+�%$�����ܮ=����1Vh���E{���B����=�?��{-lz�����K��f�t��.�K̞�h���0C�Xs#z����cdN���l��#&v�lp0[7�l
^e�L@ݬ��;�qt�,d�O�y����p/yυǍl�k�R�kgH�0&:?.�f2�zq��4��ZYj@�2�tLЩ%�v]ڐ������s{�����S>g�<Ό�l���V�����l�8�����m0��b�6��=ˆ�N���~�����=�4C�9�t]u����D,l�)�ʁu���!Q���p-t:w��]��=��OV �`���$Nش኶Ov!n�\L����l�g�Q����E)ǚ0�fL�O�S�����Y�($u
�h'�k���I{t��j�z;�v��X%ec���у��\�{�.n��7��W�&���{���O1����������!�y.�6:#��~VW�H�7<�}x�/������� ���(�I�(�8q�8S���`��q��Ocz��M,'Uő���g�cM��bmɵ�`8ʏ��|�����x��r�Q?D-_(9���+�п�r��6oq�n�x���� .�hS�Tf��YǊ��?	���� �yS�lʖA��f6Ȍj��|ٗ]���>��O��F�0��r���=���9�ԭ��/�_\�y��Q|/L���r k��@r�}b��?{o�+Iv��}7����^����ޛ�V�w�5�F�F�!����?��6�0,�l@#�3#��H�ɮ�j{��=3��s΍���\ޫz��f�<du���nD޼�Y��6�4�8OȒM�BN�7�����Zb�C�8!V�6��%��*ɸg�a�$���K[���x��_`�qz���=�o��ʒ�8�;��,�]�����N�5�p��&�}�k8����3����'�[�n����`w��n���hc�����}�ݹ�ĵ$я��֙��K�F���DJcwSR�*�PWZ����-�t)+� %���2Uj:1-Mm�y��֥P�w�gDLC/6���R����(EӺ٩5���y�����T�!̊���^p�Wûd��TV�I�\@V:���p>�Vk{ݜ�s&�n`β�k"�&��U*��lQ�X��l�8���QX /3wq�pNc~q�iR���x���.^M	`�ts���	�vuô�Tb�8h �z=�[�لM;be��u0[����ex��vٍ�&��*�V6�j�vOsG��/�T8Q��"�^6&N*�i�����Grօ�u.ME��y����q�������>�>�[��ڦ�����2���@�y��w���zo�a7�#L��h�3D+Lt����6���߇��]t��h��w�F���1�s;��O�I����C\�u��Y Iy�x0m���;������o�5>�яq(�m1��/��o�i,�n#i��q'z)~��͝M�X��k�/�$�lR�<'�.&��Xx�����7�~�d����O�я�kyd�ے�g�Rऎ�?ϼ+q�a�j�i�	��:k�2��Qɑ�Ԯ�p�O��o����v��6Ɂ���#�n��V"bM�-ֶ�>�З���;�ܚ�D�:���s�E��g�������;��.�_�|������K���lr��9[�I=��#:Rc��wNM6��V���/K���ڙUΧL��m��.Y�MS/�I�6_ұ�Y$q����l1�]��1�;�_��5���1��I��p����X�1&�1T#�\�4�(�U�,�I��IL��r��_�����s��,���"|^]Jޒ�'��M��"�����û�5[!`���5��l0����
�J���Yh�ۡ�Y�n��]�#�}3q��Z���ư��B4��o�n9��o@�~��)o#��uc�ِ�y~6������F�1�[�����NgA�mH�T~~��:�G�q���c�'�:|��M�ǁ w���)'�XY)�9�b-^	��5χ�	�K�l��e��|�a�d(Ϝ�-���v���)3��l�x=8�2�3����d�>��Q2ݚKS�&�u�V��+��c-���/X��5�_sao3 -��-���Y�6Y����ų�0΀y%Sx)��IM*�+7�f�Q�Sܕ\�D�0" �rh+k	�hc��d�Y�d�b�[l��D�jMڔf��(�X�Eck8Y��,<e�7�u�f�K�8�{�� �7ep�;����f��~�5OI�8 �vk4v:'wR����Z#i�v�8?<���?��7�n�AqY��dY3G��j���&�cl��:=�pD� aM$�o��*t�{���XZh�E�Rw��4��]-���7���{x��0�m�ǃ0��p�s9Z����g:'��M_��5	�&����\}����O��\��ｏ7^{C�p}�I����p���Hr�#<􆍭<ͪ^rU��g���w�Q
	��U��Ȁ]O+'$�
�L��n�����	�
*��'~'mU
�hci1�XB���cE����K/����\Q>S@�uL2�"KS�r"ێM���ZI�&+���f��mZ�t�ҩ�˶+���O���%c�.�Sm �����#.���� U��m-��%�k=M�/�P�92�6��IY�]��I?��P�r�9��M�R#�]��C����K@O��y�!�7o�Q7a�ژ�Њ�Tl�8�;��u�8 虺�mn�	��=>%���7H���A
�`B�4v�D�.�p��' `L��͛J�1m�Gd�'�	��	Y���f�a�n���w0�Q����E��@w2�.q5z΍z]������=�1�Gcc���㏰ww_����F6� p����Mc��:HI��H���C�H�ܨ�O�3�߭-�ε��3K_�Tä�Թ���Y���<J�ycȁ����lK�C憷�nN����I=�4[��lq~�$JZ\�o����/Y�-��ge���p� �[���R0�+�їdK���ma��i���/�|����ϗ��mZ����˸u#�i�	��-�ɐy��ȉc����<�Z����U�:������L\=�v�l.�b��D��mp��a?�2.��,��V�e\�SZ[��s�<% ��1l�&L�����SX8I�p�c��7K�=��?��헄�\���nm0��9��c�\��Ԩ��w-znt+l���G<DH �ڭ;�8r����v���7h����n�#�eφ��֜t~��}��&9�R
6,��mt��1qN��KL�{B���ۻ�Ɔ�n���E\n5$��n4a���1�y���p�Zw��Z7w1�1�}$���Y}H�G�?=�7id��4>2�w���Σ�N$���vݗְ#�}�CK��l�6��P�רK_hiK��`Q;��qv��Vz��b����CP>)4ܜF�i8�ٻ I��? \��
#��XIoWF���������NHkY�s����E�K�DR��RS�Uj�0��j��y� ��i�5c0I"[��2�Z �V	`uN��e1s�\��Nd���d4�e��q�(B݅�fB@����%��{2���ɍV�ҍ�#�f1c+3�1kgf�Y����|DV:��C����I�(w��Zm���G#h��w�[`4�9��FD FV<�o�sj�v5��JV.�e�|Q��6�h	�0�Ԥ����C��P���v�t���h�m���%��c�������	*'���]�jaBו�{��i[��g��	\�ѐ�C���ᮿw�%�����1�~�����'����p���r\�푢H�����c��C.׋BR�)pu��]yṆ���M�����������4o��e�+'�} L�|:K�_/K��$>:(!�H����-��!ɉ�o��S��Y	�.l�����7ߗz���j:	�k�Z�,�I�E�e]eq��*��"��q)K��,�B���C}s�(�Ά2�q���-r֡g�l&?a+[��y?m��˴��o�e�����	���Z�6'�J�ɧ4���)6� l6���K�����dc<	ɒOP�k	��[�HQw�O�:wt{hp��F��,$ �ݿ+�v%���%h�(���EV1���'h�Waw���|�B��G�龽�1��jZ|RX	�0"I�c�M�6�8m�U��jC��HY�sN 9Ɲ�ׁh"����'F����Fޯ7�:)p�nO��P�Ho4}ɢ?��vQw&��$�q:x��Fs��F=C	K�O��k�}L�Qo0�,):Ca���jc۩���<��EO��d�*���R�S����-ˆ��\]Ц\��C�;;>ц���<%���R>��}����r59�����I�d�4�Q�*��*\��V5���+�п�b�c����Iǚ�K�ak��}z�`B����vF��ed��- �ˀy�M�,�=�k�EB�I�s�Zv;NF_�Ɨ+ݝm�:��O�J�������|���N�n0;.u��=ÊR���� Lj�mL���yM���n����-ن"@' M��ڛ�G�7����ED������d�O��
g�k.+���{�����;�\�[&���o`4��%�k���t�?>�V{7ɚ>9���C���pF�r���wo�ox��$�8!���L�7m��IA e"�W&�	�ϑ�Ǩ���6���C<���a����=��9Io0��#�vݓ�������ҊUK"�%�[<�[�rt���O���d�;dݓ�~p���y�nCyFhq�Ye�nU�z>�.��7wٛ痗d
�/��9i��*1$��^"����t����7��LT~~~vcRl8��5���[�p�@F�\���Sm[޺}-W�5�_cye8L?$ۣGV��~��]3�_#����7��Ǉ�=&��Y�t�+�o�Jت,$��5.��:u��-Y�P�!,�IBO��nk
��c)D+5�I����s*_�ɲ�Z�:����1xm�����~[d��ހ�GY�-������ͪMR]p|��3�j�o��jb����G�5���A��Ï?Ĩ���w1�X8{��X�M��z�0:<�53�9H	�{h��7�t6��yG8Ĺ���C�>�a��G����؟���?D���wQ�n����-�^���7��9���F�(������|��|��1��=�����o�܁�mc`�tp+�c���~4�1����k[m��?,7x�

�Jf�O@�^��c�ۥzG��.>y��X��z��]t��q���B�J^��s/t5�}nNA}.�R6����/���%�M���;�sDώ)y9�ͶL�#q����aO�2l+�}���$�镰U�Ý�:�u��Z�,k@��2��$�Ǐ�[~S�\�\�T�ͺЄ��_�����Ǉhr5�p2��䄯X_�Fsa���+[B��Օ.'�������|q^��s�����1��tۚ,�Z�k6��b�$���2u+�M�X�\����K�,&�I"z)��^d\�����|�$�	\���������xB���1)R�h��������:w}�R��DZ��ΐ@xOzn��л20���J��cL� x�u��K�p�����Sb�͝=:��d�w~��r��˯��\�N1�{��MR0��F�q�Y��c�U������ĭ�n�G8��O�	�U��t0v���(U5��M�:)bmv�K�_<��!Ť�qzR��� ��K<2�ՓjU"�����j:��s�E
��.���E4�8t0���o��n6��S�=9��-w��!5-d������}2� 8�0��L���3wsS;����\Yր~�����=|�0}m�%�|�z&)Lf���ƍ=�[Rkq�%ŵ�0�~�����'ə#Ju�Z���|�B	���1����l����ҕ2����SK.�
h��h�愰���!뫦��-
�SJ��&~:&+u|��9�y�l=߇��R瓲ĉ}�}(1�t4�����s�� ���	i�6tϏ0�b2�氏��[��\Òs����Q9�*�:# ��	O?�E`�c4������ �>8��?�a{�,�[h�Z�l40"�Ud�;���	���K�[��O�{D�9�ߏ�P5�'�H�Y�V��'4O�~,�#[d���\H�%�)��<9�X�O��s�1�g'�]����ovշ�s��L�_ڼWZJ�*�2�k�7��uo�X�V�*�������t&��1��'ҷ_'�g{�,V�%hi� �D�����a�{�(q�U�N�3y
g���GGh�We-_h��J�׀�rM�߯�8�<bR�p8�r'v��d��'5�4I6��SX�J��C����i|q�ڴ��$ͭ)��~ع,���g��ϋq���;��1y���	���&Fd]q� ����X��s�pK
�u�;`e��bUs�_���(P�:�f��d�ZA�#�@�뮙�5��w��96��4b|�),m��c<�к�����R�P�dQsr�Lh�n50@�bpt�6Y�L?C�NN�ڢcGQ���cd�8��ؽ}���Ǹ��!Y־��6)sAw�'�x}F>V6�4��i��zq.��=������0���%{��q�	y���K�g��V�#A�;!E�[Ɏ�}}~΍,��=��]O{��lX�f���-)t�b��`��?������?�oP�:�|�-���Z��2#SbH��2�'N��*U� R��J�����Qj��p�>�Y}�k@g��?%�y�,�uǳ��&d"�U�d��� ��&��z���J2}���eF/��g������\u�ZNQ氙�����U)���u�m0�;�z@��e�V���&'X浢>Y���8��7=�� ����&���AxL �G���]n|"�N[*-l�5�V=�8ڔӱ���#�; ��𿇟 �^扒xt��v��%�L������}�98>��J�	��Lу��9���OV$����%r�����O6�NB�{*wW�5�A�#�cӵ��ֵ0�N���,s�%��F�����zJS���r_�a8����:�C�֢\5���5��<˔��%)c�*��;f)+v�!Qu�N�y&���р�M�3o�������Y����bҽ�st�m4��E���sG���_G�^��0�A_/.�kjD}ڲ�k,�SS���-�1Yla�ͺ�#Z������Ң��ƭI?�D�f��?ʕ�ς}I��e��*J�2Z�jv󒅟=Qև�Z�A������9�V�#q\���=�3��:Cn"�w�$�y��f��M���Aje|���Td�����O�A���6�N�����Z�Ջ��$ٲSt|�@A�Íz����YI ���eK_���2T�h3�ඥLt½�E1��d5o�릜�>���v-Ò����Ѿ\��`;!P��.j��"0o��\����D
y�cZXӱ���мJ��e���S\O/��!��J�.ES��z�2Wr���,S�GI�F-l�g7n�{�l�J�iO��B���a �^8� ��Rß0�}?>'82��x��h�k%k0�Td��X�8Мp�{��JR��0�i��.Q�@j͖��0�h+O%2-3�"1g��V�&Ϗ���ԕ�t��D���{�������{CWk�j�P�rfv޵K,h��`u^�l�p1 yd%;ڒ}䩰k���NBV3�("KՁ�d�8�O?�q��ω�y쟓�TƞggϦFǎ黉88�ό}�2-9���'z��D���2o��/ceA:�i��y]i�m�̄�ʱ%#��S�2���f������%���GL��w�rK�H���i[�Tu6T���33mN��6ϒ��z���5� ����_ͱ�C��jn��s��ժ,K��Q���<䐉(���0�	bzF�o�VT�%Q�d�$1�`�� E�;�0+B����3�7����:��Z�KZ�Z.'k@���J|WZ��Tʝ���*'r%L|�H�.����]��m�}��YaZɸ\k��4i-��)��'5'�+�*�3���g��*[ʏ-b��,{��.m��`E�n�Xo~Z��r![`L�^�2���ȅ��m�:~2Vi;��gI_r���j�E����{�0���W���=K.7�-p75�����+ӇF���0 �b��XB3>�����6������_+R8��^"���\g��+�W��:�M�d7^�-ɧ;�$��@��y0.f:���=2O+H����Ф�*+ӆ�c)3���\�j/g���ѾT�s��.��z������pd��T͓���GB$���ܢ���67M�WfÓ��-t������YoH�°ەH�;�
C0I��	�2ס���Y�/I�_˯�|���5�_gy�(�R6�~|���wN�����H@n�����z���P�Ay�0*>2�2����͂)��Y8���9h��]�µ�Y��,@�ujVe�Q���2es*�F.4�l�օ�0�t^�,�^MJL��4��XEY��z���ñ\'��IN�@$g2�n�I�/�e���w��%kYkM����+%TuVX'��2��<Ge�L��]����m�͋�����F)I��X���Ja�� /!��΀��Ϳ�� �'vM�>�y�t3�2��"&��ӂ��+�9�L<_hW�4w"I�ȵ*�/+�ĳ�QL����c�f��h��{)q��k�ONK�_���P��M���,I9�����;�b��-!���J'�mAGB���J'p�,������P�t������ܞ6���п����ր~��w������߈�"���Yok�82yZu��
>��G�1Z�K����,�)K�:�B�5���+��U��<s�ԥ^��T�\�V���B�sNG��}˾�2W8�@���pwJ�ʷ�]3;^���d?k����;sx�mWf��5��)�(Zυ4U?��i���7(>��8U`J܂�NeU�I�ȟ��_y�J@{���K��o�в{�^�J��w�5�l6��(���]c��I͡	]�.zn�-�	)�L�[G[�MR�N�?��8�`rp �y� �ӵ�D��xgg�_��z}U^˕e��Y��kV��8�l6F�����[[�Ju�$���GmOa�͗���M���YcK5K�%/�J�|Tvk
`�q�����)���k�XK�������$-ޮs�qv�gI�Z�o���*TyM�Rx��Lf<�\0���T��+���cf��gt�8�?��R4~�&�m�<M�d�%�<�A�x���4����2{6�8'�%���7u���R���Cp�<.a5U�r���.�ͶNk�u}-W�5�_cy�Ⱥ{8a���k�/��p��-�on�񁄻l��G!�[7��&��BR�Q�V�s�-�<Y-u`.�/�U�*��-�e�xn�^$3��b�c�S�%.M[��c+��R��ͨ���ZZ�U:Fa�5W�c�~�=_y+��Vx.�P�[�@L��e5��2mO�i�b,�4Kp3�{9q���]2�{n�����_�8?'���ǥ���%@oz5tz��co��p�P���fD�>� ��yc�v}�e-W�5�_c񏷬�٣���'�'����[_�
��v�
�� R��Dg����x�����b%N$%��:��~� W�cϭ"0fK��za\p�W���^�9_�*M���Ꜿ΃a՚�����<���ʢc��߅�,y2�*���Ye���k=�o��
U���[��Z��*P6H�G�3����dBiDd#&�vµ�;����w�f]j�'��r������z�O~�K���Ɏǚ���(P�	.kkr�X��ؒ����\Mր~���<B�I����aO�G�N8SLڎJ�H^�h��� �wn�#Zz�i���s��f���C_�ޖ�1��ʖ�E��C/k}.9c��b��l�߄���f/]i�¯�֖y���/:��k-QB��������Z�$-������,U��ed�s�ϵJ�Z*Y�d�KV�q��������й�!��[�c�+o��,�hb���`k���H�w�ݰ'E�J���D=����\�I��hۉi���<�T��k@��b���e۶5�XnK&���L�|�+���"��&dyܸw���bSR m!��53��UN�2��.%we�.��w��S/c�< ̾/V�~/qqR�kS��Qn�,h��-�ʹ/�U�t7+����0IE��MH����S>J��Z���<�ʅ�iuD)T�\�+WvL��oc���!��Xz�H1#���p��Yn��i+���_�=B�0V:�ڕ�c��g�^�::���ֲ��Keگ���mY��"�Gh�|�.�^��LbG	�I�u�u�.������I���6��MHQi^�*m��\��_�q���>f�~�oQ����]�V�E�vZUd�?���܂�Ʌ��J�[�,�%���S��<�,�\`���K�R W��wsY}�=`��0����ke�INꓟ�)��D8�=�ۛ�x��Ll.��s׻!7��`�!&�=��!T��w�+�QiV�(i��ɉ�߼u����\{Y���[�G�JU���uZ�G������=D� ��u��ݷ���Oj�����.����%��*T���d(�ܝ�gMÀGN�RM*��PI6�7U��reb�����5��򷙆�����ƿ�Q=/XE��6�'����f�[���C3�6����K���h�eu�x�U/A�j ��M�|r~5�1�_�Amf�����Tm�BV�oi���r�L�k�����i�y,S�/��]�<�T��ma���<L�����{�<}B�y*߭-�y��-�rl06��V����{��jkY�e��X�Z���NL���p%�Mֆ~�v�e2�}Z���������>ܭmO��%3�Y�Έ>0�ΰil���Xu'�]F.�Wn��M�"�e�q���(�Z�ŀ���-?�H�be���t$e�_����ÂP��x�±_�,Vf�	�X���2�s�g���NU>�3Z���S��|1H��:�lm/�$b�vN�;=�"����a��J?CB�#��?;SJ�l�)xمϜ��4��έ;�DX�Z�(��+�k1b�V캱�ׄ�F�Ht|����ܻ��F�ÄL	����\�a��h�����,gw`HF���꨼�.��=WM +:weg�O�����U�A[���)�M�/��	R�QO]=��w��o-�4��(�j�y�9S��irO��g�S����˲�e�
��\��܁�~� >s2��&˛���$���}���;@��8�H�DdeGR��T�����~�����Ͻ�8�I�3��y��ww]��|�;�q���|��ą��_�/�E��������.]qo���O�~�M4w�`�
�<�WjSk���������\�-��q]��E%��eeY�օǠ���Rb�b1?�"�^��^ňg��~�`Y�����:�3�*#3����?=���y�|5G�����m>��*U7{5'b�D�,<C�1Y�<�&��N<��B`��=�G�Ы��m��%\�f!�v���4�Cl�l!�j��sbW>w*d@ߡ��a�l��˟�`-��|q�z �Z�
-NI�	7�h�k����>=@��c�޸�ma̜�ܴ�����7_�?�|t��4j�s��Rfz����	�gU�Ϲ��-�M���Y|Ӥ7�z�׳���.�U�!�yV��>PQh��\C���C~�ʹ�b�����]���ߞũK/���b�{��¸��g�g���0��T1��B�����ƽo}���:�D�0I�� ����3��%h���87��R�u���_��v�w�N�~E_�Zֲ�k&�x�V�GvD�!��bۖ#��ggP���%��֞Hܬ��`�嗱�ƫ���g�%K��u�ؤ���o`^D��\s�9.>�j��l[qLy�eu��c��<��ؔƱ:����:E�Cv��2 _�z`Yܽ��^���Es�s���q=���(e�	\7�g��6�~�K�3�6�d�(D4!!�\O&��?�ۃÿ�$)�#�:���%pR���)қ7�h4B�e-W�5���ɕ�>��ڲ�����jq�J�
ڣ�F�О/n�D���~�,
goo������Mw2�X��t�*O\�9�|z	�����bU�s�Tݵūҗ��������.�/�(y�^�<��b�Ҷ��YA�����u��]&^~����~9I3τ�D��#�pMd]�q�׀��!���rژ��)�F��:=�	��h�t���rV

�Z�9��q����No�۞��j��-_����Nր��&/��G-2\ǵ���斚������p�:\�"q���B��F=���u��7�	����S%�w�8��5���]���Z�lU�̖��Y��kua�]�Se`�"^V�Iq��+���˾�盏%�eY�x9���Yٚ��C����e_�%Ԓ�ރ����y9�*�L�Ϯ�,;���V�׋��l1;���J��cecL
���p�k��o�&�����2���dp64�Z������롞�ҬM�/Y(
��!۬%��̽��9Թ�Z�/����ӗ5�_cQ��6v7#��ZQ��m��%
6�v0|�#춷��ub�*��I�d�M ��7�����	�	��8�&-�67��\k��cSm�s'SӋ~�P�֣E�����b���p��}��rE+���\��e�S�����k5)ή�EzA���|�:ߖ�W�ҾbЙTA<-k�!��b�uz�c�)#ew��A�Z�f��R�� ���~%%�b�/ �K(���蔕���`���TT� i��b^p�l�dsH%&��|e�8I���(v�4�# �5kx��~+��~B�:z�}��5��8{�>����'�h�7V�7���4�S�����m,�V�Fۻ{Q�n_����]ր������쁬1~�S�gK��on��a��?����-�i��&��ذj5��M������� �,�=n�BY���r�nv���f[�"�<~F]�m9C�j�3ww����S���Uɣ�B�]ʲ���L��/7g�<�!��0,�gaXf����6�S��u��5YNL��>�b!�n��`��������շ�I���p,ꈎ����M�Cg4�����5�x�2�KJ�0L�ʀD�fX���[��t�*l�]-z��\b����?u�����B����&L�f��$�)�G�p��S�y�U�d�$n$�EE�EJW��;x�[��{��p��;�� ,�L'�D�!�D�|Ē�+ud��<M<���[������ԥ���_$���2p�$�-9�2��g`9�*~�`�g����`��e��Cww���\O�C�����V#�v� ��HȺ���n�7緁��d�'��rOb��3��?�Eǈh���I ���Ag�ك�G4�=��.����\?�z���q��+�Я��a=��$	�P,��tŋ��;��]� �3!$�]ԶG�^���^��o��G�����p]S�SNv�E��R�b1K��r^$U♹ϖ���|g��c^�\��u�t��O��z�|�~�������I\�`=��*�*��������|vi�j9α�f�	Z_��;��y��I0fk�v�&C�NY�n�w����mR�d�ۡ�~a^��M�ga
V��7�a��դ ������;�Z�rEY����r#�aq�[,��Z=B�:��w_;;�km�s�ڨ3�;��!�@���x������p�����HV�) ���y��d�'�d0S}5���o���,�E��5չ뿜�������� �,�I�A-���M�kMc��ٗ�sYY���f��m/�U�Rd����.zx�(H�T�^_gaqsF;�MeP��6o�_�2�q0��&tnu�`�L�` �&ύf[n惇�uo;Ƴ�,	�&�@�$K84��wE��ɢ��V]ѹ���>�}-���
��[�.BV��I��[�h�i%�-�\�6:8D��e��j�0gqَ�#�g�n|�m��?>FG����)����,h��xy�T��K�;_�l8ϫY�eW���\���L���m�L����cѵV<f��j��e��.�
_��){q#/�,��Uv���6i�MC@�1�A0���;��}�����]����c��@���F��arx���Ö�ÊC�m���ι�cRz�p���Y8���G�-��ݞ�N�k��Z�,�B@_���Z4�T�L,�A���Ս3��(>���9���ϱS�acsp}�@��0f+1�;[x�;������MZI�l���P_���R�P_2ƅ�>�=V���-<N���y������ܣ�����_�!_}�k������+d��<�SYf��d9���Y����+ϔ�W���3A����W�l��.���/z�'�~��9&��|�ӟ��x�F�N�%^.�VH-[�LDr�ey*l�#J�~��I�k�P�f�jY�ܯ�褭�� %�\~#�'��8��V҄b��)�w��5��	���i[D�GX�q�7�����#�O��e_�hQK�5+������
+�MϾ_��/�6��u�<�>uO/.m����xN���)��k��t�]JY&	)�p�&��o��~I��!)�l_ǃ j�vf�#0��;8����[���d�v�&
l�M�����R����]q�Q$8�ÿ9ϱ�8�����ղ�D�X�քVm��������g�A �]���>����!�({n�!��;c�u�?�c�$L�������Bw�5��$�5�Χh5�	蛴�]�?�EV[�]��MMT	'�xUf��f7ΐݔ�
P\y}��*-A��Z�E(]/ͳ��q��03%kK3�i�`~L�N�Un�S���H���<6U�0X�I0����8�R�^s�
!ϼ4���D>u���bE4��M���f��8e�[���o �o�GstDV�5L����6m�aG,r��O��9��	��{pB�e�p�2y#9�����a[��~F��r�����bs�.,��� >]Y�5{�[�ѸI ns�-T:���ق	���G����Z$�%"��$P�t��b��t���u<x珏Ъ70!��[�r�y��E��6h��_��p�WeUL����e�[ԁl�5�lY���Ϫ�h��.��d����3ӗ�{r�����|7����yq+kNS[i��2{�-ٗQ��� �a���pBs2��������1�c֨�כ�'����2�5"0'v��P��F��tl;;w�t�H��f,yf�+y&!TH�Ȃ�v{��E���~.���Я�X�����M��d��
�;�E�NO~�4nކ�<�Y�w=ĜLdJWM������w����u�XX|:��$ 6��U�%;a.L*[T��HT�H%�9Z��yҌ����3y��%��;ݟ�g���m��K���Eu�In���',.B��!n)�빿W��QԞ�_��,cޔ?]	3��2W�cByJ�~D@>rj�b��7��{?�����d�d����;Rt?Et|B����=���O��h����|�?�e�kH�a�cK�o�SL4�nw&�aw����s]'׀�u-�����ތu���0�(�-����K��L�v%������O��jA��q�	ocw�,���;�x�w���ǟ����$��b�-B"���о��WWe<_�^.��s��+n��ܨ�c��]ZΦ����>��+�����@�r�]������	ts���3���M��Zp�u�R���-ń@��V��]��;�wnc<��vd�7}G�g8���ku�}�h��?A��£�y76ʫ9��2@W���@n%t�X��q]K���Z�rEY�"���Z^��R�r��d/�y$S�iэL2siQ�R��ÓS�� zB�bo�o"���G���_~o����8M�
�x:�lpܒ݌!-�N֗�ܬe�V�d�>_Dr�H�-�7@,��n����������֬	�O�@�@��5�p�
],�y���K�@��s���hb�����Tו&eEL>���i���v�����]q������_zx���a0�!���p;Ա����p���m�����C�Y�����m8\�6�=L=8��o^r�q��tf\���V�~v���劲�E�ys�8��`��Q�xq"^ld�x��E�H���u�u�o�'B��z.z�u��0b=-���}������M��O��ÈV�Hʀ�JS���b��U\B�e�����y�K�U�̖���ˤ
��b��k����|�x������l��\��7������\w^=�%w,��BV"i�Y�m+���Y�w��5nh� $�36�45�Ο~� [���WC2�1Ƈ�h�<�ܳ��1Y��bB&$Sp&�nF�h4P�q#�[[ֲ�+�Я�$�0�(�X�$�%#+�B�3l)�ы�8q�a���>��V�����7(\�}%�cH
���=|��~��tq���-�w83��	��E+�*�eK�.r�.�*�������u�*��^�:�b��}�����{���-X���]��������(K^�^�b0�C�9��8M$�Ӣ9:I"��`�����Z_����GA �E�8@������5[蝞���!b��{���{jI���#F��q鴑���1��b"���_����6`-�@ր~�e�0򞒡쨘=a�PRV#��,Df����qG����>���ۨ�{	g�s�u�-�!mK������n��{8���{�t�&-�Jb�V�1}�^Fڡj�N�!Ec��Eekx��E����g�^=��1aa«��g���5�#����J�.�����������x����b��0�����r'�EմZ��"��V����hTP[��]�p¡�z�{������v�ѐ�gI��?B����g��:�	Ξ>���	��M �Tn�%��FѱH��ٞN����:٣�#4�l�Q�7���\Qր~��i��Qk��s��(D���8Y�/ץ�&�~G����>F�o��^�5�����<��\�F ����|�>���ca�ڳ4�<����=/�	�lu��3[��;c&�P�Ļi&��0(XEs�JDu�3���.[�feY������zw�|A.�ȮWd��X�<����Ў�ƛŀ�J`���*�]�t	Hs�c�^�٫W]�f>/_��& O���>�5�ҧy�~N͚'�?�>E�+<�Mu
%β�{�x�$
E�T�\��N�F��U߶�	Bt�N���o���p��n<�8	���O���@�o`���HG�G�h�DL�6������Y�����\�?����s4���,a��Hm���ɉ�|����C_�Z��k-�77�ࣔ�ՒDbڦ�$� �IP\j��g��D�G�?�Ų��#�Gލ]�{@���i)��v7�?�S������G���y�� �>���ifQ��d}k� ��LّY�gA�����9\�Ό�v
p��\����ؙ��_>��dQ���⎸�N~�$�'B/8�±��_Vy&���#͒��]e�̼	��Y�D	b�������?�#��p1 ��S���!P'����9!�6���5:=A|v;@�����D���*\S�|HBe{d<m���Վ�X�Z�(k@����mŌ����܇w�=%�V�M3	��ה��`��>Aݭcks��&�Ҏ_�O<:G�Amw��|oӢ���������;����%9c$�3�S�R�[Nb�^g�p�ga�Y@�%O䪂�l�y
���X͞����E�dq��iq[a�W��u�gp�&<
F�!-�/^e���N��b�[xBVx�����w�vO���+�� 	9�����8��?As<A�����X�7Wq�ZV|�p��B�i�:���]��ߍ���+�З�lF�Wύj����mF]]�M���{2��m�.}����?z�N�dk�K��I��AB��K�u��?�6�<����ﰕ���l�}�����2�0�t�R���hY7����\�ӱ>����v��].��Բp;ԜR0gvܯh�]��\��/�.�����_��sZ�n�<�Y�4OIC<����ob�{��-����w@Gao�h#�t%�c�^�9����E���%+޷-�$�d��˨�R�Vp d�V��w��Iҏk�徖��z-�� �p&�X��65�3+��i�w��UB%)j��-���?|����S���oָ5+�I��N�?����������r���A��ReܿӺ�c��y/��y��M��Y��Z�e]d�YJX��2�O��__D�"ձ/�����l�υ!�B)��y� �zN.uN5ec�J��)�\w�(��Cs���[������H�d@�I��9?���"ؤ�F�Z�,:���)� B��I�����Tg��,b=����ۢ�p��ٙ���k��Z�,����j�V�e�F��3�@(�K�S�yw�ٝή��L����798��k���ژ���-��=qջ^���1�����[x��'�}�'��c�Zy���pnV=ǒHR���q���@[�Y�+D����sU��Y\���j�,��ڿ�1e`Ϗ_�ٞB�rUT�����X9.�?_�^qL�<���'K�T��+cڧC�=�yx���ė����}�u�A�'̈5���!d@'`�o6Ix���>��O��<�	�]Wڡ�B˱���=-�e��	�L�38aO*:8y/��A��w�r_˕� }�_0�}���D2��L��)X�t�2 ˠ��-���Bfp�i��st��[�h�ZR�������d��*���`Fhܻ�7���/�#��RҰ��^j�,���D�E��
��eA~U��e������Z2��m�0n*9��3����gn�_0΋��	j�
�E�^ާ�/�zL�je�'�[N��g]�B�[_z_��?����H����a�Oʢ�q����	���� w��k4��O~����Ms�{x|n�
�V�s�
�D:�(�����Ω_���3+��plx�ýް��\U�.�k.I�:	�g�n���ĲaH1��62��4mxA�� 5��8��?>�Nc��0���#�ک%[�`ތQ2���[x���u�������D�UI�6m���ژ[501Kd�c��VK�E�W��Y�U`.	}�j�r�/��.r�O������U { ���!�~�l�����[�e/�L++WK�]�8�}@���n��;�޿�3�+�ʾ�QO� �i!�H���`�o���k��{rz{<D����AX��)cUy��rnc)��0��>Q��pc����x�����reY�u���T�Vl��D-�
-�G��&��6��n�/^��>5� 1<ڡ��'?�)���hݾ���?��Ly:��j�ā1YM�{x�;��C������E�9�k�-�5B6�N=BF��Z9�>���/j�լ՜k.y�|.	3�U�����L�r�W~�1�T�u�*��('��^�&,:O��"�]������v)�\M �J5.�E�f��?/�ʲ���a�9g-��>�Mr��N����|�}��]�z��;�&�y�>Psp6b%�٤�C�c���9R����v�v�<���H{}4軩q(�q�Xr��&�}q�g94��0@y1xGq��Ҭa?R"R����u�tǞ�[��Z�,k@������wn�J��ήJ��3��4a
�	�ş�Ǵo��0����1�6��o��ф&t{h�nТKV:-��p"�p��������7��??@0q�A��Ƭ$�3�;"�Y���
yaU�*�O�BQ�V�\���/���r�����E\{��ռ�z�Q0��*+<�V���˒1�t_���f	��m7�:FI��fD���n��[��h}��������<�F���#�AHָ�h@V:Y�~���?D��ŀns>�^�,X���cE���me���|S�R��Zͦ����
���u-W�5���9�*�NX�[��d�����Z(\ݲf1��M�`a#&���Opn�h����o"  OFCD]Z�6��cZ�6�����~�9��+��9��	Y/�%Kg�J�eu�K���9!�Q6t�\�Y��ϖ���=]i:�Y�3q�
�U���<O�w�/sd�a-\�|z)P��̗f�/y��~YY����'<�O�Z�� �w^��}U���&}�'���h������w<�~�	_Y�ON09:@r~
E���tv�x����S�*����Rݫ�ӿj������Xh7[2��`���h��W��$�,�s�,J+[Y��Ł%�CS�Z%˘� v�Y�$.Ƚ'|��u��𼃃�[�	n��tz�#�xv�r�	��	�_{�%�c:ѣ�~)T�7�4YKnH��;چ�]�f$F]���;d�X�Ly������%�Y�DH?��%_��O�k>v>=ǳ]�9Vzf�򫒥�t���\�6��}z��z;_zo���d��`����"�z]أ u:�k$�3l�9�d�=x�I����'ڰ��Ue��������`n���iy%s�����Ro�x;i��6��k"W����Z����T:%ۣT�m��L���l��5�,i�H�&��# N��I*B��!N=���}شp�����e�u��!P'˥ըc�w��wk.������`���.�A�2�0%�4i���]����N�oUf{��z���W��i����Y��g�%K�Z�Y���q�����R���\�0�$���O� {d�������;��1�	�5)��@�?Vp���Bxz�����ǈ�O�T'0���A)U-Efi����]�_dn{eXmkѼ�Iiev��pl�a�^��reYO��-�Z*�J��$yM 7�Z����s�.�I��F�x�$���'$1d��"���������`{6���m�ul�k�j0����_��/�����8�������E^�\�g�,�<Ikh,=f��y��J�S cZ�r_e�/��9f�+�W��iX���}
�y�<'���^��7_�[���o��(�H��d4ƨ{��?��d�{�Ft6D|z����brx�6�ǧm5:u���q)3Sm���9���Ee^ 	e�rk��8�3��u��яB��f���e-�!k@��Bk����X9�+;�mZ�"n�`m����������-��,ZH�c� F@��u%Q��&�m�?r�`2�n��K?�&�4�����?A#M�	jed'JX����j\I��Z�IMew�����k\��*�{&���k��[�E(yU0����x	r���gY0�A���g�UJ+��x�q����/�?�Cl}��$FY�a�t�0OB����o=
�#%�\Ӽ��gC�l��c�#+kd���-�|[NrS���C!�)o�ʻ%)l�=w����k+G9�B��\Yր~���4���ylY*慥�r�3ڗ������l��q���T�B�����X�5�"W;�d5�����6j^#'��S��N���� ��U���_���1�닕_��0٢ȶ�҆ܦ�:(���������A99lI-�E�����5������@u$�q�Wƣ�l������Y�f/?;��2SKfK��yZ|ncG� �KٗVv���0Ɯ�F�#��)M���.��g�5���&��E<Ow�?=�&�6! ;]���8�PУ��I��$fBC�q�4Ѐ�-ӷ<ʋ����+�����,͟I�w��s��'������m[W��ֲ��ڋ�aE!'��̇I*���J�rL-�܂+35$�\#�M[HW��gP5�_��f/�����R��5߂��$K���8$������=�����_��ɒ��x�
#��6[s�|B@oɢk�8m�G����1#́C�P]4~a�����*�EV� �4(��}^rV0�6�Q�8�:���g�]ESV(f?��p/����S�$�@�}ʧʈ*'Qd�T�a:^�)?m�3U/L���##�prXjɳ�#���W�
�	&T���fF+߶�m��Oi,�������O��*"���q�E|�%�|���uQ�F+x�&��_���C��`��U�RLiL��@�Q�c]��$�5UҦɢ��6MUY�伂D�������/��I�9~����v���ʲ�k.�h�"ZT��"�Ԡs�NN��u�r(�X�ڴ9�WY�ac��k�1Y�z8"눖��SZi�܂ϱJ�%ŢF��B�M����ş޺�O��o����p��#R��E�wKq�3-��N�&��*�B.��U�s��b�|��(Qo��+ƳЫPv��P.#S���g�1O�
	�.A����gI������ơy�sD@2�SE�=�[�ܳ��pDstLvi>�[>j���w���Ko��XC��"���=ă���S�6�I'�&����	N���z��t�Z��	)������\\A�q���Y�i�l��J����_�v	w'��X���F���Iza-k������+MTRc|�)V��YW$_����3�0���{7I�'HIy>}
V"�2獜���&�G�p'�ȵP{������}����;�Ǵ0�7c���R�W̠��3oF�)Q>^�'���"�x�p^N�օ�Ȥ�e��z岺Uy�}�oe���5)�M������g,
�	��,$9�{��w����b0+.�s0\�j�Њ�k�H��^��?n�#�,��>4���f���N&�>=�@FH�=�j<W�������!Ϳ���J�.�'��«S�m��,<!	�T���M��'�� QI�q����«�c�6�d���Я��l*H:KάƢ�qO5ku�������U@�dNI�t��	/�8�1��@�g9G\���C�]L��`L`�Q���7����������8��/�OJ��	�}m��R+��V�;4�Q,��gc߫�}>-`ͥڄ��a��j�����}^�Eu��}f�Ԕ�<� OeC��,�aʻok+/�@�cy_#E.I�/S�dIK]�`;Y6�t��������0$�|8# 0����[��J�|��<y�:�K���"<?��v����%]	`����&D��
�zlf�kg�#<L�S(�q�Lߧ�CA�������:]S������Yր~�%N]�Ô��l1����^��s'k�s�����0��u�$1*NФ�;��B�?�aw��/�k�G�T�F�G�\-"K������yi_ڬ�ɭ�����|D��+�P���Ħ���o�na�H������jҗ��U9�/,�[b�粬�|��t�+�,�Wg��y�\�oy��7���X�g�qb���vB;��B�˯��o|o����_���1H@H|<N0��E	�z	���v���РstO��1[d�m)[�2�<�<k���3�%T�f�D�g������x����2������~��Ȣ߄���劲��.��:�m;��9�<����&i�*ӅŲ��2�(�W��/!���L9��0�U������6Y)�d÷mD�{m����Z��1Z���]ܾ�2~��K|4�k�����c�&�n�J֐�y���ŘL�ׂ�&�=g�yU��l_�t���"�Q�Ώ�?���g����	�K)\��柦%��L�"^��j�$ũ�N2����G��]8/��[��C����I�sq~r����a��y��4�q���	�y{nM��'<�,w7i����G~���������]�>s���9{��2;V����3�^j�-?/�㒴���劲�k,���+�u�6֊�����]���ʸ"�J��1x:&^�$���v�}p�^�IguZ�'>�s��6s��,8�:F!�)�n���/����_����)Q@�9mn����l噬伝fd���=^:Sg=��;�2��n��X�J��S����e��3�X`y���-<_)��,lw9�NΩ�����Mv\�}๹��v
 H�M�����%K
I3�Є>��|���?��i;��r��P�V��v��n� ���%��;�{o��$D�:�n�m�ܼ�ug?�^l��`��N���|�~AmGϸzJ/�c�Q�*��{߀�����������@ƏQ?�|�B:�C�'�S��<$�(�`����]��l�Op||ľ�a��Z#�f�PK'�K�Z��5�|�f�ϲ6��R锽J�{cɼQ�}eF-᛾K�D��hI?���q	��hx��G��npٯ���ͭ很�?�HF�5Y�t����ŭP���l�ISt�
�ɣ�&x}VWW��kx:�����>�pAIc+B�>.�e���o��
?���Y� Mj��Pexe�L�:0�l�SIA��/��G����vJ�S�g�ٝ)�t�Zw���y����]/ʡ~�_�K�j(��pk$�f�=�x���mx�O����+'-�
����!�U���#�C9����}��}�����Ǐ@yx���t���A��j��`<��o����*Z!�#�-~�';׵�$Nص�m�a�Y5�V��p�
�'Aq���$t!�.��j��T�CW�0���"=�Ԙ���u)Ci��ҭ��Z�E[���F�T�}�)�]+�QE��
��S"���Z�
a���%~x�8��o�	C2���VFp�&�]y0������	��?�>��� �H�:��ב�E�n
�!L�Tm���jcm��y������"�i�ٔ�Zm�[�v������KqciΏpc��V{{����p���:@J4��?�ؼ�5K�N��6�R���Ai%-��~��q/��p ��o������я@�M���ti�s=���!���#:�ln�̎��98�=���FM>J2ȑ�|�"g�)���1%���oʂ�����y��Wz�i��`�ӷ�-�kMʊ ��#��
/Q@h���(C���W��A xI\ABt�TMVS�M�!�¬�r���r��xz����>�)�Թ�ws�%P�Ն<�<I�x\�aT� y����xm��>Tx�hgw`�G߇���0ؾ��K���3�x��p�qm��"\b��}�|�|H+.��5��:�}�I��m.�y�����/���.�]ԏ\A۟^�8
�� ��x���7�P���'
���f����(���~~�W	�;w���i�z����>����1�ټk~�B��{0�c�Y[�������Ĥ���\>�tt��	��	Xpv^O\�r�%��Y���(��g��,4(����F3���c8l^Ad��J@��5�v1q�ċ��y�C)I�%�]�\~d���_E�`�ͪ��P���1��a�u̺�w���o߁k�oA��@2�qu\�܄���xn�{��_�W����	�������AX �%���B�����U��a[���[�rǧ�2x�b2�}��ǟZ�8�o�^�rf���>an�M�0G�E@���~�<�)��Y��&�"P~��������������>x7�a��CVS���;�eI��>�Yc<F�0���ل��!�c3��ѳ����G���[h���j��89{g�M��u�-T���t�������Gi��,>w��4����^B�W{�=Ϛ[M\��$p: ���Z�^��I���'R}HS0F�+l%.�А�Q��\�߇0EB8��c��ևC���E0�a��A��!��C��xj$��_�vg	���.�+H,���d_{��]k�'W���/�"1ϋ�8ݍ��c��?S����>����~�8<+Q\��o�������4 P�M?�(�fApCJE{�rx�6@χ�q2oLjcR@9�As<�g�܃�n܂�$O�����p}8F�-�Ç{p���P@H��P��,h�
N����i6p������g8��w&�v����h�'渶���1�ُ��)��A���Y�@�Ԅ.�m/����Z-�ާ���,P����v1;c�7/\�M��4�<�*����'$��#GC�6���|km���<����X����戽��@��5��W@��������>
�����Ƀ'�w4��0���ꍍ�Sg-�I΍������N-Ξ���<]��pq���izN��D�"��ٶ�A�]�ygrU�.G�S=z�����6��g߀J��>LP�N��"���R���7�������~��&�O�؏�!��u*<��l{��[ׯ��hz(�����������S�v�ԻO���X��������W&I�ϣyY$Yv�����ߢ��y�;�}׷��q��٩������G�h凑�������Y��&t!�E��uέ�����B����w���iBp��g9�m��~V�\��� )Z\��&���#�Fk����߇[���&��׸XOp�&b2�_ۂ�C�'��+���-����p����ݿ�����=x�ڇk����%K��Q��Tu��E��������m����yl�x��;�UU��,p��n��@C�qm�y]AIy㡆#�"�4ԛ���w����?���)���)��1J9Oa\�p��=������:�Q@8��  	}XR��<A�|����a�M=���S���(��q{��v4��~�^?�jr���9�ٿ��Z�)��)' �%�1�>�UU�y�Js���ydN�Ԅ.xyD*�Ukn_�ܭK��\���b�Z��u��aaU��i�A�5�k���O�1�ԫ�cH�d�w�h��7���u8�*���'�o������!�8�jy5�ó,E�݇�q��o߼��n���o��׿��0�Aq+W��������0�����͞(��<�w{����nP/���ӟ�ƙ�ϻ��/N��������9��.����{�m�������[ ۨ����%s��B�- Os&sHJHPpS�n�+�F����f6�hN�C���%S�	�7�Դq���¤�S����Ցg�x{����wy� ��{�㌦����4�I�<Aϱ"(�����%A�7Ey�`�q��)xq\B����<(O��U>���&Lm�������§L����(�Xw;[����@$�&HN�2�LT&�rx���y����ߠz}����@L��pa��)���Q���!Mr(���I�V=���M��7����~ ���.�g��ZWCzxn����a+�R���V���3c����`/��k�8�*p�,���s~9_�_�K/�"����3��E���:��˄����B�s9�mfx_�)���6���o���\��|L��$U��}�>�|��>K��H�A����MP�5��{M2����d
O?ey\�+R����F���ŧ}&n���҇��]�h�G�R߸�C����Z�]�;��ɾ��<��Q:%�������|�������'��H��m��ey��s�M.qcVi��KR���5��$c�����m3��זLv�o���~��}o�Pڿ��yTx��EЇ�|U�³���Ĩ��ą1�ϡ��̐���ېQ���>+#�%��#&ރ����2�͟����7a��1<�͇�O�x�t�����5�|�G�����nPb���,̱C��FJ5��>���Q�!kdUS�
��e[�ۮY�9rsi̵zQ��3�n���h��pB�3�t,�ɉtB��?��@�K��⡴*�w��G)_A�����8��l��-%D%�ȩ�@Z����1^�n���o����Oa���Q�}�;<Q�L�HԬQ �+��U���S�3_c�V����H����{=�̄'�n̧��)7u	����!����=m��i�⠜�B���~t�Ns+(ٞ����r>�= K �y6��T�s7�<=�t���3YHi������Ë���r�#� iգ�S�d*1�j\�7�s�E̙�5ԭY������O�=m����G��C8�\�(`��c��}��q��>L�a��M��p*��x���#�!9� �!���P�2��#�U�F#67`��[���o��7߃�����d=��!�C�`�(ac�g2��)��2����i�Z��B�s�����U<�q+��G�y�Q�ۺ��8�� -8) 9!�i����	"vVؠԢ5��z��n�|�B��DeH��7lm�g�/I�B��e���"+a�G�̐ďi�� ��u�v���ß�*�mĐQ7=�֥�H��#��BC>�@UD��k�Ϗ�53xce�����O�@M|���,��`R���}�;z��g	���m�>�6p���P;���)ܽЋ����v7���C*�LgVPF�Z:RzA�ه��X�~,�.xi|A��eT��R��'�>�A/��p�Q��Z�"x�c~�W7*�� [w�ɃȁRy���-�2�"��vr�2I���#(f	D�1����z��c�=����#�=<���$�L�Ĩɯ���ECt�l#�o��{�濽����_�
>z�Ƹ��xi�m\ǔ�NdF�Ҳ� ��f�0�pq�)��TR)�#lM��Z�@���G��y�����m��U�M�6�^�:�L�~aK�m�rFaClMm��Tl������9�#�����>�� -�4��y���nl���������[7�	��lnL˨�j$l%ju:���6x���b�C�����`H>�	?����d�Z��<�z��4�}ػ�F����on������w���H�t1&�Y���85P*,��:��$�]�����.d�,(�Z��8}��-1/��b�*�]��T�@j�ݴQ�`�K2��,���AG�M�/�D[�17�8��P/ae]��[�<a|P����&$�����_��ݏ9yz<c_��*^jI�A`݇xc�y�-����������.���(0��L�
�V$7$��kX��v�;�X.#ϗ�CrԵnC�֪a��U�睚]����ܝc�ˑ��_y&��}o�o�M�:ف�\�Oy����g��?�8>��9*�����ŕH���� �6���߄�;п���� \[G<��'O؍Sf9�dN�y�x�b�H�g�_o�D��h����P�p��Y
(��t:���=�B��#�p�����@�����)��4�Q��`���>O��+w|:������bSȧN���LWy��#^����dGڧ
^W#(Np!T��TP{���s���fZ���-������T�Lm��V�p5�Ћ���y|�X3D�$S-��<����%�H���k0������VQ��F��	���7����S}\*�Qϐ`zQ̑�����_�%\�������8��S ���>���¶�(�19ȂQhm<<v�oJ�j6e�p?�c�]]'��&ɽ���H�`��[_La�!������b�����ō�ֳ)Σ)c�4�^ 
�b �r$c|���Y�9������#x���!����N=�{B�n��c�X/�(�Ux�9�7��S"�C�A��t-$�<#��A?�q�C�Q`7a���C����#[�/$׆6�\u'X�<|���9g�yj{��R'l�R���@D��a��FH��܃4B�4�Я8���{A�>t��[��rq���<]�k��j�`���2MR}�݁��KDy��IKg�U���5G�s�u2��/0��'e
e�cCV��=�T�x�o܀������g��9j�נ��p���w�a��Yc�%�T�	������א�8"��!|����>z�c	 � &��(�z�H�H�9j���泮�Iqnnl�T7�bh�K���N��;��ħ۬SioAX���5���5��u��Ĉ��#�?���S��d|����Аb�7!\B��
7o���}��CM|�ȇ�7C��p+�Z�$<���j�{4�{���=A��O.<�����f������e����74����5��. ��:�����}��i��6>-MO�c:#�|~���m[ÓZ��6͏�����; ��5���<pG%/	!�+M�'������	�h�Н�g�caR�ڈ�'J4G�K�0)h���F�kknN�ٻp���F���z��vPjYD��r���N��P�]?�2O�B������]8�Ϡ���5H�p�q��X���5��.��#�&��c6�HN��Mx�/�6��&�=��� ��G���gGOQ��j��N����5�������*C�d��T���97&xΙ�ug2��6�"��F���(�kRɌ����h�w�k*�(y���ܒ`��D�Y������7߁��� ����������s�7%�$l/]j(p�懨�OS�c�W�#)H�D^T�5�e���z���ޫ8��G�� ���}�y
�D�x�?X&;"P.��HI�yϐ�X�9��آ24�y�bBf�;%N�1�g��ٌ>Sy[*ៈ���Я2~��.u�e�Z�m�[s������5�E������{�ҙ�;�ޖ���46�}W��i8��SSS>Sq$�0T�肴CU�0��H�%����ߺæ��O�C�����w`4�AZ���w�x7Q�`>7�P[T1�9�������Y�T��?��j#s7ՒGM���_��w�>��.lc���g��i�t�[=<���4P�@`-!>���Av<������T�S��E-zm�s�k��Onw�v+ka����R�����η�k�[��X�9T�ٹ�����}5�-$𞽷$x��4C���2�d6��
�8N�IJ&q�� 
J������c�)����c������<Ծ����Brt:���R���Q�O�<ն%���N1�@]��F�tqݱ{8(�Eq��
��s56"���t���F(� !׷�rݹ���qԗ��W�S�K!����]�.˸*�0
B^d�B�:�g��kc�]��t��O�ӹ�q�|�I�����7J;2�f������Nj^.�����F���|�ǩ���_���>�E�5��6�8�	 j~1j�[H��H�!�oyp=$2�WE�H�H�]�吣XR�yzuh�kH4@�q���!���7���]��1���s��C�Og���(�:,+��v����#*�n}S����9Ӡ�����&J��LN�}����
$�X�=�Rw�$�3!a�XkҴq��$@-�,T���CH��x~�g7~�S�*��F��w{H��%�<IٽA�e�L9�mzt ���0�#�q��Y�������&̈����i�ͪC�d����=������&<�<$���t@m eY�JeU�p�}F���=���s�0����Ӎv[�-��R.Ƥ�7`�ۺ-�&8Q��DGऋ{(����Hq�<W�H��W�e$s��U�x��PǪi<Ze�����n��w����Am����6\|�6�������}�\�6*���} 8���׬�R�k$i<~���?�6wv`��mX��=$$������[[p�Z�����JX���$xxxE/���)CG��ɳ^�ZVaJvHd�+�0��;��o�?Y���7�n���#��!��������{�ݯ~$���5� �k�HF�g
��O������;#���I�b���'Ԉ$
95��>lݾ�j����C�e��M(=�C�f@��t�߇"�`�d��H�6��P��%
 ��t��K*͚@I>�y�c%2
<ShX�x��*'6�I���~r�����=�t� 6�7AMSػ�!|ԲǊ�|n��)E�1�ө�<ք���eo�j�6�����0.e�u+�,�_~����<	.d"���q�T�/kX�+!�+\<G꺣� K�l�Eˍf*����醶�LU���5���P7��7��[��j�`�ˬ��b�ҸO���ӡ���XG��F|��g��<�9u��4O$� �|g0�)����P�S$���5����j���1Z�I�Q�I��qA~z��F#&0
�K�v�:b��Ք����x�o}�=�����G-}���3$�9�~�$����;=:����#�������@�`�7�6�?q�1Í�^�vm���g0@A���>�K�P�ChK���C|)P�&wH��6��q]�ʴ.��O�vS$�t>�	���r��	��l���u8:�C>�`=���
�������=��3���0q�1D��l�'����J9�'{�k*� ��ƈBD`c*�=�u-?D���pes���fX���:�y�7���c�\�Bd'�>�&��nIݳ��Uq0d�h~dj��������SEh���U��j�a��^M$�ҧ��wa��)�6��lh�M�J?f�kV�����p��T~~�˕[HO9�N�Ր�Gu� P՝WTGx���q�}$�\[oށU�k$��>E����_��V����#	�����G0@�^[[��W��0���B�D�b|"��S�XƚvX�LR�;������n���Q���j��bH�Dlx*M�ߕ&����Lb,Q�
�o�!������]lڢRv��,9�撈$�1��i���e�9	9���G%L��<�����6�֑�=h���*r���xm�	����AI-����G��$u:��ݧ,R>��4T.��F��R���.�e]��=V����뫆��s��/�cQ�ڙ��{#Jh+p�&0&6ĝ��s�F�wu	d��b;
�6�5�#^B�WǓ�C�5Ǖ��c�~^[��65�6�s��6��B������+T��|����������EQV+�������ߨι����&���7������Α������O����T�x ���n�@�Z��x[�>x��79�2)!~?@��ߑhJ�I#yN�k�ހ���EX��fL$S$����<]��Ɍs�)��Ė!5�	��7M`)$��5�^�7n�|��ܐ��|8V�]c�M�~�m�BJ�ߗ����]�p"�IDq�|���O�BdO�z��'R�Bn�x���	[޹qn��{�!n­�<��@ȵ^�xR�<w܃��3��B�7��q�?9�K@�|¬�~F�:	��p�� �2.BӉ�'�vX[r=��v�o��V��g]�W7N�M�,�s:�=da�q����$��Z�|��/!����D�u�Ђ�Ѽ����N����i͹Y��r-l�xIl?M�bJU��X��Js���}[	̜͖]�(���-�B��u��Ll@i��H��5���O�Aoc����k�=T����>B�v�IC$9a5_��0�Ι,G��"����:�ῊSݸO8��{���'?�2>q��ɜ,���6����`���t3�2� 8�J��vR�8p�b�)�=��c&B�<pnD��j�S::v]U���&{��EAvy���5u���?�!�/�����Ts�39��2�����FM^5G(��0�J�kS���3��>����5��>������H�=�;�~�dj71>;x����L1�s�e��v�?�t��{2n����H���~:��	�
�;.���~(+z��k�ɢ�/�8:?\_ x�_e��Ȉ
�jmڦ�-��sV=�ƭ��2�+�#BM�h�^Ú2k�I=�ش+����z.�S*X���\�7K����G�����4n����(⼜��of��$��V������1j�oĥb=��mG��k�SG0*oZ#A�*۞�7������"��{1�=#fS$?�<��2�)��%x�5sN9/&x�$hm��\#�@��K$[�S!��EV�F�5s#d�XS$kAQ��wPۻ���+��{hp�����[o��N�S�ڸ0;��|�=�oI�В��C�Fl���Ԙ��T��G�"��?*\W��mV�V��E�&��<~u箟~;e�Ԃp]D�I�$�S�䉪o��o]?:�'�X�j�]���%v�Hc-�l�?���I��2��%!�~���ڧ�k/���'iMaH�~gB��Yli2c�v�@��4�.���;xߘkm�����7�)�еiFz���t�6(��{�����ک]EI�=߄�ض�$e�Җ��5��q��!i�B���G��am�:l�y�t~܇���7�P@IQ{�)Ç��k"Ւk�S
�I)C�8
8g����#��H�!'�C5Kx<a3���Y�y4��xh~H��B��Z���[5�4)dL6��R��=�(%i�df��(Ӌ��i��ɗ�K]G@��H�e^�]�?g0\]���*̏Q#���CT���ӏ����w09��3�*�x���(�<s�j
H}k*��,�X��g����AQ�_�U��wgB#�w�GΥ�g�@ �l�\Кy�]�<��l/tWC�k5m�2u+жܱ+����\�r���)����P���}
�� X��-ik����UF��iT�k�*J��s�7�E��+.��,��rWRT:-Jv�l��Zx%]�L�boL�{���}�=�箴>C��{`7������0y;sg[��e�kVc��-���6l���z��'>F��!�HbG�ރ5�g>��*�����[o�pk6�#�n�!EB�@�OP��|{�������ĉ�����3a�xJ�SL�V����p{J����"������x2�2V��?�7��5����Þ��scs�>~�(��x40�P��맂���ñ������1T8������c����������3nk���m�5�+���)�! !JQW��fm\�֯$D�o�Ę�˧�P��@c�[W+�}��9�m�:m�͙�I�2(`���/���^�����K����c،������p�0��.�/N�0�_��EAN7�
���a?h��������UF��h�Q/h���5i$���ŗV�Ǚ�����Lu�@;���u�~v�z�$�����K��5�s�[������nK��cوo�d���tަ{|�TU��I�cE��,L�T��,��?|Џ`��MH���/���a��-�A���;�Gy�3>�qj��B����BЋ��X�7	(<Pl�5sr�S4�!������BU��t��y'�:P��<�}&|� ǥd���b$���Yr,+�����/��؏#ȩ
^؇���f^7%�WoW"��V���'p�w���G�A��R8�l����Dd�ݞ)իG~W�#^��v��U����;�~�U/�aؠ@v1hSΖ���i��i��	��ow�^���Bm�{�LO{Ϛ���όl�'m}���P�Ը�[����-TP���Z_���G)2z^��@� �~�ᣆxd�-X�	P�T������E[i��I�T}�49�Mm`�2.��vp�{���#a��kFm�n�o7莅�jP�j- m��r�l&����on�k4
/�5�QLbE���G���)|����[[p�֛�y}��c�^�(��h��F�I�N���L�Ԇ���.��HZsV���B�FOZ}T���i�H3&c"t2�sD�1s�V��f����x`�۪���,Aoh��P��6�y����t=K�������O0y�ǩs����Գd�Zz�=�{x�
�C�oȒ��Cek�kK��)y�u�T[|���[�!Ι�PȤh�;�K@!�ֺM]4���a��V�W�����ӻ�a��sß�(�A�S��X؊��RԸx�<�˧D�"S�O�5���QXD�YSkZ��e!�~��:�}\�G�A�D�L*$��t�9�����`�[f�9��놚�B���"Uk���:Mi듯O:-L����N<u�#��*h�=�p�E�[�(,ȼ0���ӛ������1׌Wl�Q�j`���,O��?�d|x8���}�pd��Q#�W �a8���ڑFH̫���э���#Q#��VF0^Y� ��a���=�جN!t9����\̹���qg4L�`F��ٗ^����]HH�Aa����t�Am��}>�A����v�������A]�8uL��;0B��0��Uq�R�GV�ʆryVxb���YM�kg�=��
u��(�A�;Su
���{����o}��责k}���Y�������VPT����6.���m��m*��=3v��p���@x��H���8�/!����!����J@��IVs�6B)��Ɇ�-Ⱦ��f#�y���&m{hCܶ쥱ܷ�7�:���
��tK �9UC~�������gf��h-������\ ���6��L�d��jֶ�hˊo4mҔ��J׈ȨX�B}��'.�M�T�Hm6گ�����Qx<�k�W�wn��;߀���I��2��M�@ +( �qr*~��?��ȼ>@A���O>�_8�,KM:�r)�4�l�s�ҸW�T7��M�SC�f%5�|wcgS4~���.��4'�؜ ��Ŝ�ڱtwoG�\N�E�;��6�rY���#6��խ�x�%G�߫�	���x���C������8,�kC��Ap�9l�?�G���Y~@-��mCV�a�M��G�z;f�f4e
a��� �%]��B��h����[;���$OҌk����.H��B6C�� ��?A7�����.�����ۖ������\�]K�v�.Q8߷1�/�I3o�k�J�;q&>Y��ɖ���J\3�qD�=���W9��"(5�h�����V�sJ�k�z���K����9�I�2(�����ݻ�A�oyr�IE�A��M��0@~��� ��[$���I"�UlYYP6�����N�D<$�|�c���7��
{�+u�L!.������8��WYБ����N*�@*�m�b�[��Ud�V���X�xcӹK�N��c&`rS(sv�ݫ� �B�$|j��ӫ��u'�[4
����y�O�o�o�M��	r(�f���H��5��<G@��iL*[2�P0� �t0HP��!�~���M�?����w�U���GO�88Dr�%��a8����]�K�g�������h�.��5����ƒ�vz�Ҷ��´~���5p0�U�iQg��r���a�2��1�n��Ӽ}C���\��H�r�)J�*�qmn"�T�b-����|;N�Ã�T����xW���p`\��o��Yn��(�|��wF���O�h�u�n|CMb,+	y��Y��q�O�\�|u�#I��CN����hݔ�^4%8	<w�îۂ@�U�L���0dn�&p��B��fS)޷q�긊-<NЃ�e��a7�^p��{K�V�Y�0�.���>���R�ๅ`���6+�+vO�L���x,L��Z��O�"��r�b4�]��;�-�V�5����E���1���$t�"Տz>�{^�"���A�
�i�ͣ�����l��]P۫��_���gP�Sn�Y�E��9����}Ҩ(ȧ%teH��ږ1�{&��ㆵ1��{(n��E@P��I�;/2�.߽[{��0��l���������o������#��6�V������
��:p�r��iu@�<c�ڷ�S�o�P!�Ǝ�UH��m��*�kQ�8o��$�Uc4���Y�I�q�#
(�����L�u*�!G��#��[����6Hir�k��pp�ZP=��G�q_�sU�C-����tv�0b,���K�7>��@��y3�#G�+�Z1�^D-p���:8��Xl\D�ب�ƴ���+w���m���N)g��n�b�gWg��/��ָ��c�y}�\�@s>�Z���<��@ik8�i�!0�X�`m 	]��lb�:��/ !�+
\h�'���o�*[��{0���{H�H�-&�j�@�d�&I��������9��B품���h�E;�(�����ޓMՔ��\�ң��,���>��	/z\��^*�J�%�3)�-m/�Ɣ.m��^50�q��ʺ����m�(��7np�UF���9��Щj��$�E�,��ua�6��`eY�B��(����͆�HС�Q�+��5�=i�&�ʐ����t4*Ɋ���1LWs!��~��N`�L��:���D��.G�%��z��gnk��+����n�B*h�c�k�&-8F:_�f�'S<I%4�!���:�<^�=�{Ay����T,�{B����ҫ+�C����7-s��G0��8���{0Ox|�`��2�����j�U�"��/������Rh�;	���wO\-{���%�S:��^��\'����S���OB=K����G]Br4ᒼ�;��{\uO����1�x��4Rg<<nN��)G�0��f8'y�<�Φ��%�	_KN�"�>
W�iV�J���J&0�{77PԬI�5E$�~��E �����I�"�s�2���f��79�Z����H�Ts=���M&䲨9]�-�\�	�
��k�7��g�;��>-�d}����iǜ�E�Pe5O����*^o�����H�C2mp��(e�$����`��ڢF�WY�d\[2&��+�B�M��4���������QP�H��3�o�壃c���>"�	����G�Ӏ��D=N����4�S���6�q���dQ����l����)��q�+���F���
]�Ə�=���5���cՃ���P"CaI#1rM6�=�a�2+8���Y��W�yuu�Y[[���.�7�xC�V�~Qzr<�D:�i�$MqT�J'	$��FS���EM�cHn���L7���}�(����P׸s]5�󕊣��p�z�#Uu�D�٢µ�&/2ܧ!���B�}��9UN�#��_�2ӟ��g�]�4�(�(��|��f6=n�$�!���P3��l�*���H�~ߏ�}?��t@���4�I^��Ey����/�[G�@�B�Y,9�˽���P���Џ6��R3]���:�Co��n|$/I2Tv=\NU��<\a�t
����#dY42>�`���M��I��X��Ҭ=ք�Q���y��,�5�W�è��X�ȸ~h2[;-�H���ʪN_����t�ڏU��\t�V*��@���J�~_*T^��eI�+sE�γ,ъ@��j*��V�(oຎ�\Pj.�5�ZպOF�)�3�r i�u��C7~�ZyD�ʶEcG���{�7z��p|��ʢ(Tq�#�m�Ԛg>ՕN�d�T�y� rȵ�u�:`��b��7���<���7�n��V� ��Vê�D@8�uC�{j��� ~Dz�4u9�P�OUK�B�ú�(���#"-/h"��}W��$��,Mص��UeU�Mh�Q ��AՋ��_�=����C6N�S��w�^�����i2G���C��I��X�I��p�(����^����D~Lfo��*G�QQMSБ��q��!����&M�p~Q��J�PƧ�	�
���p�M��~J�w�ԯ����(�J�5E��췩�1�a��D�,.A��yZ�(����=��i��J�Z�Aì8dE]M�"�ZGeD���7B)#F���2?�;�>Vkk���������Y,9����������_��Y5��{�~8F��MXϓ�tr�v|4���8jX�SȚ�Yey�#�A��t5;?,��K"��(Α�zOvGH��v�j�d�����n	��E�Aő��T����r���IڛeT?~�ٰ(Ҳ��qI� ���k�����k[�]�5�y�Յ��+C.�Ud9kq�oQUȷ��zMyQU"\��<{!~�������Ll]/ �FS�$KU䅟�EP0�㐃����
����)(��VA���JFM�J't��)´7�㵭���C!�����\����B�E�	����%r�_����o�>�Q��A�����]�r�Ϊ������̑eP�5�c���Ĩ�#y#������<͐�( ��rB���\Ÿ�,�ט��p1���*�~s���W��u�ϷR�-�9�TP%(tUxHص��&������g�g���Vr�]����Rt�eP+�W��xh����1�5�AppM��:
A�)�!*=j�@v�8�t����HX�1㾩=��}�f�~J�W��-�C��(x4(����`^OtB�P�(x���y������V0�o_��콿���N	_B�W��-"���	���"t��U��>LF����[��.HG�2�~�*�C e���5M[o��աw�����v��֣�V3
F����OM��y��(�c'E���mB!�a���9�'�My��'f�����u�1���9�J���A��8�2kt����.������?�Ǭ���� V��H��}�o��N��[����~�1j����S�z������v���+�W�Я�W��_�R.��/�	���)�@p�!�夾廢��j]�@ \e<�Ѕ��)�	��ĕ3�2���@ K !t�@ � B��@ ,���@ X0�K��@ �W��Я�u
�/ i�!X
\�'�k0�_QI X�>���>�]n�@ ,dE} Aq�@$N�@ \6��!s��)�ς�����@��A�)�� %g!�. �u��d,,?�� d.,?�̗B��@ ,���@ X��+�-�B���JC�\�,B�`	 ��c���7"�@�L�5f!���c���H ,d�YF��B4�@p�p)	]�Z�Wy���¥$���Ԋ���AR����R�U���W!s�@�lB�`	 �.��w�@ xQ�>W���u]���l�@�RB|&��7+��K!t��+��e�W!t��+��́@�� �.Wb,Yz��U����C] �%��@ K !t�@ � B����D:	!t��RC�\ ��@�B���8=�����% d.x] �.�@] �%��@ �Zk��m��3�A�k�r>V�@���ɜ�����׌�|��@�!�.�@]p�!>�@ `�.7��_o��%�2���B��+��kQn^2��*���[��Ȉ/��~��W	���/�R}�F,^).��"x�pI	] �˼2�4^B���9�.���@ X��@�B�`	 �.�@] ^$_@�UC�
C���A��_5�Я0d����k
ў�@�"BM!d.���@ K !t�@ ,!���R���=^�@�u�ꭶKE�Zk�xm��k;0�@ \z,���d.�W�׊�_w[ ������@���Z�Ձ��	�����'�Kɍ�n��@ x�q�	]�Q ��@ K !t�@ � B�WII|y\�p�@�� �.x%2?��g�@�@�<|�.Z������.O�@ �r���˚P����k�4}�ˌ���/��~�/�4	�e�kL�_ ��&���r���@ �(�������4
_����
!�/"$]M���A��jB] �%��@ K !t�@ � /O��-g!k����	]X�@�;�
�+�����a0����@ K !t�@ � B��@ ,^��%F ��/E�B��@ ���@ K !���\Hg/�����WY�^k����B�\ x=���n�\j�    IEND�B`�PK
     ��ZVX��<,  <,  /   images/6bfc6843-1883-4a57-a768-11efac5c5eb3.png�PNG

   IHDR  �  |   u:�,   gAMA  ���a   	pHYs  �  ��+   %tEXtdate:create 2024-06-16T02:31:32+00:00���   %tEXtdate:modify 2024-06-16T02:31:32+00:00g�JD  +|IDATx���ܗ����W%�0��
3����m&��9+9ݑt*�rH��N��
!c�&9�6�2��A�f(�"R��}Ws���������u]���Q������������w}���]I�$%ʀ%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`)��I�j�Ky�;��f>G��a�R�-�ߌ�C��H�Tt,��8~M3�Ћa!d�A���2`)f����6WЇ۹�g�$�hXʎ:�`&KV��q��B�s"Q�^�.I*��c)oҏ���E��ڭ�����?
m��$IJ�KY�Е3��,��W>�>��Z���Rn�j^E����-K)�n�BF�?������F���$�.��NB�����=�r�чn������ ��J������&�)�$U�KY�c��p!=�U��o1��}5�|������C��j1`)��8S�]9#D���`�jV�͹�_���<�$IUf�R}�.µ9���ϥ<��kܶ!��65��;]\G�T5,e�+������1/z��B��Pn�#$I*�KY��J���4���r�0|%�M���0`)��e�Md��9����r�@��H,e�.f|b����=�nsIR���7�N,Zu�3n�4� I�j��EKY�άϏw3.�na(� I�*��M��Gsq�Y�!������$IZ	���C�aP�Xg�b���80�ٌ�|�$I_c�R���>�����J|�f�&�=1�8�}�$}�K��iAiCW�H|�oH�М�]��,�ŔКQZ��Ǯ��}6��\$I2`)Wfӛ~GZ%>v3�kna�CI�Ky3�Q��-�hG���^���CI�=��h	�Bۅδ�Q�W_b�CI�/���:q's6�I|����o$I�c�R���@s8�b��Ƕ`(I�e���M�КnW�wĊ��(�G��,i�it���2�CE��B&X0���0`I_xy�4��!���v:3ʂ�$e�K��bN�P��C�`(I�g���i�4-���E��aE����$e�KZ��t�rN�[$>�CI�4��:�q�e�Y��`(IYc���d�4?�[Z��9���L$Ia���<��q'>v���f2C���H�Rπ%�{������{��]���� IR����,b\hm��Ex�4_~��^@��Z,�*��VQ0��F��]q��i%)�XRU�`8��-JR���(n�p��;o�`(Iic������&%)}XR2*
�8�s�9�WGp=!I*y,)9��`8�K�����$�����U���Y0���2`I��2��[�� I*A,�X,JRn���(6����0�-JR�2`I�7{y��<�����
�3i�P�J�K�_��^⣷�,�~IR�3`I5��ît�`(I���%մ������%)�XRm��Q��`x	c�+H�j�K�=��8�(��-JR�1`I���î����
�ӹƂ�$�,�T��[0li�P�j�K*+
�e4M|�e��)�a��T|,��T�q\�
���VQ0�B$IEd��J�|F�te%)�XR)Zʤ�,JRJ��ҵ�`؍{Y��E��`(I�3`I����V��W�*�����ҷ�`ؒ.�D��G�(v���1$I�0`Ii1����Hõ�ehNI*I	1`IiRQ0C���Q'��W�a8���$U�KJ�%���F'6H|t�0����t����������0���\�H�
f��ҫ�����L���$Ā%�۲����Z��ac�8��!����H�"��,�Io���"_bths�$E0`IY1��������a<�$iXR��(v��K|��(m*���b$I�d���g&ݸ�c�A�"��_ho2�a�A��R,)��[0�}�����g�$}�Kʮe��ũ����h�4�2�ϐ$}�KʺE-�f,��E���Kʃ��]Y0����I,)?�]0<*4��Tɀ%�˲�����m�0zE�p72�7��3`I�3�r��`�)���݌b��S,)��(cJҵ�G1�����1`Iy���b�aXQ0��˸����$�Kʻw�q$�}zq�Sn�PR��$�(6���&>z]�i��&"I9`����,zs9�s6�-��r��`^A�2΀%��>bThm��E���~���},E�2ˀ%雦�֌2Nc��Ǯ����`$ׇ8'I�d���r��M_���W��[0�K�5����9,I��	�BkM7�+�O�&���,J� ��5�Fzщ�|+�g1�Q��$e�KR��З����S�ћ3���P��$e�KR�EL��`x,��1e�M��;�IJ5���T{r]آ���lF1��HRj�$�m2��)��"�ތ�e"W�/$)�X������2��(���Q�W�b1��2,I�1�N\��tf�"�^Q0|���=$)EX���r�ҵ(���Co��j��$��KR>���v�Nd��Go�Q�Mc(�I*y,I��'��IG��MFo�X�_�xI*i,I������ҍv�I|���E��1I*Y,I�[¤�ZҙSY7���^^0�x>F�J�KR�L�q,=hU��[s�r##xI*1,I�4�Q�)Z�pSzq.P�$$���$۲����JM����O��&"I%��%�f̤7�8���T��w�:2��yI�u,I5g~�2�QƑ�K|�Bx�����0K��Zd��T��V����6L|�����\� I�Ā%�6�Do�r4�sFo�.al��e$��$ՖOZ�rD~�_Y0��P�`(���$ծ)�mNg�q�c����fr=���TcX�j�[��?�Ѓ]�0���B&P��HR�0`I*�*���Ʊ�O|�Ɣq:3�;�I*2��R2���$��;��]��`��C��$�KR�y���p��oFߎ��[�sHR�����6��9�Qh��`��/b!�û�Ɍ��B|���ZSF&>�za�2�R�],&o��2쳛��6f,��¿�����Ϋ,AR�����6�s8HU��pȚ��<��sxH��it�b:r[a��B{���"��bO���_[��7Ƣ�=v:��o#�@,���A��:�ݩS����v`��&15D��К�wy��,��'os�Л��ϐEu�!�ȃ���έ�j��B[fv����sD����8�О#��n�GZ�2��\�f4fEXV0ܝN��:��� ����P&d�ը�!�_�4M`�f�%�%!���񼆤52`Ik҄����A��Z�9&��Cp��fO��Ջ����E�5c�(F�.i�S�c;�i£�e��.�/��V�*�Vπ%�N:�xը��д�������5��r�ю�E����U�ap�~؛:�c�n�kC���LE�*��UiC/���ڑA\���r�K�7��!��ʺ��ހ�B��8>!M6�K�I�׬Ǉ6����(��K��:!X]�^5������T�Q�M�f��Vy�a7�-�譹�K���Alʙ��I?�~����&�t��΀%}ݡ�S�wk��!��Q�qi�(Vۆ�ծ�M�B�����D)�0D��"�Iޮ��\��H���e[������u=o�%ʒ�)��T:<���]Y0|�����1��'1�o��ؙ�#��t��j�KZa-��2S
6e,����\�ͤ7Wp,݊r���!`]��,�)
Z2��(��P����H%��?װ�d�b}Y���cchKGR/��7��q?�%R0\�KB�,�����'�˟齅R�RzsJ��=�W�Cru���r4ϢX�
��qzh&>z]�E�et-�V��Δ��y�+��ϑr΀%m�x~D�jœ�O9*�K��r���ܮЊ!\�X�
��#�0AE2�ҋ=9�� �Kyw 7G.~[[��yk�d*�G�
�]9�?���va2Ck|�F�1O���3���B�KyV�K�0����}�X��T�)�mK�I6J|캕�J�`$ׇ8W3v�ZQ�����K�V�e�R~��u�BZ��T~���U�2���1����0z�� qk���x/�ccҡ}i�a�Y>[*�Ky�9�4iʟ8�?��Xĸ�ZӍ��s�	e�V��a���49��8��H9d�R>5�^�#m��n�`��it���\��9�g��g�\O}��`&ю��rǀ�<ڒ?�Cb������r�Ӝʛ�?�a8�n�f�m��v"�U/��r%���З����S�ћ3���P��踽�sNj1�Oy���ٷ�;�%�{lE��(�fa�mI��J�{���:R���?�?�<��p ��#LY��Y_��Z|�i���o��6U�"&�VQ0<�g�S�Tʹ3�����F���+���8����_���X�`�cx������f}�f�ZR�y�w
�f1O�68��ZsǱY��A�ˍ��*
�=9�.lQ���mv���s�9ҩ�����n�o!q�=�
�b٦�О���ݶۆw�!�I9b�R�4�v���/0������b��'?
���W�e������>T}o30��)��"�ތ�e"W�*��3���9��CH�C�8�V�odKNq��D���CP�)7Xʓz!���[�9,��Gl1���-΢Ti���=��)(	�./����(���Q�W�*�}��L�����m�g�)ͽN����*_����/��/ ��Kyrm�_5��ǣ$�]�2���Z�5�q7��<J�4:q'ә��0zE��-F3��;��U��aNt����b�Ƕ\~U��ƙH9a�R~t��#/�� �1�K�Ϊ�R���՚y(9�0��84��b7������kT����Jg8�p3=�}�תL�-#�T.<#�X�QN��;�g�>f�|��t�FF�w�[6g4Ǡd}ν��ʙ�X�i=pTh�ʄ5�q~--��O��OR\��%D��U��p��i�0`)sG��y��̦&�������XG3)�,%�i:�3���٦��flx�ǆ���*���	��1�qK(�O���]��-p��!X�Qc+7J�Ȁ�|I��X~���:jK�ml_�vC��g��C��^Жn�Kl��/lF/zpwx���0�3W<������� ~�EN�Њ1��y,���X��ѡh�]��?i�uW�6�=l�joŲ�����ũ����k//�b<����j�g\�aM�4���L�&6-h�cx��2΀��ۊ�n�?��\W�1�����ʂΗlO?��b�A7.�X�'���*b�e����-(3��KȗpC���3|ٱ�m�C�z)�Xʾ��<<I��݁�7���,��9��'*�y����`�	�87��XZө�mS����m�'���n��S�)S��0`)�~����T.�\�n�.G���u�]#�6�ݲ�asN��i������Mڱ��j���U����!x�;2��R���m�YP��8�$�~���E�߃S����̢7WpgUi�5٭�����Y��ka� sK�z���^��9�0���|��{r8h�B���W�~D���yՔy�]9�
��&�3~Y��bN�	?����)�Xʲ��Y@ￇH���1�S}��\^��;��)�5��ӫ��Qu-��t|�Q<B������He�R�]P���+��oa�fC:����j���r4�s?rwn����P��<�wC��T�(��k�f��$ K��6�]�ٷ>=�j�'���`xD��T��a��w¿���Ku�r�kPV��]=Y;�o�����#z�S跚�WTl��)�,6.�cU��U���;�"���W���I,eզ����Z�Eh�pt���pu�Moї�Cv-�T�q-���G�?�#�vb �A� ���W�K���tJ�s�{�6�o�ppծE���t�؂&��׭dϸ.s��]Tφt�|�2`)��pft��%wq�׍�=�E�\���J�4:Г��+�G�R�s����Ⱦ�Ç�yH�c�R6=�mL��-���<ґK�ӽd��@s8�"r��t	{D��#��\�I�W�%z��Xʦ�+@�䚥�yQ�V��GQ��������4L`��/�НG�E�ހ�,2`)��!#�e����b�eӨ�X%h��kؑ�زZ��'5���A?�G�< �c_E����=u���W�J��iW30��/�R��Uke�^���9e\�1�*��n��[��rW e�KYtBd�߰���yQ�+5�p&���Ye�p7�����8�0'z��R��r.��y�K�c�R��I��~���U��oT�X%�t�W�=غ���K��ׯ>�ѯ��H�b�R��ox�n�9QwG��!����A�K�hGW�,i�+��qV���.�0��,e�K��6�גT[�y�[�&Em�><�J���c�]tB(K�k�M��~r)R���5�gT�ɼN����u�@V�4��7��y�Ǣ>��C#>F���f?D�K���b��4��w J��s�/�g�h|��׀}y)CXʚ�h��;I�������b��]�_����~cS0��LdXԄ���-,eM�ـ�R?n�
X�i��j���� �F:-�����ΕRÀ�li@�~����o�yD�}X)�oT�7x��z8*`}���)3Xʖ�"��ɤ�#Q��D�7k[�oZ�{��i��)}�K�+^�%�ˀ�-q�T���`��~-X���%�`���W�ϾuY�J]]����U���G��C�2e�k@J�G��;i�2s�h�����R�5#z��+��ߣ�!aߖ��1�Y�V����H�4�t�uatKV
ĝ�I��@�oS
����%B���-.`��!T�XRF��?R�HΗ�ĘˊU۶�����:Y)WXʟ�)��q��5_��ڷaT���s]�,���+,�ϛ�]�w`�J���z�Aڽe�R���?sI�9Q���ҷAT����!�K��>i�AT����U�D��{�KY���@,��"�^k���*��M�w Ȁ������[7�܈jW\�J�"�,�KJ�:Q�\('��h�{�KY]��1`)�_:�;7�9�4�;7�v�ϻz>U�c�R����FQ��_Vʃ�܈�[�>+e�K�7�c)���j!*}G��(����]'Ȁ����ڱ����ϝ�q�R�'�M��N*�K��5i�MT�wQ�;3�5&ݶA���g[�N��I-�z������Z�n2�F*�K����iw���J��Q��"u�jN=��1`)�Z�<`���5���W)�/]i�R�:`M���vʟ��+��z4��7�����"�ꟓ^qk]�2�3Xʖ���~���Q3y��5X��.s#�0X�]x��j��s����%�G�a�_LZ�����������ڦ8`�e�R��-q?�Ӛ'I��zy�J��Q�@�"���IT?�Ye�K��:�~��ڀU?�l��Q:<�k��ʧu=¸��x)CXʖ%<A��~�0�tjúQ�G��J5f_#�~��q�"e�KY�hT����
itbT�I�%��2�� ��	)X[G�s���),eM܏�:Gҧ!����h�o�ϗ�y��F�;�n�KC������L1`)k�fN�ҸS��`��~��䑨��$����;�:�!e�KY���CY����H�����t�}�:�0`�9���+e�K�39*`Aw�']v���~�Fޙ���,�qD�����"��#��	�9,e�]�ZZ�h��l:��#�f���c���ᔈ~u�MGҤ9GE�[½Hc�R����Q3�ԣ'���8.��x�.��%�Lz\�Q�����Hc�R���ڰ��*i�;���*SP�<bӶ��s�I�����~$P��Ew0<jA��\���K+N��9�a�,�.��y
CRS����Q�p'R���E��}�g��ȣ���ȃ܌�g,P'�_��'��4h�	�=��#��1`)��G�:g���vm#{��%sSi&gϨ�s)uk� +X T&��M��E�܉����ք���^����Ȁ�y�����|/��,�hP6��M�3�Q�}���]h0�G�|�aj��ĭ�z~'|$(�����X]�I�d�RV�ȯ#W�1��XH�:6��
�RP���}ƕ��{:��@V�2�u#���8�L2`)�>�j�D��.��Di�>�L�b��k�G������y���w�"e�K�5��$�o��Oݥ���qt�+���'�#��Ⱦ��u��E�i_�׷�)�Xʮ��puEt��y�'(-�����{�)�\�J�HzF�JXaWn�,�������j?(�Xʲatf�Ⱦ��;Ji��:\ˑ���لRo���g�(�����]�0��k!PJ�e�R�}į�=�wS��~�B�������`�	�9�]�{��6}([�6(��(��2`)�&�����ޛ���Ȳ��"�NYf	�J�X��XL����.#��l�ClY@���)�Xʺ.<[@ѢOr��v�a =�����a*7rr��=BĮ];�`A�jQx�R���u�����
��m�� W{���ê0��Qv����K�+teð���h{q_A���f�j��Xʾ�G��7�O��NjǆL�GnӋwQv���=��8���G1�Fm1��Hg�R�}���:�.າ�����m�����-�9��;H�'<��?S�0(�S
�(<�R��KJ�Ky�zE��B��h^���	�A�]�V���Piq*����1�qi�^��u�@�W�[��SH�g�R>� �(p��C0;�����#8��q����cy����}؃�jh����>4)x�;.�K���Sص�����:�7��~x�~���~�y!*���������{����[�I�Ta�W)�U?����U9#P�5��2�bi�`��Җw2e�`�goՈ>G7�X6���Ua�E���H�`�R~������oW�.�����ğ��\^�kX��{�~�eKCP�T��D-x����;��ڄ���Ba��:x�U�a�R��ʦ_�̺t��1fvBϥ>Gr߫���9Ե3o!?gJ�o���<C�Ll�����0m��u+`�*)�Xʗ���:)gC��6���T͂�N��cx&U���ʾw8��͑�e���31�S�u.k}��A,��M�1)GXʛC�)l���j� ��~��m��� u����I	-J��z��x��E���)e��b��<Y���[ӖC�3��y�eƔТ�R�0`)o�҉�y��h�ѡU,�3�'¡k�Wӻ.[ђ�Áj��^�^�%�&�+���W�.�/��š-dj�g�
{�k��~�q�cw`���nG��į�J�K�������$.oZY��d:��.s�`����Y8P�����/�C;�D��8s_؟�k~Z�O�;�����/�j��1ۄ}�;$��.�)gXʣŜ�P�%��$|HZ��k��E��W��A�Jl���ZMJw�^)�Xʧ��e.��0iCmz>ī�Q>���!bU���ڰ��\��K,��P�p�I�'9�;s�?��І����L@�)���ffrې�9��(����+i��2)�Xʷ��7Ҏ�6�N�	P�O��c\_�ij�}t,��RR
��w��S�re	�
��f!�p'�r;�R�ӏKW;��,i)���[�C+9K��O����>\͙��W9��"�K�0�9��Y�R2�.<��M�Й�B�މR���\�<$���З;��a?J�B���箴��[�Y���aJx6��&-g����/��d�qm?���;���3��}�uxm?ޡ'�PT��K����6�zq&�k�9��K�R�W�9�Ї�k��g�xI_b���nnX�B��Ɇ5��SȽH�y0�6a�=��yׄp5I_c��Vf^:#85���k�1'q1A��)������N=⻌d���7��,iU>�������-�o1�y�z��Oٙ�Ƿ��8�3�����HZ��:���I�V��?��p�z��H�x�s8�}���r��L^A�j��5{���v��	�k�f2�.�#%mIe��<���a��,�1�7��FR���`]����v�b�p>O2)����]E6���A��=�-Uq�ٕ{�C^m%%fA����-i~�
�կd��+�^`�k����fThu��ڪr���}�a볰�a���<�RU���y����Zl�&ᐵ�h~-�:̩lo�_Rm[�ҋ����ؼr��ZM+�f!���r�}�׽*P�.�T}�y94)=����2`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR���'O-�@�    IEND�B`�PK
     ��Z��s��  �  /   images/9d204b9c-624e-42df-9128-467635275a1c.png�PNG

   IHDR   d      ���   gAMA  ���a   	pHYs  �  ��+   %tEXtdate:create 2024-06-16T02:31:32+00:00���   %tEXtdate:modify 2024-06-16T02:31:32+00:00g�JD  �IDATx��kHTQ�?�)�OP�#��
�Q��BȂ""����B��V���0����bR�z@�!�C�dDjTD�� R��f2q�j�{Fb��^�{�e���^{߱� J$�%i0!�D�q�OD L�t����S�ijd��#�#����9�-�4��Fm����s���
��p�����~����p�V;��f�I�Y�3N��f ^���W�IR)�D��WG�*�H�4�J�*�N��bUj�qHѮ�(p�~E8�g:c/i�o ��,c�8@���À������:s�6'�`�2�-�*A��{�MJ�%y^�:�J*�E`(;��h��&�]���D���~��F>qȜ�$P��fd�D��8�Y��,W��S�"�w�bFd�h�Hp=�^�zNv��	_�S�I����z���lߓj���}���2̈��,�<=�l����e�/��#s����$�mFDb��8���a,PI���Sy�ϕ�:\�\�ssS1�+��	����]欖Pz6��>Z#���=�7Z��6������fay���1	�s��^�������i�yĚ-mv�V�¥�7Yu�o�K�nˠ`hҬT�����dmA���e�{+)W����,��v�ѧ��f�J�*�*3�y�����[��%��S�%�q�/VV��o.n�3�����5"cT-�&�w�g�ʐ	��`�}fHf��/T�UX��^0/Q<:\�V�U%&D��4D�D~��I�
��    IEND�B`�PK
     ��ZP�x&�  �  /   images/9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.png�PNG

   IHDR  �   �   ���   gAMA  ���a   	pHYs  2�  2�(dZ�  tIDATx���y��g}����Ό4:��ut�,��Bb .��cKR�uRiUm�6U����,��J��zۉ�1��C�c���6f�lK��,i���ߞ�>��g���<[���������ꑫ�s�/�[����Q�1�`v�yꙁ1�
BPQl��fz��p$`&��W *AE�)%���_5�Zf[S��2GP�l���(��#�ǵ-f�p�S �LT,?%.5:j����gX"w~��r����W	� ����V�_>�Vj��d��� @!�(-JBJ�C����E���c e���D�?e�Q(����5��OvO	 �0���������l�	k,O] �DT,�w��H_�h�	��	�cNT�����&�%�CP���oZ%7ߵG���r�	���L�9'��k�~������S��R %���d���}�_��٣��RQc�EÍ��Ds�� %�����e��7xQM��;�Du�S��9�ՃZ��O�X `T��U�W�����u�֑�ɼsNXoT"O��O�b�ښ3	�e@PQҮ޹��t%���W�fr�F���Ñ�g��l7�>vtN ��*����&	�o�vg����_xP����艆"[c�x�� EBPQ6�V���n������]�^��v)���V�R�����_	 ,1���sՖ�r��z�ܰN���T�b�B��Wk�mo��
 ,���<��}��Vݣ6�(%�#�+`&��� � AEٻ�[��n���^���uJ�C����v,��D `TT��W��>�k>������W"��2�5~X#F�Ds� �" ��(�v��>�'�c6�d��sJԟڢ�4	�c"�6��L pq**Ү6���NT���c`ѱD��=��DPQ�V����޻}�1�`�x�9%�����P$�Z�m-�_ \"����a���C�$��������l�R��'�xT�Z3� �HUc۵�w�{��H�����Rs'�� �UEJ��+0�L�H�9��_�n���cɸ�$ ����*�i����-}�G���L}���Ñ�?���%���
 �APQ�6�Y�}���.��e��%E�E��Z���BPǞ�6���9Yx/��Z�׽t_+K6�  pA.X��NB��������P*�1���*�'B�`�F�<O U����!�F���}�J���D�w�+%�E>j<<�f�3M���jT���o�8�����%�V�+��H�Lĭ���DPF�!��M\��B�ld�����j5�ň�5���BP���vc���-�s#��u|h:Z}����ku��9�C T�
\��{��>�^���j�^R���UN7�Ds����T�2�y����8u*�1��߯O9�ը6t,�d ����~m��o�1��5�PIHi��p$�o"5f"�sL T�
\����z���nXg�����C�C��VՉy�'�IP1*�Hv�������1���Yy�m6_ �����ΐk7(������:
���$��1g�Ub�͙���FP�%�~�*��q�Xg���N��s�z���P$���lm�؋�=�,T`	���}�_镳G-�B�l���l]6n:����@�!�@�e��5���C��*��g��j��*�ڒ~Z ��
ɪu+�����Ho�M��j�F��Pc�_��f[s&! JA����OWb�	�%s3��sJ�cJ���� p�ް�LJ�
��EP�e�3|��n��������"��d<�mP�*���V���n�6�����sJ�NQ�[�H�6��lJ�R ��
������w|p��O��l,�-�tW�;��;�WU6k}�7# JAJ��a�۴�V�kAJ�R��DC��X��zP ,;�
��kn�:�uf8���uJ�@T�K��� ˆ�%j�U+�;v]xM�%�}S���E�~�Y��K����)Pt(q�v��>�'��kv��1�'��?	E��%/mʽb��!�@��u�&	� �G2ҕ(8���]��`T5j3�l}O A�Ȋ�Zy�{�;amp�j�@�x�9%�����P$p�6l�dS��`IT�mغZn��>I�>�]c8=����R*R�k"������;�B����!�@�vm��n�s���L��5v���`��9�E��*P攡d���3�#��j�"���Q�ֱ��y�h*P!�4����-}��cు�B��c�pc���rf��� �b�0�w��>����沅NϨ���h(�%�ֽ��T�B�q��7xww��SJŜ�jT�2�����BP�
�ru�\��^XݍKC����y"	4lm����KBP�*�\#���>�99�ufb.�Rr��Qw�O�fb퇇��p��"�߾Q����K��+8�D��*�>�+K4Y_ "�@�1j�xw�BX3�{��"T�f��K�j5jhk��[@A�Rk7��M���{n�{<>8�w�Y�ަ��Í���5�l{�� oAP�*�e�U���k�^X�.4�_TNEÑ@,�>% ��
����-ޥ��c�ԩ��l��o�R���QQ�L6Y�����W��N·���^X����sNX��~�V���0�-���r�[lܶV6~d�t�xa����T�#J�8+�jm;v�%���@ � 
�q��.��xW�X�:��h(�%����B���:C�����k�����Rt��5�m6��X"��� U���(�6����H��։�B��/�x1	|����<���� ApI�^�������]����QJ��l6��c��
P�*�˲�-�ӧ�
L�z��~'�Q���)�� ���l�֭��߿���Hf2�����SNX���m�lɴ
Pa*�+v��uާ+1��Ւ��\�9'��Q�GÍ��g��ؙ�3���A�hv�������3��f��^�k���%@ � U�y�m�����5�wN�ک���{����5�!@#� ���ͫ��+�3��~Ē���B�w�'	~M�̙���f(C��r/�x�R���>�T���lM4	Ēq���
�(��u�|X-g�Z�Z���H *�a&�R�
P&*��Y}�J��]��d�o*��R���	E�?2D��x�� %��(�M��y���ފ5;[��=Z��]�����19$��@P,�]7l���=�Z���w��A�h3��+@	"� �U]}���=�%����x�{<���=Ώ�QC�Xks��(!@Iذu��r�>I�>�����F��hёp$��\N�'_H^�EDP��m�6�_
q���J��QkGÍ�X�9�� ˌ�(9J)�����'��d�G�ω�����6����b=/�2!� J֚+��;wK_Ǩ�b����ﻜ?n<�u���w���*���y�z��q��k.k�T�T��.ܶt� EDP���7n����6Xp�Y�Ɯ��A���ZM?!@T ee��Z��};.�5#���lD�WJ���b�X���� K��(K�5r��IϩAi?��鉹��J���E��ܤ���,��;?�K-@���Y�Ŵ�m��>�Z_�9��'zO\�m�GVo������Kk�����}V� ʞQ����/�5#�����sc2���L��B�n�GV��I��BPT����?������t޹���e��>Y��vo�ZS�E�+EPT�-{��>�_���j��?��~�[��sV�k7L�+APT�=7o���oӒ�y)/m�X���Z�m\�
��կ����;��n��:dM�����P�CR�~������+�� � ���mke�G�Jwۀ�xv2�wnz��Ys��_UF� ���>�� � ��{���#�7կ{'�|qY*���ޠ�)�ڕ�ٔ�+BPT����x���,
�
��,t�Û������n@��|ӊ��r� AP��G�]��2j�]����Ũ=��{� Enr`�j�׷]��~dˁG?q9�o��I\V� ��Pzb��_��9���f�7ۮ_�	�APVf&�NH-�n\`R��Z��x�	���(���쑌䲶��Ί4n�+@T %��c�������	�k�Ui����(Y�3NH-ɴ���Z~�JͶ�y�	APr�8z+�s���ωV�b�x��APRR�y�w��f��|����R� �
�$g&�ݻ���`�Ui�#�O�� %��XVs�Y����M-�f2n}W�DP,���^L��9�9����tL�� ��*���������?����1���8�
�h&Gf��uf�P�W�0�ds�Y�APnH�ݻ�p��(3��J;���#�L�.x�kje�L<ۻ`u�RDP,�ѾI�r�����F_�Ebm��/(c��rw�!�l���Ӣ��'�� ��X4�YRw����B�[���jm�L�*Ap��ǼMG#�I�9��)[��ɖL� ���l�}������!�9'�'�;O�� ���,��zw�:��������Y*ApI2g��ǻ�J�h��YWWk�iw� U���(c�S^H�:F�ߢmgU��� U��𕛳��v��Ԓ�"�����B@A�mަ�٩���j�U��̄ U��x��Ը�ak�>j��ֆ�lI�&@�#� �MO�y!M���sV�m���l�	 A�9�Z��]��+|����z�m0� �A�\�/����~G�8�����Rn@�ǻ��G|���chk��[@A�2�#ݳG,9l�c0}b�X���� XA�H��A����Ĝ*}xڞ��Ǉ��� �T�
�'����}紖�[����pI*P�f&����m�L��Z����  .A*�{U���(��}���`� W��ƽ����������rf��� �b�C3r��%����_�ֱ��y�h*P洭�G�^����z�P*�ڜ�� Xt(c�ׇ�ǻ��L�G�K�� K��eh83)�G,�Y���ۆm�l�}Y ,)�
����Ҍt%��Z�m&���@QT�Lt����+���|紖����6�^�?/`QT���w�y�wG����h��R#�y"�:%qPd(Q�#3ފ�:3�?��+��X�%�� X6(AnH۝�/-cZy�=( �AJH���w�����`�|Ues�ċ�T@�T���Nz+���1�A�_Ԇ2���_
��BP�e47��B����;�Ew�6ܷ�|[ �$�
,��Ā�=byQ�e��e�F3y(��uH �A�l�{̻.�}��G����lk�$D,P�*P$Sc�^Hӧ�|����b�����lT��_��.gp����)���� (;XB��ao�����*�F]�6v���P�*�F�����u���9֗��Ϊ4�sP�*��rs�w�Q��>�A-i'��1����@P�Eҝ�b:;���sB���b�I��/��BP�+4�3�tؚ����Dj�Ui�1Pq*p���缐�N�jIjCǒ��!P�*pν�+�G2bۅ��8��U"f"��� �x��s#^HǇ���<�k�U�sV� �
����-G��G|��_i1bm��aPU*����^H��?���)�f2n}E T%�
�sr��t431�;�J�5f�3M���8 �h�-C�	/�C�q�9gU���D�:* �A.�����+S_Z���{�}� T��~G�޽��ھsZ{ߓ�� �o!��j}�G�ǻcS��Z�Y�l,��wV  ���414�4�>��话U����& UE���W{��Q��`�I �"TT���Cަ����&���_'���N������g&���o���J��MGm-�_ \"���得�}�뾧ԏiW�}O�=��DPQ�:O�;�RK�s��`���c2�6���+@PQQ�;G�ǻ����`��ֈ;O� Xard��uv�w�Y�Uڎ%㙟 ,"���熴������1mh3�d=$ �*�V�����hj������Zm�Ǜ2��O�
T����I/�]c��Z� 5�L>��� �#�(s39�����&u��f�- P$e�+��}W�F՗֟�߳�<��Q����"#�(i�c]����wO�b��♄�% Pl%��h���x�Gk}\�2��� ,#�����qc�ww��)��m0� (%ý����Խ����o��:��ᮔ @� �Xv�5��NH�:G}紖�C��f�%�CP��~���&tJkK��_ (Q%�Y�~~��Z��'�� JAE��?]�J{�	 ���Ң%��6�-֓ e���$h�s"�=���Rj� K��b�iy\l'��ӝ,��/��7a�T,gU�+���9�� @�#�(:-ҫ���X_ ���Pn�yꙁ1�
BPQT���' *A `T  ���>�9�<    IEND�B`�PK
     ��Ẓ;�  �  /   images/f39c2bb7-8598-4025-b62d-e677fac223ba.png�PNG

   IHDR   d   +   ��-�   gAMA  ���a   	pHYs  2�  2�(dZ�  dIDATx��ilTU��[f����.����%j��Q0�� ~p�f�Q	FSVk����J\������"(n�H��e���}�����uf��9��1�	���涯��ɼ�ߜ�?��;<��I��I����փ�Hd<�2 �z�f�r������əS���O�ZZJW �Ti�r�b��Ò(o�-l#0+�K��hu�cۖ9ނm3h,C ӒPu{)1X�q�_�����x�u3,s%�4��ǚ�@dY���ʅ%P\�omo�<�v�V����8|��kI�W]S�}p��a`d�Y� BB& 
�ͷ���B��RW�ww�7�7Xr,Ǩ�,KP�t�����y�V2U�$+����`BY.�]
��h�}HE�_�1H ��ʜ���p@T���L��%y�����1���~/oG0>���.g�D�a�(�c��*�I3&䴝���m�Fy��m\�)Ø�H�Z�3��@2"������S��]P���y'�}RH
��8��X�Q�8L-� �J�F���)㡀���ࢎF���@�2��Ł���0�?N���M��J%`0͚zk�T�C�y�����Hz/�_;̀�/���8��Ȕ@e�Ś�����P6s�������8��!��v�2�##�G�y�dt�_
����i�������tG�B0���?I]RL�"M6=U��c�\X����;q(�.����f�^R�1�a�KYD����10�6���y�E�����ñ�����A�_�0/��#)뀐�i��s��g��x^�u��
Iqk*%~dg�ȈF��a��@T�4��m|�˲
�u��aa�a�{ZH����=MQb���'��@T)�0�����Y�cpqg����Cxz�,��T���٠���J�N� �?��O%M��1��bA1�"��F�c}+�1᭟�=S�t}KR� )����P�,��B^��Ɉ�T9��BW�%���N&�j�l����`�oޤG�a,�/M�r�nKYM��E@�%�C`;�\����/y%vX����pn��cs:Z`\�*6ov[��-=�m�M�!�&�_8����-Aw�MNH�9��s��iW3���B���b8QL������[S�B�����s�rr��_T�J�u�L��8�$>Vl��y����$�x�p��3�
̀��	��E�썶G</U-9r^�C��n_`�
K�!+� ��S�p8MvxP�NQ��.�����Ϡ?�����\���X4j�����6Z�6��pq<����-B|(�>���\���-^�,D�ﯻY7��0QDPF����¾x=��x{F��R�(�E0�����'<0�i��F���-pA&��Ųj0���5�il,�T"��rp0v �����I�UF���* �O�����1N�ӯ�V���Ez��7Ad�� �%{
�b���	�7Z{W�7.U�B�z�|�M����C�Ŕ���p��ptԅ��v�����0���/Bɸ�&�}"�)}$��Ic���L�|"����K�Ke4����*��u&�I7˙����ݮ�Ox�?J�L�������;L����@T�ybXO�Ot�ۄ����'�IEU>(�Q��8h���.�Q}"1��vLc�.%c�n|��x�������&8��;*Fː@X�	̖���G>��7��K�'h���;��I���OHx�B�F>���>Q�>q�|�����>��9��0@��'�����]���O	��G9�vI�	���ES��#C �T��U;��h<�ڃ'�AK��:���m@��8�L� �ё
��GŴ�2��%rt2u���%\�m�:Hw ��|���� aY}D��'Z3M7�6�j�ԓi    IEND�B`�PK
     ��ZFI��  �  /   images/3d3e563e-9ba6-48b4-a3f8-79399330dfef.png�PNG

   IHDR  �   �   ���   gAMA  ���a   	pHYs  2�  2�(dZ�  @IDATx���y��}���ӳ�[3��i!���0���N��;�/�k���W;$�J*�+��[�zp��m�ڙ���1��k�� �@�ݙ��}����;3={�N?��KŞ�V{���T�(?�����tϯ�N�I�g՛M[:� U��br)�F��ʆp�L�� �A�TX���a,��"fS*�A ��TL�"��ꣁ@�\ݜ9$ P�*��sZ��P�����fc��� �_٤���[�J�QT���^��FC$�Rie&ҹ� T����D]���&	�����#�l� @ �(S�s�?�X��4�}��W ��T�5���O�>+��P��5�( P�*���~d��ە�7�{�(�C�j�5�a6���	 ���)�<4]n�v���u;3r�{��sZ��Vzc,L�Ro6�:�
 �	���q�;�x׆�/���TL��h�ꐙh�}G �T��/�/��s���-m]Eg�R3��~;���2�Zs� �Bei��z�5�x8��i�P����R�3�<�	�\فx�5� � �(k�-��][XNX;�g�.:�D}A��H蛆�3W7K�� 0A**��Gnoޟ��?�B0�Q�d*�� �$!��3�������y����R��?�b�`Tk�L�vm �`gż�꺥�:2�f��S��R7*��!z��2��}B `�TT,����iu��L�9�䯆�@�!2��ܽ ����}���K��9��	��r�����DCQ1�x�%� ㈠�*,�]/_�z�\}����-Wj�F�m<��_�oz5�S `TT����M�r�vWF�����8a��Qg|)	�Kc*g:��1}x �BPQ�nxWH§O�/��F����`t���T�q�1"��Zs���w��|��S%>��ԻQ�5�CQð�Ɩ�V��DPQ�.�?Cn��2y�p�{1D�w��R�i��O�
�~���|�� 8C5��+掜V�ݓ-9g(�=]��H�L��� � AEM	8��?�|��k_=�]tN�������H(�EǓ)�? |TԤ%s���k��kǻ���J�^����X8�ce�xc��W ������빽Y/����3JVj�V6��f2m}M �T���Id�\'����|�9���PTiO���
 �FP�ӂ3���-:֌��(�f�D.s����|��f�%�, jA~˻Λ!��e�I���7Tj�3��3��}��ՙ�����	 Ս�%|��sG~�>c-E)��������
��DP�%7]�������9a�a�{�*��tn� �)8˂���߿��[u�ڞ/�f�a�d]C$��#ޔ� 5��g��f{���%7�����u�h�2����P�*0pɼ����;��Q��������%-�d:�F T-�
�Ѽ�u�?�Z4��}�F�t����H�Wu�0Ng[@�!��9�d�L�r��ꆵ��PtN��������1�\�|�G T�
��^9���/Wr�	�?
=��U!3њk U���hz�!��򼑰��^���,sʺ:	F������FP�*0����m�.�֣]^XOv��TS�<�51`��k�<" *A&�U��]vg��j]jRŦ��hC$O�r� �����K�|ͦ�����R3�ȷb�`TO�� ���d��:�5�x$��2���z�h�EC8��J�Dk�5P�*0�.[4ӹ�˖�֞��R�����"��r�9s��R�}� �A�����f�y�o��Cӂц�2���#�,T`
ͬ7��w��f��D�w=(�B�45��+����9�I ��
���˪,�ԑ�5����k6J��۶��p�!�'wt���@P�2�T�:��w�R�����@4	���=`�T�}��#aM)�f#j���w�5eē��S`�T�L-�]/Y<֝i�_�QJ]-���ͮ�ͦW�;��#�@��|�,�ڴ?煵o����(��(�6�Cw��Ιw��0*P!n�(4r��V�9��m�`�v�fc*�� �� ���s�Y8rx��ޢsJ�EZ�c�iu�2l3ђI L(�
T��ϐ��Is[�k�w��sZ��h�S�p���v��m�0!*P��9��i��=�҃J�f���6��Ɠ�����#�@�3�c�/_ ��ú�Xw�I5_)��X$-h;�H:�� 7���L��5K$��ㄵS�Z%ߥ���2~�	��P�ll��
�sFP�*s�Y���ޜ�5��B�+���*㉴u� 8'�R�84rx��k6�T�9�F�֦֟
�1!�@�;= ��o�HX�v�Z��K��>��Vڢͦ��� 8+�-�!�e��P�{1D�o���M���"��F ��9���V o#�@���sGN���^�Q��޶����`�1m�P ���5��P�GW,y����ld�V����hO��u�$�
Ԩ��i�g�_";�u{a=�/�f�D����"��b�M��A�;*P�޳l�wmܓ��:d���)���`<���. ��
��������p��R����X8u�k&ӹ5�CP�ͬ�/\�h$��;��*�B���!����L����8�
�w\�p�wm=h�Z'�]���sJ��������+̌�x{{�_8Վ�(���iՍ���VR�?N7����C�DKn� 5���5�ΐ�^y��m�7�{��)%�D�ñp0jkoj�=+@!� ����t��ڥ�z���ɮ��J}�P�LC$����̇[;�P*��r�;�x׆�/��Ė��PP�h,�'Rַ�r���x�|�,��E������S��w5��Qe(3ђ{R�*EP�قYurk��5�C��k6J����_���_�v�lڞ�!@�!� ��e�fzז�֞��k6NYo1�-�H讙�\��=�/@� � ���GN����~��{���"*ޔ�5	P*�q5�ސ�������=%&�
C$9�|Ո'Z�/P�*�	�b�tY����:2�f��]|�F)�q���p�a=4d&wt�P�*�	�T�:��w��������P<��}W�
CPL�O^6$�i��Z�5����X$�b��T�)*A0iή�?�,	k[�ԏ|UD���sZ�Y P0W7w�)@�#� &��gyצ�9/�}�v�9�䋶���;�Ks�5k��>0�*�)s�E������sNX��\f"�}L�2DPL�����,	�E用E��"��-v�)�Q�2BP���ϐ�uˤ�-/�vf$�;Tj�S��j��Qo�l�wP*��r��sO�t�S�ٝ-9���u����
ϋ7���`�T e�P"���#a�~��Ĥ�g(}_C$5�m6��O0E*���xN�D�^ℵG��씣�@�9���je�fU$�m&S�&AP��\2˻�ߗ��:P(�UsC��N^�㉴u� ����}��k6[�^���ph�vO�i�	&APQ�N�-�=�f�3#{;��و�K����k6J�xc��&����W6i&˳�`<\�`��Ň�ɶ��k6���k67i�n����d��Ů�}��[�=	�����~�����PT�kW�9�n�[z�&��+����d.�J~�go@ū3���$r�pXw/�fcZrޮ��n��Q�]`�T Uc��i�g�_����|�5��7dI�W�k鍒uN�C3�p�*��󞥳�k㞬���!��#�9�7���]�%�AP�~��y#���/�m���q'���j��0@Uͨ�/\�h$��;������E��%���ց9p6*��p�y3���gz/�X�+#]�ſU>��V�V���
ց�	�
 �8 � j��F%�[�o�Yx�|1&@Usߠ�����g��GI8'@�mmƣ�f0.*��3ڋ�0�*�����Ճo�]��1����s�`��"!�ځq������.�>8�����$�'T �>��Ѣ�����ߍ��m�� � *�����������x"mm����;&APQ����|i��J�d�zB�I@PT����Si�Fy?|"�C�IDP����{�����`l�'��t� ���(['�eݮN�~��9�n3�m6��O0E*������3���Lꬭ�xS:�=�APV�ۆ�`2����hy`F�6ؖ��T e�`����������vN��(#���^�y���}@i�L���	P�*�)�i΋iߠ�;���i]j�׬�� e���to���Bږ���sB��@�`�n�zS��5�
`Ҝ��B�>�5ʤNi1�d:�� ���nH�;�-�K��'��w�0��J9�Q7���ԗ��e�`&wt�P�*�	q8��t��9��3�0�T�*A0�zm/����F�ԇmQ��$@ � �͖�Ӟ�Q�[����~�Ap�v���Bz(��?��/l;`6m����T c��3䅴�-�;��~U�L��'�R��l؝�b������O�v�`�%@�#� �J���5��]�k0Zt�Nי�;�P*�3r$7��F���sd}��*��j=+@!� |ٲ�	����`��cʐx"e��T %m=hy1��mF��oό�8��-@�"� ~��S�k0�;��`�ֿVZ��V+-��=S��T #r��k0������7���L[k����lܓ�b:d�ރ�Z�N��|] �7�q;�u{!=�eR�H+�lJ�
��AP�u��B������h�J�	��*Pc�[��vfd���h�'��D��� AjȶCy�T���Ӣ������h�`pAj����J�v�6�[�ٔ�^ g��U,�_�B������٭�6i�`L*P��ߛ�u�:e����pt� 8'�2���8��N9j���8�����٘��
�sFP�*q�k�����ب��}����#���`�T���zx�=�����n��/ �A*Xs[ދi��F����^�ߖ� ���`fxf�)�5��V��H�_ ���{�མ���������k0���� �@�ش?�J��l�9�Tz��i˼C���"�@�{�D�Ҷ\������l���N0�*P�Nuz�w�G�|��-��x2�}J L�
�!7��˟΋(�-G��)GP�2�rN�nL;�ө��!*ē;��@Y �@8���B��D�����@ `�n�l e��S�w��B�y�(����V�L��G@Y"���r���30�v�]��\���EP�I��d��C�5���+0���@�#��$���B����t�*�LYO
��AP�I�aw�{V�����u�V�̷@�!��j=:�s�kp�I��u��ҝG@E"��8�^�y��g�I����Si��Q T4�
�����5�����h-ǔ3�j5
��@P�q��AˋiW�wN��;�m�n>6��@!��9�s����>�9'���ӆ�p:�*��=S ���c���B����h��k-�w���EP�1xvO֋i�.��DtH�6i���T�,�z��i{��-�Z����Fi*wP ��
��cր�׎w�6�Yi�;�����T��`A{!}nov�ѓZk�k0
��DP�^>��bj���9!�oִ:���;��.P�*�[�u�y!���;���%f2e5��GP�Ӭ���5�d�G��RZ��I* pA�3R�T�>3�s�9�� ~AEMs�����/-?V�s*MY{ � ��I��Rw�t[�h�-G�) �������u;3ޛ��8�(�9��/ p*j���]�T꾃׏��j����V� �"��z2}ީ��*������6�R�� g���ju����)���>[�xS:�� �TT�M�r�vWF����F��1m��[/��#��*o���N�m�~�A-�j�xӫ��	�sGPQNu�Z'��G���4�a��� �#����H����i��J��t�^�	@PQ�RG���v���i-�����' &AE�9���B��d�������dk�f�	FPQ1zm�����|�ևD)�u�� L������J;�gp�5�o���Y &AEY�urx�P�F�����Dk�5�)@PQ�:{�ۻ-m�����VfS��K�)DPQv6��x�R�Wi�{��ܯ�|G �T���nHOv���S'��7�-G �AŔ;���n����E?gh�lL� (3S��/�����U���j (Se�9�~'8#h��R[� @#�(S��m�I�ZE,�rGPQV���J+3��~. PA*ʂ�2h�vC�M&�Rj� ��b�i�����!&к�~�/a�TL�Ͷ�ٔ�6 T8���p�9��_�yP �JTL.��g՛M[:� U��bR%��W �A `T  ��]*�ܴ��    IEND�B`�PK
     ��Z��C��  �  /   images/89208456-78cc-4fe1-a1e6-da24e243623e.png�PNG

   IHDR   d   +   ��-�   gAMA  ���a   	pHYs  2�  2�(dZ�  oIDATx��ileǟwfv���v��UA�z G I��J�1����cD��p*x��VEc�Q?LT���Rm-��^,��ݝ�w��yv�5�D���Y��,��4;��>�o�w^	J�e�|w�n��N�ߗ�*0V8����Z�_�������⡣�5�zX��9)S+\�S�I�6�0V{D�]�hl�[u඾���5`ql$��º3 ���+/��w���{$��X��LÄƎSF��}�b �]C�[����L��wtGkLޕV����w�.1E0�5�p�*Ƅ�@HE��wÒ9�a�Y�	ۻ��G2fT}e�[���-�,�����:�X[ �!0�Q��֍��i�{��HbVs0�m(�l�wVy$�?.�g)�il//(�rr4C�.�R�'�`W�|��ь�6�%��	tN�Z���� c[ �E7��~����a�$�剎��"�ˋ�v=�Ee# �(89��S��	��p����y�_��+�f�h�!��-~]<3���Ø#��p�\4��E�����쑿:W�0�\햄�"���`]���Q@xT���+����*h���;�AΨ�c�/�������0�B1��X����䗪J�����R�q[��zc�ۭ3(�/���W��q,�ڀ�7�&o��>�`VT��&�5e²Y�_�����~�>�����q(�1�P>�ë=>�|�S�
�l��_hb��i�Y�格�P��XFۄ~و~����x�fwde�����Hp��3`�d�&?w`8}oV՟�)��������)K <�1t�I5xx�D8p,5���@8����L�Ba��s�����ea�_��_��W�y<�~���x�\�'vr���ԑ�O�J�Ӏ��mPyp�n��_$����֠_��/����7ų�kw7>��g�D����ҋ��U�*(U� �9KT�ѦX3�����Ιc�/�ۻ����;�'��z����\��+��-�,��V�Y%�s�W�	�9b��r��=���_��ӛ��B��$�!;f�<m����"��u�/.������h����pdkf⯅��Z+z�JC��b*��`�,�?[���`	��#f�P7���\���c+X7d��נTA�����x�2j-B�#��G3��	t�d~�c�'G��t)^ǌ����o�ő�^wtr���,�,Y�A:U�pB���(�&FR9�el���y<�Lmn��������.딆��nwS���b��/����<���A5<�`��J}�e�*B�_}k(M�(�s�����%�2,q(n�vH��� z��tE���NE3V����5�ȟC�P�.����l��B�.��I5_�I��9mj|��%�t�(������=�Vh���hJ}���	E����XvLY !OP����d��)�~��XY!�{	���w¢:G���"z�?�EOD��x�;�kjU�D�A�����[�#�pO���eZn*'��+x��KHșL�U4a���_�pr��2��zc���I���x�/mMu����r�R�@�`���.�a�~b7q���/��ዯm�{�p$��ġ�ެj�m�M~t��uV�Î8=��=Nk�d���xV{�^���؂�`4���^+�)�§��X�y'��}�kpx��(t����V@�'��`z�?��^3���B��i��j���?�6@�G�|���:�~*�U�����j��W� ��sl�-	q��3���M8*mDOD+]���a��wX�OH�oYl�#%$�*��z���~�dV�3�z����)9����pB��f�3�$�d��,n%�%�_B�*�    IEND�B`�PK
     ��ZP��/ǽ  ǽ  /   images/0b351edc-7875-4477-b820-546ce15be531.png�PNG

   IHDR  u  v   ��:   sBIT|d�    IDATx���}tSwz/��$۲0���Mblc0fB��3���@��0�b�!d�qN�bν'�tAgڣ�rf��i��Ճ���M�8�Ms�z��� N�`L�~��-�/��ClE�e[/{k���Y+kY��O��g?���S��ҡ�D�P�C���{HDDDDD�;����_��{�R�=�p����V)v9""""��Ή�:�t(I�R�)xZ�Q��5�cR�GBנP�@��x�1�cR��+o6I���t�|�&�I ����W��ǙM~��<>/(�^h�J""""
O����=�p���`T��F��:ix./M�8�IV�0<<,�0������ ~�}�M�Kb�J�/^:���Q��)��ӣ ]��+���!�L-[�,(q��~cP�Qx��+u>HT�*�GT�K�N�F#�0�����BN�T���@{��c�NQ9*���!�S�=�p�n�DDDDD��abg�{�aR祄W��="""""�G('v�~I�v|b��
[�M�6ן)�B�;JX�&"""�^�N�dRDO�f੅�`�b���y��A�����DF=T*~��"�bb�������_��g}� �L|v;>��f�@�|y`��6��~�PN�JU�Pث�B�GIDDD^B1��^Jx�PI�g9������~�1��y��\oo/���@�Z����80w��Y���G'Q�f
���c��	��0����'�C
���䎈��h�P�:�aLv��0�Ə��8��/�ҡ:m�Ҡ ^��٨���w��cqyX˸�˸�Ըb����q7��
B�b�J��X���Z���qu\e����MRʕP��{`<�}���R�a��A�<�,]�q��G��s"�������m>=?*v�~I��v\���H�����_�W�J�@�g�DDDDA
]1���1!����(F~�r;"""���N���);`W�*���	F~�r���`�#"""

�r�f��0e�tk�f����봯��f �S&&�ݮC�RA�R1.�2.�W,6����O�P ֋�y�q7��I��f��b�`xx `�Za��  � ��������"��<x��:�����e�?�S `||f�FGGKllRSS��!�2.�2��q�b��1:j���H��R*��?���\�e\�<n8`RG����`�Zq���ޅ��?�6�������9Z-���/��#�uB�)�o�<`�P�B�|ǟ_W*�P��D h��q�?>�v�Wg�˸�˸���B��J�9s�tA*\����xu1ʸ�˸��L���������z��c;Vcn������ݻ���|���>�����ݻHNLD�R	����	L���X`������͎/&&�y��]�����BZf&������(�k�Z���?}(��"<����8f}��6��1���F�oV�[���pa�P(`���q�q%�+�@.H]/D�q7�qCYd���fý{���ڊ�`�Ղ�y�H���%&c�}p���� ��#QJE,���0������F���`Q����b����ܩ����)lF��� 7&����q�q7Xq������˸��	���&A[k+�:��א9/��x���`��8J qJ%�J$ƨ`�����������'�=�RRR�z���.�Z��ƕ6c�MPR8.�ZZZ�~�ʕ�D�0c\�e\ƕ�J����;ר�fɒ<Q.D�q72ӟ�|U��Ʉ/._��cu��j��Q����qc
̍�A�J��]��f5z�菡/-EFF�#�"v4�=W#�x�I�ꛦ@�`
�����&�)�e\�e\�X,V�_���~�q7��"��d��_��G���I0wv`��W�1
t11xT���}�O���B{{��1"�ݎ�oa0�K4������:��d�o��a�ڄ�9��&��$�� �T���x�_���＃��nIbE"��� �&�D����(�0��r###�M}=p���`W�A(M�*H���D�u4��?��ݻ��$""""�DLꢘ�f���1|�7��SWWP�����k���gQ6��t��W��!Q4aR��Z[��#;I�� 't�X�ɱ1�{���ٳA������(0��R###�ZW�m"�;�2�r:j��qq���Z���m� !�r�a2�MY"��������(����B�sc����e��F��vxW~�kV눈���|��.
Y,�7��|�C==r�c�����~�vÜV(V��ЫE&uQ���Z�#���N��,N�D�݆�S��J�
�J���@DDD�b�@4��ݥؖ�,�Y��5O�C��`���54`�ܹ�Z���
�����s����{H�'��9?>T��A'Ʊ��ӽ~nll�!�q�qe������u			�˸�BqC�� �L����z����_H�X,�tu ���m0�X��!t~�%��^QJn
@7��C�^�N� @�MY!�q��Ұx�b�~gxxV��7H�q�qŌ+�����;V���Ì˸�+s�P��Q���/��T���/�P<�Q*�Q����,�PB��.N"%��@������D�/!!j��q�q7hqŒ��������{j�:�J�2.�7T1��2��혫���phn���cm]��~'�PB�B�����=��WU(��K/��^�1.�2.����Q����˸�x�P��Qftp�PȾ��LT
��^ht�Uj��h����^:��P(���u�J����.�			���^Mkf\�e\��5�X
E��!)�f*)�2.�70��2C�3�'�J���.���(xZεu��!�*]LLFGG���+�x�v;�2.�2�$qŢT*#���q�\1��211*����ƬT
�G��P���P��/^n
fܹ�*W /r�͆��Q��ĸ�˸���v�,�g\�e���5uDaJ�b&�F�t()X1���P�Jc�����E�ؘ�(�*Y��B��J���nΏ�ؔ�6G!""""q1�#
sBb7�Ǉ$��oʙ����(ېh��j4rcF���,��B�@A�Mِ��������])�x�P�æ(~�����w2�����:�<�������a1.�2.�J�A�<|�rیω���q7��"^9{)��C%1P�	��K��?��Ǽn����+z�իG��~��|y��	Q�-���	Ld/Ď��I����%9n����Ʉ�f~��@���ʡ
�BiP EQD3���,�+uQF����/>Gl|<F����G�v;�͐{aK���1P�Ѿ��'v،C�Û/x���ĩT�
����Qx`Re2�z|u�#h�ڐL���vL���Z�B=�O+�|Z�w쯼��ݎ(lm6�\����

{�(Q(P L�%"""����.�:�ڝ^<��>�R?O��&��		S�#Y����;�?P�v;,6;�=���P�i�Oʩݑ�8N��Z�>��  �ͷq����#"""�hƤ.����M��ۛ^=�؎՘+�ǳ`u�?�-�B�Z7f�#5�		r�h���4��� �Ä �m\���.�2��,��`�Z�����Iu46m�5�������CDD���A�{�i�3����*�P܌���۠��?�{(DS�4jԾ��-��.@��2��I5�v�PV���t�ㅙ�0���/+�'""���J]R'$ ��߃��fHU�6�s�h�j��B4E�~1����� ��q ���#;E���AY�竺=ې�Q��ݏQw���gBbW�gJ�����$�()�%i�����ꛤQ���#�����U4��`	�����I]�Z�y3>�������H�6F�6<U�W�y����6��Q�� P�w�3�[�� �a�ԕ�03�oECKǔ�7u����h����X��3Wd%��$�U��P���V�0[��kB��IΧ$�Ez$͉��B3�zM0�;Ө��ك�O���G�؁�Y}�rпk9�:6?�f4�t�� �9% Z:`�o�}��1���P����(�#'U��7�a8�i�n(5T� �T������R�π�]����Iա��է/OIn�vJ���Caf:*��(�L��A��I]�R'$������e$��b�����2a��j�!q�rV�$�؍ӈ��t�Q�|��4�q��}�^??ntK��J[`�1��[U;a�o��TI�03M�=��.�"�@W�F� �]��8V,q\��t�$/��b�����9�Iա�j�󮼐 U�_���-h�Daf:��lsܬ��.I�FyAJ�fKrq�� ��B3J�`ܽ	m�&�w�|��+�B�!$��bT�_����]��$�%yYh�ډE;O�d���1�p�ؚ<��_��B�]Q���B���)�����s~�m�&g���HҨQ��.˿CR�(ңzG)�zMh���o���AR%�rbR����p��e��Q��`�b�� ,6�J��/�"�����'��^�Ռ��x�I|��Ը��� ��+nt�>���:���˜�i��P�w����[��:��iҜx���L�<�ԫ��:	��s�*]����b�P߈���h�쁡����0�����fA����8Ū�+U�IS���ls\ؾ��(q�V���0l~ʭr"er'�o%�G0`�¸{�:{�>��ӗ/m~J��M8\+w�k~�><-J�$�U�W�����g����U��r$�6!�5�7:���F��)��5l~����`��*�^�S��*�����2�Z���|�#�%��(�����?�	]����ڂ�ؙ'&`��P��͎�+����^%vb��&�3�s����Gб�ȹ��5����h=�t�^��4���gO�	�J��=DI^�ǋ�����VSg���\����k�����f���:{P��%JL)�XP��Ǩh�pT�&�-h��ASg���sRu��v�y��1����vK��-I�vN��:��B3�o�qU�v�#BE�����b)��r;?��\q|��r{�����Ϸ���oEݞm0��$i����9��k
ڍ:�����^�O��o-��(�NH��?z	��7�@F��:����Yl6Xl6<��z}PbF#�+�l��TqgJ�H��wocw�_���6�fck*��=f��4���#p�J'֜T�E}��V���rR�n���z��
����sKĎ+�f/4;�r����V �zMn�[CKrR�S�����dm[E��9�q��b^��A��M0���V-��b��n������3��{1�}0[Q��ǎX{�IV}5�7b`Ă��U(������0[��TeMҨk7E�Ć&u�y�����������I_��yX���{�R��g���J��%vR����I��	�_b�K?F~َ��|���:bO���iHr�<����6���]mA��RwoBCK�V��X��<����C��R��e�����ݛд�nu�;J��ԕ�WjBr��Q�di�#����B3��ls�w���>V�_�;'ޙX�y�?0b�m�p�w0[a�Ќ�T�֯���j�5���0��PV�ܣS*7�a(+F�ي�3W��h)/�s~O�|�B\C� n�;oX	�_��I����Q	��N&�$�I�:*ۓ�/���(_����Hä� 8���j���~�0��+I�q��	&�
<��V�$$ub%���+�kb���5���Q/A�`�xu�t�l5ቶiH�;J���O�i��tęr���	�/��W����3WP^���-�><-�U��T �)�U�v$)��-q0�7��܀�*��.W-�u|�;���*li"�6�7����/4;�f��%VBYx��VT}x�ys	�d7w��\AҜx�t�����K�r�|��g�8���,�ñ�I���ZQ��<�B(܌��j'>����r \$�z�$�3��wl�j̍~�mƥ�%l-7��h���=Q�����0n�#&�Q���	�����{�3u%�=v�44#��[̔�(�FG���#K��ێ�1K��v/X���&i�h{mϔ��+�d��<%u{�9�	�֯Dݵ[nI�q�&$͉w�o�".�m���ׄ�w?F���:���H�`�-�3���>(���C��{��J�4'^�q�$'U7�1�	[P��3j��A����_�
	^�>/�r/l{!��TF,S���3.0��Y�~%��e=�� |�#4u��|6���,�+u�F���5�{��܌k�|Z�s���N�d�f�æV���ǲ?�C�Nn�>���1Y�&<�J��S\MW�4�����d`�"ZBmӐ�F0u{�9���0��n�6g�W9)Z�,�FI^�dӢB�1n����dO8Z:B�
�{������ӽ.�_�lǏ��P����*ؘԑGz=2~�:���q���	�qq�%%�n�atx��a�'<_H��혰�a�c:[|<����d�ȅ�{�T�gm�-���<�8����g�8�)��t��>ga�]�$_DDN����/����S��e�����`�b��4�S������9|s�"�{�C��F������v�Y,Ǹ��ݎ���1O��%6bޢEr�I�R����bb�������_��g}�߿/P+��C51Ԙ�΃�l���-�Y���ʊ�����$R�]7[�Nh�`Jw8��G�4$O�w0M6\�1���(Zp�exj�#���{cc�]|����LR������ہ�۝�u7O�뜺hQH�7�]˳�����s������ΰL�����q�g��{}&��[�M�x	ӳ�O��ݙ�����~��;�q=6�u]�S^���M������R�]7ݴ�$�ڹg��Y�S��q�X��|%U����g��d��w#�N�F~Fηv-f��'��z)��ԑ�ع2��$�Ŝ9j|��9ѹ�g��3l6qo8���0G��Wmw<�������fO��!n�(/ȃa�S���"6��tp�:�.@s�}��|+�!/?#�+� ���j/ݐ<f��'��z)���E����P�Th���x��=��B9?]U����F��U��u�~q��2�&���q��Ձ��w]!6/_��Wc߱��� q]ﾇ���b�'p���o�-y�q��E<��2<�jYT�'�ߋ�[ס��)��kr3 &�U�}]�3�P�w;��q3>��ɋ8x�d㐋R����j��s�O����R�".���_$�E%yYh���l�!eB8����$��q���|k'v�s��B�B��lE͹&�w� ���ηv:�h8O\���Z�G�6����gp���{�9g�'o:aL���:"�($T�=ڂ��J���|�ś�w�I|k���E�yM�7?#mJU�sּQ+I���ϭZ6��-���Lꈈ�����FU�WN��^�y�h�ϸ�$u{� ���,Gv�Źp�s�^
��q-�I4}/jvn��XVr�dSm���2}�պH��ʤ��H&����=�$�;0b	�F�MXrRuAm�ϸ���������}?**�b�êJ���-�[�,jΓh�^�۸��y���Bo�-z����A��8�uݴ�9��m�7��7T0�#�r�� !�}Ͼ�ix0<����q A��i2{�Ed\Wf�Ǥj��DW��+�����\�578��uT#��L���;�F��V-CG�P�.z��<����i��dRMì9ׄ-�\�.��A�h�V� &uDQ����T*��
T*�����װXş��so��I��TJ�`�"\��+H1�]����T	N �����T�����ͷe	y���,xU�h;O���z�v9���0+?8���2��ȩ��F�I]��Y>���Gg��y�wa�\uF]������סP��P�����4�Q��~�l�	���i��$g>z�� ��>���mbv�j�������Nː+n�JҨQ��9�:�TA�F��Mn�ih�@��Ge!�3��q��ͬ���nv�:�:(��z�D��n��d��|\����4�H�v)`RDm�Ch���;��G֜�ٟH>��l�|g@�a����<����<���;���6H Q    IDAT,$͉��}2I����-�v�LҨQ�g�c��ӗ�~f�oD[� rR�Ά*rOդ�s�l6/_��Ϡ��e5�=$����{hl������k{���W�'�v�8y���?�_ock��鏮-��w���Ps�	�cZ��#�:""��`ܽɹI���R��}Թ��� ��O!'U'�vEz����	����J�f�di6�:����N���e�;�1��j>B�>����?(y�h;O�����|4�~t���h����D��:""S��0[QQ�w$y~����(ң��G��K�f��f��0n���t���)z��F�EU$�on�4�h;O���F���PŤ��H���>}�Y6��۳%yY�>sE�΅I���n�lE��+n���"I�F�F͆)�N�bתe0����|#���������o��cDD<L�\\\�^4	�%8���&$Jm.SO�d�03]�ꜧ1L69��9&t��N�:[|?���X�F�,����jl""
&u!*F��J5}�>�(�ʐH�
EP^/Q��>}Y��j*���>�$/K�M�#���N$��ߢ��-ؼ|1��fmz����i��1Q�aR���P��������oJg6��9o|�	��A$�6��@ݵ[�*]��������T�_��<T�����&׺�a��ŲĖ�)ɇI]����\�+}��K]}���F��0�o�Z�aE��^�O_���%yY0^hv&�9)ZG�ˇ���y3�=���  K��L��A�(�tDD�I]���i�_���AsHT���j�JT�_9�c��FѧdV�����AT�a(+v�Y[�	��Fne �5���JN��An� ��\���D�]�����:"� 0[=�U�����-��ڂ�T�s���^��Id��f%��?�ڿ���IQDbRGD$���#^=/'U��i;ö����k�4F��i�(�]�����O��HCVr"���s]E�.���řIQ*/�C��%�f%\���3�  �]�"�u/l�MD��03Ezf�;g�q�zM����K��E��<wo���-0�7�M�2�ބ��[R}��w�֯DE�9��o�s�ٱF��n���S��L&��i{m��}�\5u�x]� 
G����d.'U��^���p�]�Q��w�àe{�9���^���Y{�#��uO@�Q56E'9���"=�w�:f��N9~I^e�(/ȋ��I&u��̕)�f�ø{��lC�ύS�����^�=�۳9)ZN|���P��U;QR}d�4.o�9��۟�^ۃ�^SD~�&�Z���qpL�du.���V�;�	n}�6���֮�%u}����)YbQ��+��(�;�a�a+���,��ن��+#�bǤ.J4u����T�(u|��8�K�P����O�]l
���v::�M��}�$/�Q�+�C�F�'͉w��Ä.��^���K7�.6E9��$�������M�=H�p�Pä.��8Od��<M�l��Aҟ����#�"I5��ls�l9}u�n9+ܳMY&""
Ur%Wf+�Vf��xS4I�v4 ���L�HN� ���p��Q�++FN�M�=0^hs�DQ������>IDDaN���x�U�W"'E����M�f^����K�ύ4L�DyA*����������﹖��VT��1eŨ(� �w����-�>}��<��M��.f딵tD�"��FE��y��Q
CY1�Qؓ+�2�7b`����Փ��-0��4"�8`R��֯D���S��D��QJSg��>�$�U����Q;�U�Q���)���g��0^hFaf:J�]e�VʊQw���QX�3��>s�g� 'U��usĂ�Ξo�"i���1��@��/sRu0�ބ$�zʖ�0[�1�><�ܾ�zG);V�������H�Ҡ�H���+��ك�w?���DD6�M����t�������$��?���+80��p���?,Gݞm+iު۳����LV���l��w?"ѳ�O��ݙυ{��ۯ�7w7Hꮶ��j��
^^����t&uDDv�K�b]3&i�0��03U��x̊"��Y$΂aR烵smXk��ܤ���VǨ#�N[�ɱ��mU�n�;۰{��!̝fBRRt��Q᫶;~�����f�˸20[�w:���7��]1f�U��B�_V�m�%$|Ez4�t����y��I��~�j��Z�q�Q�R���������!��KN��U�(EN����MҨ���P��Q��N����*F���>���	���䬘U���hܷ��ݛ`��r$q�W:�Y�E"&u^���~�slԺD�q����Ά&��#���%�F���Z���	8���T��圮�%��2s�����7w{�S(����|#w�L��4�;�W�zM(�(Z:D�j��yA�T�(��Qw�I���''P�~<ܲ�[�N	d��: """
?rW�\��������C��l&uDDDDDDޒ�b�:�L�V�(u&���� �oq���*fR��Q���h��A�ύ0^hƀي�w?v.Aj�ډ�"�dc�+uDQ���Hиw|�^���C�0.�$�3a C}�ǥ?���)��;J1`�F�>u��E��{C�J9���:(X�	s������&G�l�lE��Gg�� L��ԭ�X�#�R�{�`��ݮ��9K-D�o;��H���df+�O_�r�iܽ	%K��4+/�CE�%yY��ꮶ����.Ԯ�_�~�[�jO\�XW�(����(�c��U;a�oDCK�v:��=����F4u��j�JT���������nݼ���
�I����ԡ;'U���?���᪢H��<Y����b&��+��BҜx��MҨ��Q�/�0�#�R�rL�;U���h���PyA��BN�n�}d�d�P��h��m��9m#����^���i��䡩�Ǒ$�T�0�����6>O���7��{
�M�=HҨQ򰃢�di6�V��e�%u���h�5����L��MN��W,���q�¾�Ez��&��\���i�#T�f��૜T��>��(���sw��E��K��/����dUw�����H�r%(�LwV�\-�B���U���0-�P��hn�R��P��&A4��9�:�䡡�f���"�����)�7&'����4կ� o��#�g����-��܎���&7s�sv=��1�����%i��
�l���&W�;J���s��p͞��>���
�4�H�ހ�:""""��]mA�槜2O*��h�왶�2y/Z	chh�pTU&W�Z��2�q�a���,�v&�B�Vw�e��?�ꐓ�CÉOݎ��ҁ�<f�;�ϭ>s�y��wor����Kv��{�C (�<�j[�p�\�[ ϯz��O��b��Z'���t�i�m�&��ن�=�7$�OnL�"Шz4#�݇e"&V���sS��>�jb,�q������3c��$/u�nI:�
&L��vE�Y��Φ�H��؅����4n��U�
3��p��m�eCKJ�]�Uw��m
f��%�W�������2%U�|1��q8x�"���]O.��Gq��.��e�}��g�CG�Z��x>Ea�\[ߠ�1�.�L���+&uD��e�x��$���ĳ�p;� ��w^�,���EX���Ci�j\""�ʹ�+�C�^O����zf�_�ufBu��f;�֯DyA^@S���{la_�~%�֯t{��j�]�Ȧ�geM�
UɆ�gϵ7YCK��rVq��®���Qs�	 P{�j/����L�]W���;�]���'��|�Y�Z�b�W	��B�䛁W���	���(b}���˪N���A��;/��  ���������5.���K|��t�,y��r6Ez���9s�ʖ7rRuHҨ=&��L��Օ�e�-E����}����n��L7ƺ�-0l~
���0[��2��j��
�d�[;q�uj���}'�㍀`��}m��<�s��E2&uDL�krB����`$vL�HJ9)Zgh�!L1�JI^rRu�H�Mi,�4'~��,ꮶ�03I��4N�6�9���칾�%���.���S �����E8���:��ΔXI��1�#")��9�|�0M�x�ٱmA�S!gC[�	�~����f��$5m������kKա���?{��s����j�w�pt��$����*iN���n�ȑ�y����1a��H�����r !!a,!!!V��^zD?2fW���#���?|D�1�;����7��N�fK褊�Mb%EbǄ���TQ�G���0^h������C}#��7�:3�9m1'U��Ι��~_LO׈E��:��K@M;����w���vT��������E�>e�	d���������P(Rl6[�7�x�b���h4���[
 q
;  �_(�a�4h4J ��Ð���x��i�YG:Ψz�\V����N���n闟�������ݛ���g�J��B�W	S��+h�t44��9���2eSs_�����U.��l��p�d��:]zJRZ:`(+�j�_ݵ[���t
3�e�|���G�
�X[z�+�O���6��^�����INN����Wm�
7�Lꈈ�䒤Q��/+P��Ѩ���E��N�JK�3���,��r%"""��!l�0ymI��������������I:Ez��):peE��{
�f&tQ��:"""""�0�JQ��N�";Y+�0�����z�=�"l�s&uDDQ,?#�{�C'�P�������>�j>���.f��#J�|�0Fu:�l�)���f��A�j_������>cn]��#���hX�#�pm��A[�i����T�sASg�c�Ym�+��(/�s�Z����f��n���z0`����e��'i�0��mJ[w��������&��z�8+uDDU���c߱�rCTLꈢ��x5�t���/��S���0��03�~�|�𸡾�ou>nܽ	�ݛP�QO�e�o��
��Iա��� ��=� 8:�5u� 'U��M��a9J��` ��F�������Z��#"���5uD�rRu��Q���� ��\AҜxT�_��k�����U0^h���U��1�2�Q�~�W퓫�\AyA��P��i��03U�FSg ���C}#��l��A��7���A��ADDD~bRGe�֯D�F��ӗ=�|��I5�4j�z^�Zx��>�o�5�03��騻ڂ$����:�4'ާcE#&uDQ�$/f+Z:<�|�l������-(��Bݞmh��P�,'U���Y��03 �������LꈢLҜx�X|���<����F)��b���&)3%h���z�I��xEz������IDDD��Ѭ�VG�w?vLߜ��Y�~�Ǧ(��bʊ����T�3�ބ�Tݔ�~DDDD��:�(30b	h�����Q^��槜�T\;UΖ�yb(+FyA�����?"""�h'߮�D$��k���Q��77YyA�s����+1�7?r�ss;��/4;��4;�qwoB����x�c�}��hfLꈢL���0[QU����'o.4T)/���|��I��v��S�����?@��l�TaBGDDD�#N�$�2f+�><���{�6��SeŨZ�-Ω�M�=�>sŹ����9Ͳj�JT���EN�ι�x��G9咢Nv���Zd�$�m �67�c�\�e2[q��>���k_A�F���4�g̃N����A|��=9��u��:�(Tw�%�&GW���xSg��'��h�5�� m��q>����H��RYQ�G�F�8��8\�Y���~�(�g��L�ks3�� ����_��`ڟ5�v�\k'�o�z�=��*�F�|���f"+9q��)���i�2��8w��[�"�=��������BZF���'��t�,š�Өa��#��_]����4Ծ�Yɉhl�¾cgq��ޔ�w��d�bד˰c������w���[��6>o�k¾cg �6���uO  j/}�|�u���~��'/N;v�F��[��U���?�'/8��؂����®w��z�=d�hQ��)�O�Z�)X��~#b�J��V�|���������O�?��R�@���_��ɏ��DRQ��Ԕ(��3r !!�k�N�P���~�t7�r�(�}�5j�,r{lB��X�bUP)��o�u|jK+���bhb|O[>~���H��u�(��Κ��k�2���V�w�ηvJCj��\�-�\l^�X��w������5Ed�L���[׹%X�V-Á��ܞ����q����P�q�����p�'/�%э�](�����E�s���7p��E\��
�c<y��oLy|�����}�+�q{|��  ��������_!?c�Ǳ��c���n�����7��s��9��"��o���-n�TG���δ�����
���a��_���]n1�q�o~�L<;�����Y�7G��e���/)f��X�#""�'����p{,sI.�sf��x-!6�w����o&�P�%�ZŐ�6>ϭZ6�z�t5*�b�'$KxYɉxqm!^\[����8|x���ӨQ�s��=��������Q:n�L>W�s`Mn��&;y�X�1m�|k��Ǘdz��c ���X� ��؅�ɳ�G�5��Sn���k���@JB<�-��X,w^*�O��ޫ(Ê�#��>&uDD��AF|U� ������^��B��~��I�t��q��8��i���9�$�8f�d�}�<~v�o,
�ؕ0��d�����p������xs딤�d��d�N���*�k�s���8�ډA˨������?5q9���qJ�[���}�㞎8�E��V�c��}oʴda<��p�鷍�]n�����Z&�6�}J��쭎)cl�?�-��)�g'k����޹�N�tR")��lْ�P(*�@\\�)>>>I����}� �-�r�HU�W�_��?�el���}�G�M�&���%A�Pa|�
�Ō����A��>� �`��c�{�F�W���f�~�v<S����Á:F�?xl!��q�����_�!p$��/�������O��{�!��dMn&�� u�
:���B�~��wܞ�x���"I�ƪ��`�2��?:�������7���Y�����͆�w7���|k6<��F���.�?E��.}������څ�N�gh���X�$�[����;�L����:ׄ�'/:�ҝ�:}׻ﻍ���˨�|�ۿ�8�K���;�S����|�|kηv��>��-:�����_��?���������9�������}/t=C#h�@Y�b(
��@�q���.����Y�P(�34�m_�F�5�*�����q��&H)Z���t�����?����#.��Q��:�dU�W�PV��fﮞH�\gw{,1)���n�����I�Z@��a^�b�'L��;_��2�r�G��	SߤZ&���F�S�5w��HC���g̓%�7��%����۸zʚ2!i���63!�6g����MY;(�ף��5uDDRF'�KY�R��Xb����p��-$ν���ˠP�_��K~F��n�m��/6/_��?y�GN����D$�.��Wv��MGX��ӨQ{�\��ų���n��4�pg2[�$k�SovonŮ'���U� ޻�?+7'""�R�e#!1s��	 �զaђ����t\�R1���8�Ņ~b#�]O.ùW���N����{e�ٹa�'� ;E���
��N �G'u^�Cv���݀��Dh�����B���x�e��[皘 ������>���.��5���m�s���L�$
+uDD䗌��ߊo:�����FO����ڧ���V-s�W�dS����n�͋k����uʪ��[��(��ȹ���}�κ}>�nj��]�ۏPhb�����6���`6[1<t�c#r'(�=��3���O^�8],P�k�^EY�&t�����r��v�R��HCv��c2y<D����<u����'��X�#"��d-�.���u�:t����=$�H��]���e�}��kr8��J񼷗?��q�߻e�?�uk��!�{d2[q�ս5���,L�B�-�    IDAT�Q#?c�3�DM���P_�]Ҫ�������{���P޿|��9�2��^���������?CaSw6�!10�#""�`||f`�L`��M����3f(�\[(j�r���o��ý������5��آ_�2�d�J��N�.�׻��K7P����_�b�G��y�ٹ��9�f�k�2�=՞[�Ǜo#��oI��Wy�*�����\���Jvq�ܺ��s"0�#""�%$$  t:Gu�61�ί?C�|xL�l���mA����8 B���A�^���.}�S�⪣�_���/߀6>{�=�]��T�4��iԨ��.�vR�G��|{������qp�:Iײy�0�g��N�$���4����I�F������jo¼�Q�5)��a���m `��)F�)ڀ�E����ɋ�iWb����ɋ8x�"^\[��W�=�0�Į�bK�	����[��ֹ&<�j�o\�wr���B�k�,�:�b���'l*��1k'u�l���}�7<������{���%v\cG�bRGDDS(Uq��O��wU1j<�Y�{�����;�Q١��nj������lE͹&<yQ�QM�hm����k�:�?�]��nS}e2[q��E�6�Ry��c*��uO���B��X��=�6(�i�صj��sq�������w�\��qn]���f߱����t�cp$%�T,'�^{��hS�3�ܶ��vL3Y�����
g�B\�o��A�(j/}���8���#�pp�:d%'���7�wg?þ���{�*|��%""�hS�C��sal\<2�W  ���a}��v&�h�e��B��������~O!�Ǡe������V�<�����6>5;7x�$Ц(�ͭ�<r
��Q���+��y���[|�lj��pp�:���ܺ���.���oL����in窘�b���~}&�^1�x�mQ*�:�:��	�����	{���O^D͹&����7�:߇5��h|e��gϯzܯs���4 "� ��b�͏<�W����q�����ohԌ���qv��C��6%���KG�Qc�������K7������йjl�7j���Ϙ�ڊ-3>'��1B��yc}P:W��]���;~U�6/��)�a$l�1�����E�L*���+�� �۸�����"d�:��zq�I����J��0��Q���z��;��>�l������ߙ�L��G��;�T�o\�״�}��e*�l-��R�+~vv=�{� t��4�mד��n��7�]��hvٚ@.��Q���{}�?�u�(��k��Jr�E��W����bo��Ϙ�׺T]|�$�������3WP}�J���f��ɉ��I]��N��E?֥U9%z��@������ZC�1�c���~��z�=��(�!�;��.���f%'bד�^����'8���?G���x�m�+�bp������o8��:�2;E�5�����=V��Y�z�\�۱�����:""�Iv�q���ҍ�K�B����Pvx׻�!?#�{��U�ńN0h�.�q�Wn�ij���E~'ukr3�������T��P�,����uX�F�,�����޴9��m�;vv�ϡ�o�}�f&kr3Q�s��ݞ�˺T���nKͯ�&wLf+�:�aMnfT�8��#""�d�'|z���N�� �7>x�_	�p�*l�i	����>�إ4+9ѯ�ukr3q���۸�6��?���z�x5Á>c��]Z�Ө�ݢd�����^�[;��Z�S���߇�(�[;q��E�X�����v�|�_�ŵuaH��F9�2�#""r���e>%.Bӏp���S~��g�õ���k/:���[ס�r�����1<����)����^qͤi{��8����f�9���Em[�y�~����_7=Lf+�j>�ؽ����)Z�)���8���[o�|��H�����c���ɋ�u��G�SA[�c2[E�н�p{	O����q:�&蛗/�����]+�pv��gn����I���ǣ�S�����y�K��S�6Q	Or$vLꈈ��i�3n<<Y{�`Ht��Še�GNy����f��e�C>_���?g ��������>�o�t�pt��k��E��!f�)����yڭ'&��c���V-�Zw��ޔ��q:��<���1�#""zhMn�O��bP���%�2���ِض�N^����VwMf+�s��yc=�7�c���'١�Se���uAٻ�S�x������K7<V�}�Z[V��������N�&�n��`&vLꈈ�Z����}�!���'>���)�P�ꍎ�!���r3`ד���k{���#ܺ.��� BE�}����D��)��L�;e-ݠeT�
��)� ����{��&�O^Ĺ[�x~�㨯��J&I#X��:""��|�8��<�����s&�}����{>�/��8���4j�=鲒��F}s+NL�����P�N��n��7��^!��p3#+9ѧ�)e�\غιf�����7�!q#�cRGDD��/�߻�#	�}�>�qJ���n�''>�������OIK�6¨<2�<�n�1x�as\�u�&�����Og����2��Rh�:����DDD�|�=���A�׋��n�&����Lh����۞�^���֮���7�M~F��]=Ϸvz=�-;y�J���Nt��mV}��-"��lŁ��.�/���XG�醍��Wx�xs�xޜO7�K��{��a���*�>6�:"""������rm��E���7����h����ـ*%�u��V��͹W���g����+Q8���uR�671��]���﯆.^�s7��V5皰E��b�*������ۢ�5�tS��H��4��S����8�p��/o�k
�6$$=�;N�$""��)Oӹ�g�N���ߓ�/��r���ـ�]J���{l).�u5�u����Vv6�c��+)�����K٠��/�}+��@V�܈M��)�e(�I1�I|����w���x�N�ӹ����M#�2}.�W>�}W���u�����"B{���je0�����J]�ߚ���sq��]���lG�{Q�&2$�;&uDDD>2Y"sO����~U0"uj�/�G�ur�ٻ������y�X����5�b�]�I��k=}�&o�0��[�9G'i�����:"""r�Te����Q��Gܧac�P6�&�/�y)����1�#"""')׶E�Ó��5�vEl��W׻��I�X{�I�EJ���N�׏"���:"""��s��\�ʛ���ͭX�s#�����BY�GAY�8p�":�ݛ��1��S%y�[����]��8��m4�v���7�T2)���qK"""�g���������� �"l��c�_��&7��/��0�{����u�ZG�д��}o�Y''�J~F��s�Ө�����-&3���<r
�+�q>&��uR���[�0Y��o���F�] �0�#""�o��z��Г��V����Zq��zr�߿_�s���������4j|�ڞ���_�z�����WQ��󾍫a2[�*a����N���66/_�|,н���F�씩7|i��Өq�'/8�4��������E	;N�$""�o�n"m��6>5�6�M�Qc������ƛ�F�^_��y�`&;yj��E����|�V9�vs н��F)v�.X�a��/۠T�-t떩Ϙ�]����B�ǟ��Lꈈ� �6���H�Ey(�ٹA��ʵ�(�db�2��ٟ���^T�<%��C�r+'�ي}�>q{,н�<M���ٻ���;��H���e!"8�Xp�d0�f�T�2"����=A�dfrj5�����`������cMrƐ��(g-r	V0Nl.��E�`ld���ڒ��R_��;�����[?���r�~��<�H����<�'Q�wK�_P!ъ6��  �"�bf�y�g������+�,��mј�#X+y������ӽ:`Ц��X�t��e,�^D���'��x��We4��Eya���F�;9c���P�/��h�� �+����;k�~�"��Ƶz���*��灻�g*<r��:?ҭ	��P�7��;^xY�O�;��������|v��dT��<sf<{�S,����7|�p�$;�����=�Ԗh��Ǵ��c������"v�:  �8�L3O5�)+�k��BvݺV�xP^F�v�yh������*~�a=s�����zC>�Gό*���3򔌑:i*ܼ��3�źw�ۧυ����|5��=q����w�=֕�ЁǶ�ÿo�-�Wh��"
v�:  ����}�����0Wm���Ѝ��<pg�ih�Z��f�7��ĝ_��o�ᕤ'f��3 X�蝹f+/#ݐѺ���z��>l����9k=Z�{ׅWO���
��.p"M}mF3���c�C�?��zC����p�`G� ���'��ւ���I^F�<�=��N��h��%���myံ��i�?[^8`�3�����Ϳ�k̺�x��4'�>�A�g�q�'"�jj��oה��4�y��9}oe͠ue+�Nen�<�(�����k�`G� `�h@�����*��{]o���L�ڞ0&�u:���sa�9=m�C�Dx{�F�9����!��}�v����F�֕��3�6�,�軤����/��3��̙��W<#b���ٜ�	=3�0N$fO5�kK�|��P �4m�����i�� /}垘*]:��ㅗc�s]�
Â]����Q.	�f����HK���~L���-}�7�nH���_?6�㼌th�mT6���j�H��_?�����;��>o\S�[W�b�F��=�ˣQk���hb��hԡ�C�`G� `��_?���n]kȺ�D��;j�+��x��ԉ�K��r0����6W��z^�륦k�<=�n��~����������״��A��������"��W��{oW�_�3���N��hǈ�3gf��ٵ�`��޸Vo?�+������S���#�{�o��b!�5Uj��%=���k���*������I��
��l۷o��X,�jPzz�HFFFA�������1����n 9�ׯGn�|T?`�}ӵ:;�S�a1xx�Z5��ӵO���P�ק�O�j�>'���}�����7]�W?�X�/��$JMY�~��;��f�꺽o��_��l���u�Z=��u��Ks�tq����>�=��>�{n�TinV��nS}M������ڕ�.-TEQ��33��ժ���#�~^�޻I����-U�s>�=C���r0��ݖ����{'㪜�=�ԵEya���F�/�^V��3�uin�vݺV�k��۔�f׈�#�קue+t뵫����ڻs���s׆�{��ׯ/���G�W[�����>���<U�j׭kuནQ��a��H��?��:���Gkt�z �L<��Q����c�o�lІ�Fx�+��<B���:0k�ቾKz�翉�o�?���~�E~k�Jb��tOD5N~��g�[�f��Q��Wն�Ks���e������z=��=�]�.������R}MUܣ�������k�J�|T:��U��ը�jK��Q�o�>�/,WF�~	 @8�=��}ݳ(�h��H�+�9�;�z��Ԟ�V�+[���_ZU�btRl�fk��̜j�oP#좩�:�ξ~տ�ꢙh�4Li��x����%�k��:�I
{~���|X��a�%�<�_�Չ�~}m���Hm��REa��>����5e%:��v�}ӵ1]����O��;�j2����nԺ���gS�Go\���ᾘ]g_����1�~����L��ghT�>���rm��ڶQEyq<�קW;>�ۧ{U��PuiaT���������z��.�^��FO�:uqHwT�Ϩ����麇����;��y�1W���?����~,��-U����Θ2��{'����bj�/˾}��V�T5 ;;�l~~~l�u�<��N�R� &�̽���*SS�JjY�x�+MM����bL�,9#.����[I������g�rS�{�9�	�j��%m�6���;�~���Ж�r�++�-�W���y���:���^C�_EQ�*
��N�]ZS8�SQ��'�U}M՜"1�t����̙��-U�:��v�e�����W���[,��0B�<B�x��a;Z�=��_?jHI��l�Z�}_�'�}�b	,�M�g�ߊV��SϿ~,��Έ>z��o��C|$����3>v�'T���'�YXغ�Z��dF(
��x�xlFp�պ���|?�B)  \Ů��z��]��>������h��I�t�C�����z����W�-���
sD��(O��G��{�^:ܡ��ް�N��V��{o���^~�d�]8��> S�e�1��oI��� A��a�c����k�D�%�u�����1��U����J�7_רS�S
������v��ۧ�E=ʹ�0�J���1������^��{5��,d׭kC���	}󧇴��
U�{ȩg~�֢�����+[��L�N�]ҁ��3F�������P�%�P\�#�tך?�������望�R�����ŢQϤʬ�����������d��D�����=8��!��]�᪢0O��)?ӡue%q�6�f���L��<pgB�v:������#ij{�[V�PEa��T�6$��R�>V�uh'�.i�C��X����5}���=���?���z��	�0�/$��;!��`���4����nB��Z���2?}l�IW_��5.�<�H�J�sT�]���옟c�Xd�X�i��б��9���co{2�軤��^5<�m�*��pF�����vEy�(��at"%3�IS�58�rv�x�u"u*��f/��H����v�?��g��7�r��ict��H֬r���d�Ŀ����gҫ4�'�j�ߍ����?�G��0��A��x=��H�O�����jo|(�s;�]T]�+j}�A�U�QS�5���
2jo|HY�k~E]����}���˞�#) �,�H�W�#�u~�1�R%Q�.�^��v��FB���W�����bڠ|1y���)A��SL��(O��{�*
��o��>�k�����:�w)l��p�G5��U�r�������{����g���{���W,�=c���@@���# O�P��b�U@u��'�-�: 0������oPS�fu����S=3^o����,�W�Oތ9Ѕ��9tV�.�QFf��)�)�[|ۦՋI0�xl�)<���pGB�q�ݓ:��o�>2r;�X=���{Be���[j���Pn�Z��¼�7�Gb�^���7���?c�����ڦIϰ���~`O�UzF�����R�q���X���5�c��O���O�z�Ԝ��7�q��?���"�=[�O;�W���u�����KW���-�/<��EO�-ȵ�,�@�EJȲ3B �Hǹ�*���f~��Ӱ�35J�s���7�����k�[7��z��O���h�!m�Xm��3%I%�*��9tV}���▘��L\Y�d:�wI[^80���b��ׯݯ���}��}4{m�b�!���t�����Ӫ��im�*׉�KZW�bN@���\{tL�n]Z���]j�y����e�k�w�~߫�փ���K��&<����I��ǆ���#�4��{2d:����g���뫵c}�Z�ר�'o��~��j�'�%C ���,����j������%5�>���b�6�u `2-G;UW�F;�W�y�65��MՖ���~��F����yNN���^5�xኛ�;ߩ�K��h�u�<ˬ���w�Q���3��YО׏�dDg��Ѯ�U_S�=ܹ�G�9%5o_�������ۣ=ܩ�����-e+B����:�}�o����GN�jW��9Ӳ��{�Zo�
�W����5��jxxX��.�ᰫxE���	oC0�u���h�%�[7�q�F5l���x�`�t�����n'�k9 ������l��F_x�EO�mͳ[�,ғF�S"��)�\æ�?���͡���fW|�Z]�=���ߑ=-]EJw��n��bY>�)����ۧ{��;ݨ�����K��gm�����s�}G�����j=b������E0:���A�^~�d���=��yL��~x�ywG���،-&��	�{n�F\�P��ٕ�?|����Ј�3c����B�XW�B������p�{|�����*=q% �t�#������d�    IDATu�Z=���q{��/��F����v�QU>���!g�k>?ӡ�wԆ��{��A�=����O]��������Lӛ�Vk�Ƶ:r�wƿ/����S�?]o���3U�����\Ymv�9/�\��UPP���jY,���,;�W��zMh}�l͇ޟ�~�?�Pæ��3[��T�Ԛ����>�:��.�)c�V_|j�)5�|co�U��w�&��	�<jz�jy�>�>����o����%��b���Z��z䛼�1���̑�jU 0w���D�%��{U�n]�g�ݔ���>:������,#.���~L�wLMI��Ji�s�'��[�jM��W��Kou��;qy�tO��G�{B�5��XÕ����w�N��N�vb������{u�T��U�umQ��T�Y����_dL/��j�F\�}t&��	�軤k��gs�jm��SI�s���ܢue+f��RU�-/P���Ϩ$���\�ۯ�wԆ�o����ޫV+?ӡ]���V� �1����{�O�5��j{�Ka�W޲z�v��S-�`�
K箅��[������wy�Z���Ӧ���z���{~�8I�����ڱ�zN�kj;��G��23���w��uz�᫟��~�5�[{��~k{��.��� ��h=~*���k`DMmG�ކ��J]�N�I��^�vISB�=�_O����7̎��=���;�[�s�v�?���t���=�_{^?��~��?~C����]Љ�Kz����tʗ��`��/�����go71=��>o�u|��V�	��k�TQ�7��#��ծ0[\l�Z�-aF�wm\��53�`�e���0O�gmi����ue+tǬ���j]ي9[`��^�k>�aij�qKUy(�Mn�鰇�|^v������E8�7�5���]�=�Iψ�3.j�K�50r�"&�~"Ia��I
��;�ھ�B��������}��k������� ��*��UwcE����	M��e������}���'C0�m��ӄN�
�GZ�T���k�+o�|�e��#w��)Q/�Ow���=�I���1m����m�茜�ۇ��u8�����>����u|�J��3��{/���+����<a��=�Ԉ;�}f�]��.�uI���z��M�}��՞׏���j����[uy삡�-�t� ӡ��]�Ѱˣ����V�B`����eFH#�G2]���>�ᗿ!�{0� L��������Tæ�P��. ��Z��e~}�{R�%��ͻ&imX��>}nj-�+o���JwTMM�="���Q�軤{/��ӽ�v4.Z�~���#�u��aG�"�tO�����a�%�u�IZ��T������-/���u�	��[%L}���g��qy�ďߘq<�����;Bk�z�FC�ئ�������{d��C#d�}����ȭ��}8r�W�=���33�����I�軤�_?�-U塯���P��S��r�x�==��7B#fӧ�N�{�k�v�릿�g~�������N=�ũ_���/���J��^�k1���U$�?���)+w��3c�w*��ڎ��z��nP��݆O�����y�.Co��~�5�/�k�B �PS�fՖ������t��M5j�����%�~�?��m��Hekn��s�9��V��V�#[nט|^��F�~���p%�}��� ו���Iq��3�O��m�EX*�jN�]҉�K3ʾ�*�_���<:����S��{�vzi[�i�{�\hs�`_x���:τ=���^U��8�����K�;TQ�7�ks�+o��׏�9^��U�+[!I3B���9>��h��������R�=�{n��\)|�'�.����{|�s��~�O����zo�{ZJ�N��is���3���SZUPF����;��L���݄}���B�4��)���O��f셧Z�a��^S�����:B �L�7�]#�@��YW�&T9,�i9Z]�Qc�^��=!ɮ@�+�-���IҤU�u�O�ե�C������42�*#.Oد���wΝ����FL�;>�ߍh�'��.��ْ����K��>�Ν�@��(�`�q��ר��t��\Fp�ѷ���z�ڱ�Z�[7�ն�<���@��ŧ�O�m�X�����5u `"�������4�o�w=B2X,6��W���MZ��Z�y9r��]y�*i�my  fc��U~�t�����+��5֫��Sr|����l�E���;��`�Y	�׆G��x�Oޜ*f���@@?OŴ��F_x�%��)�: 0����?�@��Ȝ�d���Q��g�TKs�++�L9y�dO�Qzf�` H���1]g�ٵb�M��s]�kt�3y'���M\��i�[Ԗ����9�k�[7���!U�ݣ.�a�'��ymyiT�	�o��}�D{�/�$�nm��F6[pyp��|�E�b��]�:#�$t/�ͦ�K��
 �Q^����^���Y�Z]�^�44����S�P_��}v��gj}�����WN_'���������F��9uk�f�Z�-i~kTSu ��4��w���C�G�bY4��e�Q8s���>Y'G��d���2r�W^�_���r����'$���� �����ʟ��V����r��S�K���l�Z��R��oC��?Sæ�9A���)�~�ID�.gk��k����y�uF$���/6���>Ց��G�)�B� 蛿����v  ���Pqh��O�d���ҭ�Ϻ�d�ov�+���ۡ��٣���W��Ψ�y-��Nijf��A��'P���J���e���N�   ��o�98��')i�Y����T�a�@@B  @d�wnU�j9ک��|Ֆ�������8w1��A��P�  ,k�?yS��^h�W�7�*�P��Ў�Ւ����k��Eiܻ��_F;zH�  �Gp�dI���"�R� �l�:  "P����?}]���uu}���T燞o�nij�)x?D�����H]æ����Xܲ�Muf���uQ���f  ��L_s5}J��a�G]#j�߬���<�n �A�  ��~�g��f�~�G���
���T7�T�O��q�F�%*�Q�d�X�=$� p�奪-/���~Iu�kTY�0�`�z KK�*),���t�4  �*��r��O���Eu�����R5l�YpS\�K��g|<}ۂ��fǹ�Qm���P����������!� �G��5顏�'s4�cW��snN K9ʊ�A�F=�*��:q��y$��%Ip=]p���������M5j޹M�z��vD�;��F�Z��RÏ~1�܆M5��;�]T��筴���y�R�^k9�*�_W�F��?8����FT����q�5l�	�D�<j~�9�g���HS!)�`��H�9�ػc쟟jMu[$��6D}M� 0��֤���B[s��W�y��*�,����Ue��(-;��X,Y,}�y4t�du��e���r;�WOU�tyB��Z?�DM��U����d:���}3�Nנ3���6��-/Uˣ��dD����T�,�t��~��n����v��ᦢ6n�0��'o2�`Q���E�����: �~߄��㲧�H
�/�2����5��f��$I�w�*v���T���h���Kp���G���G���Q������7�	{�VY����|��TS��<�,�W��m��^z��p;=��<jj;���ҩ X�F�;��� ��X,z����JϋOu���O�m�(����R  ���:����х�?�u��ώԨě�uA뇟�x-P")���v$t~pM^A�C��6J�褩i�;~�3u$Zjp��� ����BO�ӧ[����f�ێs��?M�l��ϓ�  &��%�xro��bm��RB �X{�C����io|hΈMp�g�f�M��n��?}=��*�M���;rUZ�N�׮Sz����a���N��|m��=�(S��S��s��pU�n�}��|o���.OJ�,�{��
gӿނ���h���a��8F ���b�]9�ػ#U�ϳ[�b��u ��Ֆ��Yw�~�G͇ޟ�*����\���q�b�HF�r
oP~�-�)�VNA���t��*\q��ӭ��i���,���٦����p#n�Ey��F����:%��g��CA�#�j���f�����*kKַ�&}���o��a����z���"Q��~���`�kܺaF�hj;Z�4�XGA�#4:��r��׬Յ�:{����UPT�tG��v�,KB��l�������
����N�,9��^K������_v/xn��{�0��o�Y[���:���p2������V|S?��E��'o��TO�����$��~s���TY����#	�XlZY^��kV)?7Sc����Z�η��(]�� ,N���٬�zroA�������v��=�i�A���	̷n���E5�QS�f5�ܦ�㧴c}uhzf���W�f��y갼^��m��iF�R��T�Y�[7�
�DZ�$x�|�۫�v5��>:7}�n��,�G �.����p��Ou$�9�ػ�귶��$F� `Q���-/U��H��ܤzz������v�,�����^�ˋ{�H���¯��n���lAܫ���t��Ia�x�����)������0�E��~k{���k4��O�-��Ƌ�6YfD��u �ht}��9�/���xhZ�BO�����{I	
rd�PY�M���I�:/$�ىڛ�T�UGނ{�Iх���B�nm0�|����)\x�Jiz���BdS�fISm&�0��o���=�b{�7���{�ܧ�6�٭�E	�P �\���5������a"�k��~�&''599)[Z����,�P�z�vh�3.Ir�����}Ѕ�?�;�pQ�T��7]��eO/RM�N�mܺA�;���Xmy�Zp�)��+f7jܺA-��q��r�30[p�{��`�kz�Ii $�Ţ���{���ܧ�6D�������ܧ�ט�����~�t���cM ,ӫ_�X_ڬy�=���@װ�&�~]������5u���rTV�gs��|�	Ym��y'd���3��j�Hz�����t�i=~J�WBَ���/�r�S�5�o}�k>�~�Ѻa�G�o�*�����3^�0F0c1���G�Pˣ���8_�;���q��� `f���zW�]�O���@@����uM?���Z,�JTg�h����}�: X��S�ZP-�ާ��aGꂁ@���9����u����b�)7�B����h��#��s�5��Ž���Q�h��CV�`J��z_]�N5l�	��u��Z+9��p�u���h���צ���8wQ�����nPæ�ｩ�Z?�$��1 `&��Xt�d�;�1��$}˳�۷��j�J������>���o�$�\�g:9�Ju3�����Z��z���4��}5���Rmyi�}��nPS�fu�����9��>���F�mGB#s�jԼs�T��W"j��}�Jݔ�ٌc���O٫bzO�M�����^������ׄ{0�z�d�������  �+���"�|���u���`�����T��Ֆ��=Zc�Xd�Z����U��5�/�I�E7�jK��M  `&�_�"���7����6ը�T�Z�����2�n�������oPæ�?u�i�N_��kg;?�urT�Mv�-����z���eM_)Gza�kpBҙ�� �rE��E�k`$�^���?W��ݡ���~v�װ�35%�J�pS7���/Å�?�  @��Kk�R�5u   �ǚ:    01B    ��    L�P    &f/))Y��������8��=K_q�D�   ,Q��   ���    ��u    `b�:    01B    ��    L�P    &f�t����1U���^��>UϏDFFFaFff��?�����⾧;@�N�7�M    ���/�גnJuC��>���������z�����O�    0\    &fOu ,]��"��ޛ�f   ,i�: 	㷧�U�2��   XҘ~	    &F�    #�   ����   ��T��@C�o3�*=_�P�j��G�   `g?PqW����Oߑt�a���    ��q�u}��[
�.���wT8h�h#�   @�4nݠ�m��n)� ���   @�d:����*��P���Q]�]���P    �wn��e��ڎDu�RtA�;
�    H����j?��5e�-�@T��;�H�S�9�Q_�H]��Ҿ��6    fm������d����:B]n���Wz/|��v    �lL��P���5����:9�Nus    \�V��U���7n�G�'���>5�E����f����T��^��qѰ��F������댮R   ����1�S+W(=}n����ٳ�
������46��ʕE�?�T�~��ϝ�P   `	����a��:k���w���+Q��ΟTaav�����$���    ,~������y���|��~6湉t�R    ���   �T?�E����0R    &�H   �%��%τwƱ4�_��i�}���<�3�kKK�s%B   �%⓮:qp�q�զ��I�	X�t}����<ע�Ң�<s�s�    H ��:I��}�8,�w2��1?�2��zn@}���O    �����#8�'����3#�>���:    01B    ��    L�P   `Q�_q}���4~�M#��b��P   `Q*Z���nKu3�o����wk"=+��	u    ����t�   �"�T���N"�   0���
t�   �I,�`gd��$�!w   �$*Z-�6�\:�����ut�   ���^T�k$�͈Y�ؐ&�u    �������+�͈K��H��ʨc�XS   ��B�����r/B   �Eo)� ���   ���]���P   `�Zʁ.(�`G�   �(��~��]P��({l �k	u    ���T7!��Ƈc��P    &�>u    L�s7��]��d��o�n�:O�׻|j���F�   `j��4�tj����ύ8�=:{�W���S���u    � �ΟVaQ����!��w���+1��R��?!�   X"���;/��?��?��f�
�    ���    ��u    `b��   �d�����8�f�+==mI>W"�   X">麠���Zm*+-������熞�л   @�Y�7XI���S��ay��K⹳1R   ��>>}>��|RO�x�l��   ��1R    a��7�aS�
2�Q뇟���H����0R    !�wnS�����sU���ƭԼs[�[��0R   �p�5l�Q��Sj��/B�ZP�j��vD�.ς��_q�r����ܔ�[m)\ӵ��   0\ݍ���?	vy�z�Ԍ�2T�Z]�ݖ�."~�M'o�[�Y1]O�   �4]�Ψ�_��.�@'�    ,rK5��$B    Xj�Ψ@'Q(   @U�i����;.I�w/X<e�h���T��;	ik��$B   �j�����"THe>�`Wr��K���m0,�I�:    	�q��5���h�V~�Gu_���G�   `���5�1��g?Pq���M���.y���[}�!��P
    SX
�.���p�א{1R    a
2j�T��?Q��H�X㶍��^�a�G-G;���n)����/�]Y';B   ���-/U��� ӡ�Ag(Ե>��j�KC��U�QSQ޼k�b�2"�1�   @B�<z�$����?�$5nݠ��R��T������W�q��mTA�c�=�r�������b�    n��jU�����|����su7VH�������P���4���z?Z�.���w�=6ӵ�:    �N�l9�:V��P]�u����))4�W��1��c�Ih��5>�u�:    Iz�zRܒ��B)    7|�-I�,�m*�c}��?�������nX��6W�f�?޸�u�<�w?�4�g,���F�   `��h\��jz�*�th��ju������.�<@s:�re����F����=۫@�؉��z�l�:    ��8wQ-G;հ�&4'MU�j޹Mu�kTY��+CL    IDAT��������u���
��e��Q��[~�_�Y}����	�   @B4��Mu�h��j�<j=~*T8%8B7�����3�^����;/��?��?��FI�s��    $L���n*>���G�P��S)h��B�K    	S��PS�f�U���Z��j޹-��#u    ���T-�ާ��|Is�T競�T;�Wk�~皺勑:    	Ѽs�*��`��ޜ�+����vD�5��f�3�]�pi|Ɵ��IC��+1R    �ר����EP�����5nݠ��5qmL�I���88��jSYi������zNB�   `Y���B�B�.,��&Z�V�����wqX^��#g�z�l��   H����50�3>>}>��|ROo\�Y,ϝ��:    ���`���ω$ b.B    ����X_}�s��P�26�:    ��8wQ��O�q�5n�0�y���O��U$e9cM   ��h�ɛ�,�WS�f5l�Qǹ��tJ�*��T[^���|u�����6����m�ڏ~%�ߗ�'�Ǒ�K�T�t���,Y���[g��P��   �IA�C��6j�-7�Y_�50��?Q��i��	{}���%�<�l���ޘ�'�E�P   �'82'M�H��-�`o���~	    I:�]���Dz�N�|��vF:�P    
2Qo&��q���0�Z�3*�I�:    	Pwc�Z�/�k~��?5��K%��$B   ��8wQ͇ޏ���	����bmZ��Z�r>J��R    ,Fl>    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01{� s����5=�RZz��2?�_#���T�   0�q�8�У���T7e^�/_V mT"�  `	b�%�666����T7#�˗/���?��    ��:bllL�������������@��   $��SZZZ��2::��&    	G�ò�ZT�e�l�,G�N��   +B���4�ʍ��YRR�����a�   bE�    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &fOu��
3��ސ���C���ci�����|�c��n  �]y��+�R݌��,�zzc�k��
=���X
c�����f  `W��T7!*�:,�>cC���   bŚ:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� �P�f�Ck��_Ia���/v?    V�:,�t}�q�%9��   ă�    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� ���Kg\~����v/    �:,�~}�g¸�\2�^   @�~	    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���S�  rm�Zlܗ{aN��߳#��   ��n�������F\~C��?i��%�n�=����\B   B�2qflB����o֐O��   @�XS    &F�    #�   ���    ��u    `bT��i�|>��n��~�l6eff�b���Y   @R�`J>�O���
�$��+�׫��\�   ��_�nw(��|>MLL��E   @j�`J~�?��   �RE��)�l���   K�����)�u�oZZ����S�"    5(�S�X,������D��%�   ���e�X�p8":�������۸�|θ{   q`�%    �#u0����R݌�ݮ���T7   H(B1>>����T7c�ϧ���T7   H�_"n�5�I���S�    a�C\&���-(UAIy��2��_�Y��n   ��:�er�u����W5��    	��K    01B    ��    L�5u �����A����n  �p\��&D�P ��seU��  ����K    01B    ��    L�P    &F�    #�   ���    ��u    `bl> �jJ��o�ָ�:����g:�t/p%¡? X~u R*7=M5��r��c��e�m)l�yџ  ,?L�    #�   ��1�@T�\�*�՘˘�YΡl��������\.��*��D���ONhrx@���2�{%B�k\�?9��˗��Ŏ4��o[���CǼ^�F�n����}�I�Kc�C�>�x��  ư���r��VZ�����+*��\Y�7�\s��ۍz<�(���u�~-��-��<E7����ؤ���T7e�  a)��:��~(�m����T>0���n���oVVV�$���L�C.�K����$��ŋq?o��d�gFF�._��,� ��lY����<���'�===��'�a��7���v�r�-��?�3�p�*//Waa�$͘&8��������&&&��ե���9sF��c
&�%�,������ٳg�D ��-�PW\\����<��?�?�KA�$##Cw�}�n��v�|��r8��H�|>���kddD:y�~�����O?���"�'  0��`�C�xV�������l|��SFA���Mx������!MK�XȪU����k�ƍ��Ϗ;x,dhhH###�����~�;���Gt]���	  �Pg����r��p�je���z�r�\���]�����٣_�V2��4��U�V�G��͛����@ ��VNq�\�������~��_GF�Db��G}T_��Sڟǎ����z� ��Y�.Uk���Ҕ��-#u���x4::�����s��r:�S%�P��&�dggk���)	s��\.}��gr:�:x�;����
"�'  H�e�R���D���JKKKe3�˥��A�^�z��������'�۽dB]��n�����׾�5egg'tZ`��N�z{{500����/X$�A$��|�ǔ��C ��-�!���C���EVV�#u&�~�����y�������D��$�.q" ���z��'��C�f��t4)�á�������v[(��SPP ����ߖj�4�����	  �[�i�P�x,�Pi ������|G��r�|>_[�ժ��Y,]{�*++����Þ�� B�  H�%�6u��ru����K�>������h�|������)�á�7�>�����"�'� �d�,#��E@�mۦ��~ZYYY�	 A999���T~~��y�egg�=���R��O���b~��'F�'  �:B��E@�|�ISoϑ���믿^iii	"��\;  ��	���������T61p���ʕ+<���������Ą�_.� 2���ҙ3g499�={�h||<�y�Vq�?��O  9B]�|>edd��΄&''5>>����ϛ�������7U��4��]�V��������$�.�Ad``@���w�=/� BN����VSSӼ��  H���b Q�$���g�UVVV[����*++Sqq�{�y�N�����9՟��'  ��X�2�� z��'URRb�"�*,,T^^�jjj�iӦy�+..�Ĩs�{џS�YXXhH ��� �q�}���n[������L��k׮y}a���5�\#)��	  f"�����Z?�pؽǖ�ͦ��2����'�H�3�[�Y�&��	  �"�����򗿬���T7%irrrTRR���r�[���{/�����LX ��u B6nܨ��k�O��k����Z��G,�Oc�  �G�K �Ͷ$�X,Kv'�e-##C;w���MuS��f����D^�W�a�=�Oc�  ̏]��b�hrrrɭ��Z��X,���,��V�|>ߒ�����jݺu���HuSR���D������ׯ���G۟  `~��
Kr��|��n�+==]�E�@@~�?�-C��v��o߾,G����K###ڴi��=��Oc�  ,��0�����˗5>>.��#��*�����5�\�[n�e��"��n�q�q݇��bT ���>�/�$��jbq����+�����)������<]w�u*--��>����  ,�P��
r��r�\��wX\���USS�$�
�"??_N�S_��c����)��  W�O�H
��/�˥��IF����UWWS�押�<�|>�_�>���ϙ��O  pu�:$���._����ȝw޹��~Mg�ٔ���իW+;;;���ϙ��O  pu�:$] ��c:fj��v]{��Y����v��nݺ���?�������X��	  "CiB�������f3������:+oKQk"������J���Ѳ��u��]��Q_G�k ���R�gI;�ͦ�˃�nF�


�f͚e�A�|rrr$I7�pCT�џ��ڟ   2�:��R	vf�j�*
z�#--M���Q]C�/��  �aA�ǣ@ @�$#����p(///�k����ҟ   2�:,���<�iq�+--M>�/�>�?�K ��갨�\.��K"*5�/==]n�;�u`���b�O  ��aQ	r��
)�����jrrRn�{��&''�!   )E�â������NA   ,Z��~�=`�w���Y��X��
��b��D��P�EirrRiii���LuS   ����7�����w���?��X��m$�ٚF��,v%j��P*vQG�W�΋�焯jܽ�(�!,��=lv��E�[���L���oþp�C�2��]j_%G�nD'e,%��&��-r�^P3�(��ΐ�~���4���cZ���{� l&r���Ƃ�~�踽�b�
���Cz��I�;�Y�2�eɿza,\�/�ŗ� �@ۙq� �~��;&udZ�t��:"�K�����n�0��,�?�����x��/����u2��u�_���Ů����,��?h{��X��v���Q-�`�K2�Z:��j����Қ��Y}��E���Ç��Ԅ۷o��1���ʙ�z������.ڛ�����8��gB�Nf�g_�_�y�,c:-Jn�:�ű���Q_�	Hh�� S�d25q���ں�k��L�ϬVVV��imll�b��4G���ʙ�zu�DU�?w�/!��2z �^'s{��S�1�����WǦ�����PZ��Z$v\~I��N����Oj"i6B*�*yo'糰r�^��_�k�o����Bu���y�4I��dV���+3������X��EI�:6�rn�m�İ t��<L�X<G*���e�Ւ�d����d2Y��8�;+w>�ٕ����P��ש��@"��<�H��WǦ���Z �U�s�#e2�ZY�Y���8��鬭e�A��Ζ�8���ʝO""�j� ySǢՎ�r~,$�}<���2�,��èK�D�h�Is���U�۷��~I��|���$""�&YƵ��c!��/�%���x�A����_��IH���U������|����<�̧����=""��TF�:��cqY�|�<�wT�GI?��կx`�L&���|��Ge=�����|�t>��v� pr�β��Q�e�̈e���/�˩�1�#jp������e�iii	{��){�W<�|�t>����A���c�,��~I5A�$��P�VWW1==�g�y�t���.�H������/�z<�s�T4�fao���œ눛��<=��ن�_���{��|�'��}������� G��� 89��cO�  x.mm`:}ng\���h���'�կ{���:^ṕ�7�r��u���W�cj�����ف��_B|-�_\�������9������?r���7��Kptv�s�-�#s[����q�?�v�^Ͽ��焫�K�Z��M&n�<u�#��R��ւ$��K�/-J�=�8Z�c��QM��V��������6|uiccKKK���X]]-�y8�YXYY���|E�Y�o��#��@;:;��4k%�{�����\���y\җ��w����7�:}����������7��<�^��$wv��:  <{��mq\�]����9z��7կ��=�n�w���I�u�f�/>���|/����aDc	�[���-�,N�xsW��v�d���x����W����z�����\���Ww�#��� w�͒?�*�ukFF���K�:6�~�b��s���j�,�쀩�{��arr�����/���}��������|fi5��8:;��߮��;ث~R�5����]�(����w5�I�_K!89O�S�R�G���l�;��0p�&����V) `j~!{��G��;؋xr���G�_wtv�7�Z���:�[��(�����$��������]=��ȅ�#��QJy��d���ϏB[ө�x_[MZKQ��֊,c��w��D�I!�N�ʕ+��d2<x� ���wiT��jm��ZΧ�n�Fpr���7@T��k)����-����!����a���M���ݥ���~���A|-��{GIDɼr+j����|�X��7���U�>'³w�u�f[Y]{Ky�+�'gv\�,-ͭL�F��[+�(��l�JM4�� ࣏>���߰��!�"���I���裏��{�5l���|U�����^�g� �ހۛmE���g�l��M�/l�u;{05��pdnK��݅����b::;�Pc�9y����jUMY������E�Z����lC��mDc���BJ}�k]iε��M[5���TSA�:��������7�7�,��`qq�dR�$d}}?��Op��Q�g��_@pr���C!O�n��$ `oi*�9ów�*���)7��X��.�#sp;{v�KUh�f~����S���yy��L� ��f)	X�����u�N��o���5��K�b����Nv��A���BU��_����������uki5m�嗒(�E��u��3�������D"����w��d2��S5��9�����D���|j;�;��4!pr ��H�^%1+�r�U��H���7���F)��I�J���CM�����Dpr�`���F)J�{����եQi#���MG89�Vn�#sN��7<��q
een2�u[��۟K����L��N<u��%��zݴ]c����ӨKت-�N�ҥKX\\l�����
���055���/Χ�{颱��u��=�})���%�?+�U��(��q{�S/��ei��d�ꏲG�X�����rM�1�����-I���N醩�2��Z*۔�ن�<?�Gm���K������J[.�<�xr]�v�sn.��V�s�����J}�Gc	��b�[k�V�tR"Qݥ\�J�.���X,����A,3z8������O?��������|�'p�fիc��&8:;ؐ��'gԆ��	僃��������V�$N�����Z
���E��q�G�mk;O�S*j�+׷��
�:���E��|�':}b[�47�*�� ����RI+t]9˗�zݴ�:�	�R�0�p8���Y�����O>1z8��x<�믿��9j
�'Q��_��M�N�@���-gw���|M15��=�+����=Ww���J+��BG�7ԏ�t������a�Ȍ|���N����Y����t)	���+{v�G�($=}�]�J}����.1����䌚�z����n[Z��^�6�ba��AJ�2�#�mdY�ݻw��3�`qqKKKFIs.�}}}�Z��/̝�D"Q��jΧs�؞(�P���\  BIDAT�)���\z+[�x�Y�#_82���;7;��t�������#�N
5J�M�	��	��4��f*JI�vJL�%������<�_��]R�YS:izLh:�����;>�����^���|C�p9��1�끫7�<����׭�R���.��:u��!��j�j�8�r� @Ū6�H��X[[C[[[��666 I��կ���s����E��{wnWl�o����G^��ֆ��&���u��9���Kx����o�vyy�}�[XO����p>����
�����+�������������/!�+��b�`o���+�!Kd�[��|�'���qQm�����Q���P��w��_��V���,����hH���hii�7��M������0zH{�'��/����ʾ�\���ػw/�S'�f[v�[K���t�;jz����� "�mб��g��X�� �U��>��/�����X���Ckk+�}�Y�ٳ���T�'����Eww7~�ӟ��+�q>kH|-���f4��c������Sy%"jD�\z"�#o�`��L�	�9ܻw���>[�&3% �������B��7��>rP�6:5��{#b��߷��;RǢF���̸W J>��I���j��ޝ�����~�ݻ�������n��	s�\�����'�|�4	Ƚ{����Y�����i��ԛ��R��WΦS����g�N����v|���|�'tI���ID�a���JkP���q� ��rʤ�L�V*u+++��ں����yҠ������hjj������֭[�����\���nA�$�A���E,þ}�jv>�|���z��&�`Z����o����y�Spr��j�o �'������59H������}�`��{N�@��'{.���\zK�$ˈ�Dd.����[�n��T� &udb{��a�Z__������o���|��)��v��N����x���ҎVVV�L&100��,Q4�@<���g��r�O�WTEs;{�9�=�|�\1�ȱl��Ko!��B��	�G����F\�]�N�;Ҽپ}�Ͻ��V|��1�ȜD���s���cSՌ���G F�}<�:2-A I��àH��h4�'�|_��W��_��Tg���v�����~�3�/�$	w���|�(p��p���D4�P�y�7����BprF��g��?r��.�Ԁ��5t���ߏ����lI�k1&�� tX3b��n\�W#f˹q�(��J��I���je��ܽ{�(��v�Ν;����L&������׿�u|����/~a�X���ԇ����%s�{����;�״>>����%�k���*$v-��]VI���R���Licc��q7J�LX__/z]:���b�Ҩ�I�ڵ��bdd�H���UMF����tbqq����*��,���	�P6��;d\�����X����<G#��ڒ$���_K!�,��B��ē�L,��4�$v�s�^��b�;;�%1XiB0�#E���D#Hg2�WCWWW��'�����'�O>�sss�{��f1r555�駟�7��M<��Sx�����Q�8kkk��Tr>wo7�[ng����-�=}N ����b��U�D3t�6|��>�ݯ��H#������`/<}�-�5���ݲ�3x긚P&n����|ϥׁ�F�$"��Y%1�v����~XVW����7�����.�:2Q��5��$�i�^]�������������a�Z��"�U��455��p����~�iX,ܸq�n��h����q�=t�f�Z�900���fD"ܽ{�n�s��Gf�g�K�#��������	'g*��4D�S*e�/4ѽy��|C����9�Mb�Rj7N��1 ���.���b�<�݈�DT�C���3=A�W�|mgƽ� ���FC �F��2:t�m�Z�=�=A�N�M��/�� �J�����u��˶�6����������9Ċ������!<xP�f4� �w~�w��҂��%ܽ{���H&�XZZ����n��n��'�@WWzzz��ގ��ܾ}��_^^�.�����c_)x�Q���c��/����l���`�����a��=p���l%+pr���o��{�Ww���SO�f��ܫ&�J��WA�:<u��v�A�>'��?�������VFDD��2�ɐ���v���6:��k�xA�i��)X�#S1CB��<�;�{�H$tODdY����YEtuu���v� ��������b�ǿ������}�>��3]ǘ/�L"��m��!]$���OeNͧ�b���>|�>��ABWL��M�:GgGv��?e_�w��f�nU2{K��6�5�#sۖ*�A��Dc��؛mjsV	��A� �+~,��xM�� E%���D���nA@ �:.&ud
� `mm��a4����o�z26����ê!������qUc���C,..b5��M@�������AI���:�sS��Y	-����=�F82�m��lC���o���t@�b�v���Ec	u�`82��tD�`˾�z`D���jY�F>�c���<"2� �9A�s�q�77��*��dRG�cBg�ŧ~�O����֍5H��t&S�18���G��e?���~��}�6���#����@ =��.y���S��Ep>���n�[�89 [U�7���_�xo]n<GgGիb�+�|�yO߲����D��0����߈ʕ��e����VM�}?
��C"z$&ud�zI�������o=��-xʰ���_��aߖ�#��8���(V�W��많j�4��M�g!�X�����;5���bGg���������*B�x7��^Q�2K��7���@��k�臈�:2� �$���ՊL&����F����ެ��T1ng�#�Ԋc�A�z%t���-q�J��\U;���Tٿ�r�!��7�`oiR�\��S�LIGgG�^�Qg[*��Wy5�Y�L��,R��.�߉�1�.������S7�ă�3�7���s"x�8��?�M�n���FШ����\U;�����lSv刊\�X�n>����;ػm)s4�@pr�n^�"x�8<}N�g�����I���z�5��]��=��9�f���}�M������D��_|C���;7��*����	�8z�hL�j!�S4�LB��� D�c��fXͩڮ�&�LWw/Z�h��TZ���*�ĵ�x�����9���8�Z�J�����s�7< �� ³w����X��Q�2�ZO�#�\�~8Q଼hgG]$;��~�G�!�C`�Ɩ9v;{����K�#�gD!Z'�~��TϷ��"�{�������c6϶T��*�� x���:}���۾noi��ϩ���~���^�瑲�AY�`o�m���^1���`u�
�YH���F�n4�|O���A&n �S[�+7��Ύ���t(u4��c���j����_�6E��O�3{�����MGt��f\#*WFV���;eI�N�.��3�*,��=z�>�#�S:�j�;؋���}�u�x89�k�LIr<��R���7���^�c�ów�9�mń�ϩv�՛+?�����f&u�+�ł�����;GD�|�}��m#%		��<|C�e߈���[Yf���;���@��M�JN��Q�j�j��r�\,v���I�J�� �U�Bϭ����X�X�����v�Ճc��s14�.OL�4��� L�y\�������͹��_���S�!�֢���oX��k&L�Hs��$1�#"]){E
-G�7G�~#�v���P<�bdoڪ�߬q�H��L�]�]��>�z�S�u;���P�Z]Wx��w�S��$W��٥�:�+�/�SϑT~F(U�����ȏ�z�5�{ng|C���sh:���F��	&��z�;ث~ �,�MG�+66_�s3&uT1Q��(�2��4R�����r�����rtv pr����_���zc���ܛ&=؛m�A��.u9dprF�O����/�8�ju��FLGgǮޣ�R%�_���q�i����4�k)�.OTe�Bٓ:}b����t����^/��_|��
��]{�������h,ϥ��9�.�ԓ�G!��=puw��ݕ=Sts�|��[��}�m]�`�*�q^}�r[�֫F�A�$X,�AH��l�,�2$IB&���$.�� �J�����u�t��(b�?�����vS������>�]N�s`w)��6L��7�\�u���O�7<�h,���}⮴�w9 �7)1:�"prX���	RDc	]MSI빂��܎�
e?[�+�
=�*U�|��l��Ko�����<}N�g����U�yV�{T:�V��7w�`�_�QX�����2��٣V���H;��|�o�Om+Y���tz.��pd�����g;�uv�]��v�d+�U����N�����}Z��3"&��B3��ԃҡV�_֣��N�7��5?�^{��6ڛmp�oG���sh:�=Ba��g5��V&��z� �1�#"������P��ܮs�P�JwKe����U��[pr��5=.Wi6�׍��g/�S ��<e���/�Sa�� �����+��_���wt�˸�B^[:?�eRGDD5���;�޶?G��f���;؛Mb7�f�S����B|-���͓{�m�YO��3�:(���Q�J(dj~�>'��ܤ3�Q�I�R��=���O��~v�2n�Q:��/�����.O�庺T2�|$=T��?r��~� �h,��郒�j�`�[��N�S���g�s�<0Z��s�'�y��LUc���i�9�������Ҕݧ��Z��p�e�Z�k�܄`RGDD5J�\�$����W����-V��(�l7��	\�	���j�,����ϩ�M�!�@v��w�WӤ.K��YT^_4�@0�:���P?��՘�u�����S[�+���
θ�k��F�O� &uDDT������r�Զc�����vـ����-M[lG�%��^B]���+���[�##�#s������Mh�D24��x#bc�9�z��89�P?B��޻�˸�h�����J$�~Y�x���r|C�r@�w���c��!ttv`�� |��[����&s���e�o�_������j�é��TZ�m3"f���T��z\>���P�V���.O�t�q��J� &u�bRW�����(	�rV�B阨Wg7�X�l� ���%L�����|C��l��=�[��4�<@3P�*���qT�2n�)��L�t5??Q����F �22����+�eYF[[���ˤ��teo�e�gy]7j��r��;��٦&����S�SL�`����^�r��ۆ^�3.��j\-=*������?62<U��?��Ƥ���H�0.��z�J�&� �$""""�0�ƛq�lv���~IT3d�daRT���([\� ; �-�3h�DDDD��R:�I���2�ɐ���pq,^�Ұ�l�㎽�Gd� ��DDDD��R:�I�)�2�eɿza,\�cSǢ)   �vf�+��������L�LE�,��/�0���-_bt<�n�0��s�QG����O�����G_ȸ�˸��5J��3��w\����������x��AU�~�k_S�<�9u5��s�V�&���2��ɛ|ul��'*`��q�1( z<?Շ}ˋp����� �2���D�c���#�U������f��f�1��A�t�,�����u�$��x��饌�ƅ���*�r~,�rn�m��0;""""s�4����j���Ts+���ș4�)$�[�_�� d��XJBW��&���M1�#"""2-:�I��$�3���CF����2�H[$���|�WǦ���Z �U��DDDD��V	� Iݣ��E�~{�Y9?j?{�"���nH��t:���	��={�0.�2n����q�;��L�J�ؑ��2��\)-�ۭ���0�QdY�Ç)$�Ɋ�KE8�2�G���q��Fi�yf����5�:����O?�4�{��w[!^����R�k� .���3�>Al�8��A��bEKKKE�H�_�V�uW�D�q��Fi�yf����%=: `[F"�2~��85z�Ƃ2�0zT�_����ʸ�˸Տk�F�gƭ︕�+���B���c�4z T;��E��/P�e\ƭ��N�h�̸��\z&t@/�$2+H��7n/]��(�H"�ЮY,V,..buuuW�>���(�2.���m[��3��w�R��LꈪOF��!�J�:6�~�b�S���)���n?����q�v5�<3n}�ݭj$t �_U�,��G<��M"""�ZW��`RGTu�(��C>S&�DDDD5��	��������H3�N� &uDU��6_Ǔ�C"""�ZcDB0�#"""""҄	�����Z�p=�|�$����IQcRGTef��	����DDDD�;Lꈪ̔	� ��C """��X� Q�1Y�rn�%H�0zT[�v;���vumkk+�2.�(�Qm�����:�*��}g�=+��BF� ���5zT[Z[[q�ر��J����ʸ�˸�5J��3��w\3��K"���)������ڊ��8��V�'��˸�[y\�4�<3n}�5+&uD|�6:�0zmgƽ���v��_��r�2.�2n�q��h�̸��̸��� 6�L���u��vA�ŧ�!Bſ@6�@v��2.���(�6ό[�qk�:"��3ro]�U��JG�!�"�V+b��2.��X\�4�<3n}ǭL�$B��w'_��f�}g�=0Z͘T�dY�Ç�q�����q�;n-��:"	@�5#1:n�V̖s�.b�Z񈈈�H_L�&�k���j$v-��]VIs�%Q�`RGdJb�rnܥW�}g�=L興���`� jE��q��U��A�M�,��/�P������ͦ(�CG�����7��O����v�e\�58�Qm�����8?jH~Ťn���Q5�2�eɿz~,\���
���C�����
0*�c�K"<g�x����k2��r!\��汶�q�^��#���Q�cRGdb�����uX�c���k��0)*	��^'�� ��p� ٠Q�1�#�������G�f��DDDD��/w�ҽMDDDDDT�d׌�ͤ���i��@DDDDD&$`ʨ�L�J C="""""2��(��ͤ�˙LPF��������C�q-��+u5��X\��ݡ�DDDDDT�2��72>{啡��ũl�x"""""jd2pq�����1�RW����f�""""��&���L��sq,���ֶ��������Y��=��/+�v��|� ������d��$��αfR���q{���L�������|
 ,A
��=�|�����I
    IEND�B`�PK
     ��Z$7h�!  �!  /   images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK
     ��Z�U ��  ��  /   images/ae1d0bb1-db79-4eca-b526-eb1d648f9ad0.png�PNG

   IHDR   �  ,   G}�   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  �VIDATx^����yލ���[���+Q	� ���R)�jVq��/����|v�=�K9�c�D�-KV�%Q�DR,b�������~�g�C$!	.�>/0w�����μ�[�m��lZ�:ԡ�[�u�C? ꀮC�St���:��P�~��]�:���:ԡ0u@ס���3N7��R�'��f��h���F��lFM�BF#5uR��H(T��C�D$R����D�M�T��c�O6�٬�Y�n�yD��:�e��`u](�XT�������������ޡ��:���T�Vs�J�w4r]�&�l�����H�	a��($ �_���
�ڬ���Ԅ�d�lX�?7P��^&vuhZSt���z|��ԇ�]]��
���WT�Q�W�ba�h#j�:�k��<�|�h���M�g!�<P3���f�?H�\�M[�t�\ *�G���U�Y�m�,Y�X����Z$!c2��IY̒:OF�;�D,b�$!j=�KH��J=6��~�^1�l^�J�CӘ:���j<��d�?we��zF(���5�V�؞����		l��\�i���5e_���.\�|�%cqK������R}_#~fy����������r���]	�M_:|����MY�+k�������V(��0�w�d���)��t��׋ѝٴw�����Q���[=�c��`!f{���o�D��.�MK��P�R�>�~q �:V�Y*�ᓃ�����/~����K27!kԛt�ȻY3�]�zz�w~�?���|�U�!���#a;8P�o�E����4��Ow��hD�uKqY<&-V+[$���Y$�_��\�R��%�	K�Jƭ+���D�rф�jf������E�4��.�X����th�Rt�����Z�^��w��tlX:��;�u����W����%�T*2E�VmT�)��j��gՊ��[�˷X]�fR��4k����5�A.���� Y��PȤ�8oZ��x�p&q�^��#φ]��LO�tM��(�Mc����BqŢ�S����������A�T �#�-��W��{�g��b��tr6��N�Ns�4Ѕ��87�����.
�K�k<�� E��WŅ� N��CӒ:��@4j��E"������3D8:(����~�m޼ٙ��d�ݗ�lv7���@^�A��k�v����k5l>��&bzf�M�9u��`^B�Hԁ�V���ؘ������8q���Ƀ��������O:-Y.���t��4��.	p�f�U>Z*�H8�tww;`$�q�@�H\�a^f2K�ӧz.�d]�n�St�b��U��A�j��͛go}�[mѢEX #��^z3��[o��7Z�Zq�!�R��9u@waȩ&��5@q ��D�q��C���9Z,�}Һ��^tӜ:�� $ 5+�F3
;�E�qv~ڑ#G�<�ځ�zօ��߾��o[<wi����uh�Rt��ѐ4S�M��ܸ�ܹs]�\ �����q֬Y��f�5�#י�������.5��P�J��&��1�O����4 �l���ݶm�lÆn���L�!v@7ݩ�@�z�� � ��xৡ���Ld�X>�w�P�:�� B��-u@w��$��OW,,�YA`c�%�)h�z���)�NH�����{��-�JN#v�\��"���
E�-�q�� �\`��E&y)*�z��LV���4c��u@w!(j�Z�� V�Vl``���]wْ%K� ��Q�9�0�a�9۴i��v�mڴ)����kJ#���l�ҡiM�]8r�\P�\��{�����)M�z��~g�b~�D���Q�Mw���*��NLJ:Q>��O�q:��&?V��:O �_�j0N��Y)�B�̜��݅��Sr�� $�\�֭[g����oD+W��I:�Ι�	@�40w�Cә:��@�ղ�j ���;�í��f��#�B��^q�v�%�8-��g�8��������.�[��hjj�v���|:���ٳǆ��`���i�uh�St��P�ѴT,����b�X~�_tGz$�ȧ{��쥗^r�.�b����uT�4��.	7!z1!#",���H����MK��òe�l����x�`�A��;u@w��%�p0N�*�R�h���ΧHL	�@����-���:^ �b>���K����$ Cw2�r[�}��_�C��!��Q;��~�W^q u+DhN�ӦӜ:t��Vo���~���� ���?j�	���f����z����wj@��F�ceNs��BP�Bl�P�W-��8�����9�"g%��˗������$E	�X��5u�Q�ѰD$f�f��X����]w�e�ׯw=�gj6�� �_{�v�嗻�]�.w�=�t��4�N]0
P�l�L6����}�M�TD�����v��14�嫬HP�N�Ns�4��h�O\U�i٨T�y���ϸ�Rb�h06W?=>�Ǒ��/�����L��o���)��i�iN��@T�0/��K��.�x����w�t *P���+�_���[�x����T�`x�MvhZRt�2�p�����R,Zwwή��Ɔ�ui>��t���o�XK��K?�N�u�t�S��.��L�T�FGǝO��'lVۧ���o���=>� �y��tӜ:��@�0m+�z*!4~�1�Z{�����] �������F�3�r�St�����H�k
dl�w�u׹-�j��)sӱ=xS�)`.t $|�	+�ˠCӖ:��@���]G
.$pe2)�r�V�10�i�v�y������S{����Ҙ,}��;R�;u@w�h�Xv*	sQ*͎=n������K��<Ӝl\c���>��c{���Y�3��D�3OMn�#d��]nYLE�35���&F�y`�ST ;������J=  B��{��.�=9���6�yr���5�\�U�<{*^rӞ:�� �4b�Lt���)�˯8�(�͜[{���y�"V�ON&&����fXq;4���D�N��l���,��<���n+>z#=2�Ax���7�z:mɵ���;�崧�.5����?v��`�X��/�`i->��p��O�k=��f�0$Zm���|*���.ET���f�	a��;��}π���"�믿�MìdءP,�!A�5C�Cӕ:��@$�LbƟ���Nz!�$h��Z�͆99g�T�x^����:������f��o�w�u�)�;�*��l�z�!{��_�Ҝ�etӜ:�� $T�Ba����8��10��E4���E�� j(��G���8���
���Cng�Mc��B�L�r���S�����8��oD"15L�"!����LP��RS��/a�1ɛo���mXo�rŒ��
�e��:4���ER`�hB����~+���<��6�;�h:�#��ŋ,��c�D�T�F�nu4�4��. 5��� %��ڑ��Y���~�}�����Ӂ�w��ჿ����'�x­2Ǵ��ɔxtӜ:���ڄ���HG
�����611�yy���G߃Y,]R���J͸�h�Ms��ک.G,.�^�Z6�ex��mάY�S����X{�7��� x)a��Mo�����v��"�S)��JfNM�j��'��Zڏ��И�"�P���ج���� ��9��vQ0��!��c��(Q[˃�54��'?�){�ɧ��*����pf(�b��5u@w����9���˱?J!?ٺ$_��<Ei�v>����c�[��ʀG]���� �FF�|:�s�j���v��w;����ͭ1n|?� q��� �Oe�]�n��KF@vhZSt��:1C21陌FB���T��H`c�ߍs ��R��-���:�n�St���j�}�`�b	�r���/|��t�\�����u7���b��~�a�= �h��ŕ\���iO��@�L�CE���F�U�5���_�%�QK��IiB�4��i�=�b�l4�1Z�0\������h8\.խT,�,�H:_��.���F��q>"��g?�`A��,���	��M�
a���\/	w�Ph�E�д%7Vԡ,����Ή�ǖ�w�����Mf,$q���-?9n_��g�gV,�,�X���k���~�����̹mΜ>��
���S1n6�"�⵳3�AN����t���X^�z�\)��dl��W׭]gWm��m&�)��c4Ӿؖ��6^v���ң#F�\a|��B&9\��t��.t�r�����H�kj�b�b�j���F�&�o�T�j�� ��>�5>5n�RѪ��Œf5.)-װ�r�s��h+�MS�������D⿾rb�+u����"����E#qkʅc�"�*���,��	l!�����̪�f�p�y����?�Օ{��|��1u@wi����r���>>�;5����'��+�Ɇ���ӏB�&�l�a��O�ʊ��_�㱩 r��3u@w��7��_,��Jdu)"��pC@�hwkX��ćE#V:+u;��;�O��D���"��.0u�Ӄ�[��z�T��dZ7���8.����)���b4f��Ǎ��:tQPt���P=	UÑH�\�ZE�� n�p�c�AS�R�fa9vRv�H8�z�Cu@w�I&d=� �+�ݴ/,���Y��N5[S�P�c�ݘ��v�"��.0�B�F�Q��&�%S���\۲��3����ζ{u@w�I���F����7�@�L�)C�h@	�� �ա��:��$ �YW���
4��T
��F�i�@����ښz��~�"��	b��tV�qjT�B���ON����M���,hU�p�ˢé�:tPtӁZ�Z!w&�|�9���,�a�
���J���;��"��9�%K��Oz)#��k<h;�܏J�%I��D�Ӊr�QtӀ|��𚎭������c�0��u����S��]��4������\t�իWۿ�w�Ζ.]j�b��}�{���s�{"Ѱ[$��`�=ۡ��:��$���� t�-^��~�g~�/^�Zp��ngf
q.:Q�5�Ltu@7��p܉?6W�ʄ�/�\U��ղ۪/���-䦃E=*׮�T�.�nP���F=T��R*Z�\�F*�FC�h�-Z�[L��9
u���4+���V�h���:���D�5��P�H��yn	�����YHI�p�b�HhHW:�����i@�ӟ>r��'v>��T�&0	F�����@�X���ʊNOj;�M�e_���.Z�.�nЬl��y�������D�x�u�4��F�O�k~�re��}mq&��h下ԡ��:��&4��g����gB��p�\E��B�)-�t�k���t�fs*�H�ҝJuv����iD�d�X=*F�1i9T[í�}��C�j2�r�X"6�,�(��iDukF+�P.$��)a!4���l� '���b6S��EI�M+
1�$̚�ӽ�>"bn���.�P�:�t`�.&�n�@�fa��ϛ�u�Z��s�X\Qq�L&�t�"��5��Tـ�]�3-uEAw�g��EJ���N�l��%�vjo��"��EH�M#oA�	�hZD���w�ʋ�:��F�ر�a�421��Y7^qew�Rtӈ��`��§�ηs�Vઑ`]�C#u@7�H�b%��պ�8���j��bԤ� ]gT����QG��ܜyy��k ��C��K�M'jZ("��m`[&?�C1׫�=>��5`�.>�n�P�}d��N�	Z�՚�%�Ȭ�ts�N;t�Qtӄ [�وDB�HH~�����eX�	�:{5$;t1Qtӈ���Z�ɗV�o�zsCg�g-w�Rtӈda�J(����tt���1�2�h���D�F�R�V��1�r�N�ß;�:���KН#��f3,\Dk�F�Ro$*�z�\��J�z�X�e�j-[l���Z���~MM-(U��H���;h����� .�+����~��$*���fך�J���z$�'&�~�x����;Gp����Qpp��o���D�7��ը7�`�j��NG"��&bk�j,�Z*���O��>�1�����o��&*+$�c���wcw���4;tQtg�4Wr�RY;�}(��l�zju˥#�XѠמ%mT QG) ����Z�k�5�iւs\�'�N�وgj�pTw�kɜ������/|Ѿ���mӕW�P�l�Lfd|����2Bz����6�W�];���̦~8g����L"�r�l�*>O\+W,�"���q>s%u�c��BXל�s����B��C]�fq�CBP�V�V��,�JX�X�w��N;t�}��_��kך�M�b'KS�j]w��H�C��!i�Z�b�#�l�C�ʅB�h!oYk ���X�rBM�L��x�RI�ī��q�A�x�T�k�^=���<f�1��{#Q��y.��T<)�����r�j����k�>���z�-6g�\˗
&_���|:dZE��EFMע���['����7Z�W��U�	;v�];vؑ#G�\,H��mjr<��ǫ���}e@f�!U����n[1��lU���5��rJ�)[�Z+ۃ|���Cvզ�������a�&�+��p�6ش�f
��s�t袢�D�r��?L���
�C��5�i���������m�e�FM�e8f�h�}��l�G���3��9�� �[�6�JB��՝g'��3$W1�XTx�5��n��Z����v��+�T/[Ut�i#C�㿿2����Xl��:tqQt�o��5��7S���x�dIi����'�������3gڝw�iK-p�@h9����_(Ш3�M�,���X�/C�Q@) B=��ɘ]�f��[}���]V+U���J˙�xtf8��Y��.�P�.:�g�J��|nx��fv��o �F�1yѮ��Mv��I��?�#{�[�*�W���P޼D}�� �xgV-qØ��F�t�q�.UdbƢ1k�S�! �=��*��ʁ�?�G�gW�����t#�������^՟����X6�����}����ŏ����o���iF3Pj��,�w��z-=�K��Ѐ�<� 0���<=5�;bZ��M��ev&Vг��[�zd|셩���\10�Tz��;tqRK,��j��ND1�����a;4x��tղ��,�N����H\�'c�TZ��XCGB���D��҂�D�Bɸ�4"��^��cHǨҊ��IuY<�m�d�oc���J'ku����r�'-"�)V>{�ȧ����_2g�t w��?{Mwtl|�x8�����V+W-��������/���۟���iz���"`�RP{N�Xx<���k�f$\>�5i���Kyj�F���Ӫ0��'|ȱ���{!��H�6���z��/�b�����'����@.w��h�.r�n||�x$�����U���H.f���~������??��������ͤ��G�>y�f��<��q5�p($�K@i4#�f�}a�M�+�Z� �Cu> ��J�a��JF ��UR��������ݡ��!'����������|� n/M�7�B���?5-nͿ��ǛUE�W�'�ͱ��ƿ�oph��itB'|7៽O�J�	G��烋���}�PU7'���,���Z3܌F#�h�<١}o��t2�j,�~���|��9b(�hT�6VuOd�Q�`�:�=Rt�p5������b��ꍈ��Ռ�(l��7)>�Q�E��sv�C�;����jn���W$�&����`�@&d�p8����ס}��=�^�sW��ӵf3�dĭM��B�w�n:�1'�t�'ϑ���n��>)���TH����+��ի�|��M��F+4�ءѱ۳�3~ef<��:Q�t&a����e?��?o�W���m�T�f"6v�X~9R����L�ayw��]Z��wk+�w��HO���NmeUD�mt��z���A���O�����ǂ{��p���48����\�*C��C����_u��9�pJ���=�NN�<3���껕���o�GQ�D
�T�*�K}��ЕD$�w��/�w:�*,���7�J�/�F�B\�wPJ�F�j���ר2��u򆙟-�O�{m�)U�8QL�~�?sD|^]�Q�z��T�#�ƂL8� c�D�Q�K��;����?�����g����M*�H�kŐ��6�*]�TƱB�	���#Re��+�����S
�~ϟSΐB(�p�pږ�ފ�F�h@�i�E}��������9B��ԹR ��H��&�8�[	q���r��㚤��t~�S���q7^�L���@�̄��*\�:�ul�=ꖶ�6��b3��zŰ9���hT��7��K�矾+������]����6��
��Vv�{!�'��D�#�&�]��5����T"���w����g#�PJG��
�O��L�r"�)W�:�JO��L������[^\6b�hL�ճZ�~��~��۟�����}�CV�Ԭ�w�E�Vn6��P��w��P$�,�9�	ӻ�ᰛ])~p�0A�-r�w�ɟst ��~����� E�ݫ�7�܌$�s��5�H�H��y�;��N������"w��N�:��ݯ�o�n�������UǺ�b*1��訌��\ܠ���x���6���n[Cq�&-.���J|��*��Fd��Z��f5қ�q�g��@����#}=�1
-�K+�YꢂG����Ukz�pD�(v�k�8� �`�a�J��kw���s��3���q�|���}�h����]�תղ���%�,�	���e2)��G?j��~�>��`��G�P�X,�t�KyG��B���)��>��K���\)X�P�y���"'�E�����q�gY��3��UF���O��o��s�m��"��_]G��H��"X�V ;�q�8~��b�u��\�j7��V���h��U�E]�(�F8j�������՟�Ǉ��|�9�n�PX:�J~<
_�غU`z|պdZ�\����/��NǷ�:iե#�^���~vj���)����	�|��� .�L��į�n��l*m����m���?g)�������[]q#.쐄��;����������X���p6r���J�t8�E{�gϕ���{�sL�������$����zf�"���,!��(W�N�E��k���Zxg�\����?v��G:g�}{l������K�j)�O��޵�M�� I��,�Gm�./r�����bb�ө�H!Ij��m�j	L��x>x�� �EucH�i_�gC��W1)!����~����1')ɘ��E�]���������������w��&��Y�vy�*M�$��y-�4�K��N�{��,��0��w�I��w�8r�%/���Iu�L( /��C�n�2�)1ڈ�	��=�ܘgPγ����iՉ+��Ⱦ3��{}��ʁ_����Ƣ�]E�cA9�E���iX���	k6�b�DD��e�6���F�+�r�S��3�+�{r��`���B�:�r���?�Ϥ�IK�`��G����ԋ{-��XU�.��֬\2��9�+  �z��<�ɸ��40Cw����8���1,3���7�b.R�T�;D#��s)LE��V�:ߠ.s7��[*��}�>����a��_���&�.B�%�^n��< L=�p2I��|��!���z�t�I�5�S���3�0������y�n�J���t=?D:����:�����v��=��'8]�|�J�x�| �*-U�\��?��������h3*�[A�yV�����ˉ�,m���jV�[�d?r߻ݖoye5n�I
���<�����&J�����O��#��Zڦ�u���?��G��_���96���r٤�ҚUKe	��4�J/T�5w�IZ��m<���'�Tu8�A%C��ql�RM<`<w�g���V-�.
%�q���Ժ�0��˜U+����$!��2/s�f�I��#��g�l�_4ϔ��0�L�SV-H:��H�&D�#}�S�NY�¯͒�O�����I<�@��������SP_�+y��\J�Ft:%7��z����^J�!w[T���^�)1����ڿ������Ὲ�zR1���\OJ��k��Ty����6<1��4mr䄍9`|�[����{�RlXYi�2���|�_��f?�2=OtN�)�Ƣ��4��W�h����O��g��ǟ�k��O��>[0�#��[,q�',f�7�'���V����M��W4��E��tr%�x���zU�C��W�i�,�ՔV]�$�K$��1*�8";y�M�kV�R}���'pT*2;k�h�Պy�gR�V��ʉJ�$!%�S612��p2b���IJ�ftS/���q�T�JC%�)æE�`�d�|C%D'5�za��ݹ�F� ��3���DN͉��9��6�΅���Djg%�/���x�ѩ��'sm�ݐ�@Y�,K�Yh�t��Y��:��C9��╈�'�a��j',�#�N:@`55�$	w�@D�S��5��3�Ϗ��K�X�T� �����/S{��4e�F,k���G���?хI{��o����[���8�
���x��K�dS<}~��m�To4c�f8EE�x�����i*Mv(�Ҋ2�*��K�kR��IKj��OZJ!*-c7������D�h������P�S��qI�D�˦J�ty�(���@wz�J�_S�4)�*��S�U�)kN[���TH��1�P�¸śzZ���\���t/�r7�N[�L��Ҫ�G��KJ�8� S�8b剓�;5�V�\���V�O��&$�,Z��X-�r(_���7�7
ċ�&] �X=o���@Y�\��Dx�o����ޭ=D��B�4na�C�lA���-����@Y��L8����\q�EcJu(�g�*OIp$�K1	߈j!>�,sQm�-�O
�l�&�ԦD�&��������� )��U��GY�&]#�a�ͨ�q�b%�*R�K"��@~�챂��w'�΁�	t2�"�HX�?*(�I*aD~S�n�-�뭒���#5��>JF�2爧gd���R�/%�%mV�����PR�J����S�,��wj|lؒ�ȖTGRzP%EI�).,-���J+ŔC��)�5�e����Qzԙ#싎�����Li���3)+݆%MK%I&,�J:?0����ʩdL!ji�i&d����lF�ҵ��S}��oگ�- �W���B2&_�U!��S=�^Hȼ�+���גQ����I�&$��Rzaz�_+�TI:|d�U?�j�H<.�Ht*#�h���)bG��Z�r��':l2�2>d3�)	QAT�]��V�H���K�4���L�P���τ�z���P%�Ÿ����F��Wď�c�5��@��J��y�sy{"(�ԓ�I���\+�����z��$I�0iEi�* ���$}\"�� �0���k��{�Ӯڰ��r�5v�%�l��yv�u[lە���s�]u��qy����hl�Gh�IW �i�I�0���tJ�DBLDH�q�: (e�&�?�OS&lH�"ڔ���1�W�YY)(Oi�J^ޝ<��a�s�(M)@�%��5eǄ%���&;����:��x��׿�H\�N?��i���%T� ��W)��y�pSR^�R���BX�����Ǧ���e���<DWm�w��^D�1!�I�	d��l���4:A���i��+eWn\c~����ۯ�ڶ�����d�����7�{�u�]�n�g^i�,��%��%�#��B�����d2�d��z�[���;����8�؝���n�珂\ހT'8$΋N[�����צ��|S��Ę��V�4j`Z�bH$"I�K�ljR*_�����v��6#.- �^�q�sjW/�e[7���ׯ�4��]m���Q�bNi��L���C˨e�H0UJJ_���N��\�J��k�v\����E$/�M/������eB6�?n3���X�$gX�G*���4+ͽ�ޥA�L%BX�`�LR�Gz"E����Q�\�� x�c���$W{8uϟ�qL��I����[�:ƣ��Q	��3�
�<8�5�~���H�5enG�`(6ޭV�Y��h�V��Ρ����W8��ύ�����\�՘�?bw�t�}��{�ի�Λo�����f��m�l�֮v�|���Y:�C@��עL���M����&��,~���\�����]D���p~��@�"��La)J�	#�O�J����x�Mi"�QI��� @Òx��B~���z\w��+������mݒy6vx���޺�e-N���I���FX���E�(�ƌ��*�R�8���S�;�F�����j��xCLs��YP6������~��~���~�_صWo�	xkVG*+my.ݔ8�'��9�IJ/[S-�l4����1�&^���+�tZ����XS]T��hՊ�xM>'�9�s]w���qD�7��uLw�U�Y���K/�]W����GO����g
�����UQ�mI��{��I�sL�@�ƒ�vS�U��k��.Y4�^������%�ڑ�{�!�eɼyV�����7){ܖ.Y� UR9≄�ȋ��d�*_x��*Ւ���}]��s3S02E!��A�?'�|7tN��G�'VWr��
�e�t]�nW�����O��G��kV��~�[>�Ǭ8�*p�ȸ�T}���>��Z%���x���������,����Q�����ewӱq��l���646n��x��?2dC�����h�J{�'�_r/t�`��I��}�-��J�ē�T�'�|�5�v�ʕ�l�*+�����/�@ �֗�Ə+L��w��v�r�;n��>{��s_x�2�5��i������l��۷�v��c˖�$^�ֺ��;iz���f���N���UG��D����$^�Tz-�������KKq�ĕ��=�I������$��#b�3��Yh����J����]v��a1�D���tkV��|����u��Pi,�u��694i�#���ރ'lRu�c�>��`�=�̷푧�����he�~�g~�.[<`�8(���	WF�1OXNm�HtY=�k���n��?���w��o�_���A�*ߩX"?2U��5���<OtΠ+gs�����UU	�ݓ�y�Qۼv�݊�N�_���-�ɴk��x�-�LY!�Ћ��_~�A���}���ׁ2������[�W&��{�|�;js,���%�$���:q¾����P�[Q� �DjՆ3)������c��/�^��$�J2U��O?j�O�6(�W\a�.��}Rf����H��T�hHZ��?��z�&9l3�ۗ�����_~F�y��kb*�S�E	i�b�hW_}�۔���|�����x��� A;�YϞQ_���<s�1�W�'A�l}B�d�;�!��V�'*Y!����I�#���A�:c������я��Ƞ�#a�]u�����TIN���H)d<���<t�2]3�v1����3*R���~�&���C����/�b�n�IWBO�|w�L{q�>{��mJ<�U1#\�����._*�ы*7����.[�RQYS]�ͨՒ}��w:������M��âJ�x�����T�߯ɥ߽�y��/��/�N_�����x���Ph�L~7�8!���c���Çm��L�j�:���-�R��	�����G����%=X�����l��c�q�I��yv��c���c����_�e#�E�u��=��Nۮ{Ͽ��ܵ[�_u�*�Y\���ߢ'2%	�)�70+�r,J2s��yi����n.�ԛ�'eF�*ʹ��tY�p��Z����u�,��Y�	�I�*�B]L������e˝O�b�J�1�Ͼ���şe�lŖ,Yl��]��������>ui>~sN�<\{� aU�(�G�Jj3�����J���:G�OťK��"��|ȿ*_����ϛnPP	4��=x�=nM�M^���>m��g
�k����2%�fϞo���I�ڱ��m?|����"V��I��]:�訪LM�޽�Wv��CGmϞ�&�c���n���]{�۷_~YǃVR]7�t����-�^a�sI��E1kՙ���'�v�*SE�PՁ�C��3���ɝY`7\�ڢ2�QT��*�j������A����F�q�Fp.�H�� ��xJ����WTa�֠'J���܈��NwY4����+I;M	h8��D�j��ቼ��۔�8Z	�|�n�z(_��43�Y�� �ʘMY�vbt�^޵��9�LO;?%�K������������i��_�����K���W���?ٯ���m�nu�Zw&ee�,ۮ��~�~���o�g��������C�{�n��g~�.\��ܵw�Ť�)ݼ�x�Tp>�=r��Ю%�#���*�oAG��ڈ�d�����[��:r϶���IH����*�L �K|���9��:���C{:.-iޤ�B%mia��:�؋;w�˻w�Z���L������Ҕ-�X�4m�ذ�|�F�U�AS���Q�(7*6:�W*��C����&[m(O����	�B)���j����z�(�R���9��%z���o��C�;&:�t�	2Y&���|3�enU��Ì�HkE3V��X1�����J��
�n�h$mR^�d=._OO���@��e�*J�-�+�^S%V܊*��1wҽ(�, �3�1���Nq��M�J��~`�gT�jt|�A��GOwLcL.RS�K��ފU�-?0,�O�<���e�0t�Έ�E����V��*�S��9<2�~;���*`q��![��~�@}�����9�S�~sd�)��-W�Yh������ރ��L �ڬajU$ԊS��������,�Q���8�m¢X.�f��5�N�����c�C��T�*Z�Xpu�@�y�E�8!�* �e
V��D�'P	����3�bɬL��ԍ�����!���+�+ź-�3[V��Q<�t[8�tJ@
��i���nD��9�t����T��GV�$q�jĝy�_�ÿ���|�f��^3o�e�51}�RUq\~OS&��LJ)���K�t��81ne�8��H�A4��O�t�u�+=z��5�#,$��ňL�t�hi��s�l��EV�����_؉����|�$S�Jv��ٟ|�lfo�T�69r�FO�jq�r��L����SS
ќ-X���ݳ����{^���>�;t��"b2��ۮ��~�}�ZY@��Ƥ�~Bw �����u������59�c���N�i'TR�T  �#>]�R�i [(�.������CG����`9W��D�h.�gP��\��)�B��	�����66%��Jؖ˯�o}�M6����w���	+�e��ϯK{�Ծ����5�*-�=�0�����2���]V��|A�)j��`�U�mZ��r)�kA���,ALz�h/5I-��#e�-{܀�}w\k����X&T�UU�B<[<1U�O�s��p�':7��Th&��v��GUغ^����=��)Wn����a���=v��L؋���#��Q�udX�ö�А����҈9S��	UA5�/�|��� fP<����R�)��q_Gf�D�E�;3g[֮��{l@���'�z���F��0s�V�O��E�얛�Y�b����iSLߪ���j���_ҫ�-�X�,g<�L&'�G>���S��O:!à���sl���b:�i�V#�s�@K������G�y;F����H���ǂ[�SZ_o�͞5�B��j|Ѻ���1�x4!�&��XW.�x]�'�X@���u�c�w5�V>Wٴ�i�s�ʥ�=���! ��}�
�Ӻ�p�B[�|��Qںfαf"#@��u�\��*��Am�Ŋ@+2P*Vy t�A�:a\�I�n差��g+S�684b;���ö���96j����7Gm��۫p`p¶�_��<B��o���l��J+"�OW�Wj�J�q/}���b�5�U0���2��1p6*�����[33������֔
��W�k�=�,�o�PJ�hN�
���LF:]��V%6eJ6d�0+ Ǘ�^�D�:A5��S��O����Ii՞l�f�g-��;�S�rK�h�t:����1jON�g��Ǝ���ÁY)���F��|��ik�9����s�S���qiHf��Z�Y��C꣹Un]�^XA\赎:���L�&	:5x~���`�[�h����:k���ö}�K��s��K/����/�d����u��A;v������L��TJ���T̊��:uBu�CPn`�����$P��&�C*`fә�����ݗ���E��ņ4�_�H���e��I����@�A`F�\���<?([�W�#Ċ��%d^Fs=��[(7�"ݳ]uϕI9Ǣ�s-*^�v͔궺LV&�d3�".D����en�G:'�AQ$�$���!�kY@I ��˟���Y���m\�ք*$/疀3[X*�K�Ukug��%�0qp���I�9ۚ�]�:5�`ƹ�\���a緱,�̀liҎ�i|����/|�>�g_���mhh�u�d����`2Me^���69dC�XMK'�&I-���?c�� �q9���b~����������r�i4GZ҈����g/w�{��	9��w)}|�jW.#�6�rٴ�q1x�9|Іeu�.x�$sD[�Y���	<91f�#C�g�N��f�KͳY3\\&赂>���m!(���������"y*b��=�W��%���>k���?�_��?!��N�?��{jy���L��S�7兯^�p�U侦$�	s�����:%�>V�e"~�,ʜ-��s�s=�%�VQi0��C "�خ[�)�F����7��@��&:�
R����TDU�*�*�\(�YR6��b�����"р�D���l�H���j~]�w+�_	�t��������'�t��T���?j�~�~{���3O?a�}����l�k4�~@FLb�2�#��D�5� �_���qS���)�a�XGS#��RA��@��'�Nk%�2{���0C5��+?�����:�
;~��'�_�n�gPw��ȟ��������c�\~h<�NHsCߙFP���p�w�W��TY��N��{؞x�{���m��OK�M8�Z(y?����߽?�J~��u�0����X:`7�j�]Y5����;pUX���:0q�E�n���A��U�s�C�5��i>q&��t���-�D�tj��������(z����-���۷^b��]��O���/��6{�[m��ٖ�2�=*I�������e����w'-U�a:^*̳L����q1ƫ` :_0Y�bz&1�%��UaY�m�����܊v������dF	m+Q�e�IM��E�&s�Bj\y�҂1gV3-��I��cJ[��NJD�;C��&�����\��_/��e%[�(�32�s2�zz�e���K�1./�%�i�% .�chK�w&��aY�����Jz���2�K2�zgX�L/��z uD�p�3�H��%�`p�A��DC�%,˥^V�T�ݹ��.��Y�g �Ӛ��SU�ū=ɒJ�j�ť͑�RCUH␏4\I��͢ c\��bͲL�H��n�����G޼�~�޷�Ͻ��޷�dkV�S�I��>Ȓ4��ΐ�����T�r^��?'r��p��_�D�C�V�5���ݷ]o?r�����W�[�^go�~�}��[�G��n�z��#,,d����`q
����Ǩ«�Rd�o����1��[��S�P4ϡi��,ʦ%��!H�d
�1�@�5@T�_I� �,��i+AGCBf{^�N�ƀ4��I�0�gZ ����9�zx�^�oH��@4�����1c�Ӫ�d�ˮ�W�g��5B��F�X<s��5�cV�9�8s�̙�4e ��N��-R��H�Y�pAL� �|>�s�]q����}�F\�}SA�j��&�$��nIQ��ͪL���]&�x��mó�����R홬�ۮ��z���]m�n���ڵ��k7�O}����`�Y�	�@)�y=�V�(�3\���ΉKȴ)1�`I�~�k�g\�7)-�����>{�;�[��dss1��Q��Yhr�z#y�b�L���l�ҹV;)����G(��G�J�buU4���L���V�#L�X%?nS��:N"����A^&`B&{WZi2_�Fl�ɡ�*d~4�1�@�vL0 Q"1�1��c��+�z��$���ԙ�8O��=������^b���K0$i{f���q���Ԕ�����\΁�ŝ~� T �|�����L9�&�� ��W05�A珯GN5(��σ��%i�0�O�e���<i�LΥ����,�ٟ��
h��Q��'�Q���ذ�gXVU�J���Bd'*a^�_�˪��1�����[W�%����[�0d�f��"U[ї����a�j뉳~��ڟzq�ɐ����eu"F��w���ݍ۸$�Y9_�V�[�̿KW.��XL��K���>5(�3e����g�����ތL��e�H�����]�V����Ǯ��R۸|��]>���貫6����|��y�Ͷn�
�J�*CRғ����UL��̜g�3f����m�ܹp�|Nz�-��pL��=%�-	s�lܸ��*�w^K`���	Kf�T�N�ə]���6�AQ���n����q�2�͛7�i&�����@H�GZ �w M��>X�FzÅ��=��v&и�F��T3�� ���fϱLW�%�z->c�	*��.�r�(OC�n���%6�+c��Y-�]s�����gK�ϲ93��[n����6��2_ezv��61>h�֭���~��O�x�Q��@S�?�5���Y��m����g�=V���@gQ|%�E�	#��S��R�$�dd�R;I��wR�e���.�o=f�2!�"gUR�81f͒�v�(&m51i+ϱ�3{��F�)Mr��u҂7Z]0Y����&��m������m[���6��s�Mۮ��3��$d�0 =NT���k�z����w�{��~���-۝Q�A4�3̈́�d"��]U�
S��a��;!�a�:uRɌa\G`oIC��Yj��'~�co��O�t��\���ɥ��r�v}��8�l=��t  s 9�#��\�䜜�t�q������n�<d�^���~��v�{�g��'����wXO�)<���#֚FG[��,����6�r�%�e�*7!���x��8��⡪�v�6[�j�����n�I�\>�fkV,�.Y1��Q�W�Vӗ�5GF�įUK�\����^��x�Y�2�]����7IR���;��.�':��tBW ި�����k2Rb�Esf	|!��eYF/���a�&�+s�{%��{�ݯ�gC_�r��x�y;�o�-�v?��f�w��K��W�؄*닟�G��0g��$������R9��T�,Yfk7^f+W]��`ry��6K
!?����؜͘9�Ғ��i+�VCa��1��X���X^�ͺ�fY�Y��$��\��k�	M��B&Ǆ0��Ô���	G\���#, ��1G�1=4?�МԋkK>@B�Z�4��������1�ee�ۂE�m�����֧z���4=�>e��w$�CwMW*a�7�w���\"j�/��5i��͛3Ӻ��v��aw?؆"b3�;)e�:G|�IYS�g�S>I��%.�;G>]0S�N7�W�pi�yh�WSP��B*Rۜ
�LAWkغ�9�����w��e6��&��P� 2�W�3�Z3�b �"��W]~�4h�v����X�TdZ3A2�������c�0/���<`�|�[���=�hkl���qi��S�	�w��YK,�=�j��17�S�
���GFӖ�p�,�헖U�����DM}Dy�2 ��`M�7��D��#�xME�~��?��x�bw���8���i�� �/t�����4�pb���2Am Ht�}}�	7g�.�b)�pi��;^~ɍ����|��'��~�Wm�\����-�����}�S��[n��.߼�22��E7/�b/��x�ty���|:���0�+�:��rG���_[^��	����@�=�Yprh�>d��^��R~Rw���4@7wKZb&E%��&��'���G�|�6l��-R����+���*M�8������*�lǮ�*B�
j�	E�O)s��F%=f'�#�����5� UW�\$%ƪY��d�l���2���	]�(��z����x�͜��©.iְUF�vjQ^�ˋ�
D��O0~��'�	`qɍ�;|���߿�����|1LG�8p��Fٱc��޽����c�rϡ���� �{ b�:�r�Ŕ���PB�L:�yЉB�쮝{lT����`ZV�2��<�ˮ}�՞Gt�5�ۛ��v+�����v��^��N�XY�����$��Z���=)6Z���j%��D6�T6)�'�G�;zR��.Q�03�Ԋs^#�{^���~���V1 FH�2s�����}vT��XA�����f��ۜ�9���0���������L�J(n5��/�;b���?m_z�)��}�3��K��c��������ů|����g���g�m�m�G?jQ�'�H� K�+�`���$�%�Rb$f=���v��X<c�X֢�R}}��]`��o��W�h���6�x�e�ڲK���E�,�5�"�M��Y8�Ъ�T2!�" R��;yM�Z�s� x��9��&�����F���
��a2����>i����nE{L�r��gb����K�s=����'��9JΧ�7�&O��~=}ꐿ�s����$�(]�-���s��)��/�`Oo�n_��C�~��m�᣶c���?}�>�O_���m�����O���Ӗ�@8lR��'��=lW.i�fչ<g����v2�H�|e�AYGG�\c<T�[|U����3&b�dM����s��<Z(�%Swe��>� ��OJ�~����������r~�|9��LVŕ�M�x�h!1h�{�=����?�U�}|�*�4��QiƊ���62&I���.��'�̐��1+�J��"2�����⡊|�~[0[&�>�t�y�Y��/��2MVX_����/��8j��ja�>i��v`�Qۻ�[�����ؾ����[�a��C�����Wv�|P�>��̚)�ݖ-]b�_�A��J�'�v��N�b���a&�)`L�؀������0!	���` ��t��9�'�D�a���>o&�{��3��#�L���O���Z�Y�1���Ȩ=���7h�`�[.K�\Y-���2B�@��Y7�G��s�������xRmw��I�s`��!ök�i�Qe����v�M�f]�7{��ky��z�$�N�!���r}6.k��Д�ͧ�l/�=��U-NM������+WʄCۆ��6'��o�Jľ�:9o��
{�;4re���o���BV���~�>a�?��͜�g�����u[��U�6ڬޙ֛��u�_�s���������VK�Z1�6�}�Z%%hٕ��"�{$ƅ��;&�L�F�
j����L�떨L��)�~�2�WmV2f����箛=/��t�Mn�ࡇ����G:��C;P�q��b
�����B̣�s�N�v�5���e���?�[�|���޻���+Z#��@t���A�̜�@۵k��C4@�~���7!<x\����&!��������y)=�|�Ew�w�𮘴�4����>5�||��V��1��_e2߰믻�n{�;,�P�D�m�x�ya��������t�Β��'�q�P(C�J��m���i�yu��2-�\�FѬp��qӕv���l�7g7d�Դ=���kO�`_�֋�����*������~�V�).��
������+�˲��<�9�.��#ЅЩb^7����c��s;�L��mc���KVڂ9��X��Ͽ�ӭ��e�$�T���&�1�8����OI�9 ]�2 ��L/c2��V�)�[�Y�e3�v��9�,�[TfQ~dȾ�8-J��UW]e��-us݌��1%� �6�����C ��Z
���3���!�y��1���_���t���=��A��z���kջ��O�FJ�sᓑ���Y��I�l:� \0���,������G�>_���n ��t��1�oH,"�q_tǤ� �T��|bv�eWؖ��q�uX�;8)_��v|� +'��E��@3�+�W�T�5�u�(��7jM��
���ss(i��H�ٙ�$��$���������,��wb�^�v;1��b]f
AE���#w�l��7Z."�Jm<J�OkC.yA@�U��_���Cb��n��?���˞x�%��V�z�M%�>��&3�Q��ujLR�l(�6�J�(=cL��i���k<�6�.Vcz�
�_4�SFҌ�<T1���B�Ue����1�4�&S��b���A7�f`��̙�NK�7��y����Ϫ��'O�Ƈ�Sy7F� ���9rȶm��>��(/1Zг��3�?B�U�>�[�j��
��ɻR^@�;��(3�
�f~F�7��3�_��9D|�����:t7 |:t��>^tlL�{��G2�K���[M�����ƛ�w/0�-'�[Tu-�B/�tj2����GWV�:`�c p��-
nV��������������Dʀ��u�+B���ѻ4�nk}��}���?��[�΄�>�-����]P��HT�[S'~�?�Iw2/f�˲��x�&u�e�h��W��g��DΚ�>�l���I)H:E����&n(A�Ѓ�H��P��b&e�I�:vDŻm	ؽYL�*Y� 6c�5���갤��CG��N�/&�$#�nҎ�8l�#����#��v`�^�v{t�o�ԵCv���(��ǎTz�g��<���0ß�3�� ���S�Й@���f  �t8R����y�'N�pG|4�2���>?����<���5�#u�8�~�s�G0��w ��A��2�U�#�[sU�� �8�� ��Ä�r5"*�e)���+��
�&6.��Y�P�{��uJϖQYe+K��������0ď��$��:N��1I��
�
���H���H�%��=3Y��]���l���a��9뚵�"Ո'�R逇�M�4��&��RY��*����vݹa�EO���D:X���(�I��L���A�P�l���j�rѺeJ�������}�BM��T��,�co~�֝��=:;`�}`�	��?л8����&��� .���Ԥ�X�d��$�$�]۝+�Ԭ�lɒ%�ɦm�����`�(�z�G]Ru�2I�{'=w&pO������j�˘Z�n� ���@ӝ�_��߲�� .��	�I�����r�q��}K�}�-�m�Y�Q���0��,|~���j����k��@�8��Ji&��=텥� �*�t*cY*iYc!�ר0h��&������)��T��~}}.��/��;EzqT�T�hٮ]��+���t*斿T�,��5*�8���`FEL�4�2abU�cl�/��CN
�*C�unꙊ�\�ȼL��t�je�2�v :Cd��> �5k�]q�[�j�]�a�mڸ�6o
�u�R��x�u����v�uv�lӥ�lӦ�v٥�2��6��K���͛o��[�֮�b��X��&&ƝY��L��z�,	=�LNs]i�,�YqLv�r��vaV!x���J�I�� �_&�����f��e8Qf��v����"�rts[�T��:�y��|HF�,Q|�b�[b-�1멡��,���g��~ P��I��f��&��S��79:T-X����S�ͤ���:��J�}KA�3�m���8OtΠc�5�vL�!T��|94��L�
cG��m�@�nݺ�n��R�����h��XA~J�����:\c:�Y�biHL"M��㒒HX@��V�QT)������3Ў�+�wRM]��}% tV���1�.��K�)5V�J�)�O�[A�P*KX�B���}&�m�8���6%���Z�rAڴh�¸c(�r\L��OO�q=�33�J"���vu�����b�����e;�� ꘉ�u5�US=�q=�J���`bV�#�\����{�.M�g���̀6���]��=0��:�h/��X����W9��KpF���	Y�8�|���bEY#h�dW��Q�������yS�!Z������-K'ҨC�u HWo�J��S�^����h����mW�ۯ�ܶ�_h�Ɇ@��x
W&�r�du�u����]��It���"��]7N�쏈�a�/=�:1b3�gZ�0a�H���F��-o�۶m������kV8�2o�,;~���8n�tJ�H� �BR���@��w��z�b�����I�r�ߢFpc:b������f�����N9M@wz>?��a��sl�e�O�V���{����}�R v_n�����_�
�G����w���[D�����r:�uL��{���b�ab�HiWf�c#�֓��r\&�j���qγI�i�V:��g*��Gڔ�_:Q�G��6������\zb{ڵ a��o=)�׍J�ӝ��˗Y�w�%�,�;�j�w��c2�F�F,'����l�KO.#5���bɸ�iKf���/WV����1�7��U	�X�h�n^o?����;n�Ү\�ʮ�|���d����6&�w��Ch��s=ok�϶m[V�d�+�ES��7��Ì)�':'Ѝ	t�6�a��~�E;|l���	�z�v���잌�e�'-ڬYO:n�̰�ء��$��:�?���Z2�SC20���`�%0��x~lLڎ���'�IH4-#)�z�t��Pٖ/�k���6����-�m����P�+n�f�ۖ�/�yI���8E0�LE���oU����\g`��o!�kK�;��FMڈ�k�8���� 1�9��@o#�f��mf�p�q$>����������%��^D ���OՉSzo����!{���T2su�����![��r���m���m�(ޚ/H��&���sg�n\�%�Ҫ��(�NX8��$���Lհ,���dݨYUAJ�jv��k��w�nKft[JB)��Ed������.\`���6>:�|�ƄmX���ۼZ��%&���+�������t����\f�A��dҊEs얫�XV/�N��LYO�`�°edO_�a�ݰ�J��>��HO�(��Mv��u��t"�̊F�b}ٜ�m�#���t��5>b��x�̔�4!��Y�t1�I0o;c8�9�|�7
���7Q�:�������s�䩽,\�y������4��4 #�	�$>����M럁��=Qi�uU�^Yh�p���X�(��}�������F�B�1�)&b������t����Vʏ�v�;��>X�G#�2IOV���21>�ɘ�@O�����m��^�U���23�Rڍq�I[=���e�e���cr���#��n��oX�9�����t5��=��9v�f����K�6z�}��l�����[��Zº�����l��a2d5����mW�u�\�c�JV�A�^I���ڮں��RئxH��˖٥�n�g���L)���#�v	�i�ؕ.���zR�2�|``�m�l��wQK괪Ur���ngnr�s�����S���Q�9u�i<wvv:���3ɧ��`(���4@0�|T@�p��JL���Aw�>C
@	� �*Y� ����-G�����o�t\Cc���#�<fe�����[�ؖ�\c㥆����=���4���DR�l�/���-�؊��lÚ�6cf��d�[o�Esg���c����uk���ظ�v���|�mذ��F����p�4��m�o�;��d��'ܜXVLJ���5�8��Ƚ�9g����N?�:\6�^a�]�J|$^�;�B�f˼|�|�����9���Y��>	��\o���&�ֺr�e�Yܞ���	�q듩���џ�Z_w�M��|����౽6�7)����%K��2���{vXNy�Rq�ͤl�҅v���j���.�$f�U i�C�v��I<,�D0-����L�N���$��1R��S���^/�F�
� x�E ���o��
ӛs�H�!�">檟SI}`�R'<q�[	�����'�A���!,K\:%<�!�R�i���W[1��Zd�(_vX(���w����t�V[:�=��6oF����
��^|���m�Υ�q;v���eMYNlV��Y�}�AX� �o�",Jc�Ѧ���zT)�o�ҥ2�뀒K��t#g=;c|�tΠs��!x^a�I����@1y���؝+�ƭɹeC���dF ����c����MY�]��M�sSv��I�3#%GxTi��Rc�������ӽ�w�F>�+����u3�iP:T*�^�穢eʈ�ĩ��`.v�bG1�!�1<g��)0H�s�q�ϕ��M������:=[`��BQ^0>�q ��
�)�ZF^h$��-ӓktJ���>h#��$���k�s+�ݸ%���J�
��с (�!x-�FDPV!���d`��M���*��ҤC��I	�����G����^xѾ��Oٶ�W	�����;p���;�&�ܧ�Y���M:�6������Y>ZL��QflF�UB���JL��
+�:��M{���U?���p�]���� 1�ҍ�U�$�F�bC"�"�t ɻ���y�%[8���YV�,-s�'�ew����붌̈d2�L%zw�خ��=�Fr�,W�1�G��	L���7- ȼ�����Y�=O�����������٘��Ü�� �8�I�Rϔ�g��;�����o�<�ѧ�
����H���T�}��q|g#���\��5T���֬Z���z��Go0�y��=3���?`�vﳉ����y�}���3��$i|�߭Z��V�ZeK/s�S�b��{�cc��zA�1�θ�t�u��%_C� s3����+������Q=������
������A'��ʬ+{>Ԁ��bPaUbUP���m<2&�AfE*k]rx����r��JH�I������q�|���޼0�}���/~����~���ɼˏ1���g��=�����~�x���!�GeRH���Μe[/���Ϛ�6Lu@�gB,C�0a
���U� ي��0+����O�1�Hӧ����>__�qq�u�K@�ی�e��z�%�`2�'�/�zb,�4)��{��=��#���pqζhR�N����a�H"_~���ig�A9'>����|j�m;0����+�[m<�طl��Q{A>�W��M��W�w+I>�����ڪ��l�޽��/|�u�Q9<b�tN<u�S�KM�>��������ؠ5+๽P%�ѣ��к�������AYL�(9?�b�f����z��
�s�H)4��wf¡>)���ן���I����-^0��/�+&)ۤ4X�l��TmZߜ�vl�d�~�{��W,.�ʠ(��d����:fS%Ij��~�%��YQ*L��}{m���np��������hK&N'd�VFm��a:.�{�v��)�*������vŖ-b
����H�a$U�x작 �0+cs\g/L~{&���1������@<����O:\#�35�!R�.}4��P 8N�Y�wߗ� ɗ@y0���6ħ���>OO>�O���z�� H>SJ���?.W�Z��VXgwB��c����I;&����>)��e&����j�CCj�}��.���w䨽�[���~rr�^ޱ�^ٳ�F�&�BY$N�ǎZ�@�z�2K�2n~p6+V��=�`��O}�a{��;uM�C��q�R�v�ji�^'��*��fţ�ӝ���'�3�T�R]XY�{��z�����cÖ�v����<�RKV��tW��(-�l�D�^�w��ꓟ��z����W�2��/���*31��)�~�<��-���T9�|�@^o��ʷ�6+v��n���ö�g���t���%�P�!��4\G��E�0	���xG �y��B|� �q��| LO�xHP���rHѭV��uN�;O=���P��`�v���i=S��\ �G��q�'��P���"�<fq� ��/JhP ��}u�����r�cq����T�a��'�ԓ�4z��ٳ۞�o���/�ޣ�VS['s=�m�X�8Yך�t�K�cvV�WXn�w�N�W�x+/-����V�nt�ibL�۷g�%3Y�̶��q�h�q�P̎O��3>m_z�Y.��şly��v��1Sf�]��pkp����Jޕ�"���*�ܓ/�{[8�t�C����ni��C�vD��w���ȷ�_���t��Ub�m�Z���2W�:�YGكR ���ي:�e�Ё�fO�:S�B1�*Z@eڑ��7T��İՆ�����<?O���$��!�+��¥h %�b*@#y�s�<�Z��̋V$@�:gH��U���u�?A;9fmi���z�?���k�S,�*i�B:Z(�(#q}�����{9�XE�I	!��-�p&���H׃����nL>��zRmP7>b����g+>��(m4㖜9GV��V���RmH˙��\b��Ln���{��,���t�y���	S�t�@�Vq�����m�^صώ�N��c'�����������=���v2/��P�NKSv��Uv��%�`���{�|���V�\�V��3��e11_��3�G!��}��g��o����%�b���#'m�$����!U| �(����:RK�#g�l$��a�� ƻGՈ�g�����ۭ`W@�K�^���HyD�᠕�b�Ҙ���e1 �5x�.�t�}�#Q�`��̐�b�&Ī�vfb�+�`?��5�F��- ���0=@sz&�@<_(��t�����ÁT�q@���ۆx�ۙ���d�ӁD����y+M�	�Ӓg��QV���29�v"�'�J,��"���S9���/���66<f��^�A���m���rn�喬�F�W�I��A�M�����ZAi˂��ɑ4���[��8+��pM\c[�D&!R�@z(+�	�}%Tel��^)�&Pn�xY�x�5�9�O���d��Ȼ�����-�Z0�j�&
��.����*�<���,��{�Ǣ�5n����6^Q�l�u�Yj����֓6f��䬘�j�E�q��*1��	���0�0E�ޮ`M���=��๊l̆�X3�1��>f6��DӖ�ܘ�:`� zN����!ۙ��!��
��a��pj(B̂�a��X�IX�b��G����0	�O�+���`d�v����isDC1ݍݾ����F�H���$0ٺ�����y;r�+�������Q{9^�������I����ɺ�����)��'����|>��Py!I\75�#�B7c*&|�}���b�(a%a$�Ԣb�T֭T/7Sn�g�r6V�[3;�j2)�������Q��T�S�|��K�:4����ܧk,vv*�+q�i��U�CLڏ���^|��I*�M`e'��*�Y�v���*2���l�BQ��Y��T�!WE�eʒ]?ƁP�%۟��:;7�T��z��B`а0L}&Ӹ{���3�g �fe���\�Q���'���}��� �ᙎg�G �9�p�	��k�3ɗ�����Plt� &������Ð/�����6}�2��.>�����'�I>�s%7A]ϐ�0`f����O 0��e_
��ᯤLz�A,.��k4��E���ʣ�		lw]`L��eu噜! �2�҂i���"O�"B����A����H8-�ʭ����[f����PX��^T�������&���	t#��Z���jw�����q�X����h"?)�_qˊӔ6k(K@�j�?��:�k�X*� L'��N�U$��f_B~c�x�]��,p�����Ys��57�`[�m�7�r�mڴ��Ȍ�����$�i�X.`,�y3�w, ��+�3%�
���}�s�k<K^���e<�2���	t�x킁<��o��s�C�I�D��`!�Q&���ƻ�V{��k�ӓ��FD52�άڋN�E���֫��k��Ѷ]�m�9��Rt����rT��Ħ���Bb�~��y��[Hq?X�	�Qw�F`r�TZm&�����傴��k�fd)T\*��ސL�pC�@L��s�]A��ߤs��7�+:��zݮ��@?��%5��	i)�Q�q�a���{\��ebz��$�0C��&��uI�&��j�O�֚z^\㪱��luiGէJ�
���9�/������*�|ޒUv���k���{�=�;�x���~I�J�'�4�����k �ip��"6L]�i(4@	L!ʁ��F��J��T&mݽ=N�3��7��ҳ`z zc�^�up��c+9f�SB�Hp�Z`���H���R�,��x�(�瞸�4�B�u��@��k'?�r|�:H~�ӂ�	Gi�&���xK�������v�]w���~�� �����veOaE�BT�sc���|ڸZ��9��*U���ã��ri�X9�
ME߀��eT7iH�jՂ��p]�{����ټ�9˦��`M�P����g�J��NI�ё#Np�!r��:?/tn��j�;`	׀�W�H�倆lݲ��c��~������Ƚ�s?�^����n�j�-�W�N�9�"�Y�_�yt�ĭP�:�CZ3]��`S!V�5�h|M����
_z�=aϽ��F&K69�v8���$=϶�r������	��+��Ʊ�g�g\�Tv�:0�F� ��`Bb6A>/������5�e39@����v@pε3�ךg�������<G��_�� �ǖ��\�5���:t��ڽ_�5k��!V��-���+-'K�&��I��b�r��ښ�$���b2����)'x�#��0��L���^8��|�V��{�f?���ؿ���ٿ��{��H�̙eSr�-M	��/�JbN�9��<�9��Ό"S
ף�VHSQ��^Z������o�ۯ�`[�ۖ��m���._h������l�̬���dj���L���҅�،���Dq��<�ä�h:��(L��`����h��C.Fd�OL��؞��e��]x�a�p��<^�����y�iX0++���	�(=�0-�>�#e%�r���|!}|?Ҧ\��f陠���$�u��)3���������=�,��ξ4!YA􅨡�,$��|y�n۹w�� .�X����s]b���I�1��LB���/g"K-�fZ�a.%w��:�T��?�HW6#�U�y=i��-7����&�鲕�e�L[=#a[Vβ���
�M�h�l�6�s�����@��SX��ԏ�E���Y�r�s�Xu|�[פ�Λi��z�f�B��)M�-����Q˕�lYwܮݰ®�b���dvH����bɄH٬�����؄eU����;�_��4��$3`�v�B�y�b)V2�@������D� Acr#Ҡ��:���A�o���ɫ��Is����H)/�r����8� ���<�ځ���??�����!5�k_����o�o|��
j��C���n��{_�eJ{%�����N�I��(���;k�c��g1's�(M[T���s6�e��'�����q�R�	K����\�l}ºk���5����7ns{��F�1id)V%�����:7�5��HC�� ��RQ�{>˴,�U�^b��YT/��NY�V���[dj�ҕ���$�K7؀��ެH��v�%K�_����7o���2	��}w�Ůٲ�֬\do��F��?���+�P������ۇ�͚,�}�̀�afO0��ىz�	K��������Ѐ�y���A�Ą�K���3h@�{�@#@���k��4ȏ{>����H��9xޛb�|�������#n�lF�_K��۳��w���S�P����n��kl�%��֫/���,�{�q�}���ڼ�>�b�z��m��{�|�-��g�o��~�#���t���Q����m��_%���RrK��q�T�4x��ǭ/�k�Q���ٰ�V.Y�x���J����<]���]���(@��}�Y[�`�[��J4e���6gمL�¸%e�g���9�6#����[q��6�������W�K�5K�:Uh.�#�ڡ}��f@������X �N\/��Ǒ������.�իV:3&r�9hIu4L ���:�3*��0�]��5gh&��BڤA�0l �<��x�	�'ڐt��yI7?�#,��K���y�8<�ɗ"�/�&.む�@�0&��_#�n>����~���b��Q	M��_s�%A{`��}���t�V{����MR<���lV_�F��7�`�W/���ߺM�v�F>��V/[l�Xqr�܇z�y[�p@�R��Q+���l	Ͳ,$i���������.��K繥d�F����(���q�';C�����^'�e/S ���,�sD=,b�V+I�W����W��
EK��9��֟�Y�Tt��ȏ�uWl���q{���G�ޮ�]&�Ȳ���Ygu��o�1ε���nȤ�c��۝Q̲�LZ�l'
J����ȧ�k�u�� . �<�W�I	0'�"=�����z�s� ���ci��@��z���
��4#�� | ˽�����f���g��1`?߅ŋ��h���8�<��嫭��{=K�܈�{ޕ�p���8���,͚O^9	7�Zsk����/_��9z��y�9ۿ�e:z�>��O8��~�f�|�
�Δ}�o���ؾl�\���C�	��])KK��7OL�����ߢ�g-�*�eţ=QY)g2$����@>�"�<�|_tN�k�:��F���c�ˈ� �����f��@�9�H_f�'�K>Y~��^�,�*�ܹ���t�����#��3���k�v�`F�s����hH��ah>>���i|�K�w�7�������o|�{��9�0�?�䙛����0�ͻ��Hg� h��D �x= �h9�������kM_._~�,���ҥK��`���k�G^S��/�&�^�����G>���&��9cV)V��m_�̧������'>�W���l'��L�;d]��2�?��ϸ��sl��e6C��o�����q�Z�3{@nF���V	�>g���L%�66:h���y�s�K{�e!d��n-]S|@��1�V�����6r�Z���M�)W��8UI"xB~0n�$k��<���;e�h�\Jx�[W6i�]�,LYUwb��)`l$Tj����a���3;���ҕ���mӕW�C�|Ԏ�T��}��������Ba�b��IB�w)�9|�=�����x��Q{�'Ni8���q�����C����73���5��$�@��`T� ip�3��L�9�c�Af��s��mJz�|�\���v�E萁  D@�2r�EK��ɬ?��L�:�y�v"�s	��o4K���%�%�8x�=��#�췾i�<��~�	�?i�Rp�'�>�s���k���{�u�����w�,[�r���t��y��m����/}�v��o[���v�?�zBٮ�=Yῗv춊�d~oU�V<�c�xF���lO����e�ltl�:�\�Q ��Ўg�:�U�&'W�3�{s�@Q�u,��⃏�����!�����Y3m���nJ����D�LɬLf{l�qK{��7�y�T�K6�aH��ʮ���c��]�̳O�����И����а�� ���]LBh�%�6V/��&d*4�\�1����"���\��-��'1`�@E��0��=�8�E�L01�5�����F�y�]Ϲ[A�ʄ<�516��
���L��V�\�ܗ�]W�� <�l���"\�z`RV@X
\��#����9���<C<���ܧl��j�S�=��G{ʭa�9.���M}�u�o[�z�,�b���|���q;)�O*�o�~{���o?o/��c{��G}ܾ�kãc��+;��^���	�(�x����Ɔl��[�p�%d�N�r�.7��R����5�u���}]�Xb������D�W����-�"͉R��x�HX�<ѹk:12��J�x�M�ʫ��V{�����{a�1�fB�NVrL���|��}��G�K�<,[3m5i�Xw�5��a�p<�gbV��a"��Ĕ��+���8M�P f�$���������;s����Ǉ)y�A`^���YZ㨉�LBo��� ��ܧǑ@0���J�8�7C9��|��0j� b�3��w.�����g�fȼ�W|��8,`��ƺ�LM��6��y��Q�ԗ��nNՑ�����~�{6Z�iW�nn2��k	i���dv�č��>^��f؈�1Q���BC&�4�T=lE6|LvY�k�%��o����@T'-ߐU!>�l���j���'�.�Q;
|��7�Ż_y�E������	���.+ԙ�U9P�-�b*�1���s��Fe8]�����99��$a�H�z�e��O~ξ���vx�l��vF+�����>�O����n�$]+Ҙ���|��[��g�(�G1m�&�]2'e~2)Zf
ӥ�N�`�� &(L��0��&|G�8�����B�9"�!��<� �O�{��7����	X�����ǃ�=0}>�O\甇t��bb��a>���Cc�����ג�y�D9��o�g ����}y��I����i��O�I�HV����_��W0��� &�a	id�fjWT!��\�K3�
p�dN���P����8/�����Zn�7����?&ki�d�e�}��oڟ⋶�ؘ��<���-�9;�eJ����_�{�sZO���oOϘ��\^�i�����a_�e��%	6�kC���d�6�;SNmR.3fdȆ��U0+��JȺhʩt|�j���$�*&`F:����L/�Y��.���}�O���y��-4q�ҡ���N��޽�U�������؏��Gd��NhI��i��c|���q�9��| �Ã���4za���g����}�/�F$�z��9B���r*7ѵ�@! DwOZ��s�s�S� �r�K
`!�N�9�Hޑ���mDuV���N����U�������M�Θ+�ד�^�S�f�&Ci��t��H�e<񥧒��+�t~���W*E'�Gc�K�ܖ���qUY}�OJ���Z��ŞY��w�Fw"j�g��Q�bц�5�fm�rV5�	�銣���b?��[,*W�:����Gǧ~}C.���H$����ɧ;>>�*�IߗU�Gh`1�I����xҎ	l��*B�^��$��^n���+d"ԥދb��*+�!��Y�ߧ&t� �xT��ŧ�(���<H<>LO�%��a���c��27�Ya����|��d�*�=0�cɟc|V�o�|�����ivo�)�7�`Z4�q�p��Ayp�����	
3PҨ�@h=��4���|�AE뢵�(���"�%.qо��+���9�`t��N@>^@�R8]c.���j�o�톥����N�����M��n�����l����d�	���G�!C��}�G)��:=�~:z"��[ڨP���3����z����{`A��
�jJ��Ф��)Ygl��YR��.��,�ʔm\6Ƕm^m��W#�F�,�.�O��tN���诤sB��
|�d�z�ш��6U�z����e�\��3-,�V��]���У��8�)IƜL
���u��a�8EzG廸��b�L���Hu�
��D*��k!7�G!&�t�D��G"�<�I��ژ����
�(Z�����e�>�J����,z��ϛ{>�����)�|zޔ�7����u~sD�2懩Iy�=�&M�I����g�K?A�@9�;�������ٮ��$ ٢����+�C���w�۪�);D�T(��ym�]`�
G�bqj���(�v�@|��Ϭ�U�S���f㖌�,�PZ�h�`��A�.�t �X)=`������붢��/%�)��;�̠jV�nj�[7*N׻���~�tN�k)�6уG2૗t��E��P���X!���um�KN���䬆<�����6푤g�OY�sS�H�*�a�ߠ+�df�^S���E��ʪ$����G�����y�9���T`�p��P�9�Y��7L聅V���JZ���_��	�w ˃�32���. ��U>�x���i j��"��}$ t�����M <`��t$.��(+�I��>�ף�՝'V}����Eqk�$d�����m߽�|�q���L��p�|�!�a;�d"�V��z��d6���W�$`���+�J4Yo'W�%_J�]�c�\�%���rI�{LZ�8& ������\'!Ew��it��@��W�Q)B={ N����t��Q-Z\�+KRHb��y�OH
�#��Ś��l��#� Ve�`|O��(�>]Ur��t�/��A�E��8>�*+�E`5>�ES�+��n�6C�>2h����cL.4"�#�(ظ�l�.�=a^�c�A�9�����S��0����dmΜ��*��.sl��9���V�`��Y΄Fh$@F��+�&��VA��i�q�ԙ[=�Q�@�B�)�H��XE���?qԎ;l�cç ���L�����:ϭ�k��"�yA��s'(T�X�5Uf�-�h�C���'F�njjq�7��;,���2��䥵�o�sN+҂��C ~:�q�OS���l�X����|?�l=iř�X�l�i=��}6�eI����2�yR�.����]�[�=���j�+�{�s��XQ8$ ����O����f��fq�r��[6�O��^��x���wٻn���/]`U5*����Uբ����3�0�`���#��(�iL��mq�(I�p��l��&8�މbJI£�OZ���`
�@nB���G����9� `@�A�PN�$A�UbL<�c�1�&�7q}���>��<��" ��_V���g���ƻq��s�r�6�9���,�C�4(��'��s�&׈ �4� �g&l�aX��?Ơ5z�o"��\I����)�;��O:�U�������=��,�DXn��e_�ڕ]q�25K�'l˚���w�a~�[���C��w�bVε�Ԩ��u�Q�JGW2��C�`���y�s��G��E5U&k�p\�zɉ�c�|�l����f?��w��Wo���X��2}�m7�w��[�X2�g$��ٌ^TI���D�������J3>�w�I��A��3]YN��?+3&j�cEI%��)�ʦl��%6o�l�0��iH�K�y�jP�� �jR=ó��	C����g<��`��s�C���s>Ήϳ�M�L��iS&�� ��Ep�U6�&`b�סQI��0)ɛx�����!ι����/�.+�/+�n�2����>e�����6F:�<5��;%��`	����!\ �����7��؎�q8�gK'R�% }��wؿ�~���Z�~�r�v�"{��[��}����[n�\&my�Ied�pWTv���A�^�5�9�i�Os{J�l�$N6i�����5���09h���K��(�ڲ��}�]w���K��[�K��q����`Q��c�l��Q���2Odf��N������u����+J/��z]9�4��7޴������gJ��07yyF�q߈<�?���8�L0�7�(?��k~%�an��x��M$�M����Ngr*䙘g|y�P�0/��?C�<�4!_���σ{��.��Jx:P "e"m��	8o��c{p�D��S�������x��z٥6o�ť�%�$$�e�%s1����ЈM��-�=a���Ĥk{&@(�s�L����܌t�뮶�o�������e��(Yw�`{����n�+6�qf�sSd�5����S�a���#�#�(
� �ax,X%ͥk�]��6�Xh���6#-Q���EO��%�rv���� ��|��|i���g��K�ۚ���'�eK�j������L��E�����=+N�؆�+m�UJBP��x�!`V��g�?��������o}��E��g�����3x" `�yp�����}��
`E���0I131Cy���{r��ty�k$��u4�x�r�A��C��q�g)7qHa ����O��wz�@�g�.??��T�NѸ��I۵c��������;����I��z�u�	��C?"Ss��Ev�6of��&�l�o��zsi�U�U{�Z�̙�h�L"�:V�,_b��F�2��'�Z�:n�F���)K�Ƭ>|�z��۶ڲ��ܷ��Ŭ�<�`����m����p2q_
Nҫ!'��T���sr҇�e�^�Ŗ��Py�z!;y�F��1�q����)�7`;�C'�\�'�����[�+.�-�mp�4��E�C�u�1�M۶	d���9�l�@��_�ʮ��*7>��g�����%e;�{�=���g��W������Yɀc��7]z)m눺�|�ZR\��9	�`h��{4��B�
��`qߛ�4�
�s�̉�s��K�����o@��de�a:���{%phD�M6=✹���/#y�S3@���/�;���u&�F��<����3n߱ݞ|�){Z�w�>hE����e�����X5&+�+.�w��-ⷚ�8rخ��
���w��ҡ�횫m��Ŋ�~UU�����7�t�m^6�j�Ǭ/'��<ac�G�^����,æFY]���Q;r䀅+[�|�]{�Z�K�|*QE�M�\}pV2���y41�IӉ�#ҳ�)d����&;�J�$�r2����M�u	c� �Fej�zIvtR~ ]����v_r�%���O~�����7�s�|�l�aO<�u�D%u%���cb���t�F�:`#�wە������Gf,+��2}��0��f���0x�6���)`��D> ��I�8@��ɂg}|�@���=4����Y�I��ϛ���<D|��׶�� `�d;���rȼs0�fۛ� �w���/��{��z��C�oL4zO٫�<�	+.JŢ��_�t��ˣ�L�t�3�(ȵb�f���M���|�����/����w�׮Xb��1?q���V���}�_Sa˄�����jy�����2�,̘a�h�q�L�i3�ˆXq^�u����UzgY:�w��@�&	��{<0]Ԗ��0!��GI������4�78�����;G��^��� �4<7�@����|�/�%�M�8t��c��T���A�͊�X2צ�OZEדQ���$��<�Ѻ$�z��O1"LJ�S&Q���{��&.G@�r��!��0�O�"o��N�H��\�� 5��3y{Y����I���, �ݜw���~�%�a\�'�#?� B��'_7>���|Y^+��p�u>�L�@2�U;��ۡ<�U@���0t�k������d�/�w�����xh֌Y@d��5��˶��J���u��agf�Y,\�baB�����_��	�~�rcAkU �s��Ô�A�]z#ؿy^�wN���Pf и���Ą���L`6	_��u�IO�]�>��'s 6��40�_q��q���W�j��^�_�n�3S��w�y�=~ܞ�yB8́��5�Q.7�.&��8��ܧ�ܧ��n'�s�@y8�gyO���I��"�`�'mޏsW��~p����0�DZ�����gx�|:�e&�|H� a>s�@>�)����,�צ��9߸��?ȗ�gϬ��"��G���20	�4����tBT�sB��('q�� ϱ>M�u��s�=g�7o����-6o�<7��駟��.�̙۔��8$���R�|���z@Z�M|��~�>�/w��R��+�s��&VG�{��K��	�F�k?a'��%���V���ٌ����h�=N7w���#���O�O�d��+�]�wȾS��c��_zy�=6�v�ݽg��K{n߱����o���#��˯X�X�C����/Y�T��JJ:6lbd��q�հHQa�U ���rI��L۬F��3���sG����	���Ѹ��Z�Fp��t�`)���|�L����)'�8w���`L�r����ע0 L�E   �8r��!<a��� �C�S�D�LM����~��qxΝw�3�3>>!��3Ք��(pR�j�Pܪ��E��~����[YP�I�ґFC!�cq�\�'�������Ĥ�O���cv����q�w��i��*�M����}�9*>��>=}u�=&,��o��˾��S62�7�e�]�Ԯ�l��&i�,������J��ӽ[�'���	ב�X�j��@�/=����������a1@�z�p�%y�c�&�	&Ҷ��	�������ֈ�r�cpx|�`GOY^<�>�,fܹ�5�1��#�g�!�[<�e���ѩ���L�א̗����ꕋ��)�-]�&<��A��|�g��>�}:�c���U�HO@�o<04�������G�`@�D0�P�kć�y>*��׈��$�3u8��*G����к����MY���|� <K����E�����'����N�����{ �.1�[��O[����s�ںl���6w�*럿������j��`|��"���Ę9qR�:f�L��s+ď���)�����r��x�hB ��R��La;���ʕ���Ն���h��I�v=3l��)��7��g���OyJi,_hWnXi��2X�K4��óS����XeI$��(_V4����{ڎ�T�Ꞛwdg�d*gY�T���o>��>�ůً�OX3��c+&��N��j1b2c5&���*���J7�I*�u��t`ש��Y��D���2_ �q����+mْvɲe������YD�?
��Gÿ����Ń	�gЃ�<��@ �g�Bh9����&��+����7�<�'K[ �֨�'=�����]��= �Aa~�s�}����l��״�K|�=|_��M�<��H�՟4U(�cO<%�9��֬]m7�t�-^���Xc��vR @�b�a��\��T6��"[+�$�'��U���h:�WX@a�ʘx�R��E�,�A�F�;q��;�V����\�0��=����W�G_�i��Ҫ�mê�vͥ+,�VT��F�\}xv2���\epΠ���u�V.��bþ�싶���R�q)&�˒L'd
��_�m�w���z�%�}l�"�>YbJ����V�yӅ$!+�奛��zq
���^s�'���;�Jݙ��DT:c�z����Qv?�c`��=t^�8]�\���p��f��w���:S;x��|��gj�\P����V">��*F�y ��Z{9Iۃ5��K��"Ҡ��A9�G>�sp�����/�A�G��z#�e&]���?&!��S��0�}�%k��ڨ��]�G��Є�L�����a��׻OH��/OH�a�PY7��R �5�ߡ"Y������	`���?�����/mw�;<��v����W���HY~��ۈ~�4n[�.���9W��K֢� t���?��=�[
�q�SI�+b�z\v�@Q�fl��o�=n�|{�^�Q���W쩽'�d1f���L�?�,����eI)*��#o&VPe��o$�������.f>,1U�R����L|,_�'���{�}�a8�3����k�R��A�W�9�h���f5�6��o�$��$���B�� �O��4y�#���`J�]��˗��oZx�8�����U�	��q߿��/e�u�z�ә�ܹ�Pca+ʗ��B<�������
��qU��iM�˺�F�l��J� �'����ʹ�L+�c"^������0��qln��|dؾ��K��o>o�?��}��6R��궔ܠ0S�$����5I��ćB��=��+�?�VC��쩫*0��<U>e�s.M�m��L+�{-�3ߚ��l"�m#%�ԥ�l����!���Cg�SH|�13���l3�;.�2��W�Kl�RY�j-I�5,���/���,�!��V�|4�g$�3F;y��4 ��0"�P08��{�m�ɇDw>��~��c�V9H�<Hۃ���9'.y�<��,f. �F�L�Fˑq9R�E�Rv:����=�D��.� ��6�qm�w����&e.J�Fc�\Ԧ�)�qt~QNʞ/Hk���]7$�����&Sa��&=m/%P�sX�	���f͊��	�Y��3��T��ʙYf��lL�I��<_�w2o2�,��-����QJe�N��>�k��6lq�4.f��A���Q��b�<*K�v���^����HV�S��ǔ�rZ�4\>�0��5���@:�>��s����"F�DE#J�	��%-���a:_ �1a6�-���y`ޏ�u �B���Q7̌OG� ���CY`h�130N\?A����Eh[����26�������sy_���4I"nP'�A�9��=�`Z���Lӭ��UʖU]�dSjs�/*���.�N9��+�k8�e�O���nY��&]*�i>f�:`����4��:�`ߜd�&krOL�g,��{�17	ۭ.S���)i��
8�\k�u��e�5T�zU��&�n@:�
az�vT�,����n,��g(Hcxe�K��)=��V�Br��
��r�<�׈A�t[���iTV: .�ؑn�.۴��Β��� �j-׸G�f��-��ѹ��H¤��,*��}�/��k�Ɠ����,�'���������G��.� ����M��aJ��֝�����"L����R����?Z�~����%k�ْ�˭�o�͘9�z���T�������E�4�1�0�+������A��	���;��*�}��w
����l�c|�c
���Ղm��z�y)�����lJPG�	狕Tgpߌs���4A��N�b0	�:6�l����f'9�o�zO�Ҕ޷ac��T�	5Q�.��ׅ����H_��8Ƚ�{��H����\yU$E��H5����N%?&��l��n�f�z���+l�+���-�[uj��&`�gf��:@��9�`c�"�1�Ό@#&cB��2���.�arQ�i��=�ӛ��
Y�g# ��g���i���{�;G��eHX4
�h���h3�m�}:�m|�7e ]�C9H�߾N�Š8,�嚿N\G���^Y��q�9��I�.��Y��7��=�^�׍�/f�!m[R~W_�֝MXo&a�/]+^� �s7����`�$��xt�P>>�fDi,�6�f�\�!<���&��4T��ZT��-*٥���M[��-[7��V�����R�sS� ������6k�P7"�x^�w���B�ةq:��NLU푧���GN�ɺ,R��/�l��2�y���m�ۖ�+l݊���6��j��1�=�֗4boD&��!��b?Ƅ[J��Vޗ�|$�X��dLH:��!����	<���8�a�_U%;����~��}��^��뽼l�&:`l���g ��$���L<3|�`n���@��o�� ��Ѩ�I��R)���1!4N0�|����g��-I0�6e P �.zWF1��r�����Wi�׽+���]|��G$K>}N`F��T�Mnf�0�Ԩ�mxh��8d��?h/�;b�UՇ�h�I	۴4�<��v,*J�6)R�ʪ�[?�]X���abz��r+�"��b�	�q�Z��-���n�Ҷ]��6_���.gw��jC�e ȺP��q����U��
��k,Q+�kߘ�N2���+� ��	S�J�~�T,��$��5P\�ܕ�W�[��kZ6<i�ʰ�I�ly�n�r���M��1LB&D:��������儳�1�BJ�(�-;�2���c�ގFA"�����{`�=v�����|0.�4�!�o��3�3�?G{*���v��1�}'�a�@7�%>q ꊴ��;c��Y��ک=�����y��?�t����'>��!�� �H/&�%�B\ʀ&�t�rμ��"��cT D6��~�a�}���>��ƃ�w�� �M����
zi\\�ai`B��|'�e��C��+/����zYZm��}�q��jLX�:n]�	[&��Vۻn��6�^�/$����)`�Ƀw9՛r~��@'�4���x����0�̄5K��M֢^�G,gK7��1���F�6�Xl[7�S��a4%;��
;n}�[�j�-�;�����볅�l�$R���2?�\-�������@L��%љmB�vgs�&�f��1aR�wo{��F��i�V�K�eeR*(��L^i��	���' ]��9�=�7:��#=@��qe4�E�\��!@��Ǒ�<�;A0m�>����]�#���C�\#ݾ�3l��Y6{�\�9���������^7LB�f�t�>�Bg��~?aC�U%7�Y����˷٣�T�����s�"����Nۊs݊�t"bsf��/�,�3`�P���1۲~��W��ۢ��mْ�֥vo��Y_W��P�[o�b+�v��P��)K5��&�:x���l��v��M�S�x��΀
��cS@I�)�
d����kl���-�ZFrid��ǭ8t\/,G�0f)��U�o�Y��K/�d(�����m���yۛ�k��Y����mW^fKf��[�t��{�[�:���z�����]!�d��e��s���|�᥾��T&]؀�<3�������I ���9��0:D�h8�c���8�Y����T����χ �t��� &������1�dg� N�,> ��~��2�ڎ@���� �����x����z~�w����Xc"�/�ʗ��T�n��M��7�nw��F	�^���+���-�(#_l��u�Ͷm˥΅Y�t���w�<	g>�澼S)X\��e�J[<�Ǣ�)7a"$`�ɊB�w�#��U�̏�ƕ�lŢ�r���.Ca�8�p��n�NZ�iW�2�`:��K�)0��V�<�z��Œ�
e֓XR���JV�ٹt�z��J�n��|��-��o/?���=`7l�܎��c�A>�O�L�z�����m��9�X =~���fq�I�$_�d�P�[%/�@�����B��!��>x�_�!`j�㜊���:r���4�Q<L�`洧M�O@ F_4�B ����L|&�}&>�!.�L͐L߄�)_g|l�Ș��"��� BLJ�E�`���/����Q�B½�x��W�L��*&�! �tU~�!]y��g���m�>۷�e�̠M�8h�\��*�G���n��2����2IYV��PE�C|��A�`�W��V~�27�7&���K�d�L�R�v*gI㊇�G"��U�4��)���=�9�N�v���F#��|��J����25T�>��<�ԧd����7�,�T5�X.MZ�\�C��ZJ�352*�t҆������?~䠽�ⷭ05�C4�[�!U׌���b�
[�b��]��1�7� �� ��C����j���&-��#�Hσ�s�g<�N<�A�p��Y05}وC|���{<�=�$ a@�Wb��!.�A\����<@I�9�=��sZG�yG�-��3��k��Fy��3�6+m��նx�*�9`��ī*�f��}��\��M����	;|h�u��6t�?�߭طk�}�s����.�����$�%�C��"VLX���v
�ƭ��g�)�,+�k⹌����m���yW������|�9���Bô3�F�7;sqƤ���C���0K�(�t'����[n�'�|�.�|��۰���w�_Wv�y~9wD$ F�a83r�&��0IS.��.������r�*�j��u�T�l˶d[�gF�&p��Ð"� 	�A���~9�~?��^w�����vU��������sO����4�>���_qLH���}���cT���뒒Mg� �i�6��_��}��_��w=���M �r��l|�/J5	�s=��@�l��}�M�`��/@�0 !�x�`�>��>����k:L.H����ob�)i	��G�x5x�Gg'�x���$S�B�k�������0HC HG���ϙ�́��o۱�>��/���e��GI�W�_�W�JPwu��s�n>�z��;{��"�����|L��{���vn��/��˄L��O������L�����9�v�7�$-f�Sޣ�a݈;u��ե�G�E1��<���P��$"���q?��V�	��#_��KZ�l�UƉ(�z�ҙ�]��)��L˴���po8�<&�?m��߯�̞y�E;���vql�^}�M;�Fx���lR&�[�cO��y�)��9s��E�)��0Q��L_�'H f� CB�Z =1��\��&���a6*���M�Y�g��NXV~��L:�@�-	��d7nt��w��7�C =�SW����H�a�f�{�@;���4�dX� bL:�"<v�b��-����|e5
���6iD&/�n�����O?gG����}������{��!+�Z���~ �&f��^{�ɧ읣�[���̓��nj�+�vF�g�+ǚ�.�r>LP��3����Q�׺�o!|I �+Y�'�İ�q����A�j_7\iً��s��[�U,��VPc�y��d�w���3��
;=R�o��9{����f�66Y�\:��:���<n�\���=#D�#�6U�ۻ�S���&G��ԅ!;��I��5��J�ݐ�Jъx���S���o�w,ˬm��V�;<���	U�%Ƨ�/�H�� � �D����y��⃁ ~��ȓ �y�A)�qho���1AI�:?�ߔ�����FT��@>[��x�Ҡ�� s���P����ĘpV���*���j�Wf!��Cy�Ku{���x�z�t�u�.+J�9}���}��R�u1�
�ݑ�޳���JxNYIm{����M�d+��S�쵷[Yy���>rⴝ9?�R`���/+ϟ�U]Y۽s���'Fm���}�b�l�B���~��?x�w���>�����o�j�J�Xb��l?�:��0N'�~K��w�F�@�H�t��.�N�w�z���-1K�a㵆%{����Y-��#g��ۏ��:j�4{�$��o�줤��!�'���s���ή>k�2,���U�-�0߻�>#�%rҤα�{�U�
r�9�spd��^ ('�΂R��R���a��E��&X�~�o L�Ϲ�c�a�SF�5?ߚ�l�hN�Cs�s	��ӅL�;0$Z�y����F�7[�A�@@W-�� �� XN'
�o�7��8OX&_�١;�ve�$��3j��57�xYZ(�m�_�����z]���H���11�8�d��O��=��glx�b9��tE�lS�0S��ɲ�Տ~b/���n��[K'�LaYk3��yuq	a�+�w�bqi:�PQ�"�=��KvQ�sd�ONۉ�j��I�4�4�11�GN�������5b9k�9�bi�`YOZ��Uz�X���K�2'YK����䔈�����*k��x�&�!M˄��b�ĕ]�]�w�l����[��PhIa	��8D��.v����V�F+�,H��݉%���\�w���0q�Oa&b:S���$Dӱ���bUt��2����0�.3ļ�G ��HOO-Ke����3"J@c��j���1�����~��U �FP^�kz�l�����EgF�֭^c[�n������b�ܲ�ڮ*|zgG�&|t��2�e��2CU���"[�0.��T41��'.�"��x=�F��hJ陫�3��nz�]iB�=����	��ç��O<��a�*��L���O�k�VkU�R(��b�v�9�ܚ\fI�kX����a���i��~�H�ץ��O�S/�m������?�7����m���z�^:tܪ�$VZ��2	Z���ɪL�Z��cr���L5��od���#ӡ�4���� I�T7��+�!�R�6o��}��Z	bD �0\C�!��B�~hs�������\���g���k��o Ԁa��^�0[xp?ia:xh��OZ��f���#O��f���7����zŕ�J���n۵s��*N���|�vf���\�d:8���4QM���Zh3�q���Ov�����A�h���5V�v�o���߷������������_�O�h]����hH��P	k6I�錷���G�Ea�/;��  �@�F������D֒�6m+G{���`��z�5���)�r
�#��NE�V��a ?iEH���������Ji�X������(�����|�v�ΈH�ukȗÏ��.؍;�ۖ��a��oBB �0̿+�϶a���{��������U�"*�Y�<C�ѓ��������A(�l�%Pz)����}X�{�`!o�w0_éb�WY���������S+ze��H��b ��� P�@X�/ho�}aìf����:>I�0e�}�?'W�b�_yj�c��$cU?S�b��)aL?�LN��N��j�$w�ۦ�T2rG�7Z1��[]6�\e3+�Zt�&k���0n�ﲕ�q����yk�uYjX�A��zNZ
��2&���s3n&�8eL� 0]�fd$cS�j��(�RY�2Lj�w:�7 ���Y�(�º���
���d+���Ό��f՚b⣇؋��w|�;}�d�ê��N ��W
�`�J����X��51�||�+��߉�O~���=�!vޡ\�	M���ތ�c	��zC�N�y�wa
p������z�"!	��*�څ�L�zz}/P��E���֭�I+�ͫՕx>��Ĕ5���&�����7�}��A{��A}��l� ?Q��,��P*W�<�$I�c*�"
��B�ԋ�o�z��0^mT}ZۦZ��FJS<oK�D�i�e}
#�_�]�K���ǅ�r�	~IaQL�5ַ�,�`��T}F�L�!W�|�a�&d4���$y���L���
��ef�[b��)�x���"`!�Y.iK��C�01c"Ρk�)E��YX�3)�Ӗl��c����~Ӟ}�q{��'�'��I	�F����,c)�D���~$��|�5~3���!M�5u\�1�=m'&`Rs���W��%_��[|�P��uMo_�u:�1�w�"�����luH ��X���ŭ����6����=,�)�!C!0	ڑqC�����%(7i���F/��G%��5�;v���_�3O?i���o�K�>���.���n¥�谋d���i��j6)�@��_��jONs���Cl
�p,�zs��x&&�n��Ye���&h*!Z��*2)�o)-�RK�ba����d�K�v�Q��i&"�� S�����lVK�6Ӗ��l�@�﮴qU�ugT�ڴE��.i&*�FC��bs"$W(�����`���U%�
�ni���%fVk����`��%k��m�/<A8�Jr����)$>�8��B(����q����]�t�!�@c%4s)�3�xNg es�*�������"=�K�P;���i�v܈U2�KNl����H �hÐ9W�X,���qt5�an�F�O`���
~�n�(a��P([8pM]+U��ȓ�o�O'�k#�C���A�l�xQ1�Lj��)1+�����i�l�mMO�nٱ�nں��v�,Z�����20�k���ڭ!��b�M�D!hϥ�E1����#�	�fgdKg�L�V9i�}��ؗ>u�}�K������?��W�o�����;n��9I�1I7	�Z��Y�kU?���=3蝒�Q����帕�5'��|FNj��"1�Bc�xԶ:�J��!�֙��p�Rߡ!!R��s� ����J䀊T<? 0X����D<i�\�R����K�;ދ�4�
�o��M�/O���&�^]B�4�kH��zQ���z�w8Lqb�h�Jǜ���~����^B�q�Rї�y���y���ĳQU��@�,��k�XMr�VO�ؒoޖ�����R�&sR�G�0�8=�Uo�#���-:��z!V��-�i�����o�����q��_}�����E����}k'�.�c���A0*>�����E1�>	��0�,���n^�t�,�v��i�=��O��?~��۱�6���M�������~�!{����$���tF��_�a$ͦ��t�(ҍ��,�,0�!.����j��
��b�)��Қ�U��7(R��ĥ���p�K`�ف@�- '��ǳ[t��ء�x�w��脰��H:H\�	BmE��\��)̃��>�2�S )��t��7�7����Ĝ�t�����W;|��1{iك���ޗ��ȅ�څ��t��▅��3�0i�8�K��d�wIX�=�J��1�	��c~oW>�6�{�e�V�u]r�/���ڢ�Vt�o~�a1�}�wC��Z���ɚ�H�/=r���g?i;6���S����2B#�3u��.1����K�&��� ��d���W����m7oZc���YuĪ�g�9z���Q��[�O�y�=p�^_nі���fV����/�Ic�Y*N�/�^��	��zY���Pm*X��r{:Y�2��,�i�!��d�� �wF�εt�H�P���8#),"vT:!vbx@�B3�1�G�L޶ܰ�V�����>�¢Lҵ"-�.&`��B��z{�m���q��w�ɱʞ20A�̀�!*L���������,k�l�Z�e�Ĥ�v	8�[P��L�&���=�!����J�:0�1)��U�]M���Y/��3��C�E�?c�gN�*[R~��Ƞ�"�jIڿh��xV�15h%�z���I���U����o}���s������E˷��/V����dm��u�}��o�����_�HXX�І�����Wh	a������׳�+&��,�Z�^z��]Ve#��=���}7���Vu\H�]-�6!�w�wa�OK���]i�uY���Ysݳo�}�c�����ٓ�햛w�ß��ݰq�]<o{o��>��0��bU{��Oچ�l|b�J��
Y�����Y�m���j�V��m[lݚ�6!��'���+W��7�A��q:�A�0`�����R��\^�y�4��������<�/Q�� DO����7��hAb�l"��m�l��. uD{�!Ԕ�&�|�|x�<ю^7�KX���4W� �3u��Sj�o���p����릛��;l��]ֽig�W��ں����^{�_�]�w�W��>_��#�o�ͮ����/U�i��^���>��'m��;w�L1)�aS�pמ����7[srȧa�Q��gY߹[�\���[aG�?f��bnk���7�-;�YF���fkQ�	�yzM>�bt	��tH�� �
�!���WZ�e<���m߸�f��u˨���1UfrD����$H\�c5���~�%G]u�ļ{�	���g����~�����A��l�6�����f��[�l�]�7ڙ�G�cҪ7޸E�ZE&�\9X����s�}��|���+�/
]�D��f���z��i�=\��|F� p�Y��0:�.)i�Gzʭ�����I	"��L��ob֣�|b� 1'.��3gNK�1���?L^�Ѳ�1���K����rL�,��2/�����u'��ҳ��q1�f����O�����=b�rTm��0Y'b{���y[�Oz'�΍��(k����� ܺn��Sm]��O�ݷg��-	#�4��Ϊv�έ6���_sN��ؤ�;����L�P�&]�W����-��;Ⱥ�c� D�?m����E1]H���M�΄TzZ�ę`�TL���2n���t*aIє')G�*	��e�pN��)(S��Ǐ�kO��q[��W�:h��|�ΞzOZtF�����@&X�.^<mo��ߎ�wX�T�z��IF�1��Sv��Ii@�I2; �&��!d~C�U�����k��IK9�f��H�_�.z�N��ߤ% \��1y7�fe���\�~��̬����#@Z4-���འ^pM5�\Z~E�u|n���g!`����v��Y{�7}��}�����ݿ~Lnäo�p��{������i[��Ϟx���ǿc���aw�v�]�9:t�̈��5џ8���/��/�｛�?���`W�����~­���J�̰�3h1�(}�Y�C0�	����@!A�hEf�obF ��3�t�����[�2.�M����;}JS6���ҜH���j�g�Ng���o|�^�o�m=�}*���Zӆ�'��v��1t&0����~QF�M��z �����8�?C`�On��I.��=|��|Y�<b�6E,\����ChP��{av.z�;AF����+o�N=T��;�Gj�y���I���6�<CX^�?��ⷧQ>l}����!6�.}��|��#v��9+1CEߢ�3���`���ҝ�̤�����d)�9]�t�޹��~����^C፭�=s�J��Gb�Ù?\C'~^:ڎꃣ%�E3]!�zϢ�npp����R�.� ۡQ�`][Uҕ+��+lLf��Ș��,\��N�='�p�EY_3�m�n}(j[�l�J�"�6l���1{��w|haͺ"Ԍ�e��6&"nZ2��uu3���ʜ��Y�&� u�pt2�_�{�MxvdSb��Y��S��%�5�l��/������	ǊCM3?=�B��ZA):�����1��ς� ��ͥE��ć�tN h[ӷ\-9��lh@,fm�a��U>�v_�a������k�۳?y���q�mؼ;��������=�����;GlZL6]�Z��%혬��#t��Y��ˤ���D�-	z�y�:?�3�ʕ���4Wf� �D�����Ho�>��E�XWA0��Y;SI�������?p����l�@������m�e2ʩG�7c�\�/n�͸}��w��o�ޕnj0�ң�b��)K"�|.k� ̀�t���9�:)7Ǆ0��T����0��-���-�*پ-k���lzt������&����n�i���o��$3h�����ge -���wU`ro��д���}�{�j���ĝ�B�}��[X���^N���#���3顄�=��i�x��6Zl�G��{#5k�
ކ�ڏjT;3Wd�!�����,N��V/�E3Q_�̒-���$M�%ga���T��~�A�K>�2-�F�����nĬ�[i���}��g}��Ly�~�����/ZD�#Ѷ�3�r������:���K!�} �(@�w:��,���0aʎ��`?����?8jEi�t�ߗM��9k&�vn�hϾ���Ŕ~j�l�l�@��*-���I�����3�'�X$���rÎ?#{�GfdۦJ��!�:Y�u��$ە�]�w������rlH��C�Ks��: $� �qb�����G�=q-]��MŮI�d=cH �F�נ�>�Z�]-0��05`�����7dD<;̡k&'0q3��,�ڨW%�fl�lӦ�����$H'�e�8����5;]��I	�V,X+W��7��m��dQ���E(�;AM�����^�����=���3[�h,�n��_V��/�.Z���V���2��=�5�)d�?U- �%�E1��nRAB��n���b�T�^>��=&���OߴC'.�Pi�NMT��7�w_������vN��L,-D%%E�m�eI*5`"��YؒI���k��&%�L���Ya�Se���Y�����g�[�aB�ٹ]Z_#"�U�"�-��%ܧ��~Ǘ`�Qb	���C��3�G�g�K�6_��\;#��R��>#}{^���c6]z}�4�G�y������e����B���P�2O��,)�z��t�:	D�*��"�=����]�V�<U��9��B�hDB��b���dE�Y\���`o�a&M�:��9o��Gn��߷׏���e;3Y��?��S������0j�L��ʗ5.L�/�9�D��l�%e8`���ه����L !��;UJؿ�wj/<��wY6ڲ�Đug㖑Y�A��p�Y�##V��D�%r2�Ү!�z;+��c���^iv�] &��h5��%�stb܉3!�ӳ]+�i-��ʸ�4�{�3�~��IISf�4���`۶lvS���pR��?��ó%��n�� Ӓ��A��9Ӭqi�\=�^��c�����~ ��w\#�`�#G��zL�=ݶv��G�VN�m*�gr7�3	��Ba��I&�Z �]��x8��M��1������:�b�Q��E����D�82h+��ϱ];�	ќ�%�p���YbU�/GG��9�����ޣ���L�W�d'�3��o���F�p�b��Sb�'W�[%�m
i��i�'��?���s-��%�&��ʴl�(�(c�VU1\ݏ�m2������2wl骭��~�� ��!=��;�f��Ф�F�@�-=P�z��m����ïX!����R���.A����'m�p L6�11�y�>
0^�G+�mLV����J2�ܣ}/��Q�����%����`�Y��aB����a]��E���0��>&S�,<�Ħﱁ�����oN�΍F�sP��xGm.넉�t����x�89*-�l�y���n�3V+4�ҹ�/p������|?zɋ��w���>nGgV^�:u�����~�s��*�:�lf�63�;{W��=��3�"!h�aw1�8�����=U$�0Fdc�$���hu�߬��YE���LX�JWz��+K�1��Se}��B`ƶ�	S�L��1���R�Z����Y����ɤZAt4���ů��Y3���vf	RЇ�rΙ(����x�Z�vNf�{��G׿o�R9��Y�Ib7EU.�&�7���A`s^Bn���)A�Kc��G�A�^1������}����c2�o��3�]'��>1�pa{x)�ejr\�$�}�����s�Ɉ�w�]0&Y,�����JE'U�v�E$MǪ0�V.�尔��)�n�F�_,˝IuY3�e�b�i���o��vnӧ���;��[�˵ZB��t��-
1ߤ�� �xo���l�l�*��J�����d��$"��4]�U�z_�l0�i5���4�н���,.�KQ�F%���*���,�*��L���4>�qSN�şSѼ�������ѽ� ���ix$!C�o��7�	��>_�Ο1�Hͥj:P��E����D�ܷ�Z���4E���P�ؚ�N?���wm����'�ڬ����R=��>����>2i$�<����]��}}��o��� Bf�����S�h'��&_��x����U�^-	g���J��K�,K��5�1� g� �M����L�=Zպ�LF�lR������3�vi#}�C0� ������6��p��Z�_��˴�=��З[���i��Q�,L�(o�A�_�Z��Ǩ���gs��6����D��ƬqC�:i�cC2IՌ�YU���r��h7���h	I>6��]�|Ii-�)af9�k�c]��߻��tJ��ly0`E�`%_��r���*3f�5Q�a#|{p�s^`5{w��up��w;��3+v�U��d1��T�s	P%�)̇�H�>���!��-�
�/;��{l	���ZT�Y`+t��A������c�k���a���6j@т���,���N��g3-��`�4-�)%���ԅ���C�Ppfn
�<g�8Z0�$z�쌬"	�vq�b��hQ�U���+0L*����}�G�,9�-j������Zs�׳l5%�f���Z�~��;y~��L�UF�[Q���{v�����k�����-��I+M�Ik�Ʉ5_�#�F$���eM	� 5VC��i��BNĩI�F�;�s1,c2L��*�ct�Ȭ(�O��p0f�
��~1R��k�[qT�!�6iɿ�|6�}��<Z�-��rv��N��NX�s������Il�g���z�w6�S�
�_g{'�@H@��]�O��~|���Ӹ�cQ�����q
���'�M<?0����W��@:�f��`nVL��|��d�y����Đ�鵈La)J�$��#)���mdP�9�=�cU�Y���@(�$�J���������V��V؃�v��ݲ��y�m�a�h���U�)��񒖒صi��y�_z��L$K��3�s�W�����:R�=���J��	a�����6��;����ֱ���o��1۹y��+f۳{�w�sȟ�:J��8;hϼ�����a�,rE�,����{5_�Ȱb3Yf�W|����Ϭ,�*�� aV�˄⭒�T�`c�N
iUG"D�u�8��P���ɼ8$G q�{�a_��|<b�ҽ�%�&As;��% �8��H�&:vİ"�/�!��F<
��oqcr�D�.�;�ɔ/f�_��'`��u���T�HA���T�הG�P�N�ಡ6�{H����a�%��ݬF�`~����q�[0�-���5$:a+Vny��� ȱ���Ț}�;�[n����;�B��)5���_�K��2�!����k�˟�x[ZQ����Gc�|�����J,,��F��ģ�(L����j�����{��y���-�������u�nIm��9�Q��lrw�僝������k��#]p۟}/07��lL�dw�k�,Hy�>�`V���c�,Hg�s2��fG�h�h��A+�]�.cV?�4�|�ڵ� m 6s��v)�Aȁ�D�-����R:�_��;!S��4+4W�|`$H S)s����;�ahF�VB��0��! r�_��=>��}JW��S��{3��K���a
jt�ا�ׂ��^51B�-��g���]VX��"��j�Q�%f�m,��*������ǅ�d�TJ��~3k:m�A����Nد<t�=r�>��fy�V��%3�"ٽچ�)�֓�۳���?=b_����[�􈬶)��a�X<�޼��?Q���E1��3��5~�2�EU����dq��տ�c{��{�#t�ޛ��O�z�Q+N��:/z�2j{TyeF��o�=�3�xUv�>�O�$�z� H̉��W٪�+%զ�����v�6l�#G��s����Z˯��a�1>��"�KJZ��yxpy�dF*"�¿�2'�����LxZ�K�߂�|��f�c)�j��^)�60Y��=�K�ғ�_���>�r�q��ls~�O��.���/r7Ԥ8�t=?B��_{ FsSW�e"+�0�ƫ���.�\�k��Q�T:!:�J1۶e��[��Ξ<ii������
�c؀����	��u|��f��o]�c��k������E�	�5uYN���+��c�E��?�3�1f	�z_��]�~�6Sg�1]�P<��?����àVK����ӕ����J�F�a�*3	��W^���[%��؝7۶u�6S��i�ҏsߴ��ec���+�J���ਝ�8,�&�\��C��c�֯��[7YD�a�Z�/}�S��̤�~��}���`�l��бr�؅�Aw�GOTD�Ì�j3�v��J(�n%�.�ۉ�~g}̑!�f<'ӃXRS��]!�{a>J�׌���TFi	y�\�=kz�u\���[�+f��j���U������z���q�Lȩ��ʗg�C��S��ޣ��{~�kb�WS\S:�L�)�����=3�7um��$�v�c�/���PO�KL�M�A~�y'�oΨ���l��4�̌����j�;nޥv�������){�s�}l�u�{n�i�7�`+Ew�֮���!?�+�4,��o�c�ˏ�M��v鎈N857����tޙ庺�Թ�64x^>o�nܺ����%�e@"�x���4���@(��	�f�<$U$S�i=Hj���͉TXN�lK�T��֝��K#�_�ԫYO>���|@�W��P K�_}�y{��g��f��}��?j�O�/�L:CL��c�
�ŔS�#�ݼO�;d��IZN�,��?��1+ь�Z,uY\S\W����.�B�<�:���U�XIR�2���|��B�~U��W�&������4�%߄1˺��a ��1#�B�j�`P��QQ�j;i��6�P���;k%�S��<��wN>�|�V��R��	m�8X���2�	�jͦku+J��Jʻb	�O�RV�(/I�g��*ktO��<�ң���@�<Hs]�r�mJ���p9��!_�����!�Ї�GD��D�[��F��EMFm��땟�i�J��$lr��=�����m�:��S��x�6�[����l&�vb�m 1�c��<[��H�oZ���I����3��^���aQL��W����4�E��Ӿ���+�:!do3���ZU�(&a�]��%/��%�a`;�J�~��VXY����t�$��~��xL#JI��8����S�u�f?��df[��)x�%@`�ja<?ЯrIE���1�>iU���T��=z�B���bҵ�^��O��0B�ӕK�={wڮM2���uU�6�Glǚ�mY��M��m��s���x'�%��Bz�VfTD��^�ߣt��歫m�@¶�m���m_��]Y۵���i�ݶ{�� �vq�-�!`�� ��\I��\�й�i煠�s�9S���b�����	L�`H$	i��LJ��R�����ׇ��}���	l�N���.�e$\K%��E���[��[Äxv����w hl�,za�����'�w��E�N����E��'�6�Z�_ω��E���e{�#6<6a�l�6I�o\�¢b���<mqj\�&f��)K��醽���6V*[&�s6l�޽���,)Dx󐯱{���������Q_c�k�;~����ݢɌ�;w����T�� &i
�Mgx��B��\{�N䄢��N,b��q2���;h�:��OV����+B�Ͳ̥����<l[2�k���)۲*o�{s���`7n�j�ɼM��	�0c�)�e�g�(3F�t�������~�6�L[o�*�M���=ʯG��m�@����(!��Ο=+b*I�!��	�FQ9�P�'<�^Qƾ����T1�=��s�\�ͅ8���@
z<�߈eRq�	@���M�Y�}ᚎ��;���-��ןr�|���';D��7m���{��]�;�4��r���m����d�_��<`f@e��6Qm�v~�̓v��iw�{��U�/*SS��)�,�wyfu>��v�`q>�����	h1���7�����V��fM�l�]y���e������L�x����u�^y��̩`��Uϟ���Q{�����[�X��c�x��'S�:w���{���MeI�c�Oر�'�!d�=���*Ӂج5��Zt.��M�7.��]_-̥��dt��T�i���xC�=|�NK��X��a�i�X_�dٶ��V��"��k|g����S���'Ǔ �T�l�a�ƴݶu��޽��c'�|�u�'-��|k�2z�Oq*�N�ʬ|�ͷlB�LLma�^�*����:���1]{�;�˙��0�3��܄��!�G�-�F��� -�d""奲���q��G�6x�^&�6::n.��م�/���3��h���S���vah��s��'�b$��rq��uYV�6����]"	�g�~�8-"7(�u����ځc��'��m㥊oF�g�b�j����d��ğӽ�.�f �|!����}K�a�&�U��Wߴ�rݺV��iI:5�;���xa����{慗}�;c*1�pJ>ȁw�ڙ�I����b�B�����v�C#������d��<q�L�<��;�=���W{�;�Ü���o��悮тj8��y��(�C(sXL�i�[��b�DC�F]��<?v�bpB��0�1X�����,������-DET3e��3#�-�4bZ	��rZ3&�ƶ�l�Yl
ޮ�w���X�ʁI��8�K�~X�ފ� ��%$=��h2uU?I�� h9!�)Hځ�G�(}jh�;�FE_�F&�,���g%�g,߽ҪM��u� ���8f�~�)YuK�e��,�풖��Z�%$�<*A������شE�}�U/�dPQ�Ѭ�C*��¢��r�� �)����Dtb0$���/�cO>o'.N�L��ڙ>��5vN�����/�����0bMe�:z�*̥�&s]��L�����%{Ĩ]�6,3�ްt�
}#�	�蝴�[�U��|rf��z�'a��'�}�u����g���i�{�gkf#��it����<��j<VK�DD��V�b\�e=���C	��n�u�	�["%&���o��"��|u��S��Ku�h,-���EP)	��e����i�?�9��܌:qfr����v?VL�%ù����q���A�&*�_迹&�hKך�Ø>~4�N2�>��Vl�橌/jm�q"�J<%Ry�6��9mf�(��Y{��s��������c��6&7��,X#�k��ٟ���v��	����cJ���L	g���%Xr��?���3.W�XM��$/���������wO��db-�=��%m����2�XNQ���̅1;74ic�e����8/��?��Ü7��=b��|>+DN��48��Ä��!&cz�"��u���ˀ:Ӆ�&�2f 1b>p-�꾊�>��~_m慃�DB���@c���(o�-��R��]W�'��c���6y��������[n�-�������3/�풝Ż�<R��ʛ��x�h�l]kwʯ�M2縥E�lxDU��t���v������lH��I��h}�'i�M3c$P#��Y���|0�b����Iq�� ��&�t5e���At	(m@{|C1v'�Q$6��u��@발���dA�W�,������N������(�Ȣڰ�ߧ"2���3���X���~J槄OL������о�eA��j���h<������3R�>u�c��~�*&�j7�t9;U�ٿ��������@U4-KK�U��}[>Y���j�DNRk��#��F���P��_�`�jZHdژ�e��uΦ�y*s��`Z� %Ee>F�}i[�Y%B���t���OA�C$L�Iʡs>�'�������}ރ��k�U��ZIμn�&��"�FI�Z.Y�h"�᥶p&B��H[(4����P��Bf�iF�XLffN~��	�
32@ab}_�@�,F�$ӌqB���nVbr*	y(?X-�OPf���w����0|�J���M�<W��M��\��`�,��@%l���+��ZQ4�*��葖�#&d&=��T�B��s��X�*�+�I�u��"X	��Dsz�������Q)3�	��C?g_�҃��TT>Yo���D2�O��Y}�g�9��3��?X��3���?S�ؿ��o�O�x�Ry�K2}'���7���F׷L�������fAw�4����r��1����+|쉕��4S��9|���`:7��dH>��`J&�r�Q��u#����'����� ��Xi<���T��a3��	I�2LhfL�-.�4+Np̢G맺z�����B���`z��������IY�Z2v�N	͜��j��.�8�iGڴ��e�aBM��`��ލ���Ƞԍ�q�NO�o��]	:��,\���Z��?�R��\�X'Ѓ_�*+�4�ͱ
pkG��9nѸ��i�)�`�BNע����h��<`�h���&�'��$ ��E��?��{���W�:=�hh���s��?�e����Ǘ�t����O���S�V쉲W�ZlZ���;��{�.H�,��W��D"6��<7��
��baC�f�eX����pY�d�g�������0B��2ۂ"��������q"���9��5�) �@���U�G�� �|�N>F���|���:~��~��������q�FE��b�R<��2��B���� ���^�b���
��}?N�]Kw�1u��f��5�vˎ��g�6�nJd�D�������+�&xci`QL|��7�p�w��F͘�ڒ��s�BK�L �0��Ml�$(��u�\��o�sf���?(��w�b�5;-�1�4�Ůp��5��]�}�������k=�\��׎���P�,�Iz����q�cY>#DD�Ֆ�*<��jJŢ�-D2�eQ�^����L�ب�p��U�{>w��������sn���?]�׳+À�*CoZC��O�e�w�{�0��ha^L1s�ݤ����}�xa�c6ɽ���ﻦ���x!�^�#��Z�Zp�հ �|	�t������ʁ�v��&
�������4��fa��:�����Y8G�-͇�ѐPJ�t�f��m6<扖�t�kG�=zar�wV���gP�V���[R��$�v���F$W�������C<�L�рs���%1LM|%3���Y�/� ��6�FK\>�|�y�?�`��5�_��-򵛢Yi��c2`��Z<r��n�����D,F���b:୓�>q��������N&Vf�I�銟��J&'#��L¢�hC�h1���SA����]�wј��ye�v�%�y�{0!Y^����\r�/��K��P����N�f�F�C��S�/d*b��|��~�x 
]����/Gj)��@�f�������a1�R�f"������0(I�c&���3��ݰN���`���g�ee��{����<��WJ�!�2 !Q�h"i)f�����j��n6��˝���u6����K��z��>uqh����J���@Ή��!�X��l�S�6�xG�jK�A^Po��Ɍ�4(�/�:��
� f����z9�/Ѓίk�ӱr�"z>A+��,�:*R��;�C�τ)bk.f^�����Y�b'ߠ�07��>��x�}��3�X����#P���ς��'r���_�%��]��c�B�N�������D���L.�����a��CPN�^�w��}�<�t~�����z��t ���yٳ+B�����s˧�y�uOaۏZCz-�Kb6���`_>�ֆ��W{����O@�u~�� fL�6n�堒��! �pv���R0���e��e�/�J{\	���s���J�0͵���	���a���`�a�#,3�2,�u�e�[�e�ΰ�t˰���n��:�2�-�2\gXf�eX���L��p�a��a�3,3�2,�u�e�[�e�ΰ�t˰���n��:�2�-�2\gXf�eX���L��p�a��a�3,3�2,�u�e�[�e�ΰ�t˰���?^��(�    IEND�B`�PK
     ��ZJ��F�  �  /   images/1348d1eb-e6ae-43d4-937f-d455f2ad4bcd.png�PNG

   IHDR   �  ,   G}�   gAMA  ���a   	pHYs  �  ��o�d  �IDATx��y�\�u'v�~{}�@�$@��Nq�(Q2EQeɒ��Lkl�cg<I�)g��#���JR�+qR��8�*UM<��Y�dm)��HQ��W������������~�a�~�{�f��}�.��;��~�R�
)�����TH!��L� ]!���� ]!���� ]!���� ]!���� ]!���� ]!���� �I�$~�T)I����M��SE�a���_Ķa��aD�i�eu��M'�@��p���|�i�w�D[<��	�˯-�X�i�%�F��]Fᒣ���$��i��f@�l
)@��ҍ���^��i��߸JMՉ&L2*��a�lc���y�4��VJ�%�Z�f˲>�&��t��^�B�^
�m�DI��t����n�hk2�\6+�C"��٩Mf�)2�3<���n}z�Vo(��1��i��v����G���� ��t�Y���*ن���	k��\������t�	����Q�"o����N8a��[���a��	*d�� �X�2�g:�k´-7I�ec-f�r�%:97� 3d&[q�����K��3��w��K��_�Ӷ�W}�����6���Vh��t a���U��7���G��*=����_��:��:��PI31Ń�X�1Ӥԁ;S��>q����m��C;&��f��45L�Z��t I���coe�Hq'�r�J�s�����3ϒW�)�d����ㄭ;��mRb�������t��+��%�!ˎ9�Hk��>2�R�n�Ag�.��-���<�R�f�e��v�S�1݌�-��M�m3�d ���┵o]��k�Mǉ��P!C-�6@Xw��57�<fʚ,�r�B��̧��|���&�%�~,�c�J��&��B��㟤w�|%L5}&�A�~�
�ͥB�Z
�m�0[4��$���f��>�~������$I��5M ��A ]�tإ�A #a<9�Ci	
��&}��_���9*�<Fe7Ň)(�������{>D���N�#�N89S�L*d�� �FH��K�a����\�����`8�̴��[컁m54e�2�R�n��bh�IL���J���:}�������1�Z�>�P�rP���G覛n���>�Q��B��6��� Q��z�.Z��r��Z-��Nn��To�6)@��
̶lJ�8��V����/����t�uVF��o~����E���K�	:BQ�]A/�\
�m�0�0�-�y`YL9m˥0�(R1k���5��eZ��&U**���lQ�;T��
�n� ��c��M'i`l�m߾���>z�G?���%��4��?x2S��<�������z���,l���A7g!C)�6Ft}��2,�PH���@d��~j���K<///S�ە�A3Ơ��^�r� �H�a�l����.��.��633C�jY������2�рS�{��}쾏��}�Q;h��ҢM��K��6��Ei2մ%�v�%����eFIB�kd��I����-[�Uy�����f��z)@�1�\�P���R��]$��t~�������aG`���A�����t�u�I�@Ebt������ 1$�l1i�'��`�As9���mHk��4eLBqH2�A�v)@�A�c�4Π�V+�%�,�$�Δz�J�@@X!�r/�3A�s���~�>��_���]J�^�,֌(/���a�t$LS)ڱ�>eܹs'9�#��Sr/ek��Bh�ЮO��JU�O�<��l)@�bJj{Ҙ��(
izz�~�3���{��{�|ۗf��H��v���r��ҍ7�(�Mo'67�}C.�6Nx&*IR
��^{�5ZYY�N����_]����9����T�f�t$�V�iQ��s\:y|���H�n˖)����X{�L1d2�z%��~��������
�D:H^��6���Q�����b�Z����z�{�V��~����:���C��rH���4�y����~���ͯ}U��� vC*�j�%@���[�]�z��J$>�J�
n)@�A2��V�E���q,��u>9r�������8َM��Zn�H�dQ"ɹ�x��5ɵ�t:��o[�+��h���t�?�8���t��WQ����*v��� �	���m�a�!��R���������M�{�P���w�^ڱcG�#���Q�+d�� �*Ǳ0����z�.MLL�m��'O�c����o�p�=����H]�#�P!C-�6P �0�_*��J�x�:~�8��K�+�Z�3�<C�o���$塞yP�&z)@�A'�aۖx-���f��{�,äDi�fU�k[��j쩧���G��mw�JA/��1֍�I�E����a�]C�D4R�H70��\z�� �0��ҝ��.߷O�/�-�*�?�mP����� �h��P�B�v:4::J�����G���>$���Z\o����w�I7�|��_�֥�s�?+@7�R�n�D��$�j�Vz衇$Tse��i��Xl�W^y�.�b9e�fH*U�E��a�t$�i���b=�0�������M��e��~e���^x�^~�eq�,��%+��6TZ�nȥ �I�0�����,r���}�t��?�4��>)1k/�ﰞ+��@��ޞ={ĞC�L	��֨�B�R
�m�T,S!��dP%QH##5z�i_���?�?s�l��-�g�4��d�RK��K��"4��<�Pt�.�6H:����KV�e����"6z��K%ꅱ��ÿ~��l�h5���}��������/$YӮ�tC.�6HlK��S�ףJ�"�:�iH|v���U{�R+0Si;�9}��<�:88hP[�^��� ��3�
�c
��*z���G�~�b�0�	X��V[�.����ڵK ����-{F�6�R�n��l3H�"�t��1�\����irz�N�<�h���3������=R\���v���+�2�R�n���h���Ģ�����o|Cr/%�2_{\j��.�J�{�<M�t�^�NIb{�[Z����� )c:�G�+�_������z�G�ԁ��9�hb��{V:	1�����a�t$a��u�<���^"��'l�u�m�;��k�̥+4�[�#m�R����, 7�R�n�]S�X�T�K��� *W+��u֦�7�5�L�K�NNN��N��2����K�a�Y=���b������z�rI��n�{����c�=&C^�c�hK�+���^���QҷY�L���#2J�{�y��z��x�f�,]G�_��t�Y,	�m�e��,�� �6H�2�J�R�$�=h��O}�zE��<�?��r ����$!�HE�E~������K���1�+&�����yl��D�_׭y0l۶mTib���=����W�nȥ ��J���ZY*�ii~I�)O�:E�j������y�i�~�������S��+d�� ���^�^�ش-�� �B��5�)���/��SeKcYt��IY@)`q�E�cKp�4�b�!�t%� ��8��-Wl�g�z�bw�����>h:��;�H}�{�뮥�ףVs��X��rȥ �F	�ǳYKE������5�Ϝ���Zә�&���eHe<����Z}�ϖNb&9.�Q��5�R�nD�0����N�<�VV����]�'���2}��Vy�@�\�җ�$	ϟ�Ľ�tA:YW� ݐK��%�q�PE�A�xݱcǨ�h���i�{��(&bvif��)�n�&.�aL]�4���� �vJ�V�iaDT������g %��<B�֨��Dϲ�Ę���t$�aw�2OТ�Ȓ_��{�����Q=c���[�l!�u)�B�~�%��(bz)@��t�$�����G���t��: ��_�g��)Q��|�Y۽�����d�Vɒ`;LE*d�� �	�d坻E+lˡ?J��$wtTW��Iκ�l?�Ph�v�M���SqQ�3�R�nDnD��t;戩�֭[鳟�,=�ԓ���Ȉ�����8"��Ib�,x/�G�� U���E��!�t ��6$NL�d����ڦ�Ozl�%�^���\KY���י����� j{/ҩ���r)@�1��(U�ً���xl�-з��-��*�*�ǔ�^(`�LE�v@k;,:U�裏J=ݮ��}V\�\�o�X@d� ���F�q$>�~
��抰��8�r>I�iD���q�z���U��8�����^��� �M3h$�3��T���������������铤A]�\�����@��ߤ��aBb+LAZ�q��2�R�n��:�+�C[&F��YÅ�.�~E�#�vl�vs�������E��b�X�uzm��w��|����i�]4=="`z	�%�|�+M����t ��Y�j�G�4��j5��ے?���k�����џ�ٟI��R�DK�Җ�F�'�rbm;�T��hg��}~�c��B�Z
�m�L�k�qf��Wl���Ҽn7$�6��nR�V�Nr.ٞC&3�w�d�Jk��r�?q�-����Ŵ��ӥ���k��%*d�� ���ё�+Q���]0/���ó�IK����m���ΠI�_��=g 2Πs�9�A*L(�l�l���4ۙ[�7WM�<C����@�bj�WN�҉��|�%�Vj�d�x�����T��L����Ex�fJo�O����ɱ/��آB�^
�m��UJ��[<��6�5vX�!�C�;U�:�~��<0�N��~g��
��&�t,#��\B�� Iz�A'0�ة��ydy���	W��I�v��5�+<��H
�m�������������6��怆�H�B���0&��%pbZ�Q!�F
�m�0�L�hRT��I,E:9�4֦�?^0�Y-J����Z|I��0�$M�N���4���Pr��_mNSN%)a=��A�m�6���`��9�N,����H/��p��R��l���#YA>)�n")@7� JP9��1y��︀�@9�4ͦ�ߪG�5���*��6��A�!M��B(b]i6i�V��3�NK�8��-Y�A��,�REg��$�A�O�U� r2A1QL<��}2��j�B�m:)@7�����u��3ga}ˍl�c��c-�1�^�ۉ}.7���]�:@}M��I�6�vh͇m~�0���a���$�@��/��o�NW^y%���}�{ߥ^|�~��_��~�z�U�$�H�_���^n*)@7´�'����۳k7��?�Cz���������t�]wR�mɂ"��2�4l�B�_
��$�,���9h�nR�R"3apEL7�@Z�ix�����XI�h�W o�H�!��(M��2����%-9�p���dG	9�0Ƕ(	���t��,Qh&�5�p�I
����`�c�z�������$+��֞pP��2sJ9�e�)�K
���)m�ԙKL�c��u�<�;U�w�d/�W%B����r����ǪNv��LR�ndK��E��t���_+��K�6�y�PB<A��&&�zay�������b[���M%�D������i?c8�B/�9�I^��T�V��5�R-����JE�M(�Hʾ*1���:d�P��
�̫RY�y�8��T��lN)@7D����ԨUQ�*�=��:uYG0,ԓ��J!�R
���61U�x+u[u�bb�,%9_	�=�k����&�H�O	3N�1���A�sD���lL�P) �9� ݐ�JÔLL�￯3-u�ΔKbmR)@7L�t��V}1׽��	� ���2tx@k���	�*���Vnn)@7D"�OLi�AǏ�j&f�cuF�#�Pv�T
��(��9w4t�3iՖ0�"K�s�J�!�H���HW�Yb�4#�Y��T�h��R�n�Q��԰2�Xo�)醳�lN)@7L�Ȱ�aZ�j�0��F�k8:@Ο�Tt�Y
��HY��D�wP�+�X��|Ud�lN)@7$��*�,#�O�t�:3t�A���@��tC$��`i�H�%ԛ���%��I� �	3L3A#>ǥ$�|�lC�;E!�M+�I�T�AY%�_] ����*4ݦ�t(�V�V�%�_����%Uޜ9_��Ț�S�33���zQrń�<��7M����N�M+��!a���Q<��{�{Ub�h�R�Y��&Biʰ�����q��h���hS�����;:�[MTB�ԬZ�����I�ޞ�"~#�I�y�K�9DE۽�*��I'�B^�b:��z�-ʣQ�X�<�m�G[@ed%�Y��t�2���{���S�xK�e��;�J];JL�L)1�QL͕U\�J���+�#J<��꼉� ݀�è~(�~ׯ�~�F������61 +1�̯� $�fE�H���;�vB�$*�;Vb-e��jMX��N��:�B �?#�=rJ��=�=9C���4Z�}:d��"��U�2�)� ]&A�v{��׫�����i��N���:������-���ZHCj}$�F�iJy-�h�ٺsǔ�^Od��6���^-�b֕Aџ�ɟЏ�x�~���1m�~	�{���i�z�
ٔR�.��v�z�^���a\Q��b�3U�W�B���
���P��m��j��zqke��/M��5�S�\��f]O�nŐ��o�٠��%��o'�f���ң?x���v���T��P������ha�4g��M)�XA0����W&�l��6���(�/������O��^~�%E3�d��ئ,E|6ɣgh�=+f��(��$K0(MJĲc�F�p�:Ӓ��[���������]ӻ��X�ƊIc��Je�
ٔR���h�y����{K��&���Q����?��?���)����}�t�N�h�ҫ����/�ʉg�������$N#J+��͠�z�U{�+�Ee�N1���[�����,�/ˎӢB6��܃.�?H�.
��g�&Ky�w����B5�����?�}��ǚ/f0�YJ��C��M���n;[��xU���yn�`"�ޒ]�L1ۡ�P���Js��t�rlz��i��t�0�mo��oWU;$��ӗ��5z�����M���BKYu���;-h�Z�{,s��(����Y� �A-�$�0a�ɚ���Q�R��ՙ���[�+~���_��}vn[Ȧ��{�EqR�l��Z�����9>7ۉ���K^�LQ�K��r)�+2f�E��5��tꖙ�Рܒú�vF-��%-ҳ�͆��é"'J�8柣�nt����,���vɣe�-h�&��{�%i��q,�p@�X��e2����k@X|�|��':rz�DH�Ur�X)�L�L\�`��&��
F��w��
������)����HQa�&�B��jw��v��Ɩz�+WLO�`�V;N��g!?����-��Cs)d���؆#�٦
�V�(\(��/,=��8�﷎�>��B���6#�LSe�*__G���V�y�>�4��1k�7C�+���c���#aəll��a�fB��g#?��c�b�f�pA	��F�� 2-�"�hĶ=w���x�
)䧔�{СEBB���~w���m�?�l��|�
be*۶,��TH!�@~�A��-F��7��z.��
9Ķ�VRK���F�����Bށ�3��VF n�!ŀKRKR��c�b��6E�*C/�-Ӊ��Bށ�܃.[�M�"�	�Pk���"**��i�Q���Q!����S�.IS;H�r���K4Y����O�=y"ڣ�V�;�J�Ymd�l��F���w����W|�1&?�4u�����c�mo)6��t�J$Ԇ�����X�an;�m�eZ֣l݅��e�/�v�uT��4��)v�X%/���[�ݼˬ��2�'�TO��_3V����[�����k�����?~i�/���~Og���D*W�8�lG!��yUo�[d��&.���� ��T΁:�,�M?y۠���u{�f��W��{�m��<>]�ۣ�4J"E��K6p�/���ٶ�Wcg�8{-�T��m�\e�����U�7߲Uy||gɤ���_b{�LٖK$���X��6�VT�,y��<�_�4͹T��][[�}� �9!)�{ӱ$s�g��;�`|f*�`�����a��X"|�C�,���\���/�]]��*	ϟ�k���տ#kY�f k+�պ}��*:��h�)�9����B7p­�4����Vʔ�چ\c�YV�M��W�\��k�=����nU_m�?����*�ֺa԰.���-0��ý?;��R��C_ɔt��TNټ7��q>I��H�Կ�?y�PY+ִ����߈V�	�]��q��F�BDN�I{��T�J�G<<e 2���?�$�]۝����mM���T����Q���]�C���a}'ˁg��Z�n�4���Y�����D��V�cR)J�@r�5�#Zz�V�u�5'�t���y(��[Y����s�1|�����w*�73՟#�%b��.�]6�7S)�7dw�.D�y*�T��[i�����k��&E]�b�ۖ���R�|gK��1ϝ� y[�{����5>�/Gc����F!Y<Gؒ��1��i�Hteh�5�0��\C�9�Q���݋l�7��^$�`��{�X���Ղ��������F�MOl�zU*%�<�������Ð:AH���(�8-��N����@��,Mb�Q.�\�b��k���V��^� ��ղ!,��k�����h�yA���N���?�|B^������!<��F����q�15_���Xi��jG9�^xLS\�2�nJ^h�Jj�;���8Y;�0�ú���E��|�s�3>�;<���j|�.�����r��^ޥ��w]t|v-q�����k�`��[O>���Skp���ȇ�%��n)�	��Y�%N�R�L͞ZrkuJ�2��x X�M䯯_8�uz�M�^�64Ӂ�ٶT]k-������Ȋޡ\��y�l�g�.�<?����[��r��O�TO`��+J�� .И��^"��S��\��O�"��n&�~a�Tz�����:xd�Z���;��T�yTc&2�^!���Ĕ�S��,K_�Vz��/}�e�� Fŵ%ϒ�/����fN}�\f=���H'GfJ�w(�d�M��+43��mJtxf��>�:5�,)�o���_����!��&����V���A���g�btZY�k�6��)���
����vO�o�S*:�3�OG�O�L�ҥs3��L���(;l�쿯��K��`��T[�6�F��G6kE'�Q�����$;4���t�4a����;^-Ӗ�qRݶ�j�[���f�U�u/j����m��r��S��]=��������S/��ʹBt��&u4h����ۿ� @�$Jx�R�@�7�Զ�a��Qg���i�����/(k�����.�
�М����"�jLM�y+���R�t������k<IO��Ls�&%<���y|^(�Q����&�T~���|�؜��i"h�}Ǆ*�C@G�_BKæ}-N�گ�;�u�G��A��X�<�T��|�>d��*6p��T�ȹD�I�d�e�K�T��U��Wu�D�l,���B9���sوK:�؊�J*�O�s7����Ju��Z�Ԏ�(�|C@%��:�6��B���dv�t�GG�i|�DSc�4���aL�F�rY���)�$��&S�n��J�M���g.n@6+����&����fp�oL�*�fK=����p��Г"qBd4w��/S�Gao�ۗ������,XnR��Z̫���'�À�J�����E����Ϙ�f� ����2����y%���6���}�qՅ�4�Ȁ�<�b�#~�[���{�8���ɔ�0>xr��Aq�R0�lx�-e���l��*3�A��h��	�N���"�m��(��@�)a Z�I�E	�4giv�Zd��T!?+�Պ3���~��Gt�@�0�g�L�O,���>�ρ��LhۖQ�'��vN��K�q,�<�,�ko�El�L���W��y���Þ��%E��;(�<I�J,���n�F����+a{���|j�zrmrD��2�N�F��L)��1PIv�Lq�Mn���F�����r6�,QcqQ�̍33�{���Dk�B���=�	�A�"ހ�NQj'u"2���8;�\/: ��3�>]7���Wk<����<���F鹌�\��)�]�]pt\���s���h������-Tڶ��2�*�S̆�œn,c�b���0$����`|8e�/`Mi�	���b���}Oy������.����Dj�gү/v�~|k>�J���3��������5	˨�#����'ðFY.tI�K�%�I "�|�B/$�O���d3��� th�c��إH�E�Ϻ����G��-�Us�#�~.d��$�~l�l�U�l;�h�Rf
�,�����<SƬ�<�9
�4����aV���.k3��a��ͣ��cM��P|�ha�i��c��H�u�t)��Em�e��9����&�]��	��0�Ģ� 0�Z0�I�[ya�%��^ˬs��|���^�m��t뽽k����u��!��SV�5�Ɍ'��-�n� ��@O;0,8�X�ҏ0�@�v�7��`��X�&����7�x1�l6jyLqE)�3v��X����	2�|�o����w�d���@��92�ϑ��;C��7{]�\�R�,�2m�ٔ�i���d�5�W�-�.\�v"����1*�-�|��hi�I[ʖ��q���-e3b�d�]�Y����^�]5yP��9�!�f���Z�qxv5l̖�˩�{��$�X)e�0u��h�c�T�g�kx�����5'B�ut�ل�Bi.�f��3�0�x�~�L��Bg����3����N��ؽP�5�`�=.T��[�����V�1�}Ɉ�x�xH�.3�X'����� ���3qܥ�g���Q��3�pe��j5��a�n��Q��l0b��c<�hJ�����P119�0-�Њ1�@�)E�<�^�n�� �BHK�@��^�Z��^�
��U��`�� J��dY��I(T��m6P]�Ȇ[�����D����{�{o�)���x�5��
�앥e�y�^q�LLm���8F�<�Trc6�y��|�R�`�%�&m,U��+1��ulh�O&8MC4j�����-*.|j����1�T	h$��\�C^Y�|�n�@5�%_�3,b��%yn`
ne6ؠ5�]�#⬃zu�$J������w�Y��D�y�z��َ3��7Z�[��,QhL�6��'4�)8~�Af1�D�'�b�0%L��Z٢��G;vL�©ST6\Z�_b;l�F'�P�M�������/��`+�<�omB��o�^�)�SGԷhh.kה��mf�w�d���&��E��rA��ܹ���l�t�6��<b̠YXSuT_��f�V�Q�Lc��l��|��D�_�[o��n��Jj,�ҩ�����h|�z�ߥk���B�`������C������Yr�G�s���^�5KhH�7S����6_����-lAT�1e�45�v{b{���}f�7�5_ͥfץj����<�t��sH�Zp2��Λl��?����`�P� ��`��<���Q�����{�6�ϒ�|����7��T�QI�F����(Ww��g�q̵�@G3҇؁�l[29�9a��}1�2��<!��������cM)qݰE�_-}�Λ�������������C�����y�)��_����$N��zQ�phk���!���]��i��OX�Uhzګ��C�m�↤�Z͚{�!��ra�[7���o�J	�e�@3d��?`ש�� �����kČ�i7ٖ�A�f�\~9;�
_�tͥ�i��Q�>r]�o��5X�|�[��~�ў�;�գ�������D����������ƅWY&@��.h��žx���{��c��J�=��>��^ܢ[�?�����&�n�sH���U�����*�z�l�(�ńv���ۼw}�.�PL���Y� U���:G��=�}�t�.Ϙ�n�6�����)z�\�h��"��a`�L�}f;	Ov)��]�	}>0�X{��^��إ�w�K?9��iХ;/���^��;�Х۷S�٠�F���B����t٥;�O>FnݣQ��p�Y���+ �[ ��	�OtB�N2U�G��f�Һ���,�B���E��t����ee�G�}�Nqi�K|�p�X�� 6��Y!��4�9�h�[h��$^����*Yt����GѳН� �>3Of�I��v��N�Ex��H�V�}6�ȣm۳�v]}9���<��z��'<�ڿ?��
�0�GF&���	���\�Ŏ�4��５�}���|�j�q��6-/u�R�����χ h�'�j�NG��Ç�О����k��z�*��9��<������׃i�Yc�a�������V�:y� �1�6פk���1��d9.�,ӣ��P��M�=�vѻ���'3��N3�I�M�a�%�*Y�6���:����Z��ڷ���Mz���t�n�׎͊V����})�������l�o�.�oJ��uh]���Ȳ�,���he�n��@�uG��r�)J�u���02z�)�!��GJ>�<���b{�\؈O�.|�hsW�������|����x�ң�N�r���֝�dM�k�n:v��z�Mm�	�g�T\�����v��ڽ4�PԣS՗^z��<���1R��_r����01XKU�5l��W���
5ﺑ�7O��Ӓ��X���b�x-���<6��.��=w���4=����<I�������sҿs���l��,�軙��V�Kʳ���@e��n5��;��_X:��d��NӁ���������Iw�����(��LϠ��H����J�rN�N[�z�<����]��H�S�tใ���^z� �^�x�8���ᕣt��b�%̪P�e�W�Ь�5i�M�Fڶ���~�H�O�Vd$���`l�5����y/X�J�58΢���V)�$�OQ��d��e���p�G8C�]IRt .�t��r���ߢ�g�k?�i�O^;��}JlA� �(dޝ�Ă0��e����饣'i�x�����ۧr6�e|A-ǖ�@��|�?&���_���1E��і�:ӡ��?�xH۷M�/|�=&>�|��v��>u:�Ʒ�E��v�v^��?��;₩�;or��\�rc�	E�X:�jʣ�1�i9�g9[R���f�H���0��i@g�dgO�ʏ	�|�}ˣ�J��{I<����nH�ئ�3stp�Is+<��%�Dbt��I�4{z���C�f�ߨ�����*�GSB4��[�xJ�?&���;X&YPK8�*%/��Y���������ki'��G��b	e!�S�|�wo/tCE��6�u�4(��tK�K,y����3S��G�� �+���"�Iy�c��b�M����F�V���7\�D���:�a�ƹ��E:��:���Y5n,R�c��O�]�Ց@=��c'$M����K�c|.�N� K��|�m�E:u�ua;im�ϭ��O�ϿQ�9��rE��G��F?y�y�g�����;���;���Y��X� ߷�5��R�갇^E��S<�\}ݏ�I*��AE��'�}�^_O3̵ [=s����9�H�BBy;�eN��<��/:H�ZԵyL�e�����b��RI��K)a'�'�k�X�>V��m�_6�A��!����v�V��C�*Ip�a(�@ ^2�ro��*m����c����~W�D%�+��6�nV�._�;������~���#���IS�� O����Y��2W�y����Q����|>�%���|��@���~"=U: 4��$���+� �T+[�T��e�8�+gt��Elk&a��g��J�:�.5x�F��Jĳi�)��Ⲯ.ς�r��|��)�����7��竮�j�a��J;"t�i�k(_���ILK�c1�Aa"����i�Ӊ6��aI�Sv�k'{�
������L��"F��u�N���N�ͳf*K9�w:�Ul�<���K���aZ@�!q6�pm9[���(;y�p�8~�m<x�y��l$^u=I��_R=Ycl�0�+#2v�S L��`c���Eoir�;�P�T>Xt��Ń'���,�ǯ~�*p��G���e�G�fԁ5M���ҋo����Y$B+��Y�*+ߌʘY	#(��y�R)���x,m�M�k����� ��?4�c!��GJX����d�:\�a4��8CKg�Q�]��=��#l'4�g�e֖;w_I�-�?���(k�3����1h0A���������<���!������Ck���T��d�!�}�[���k��YUG��Ck ����d��Z�%�T;��"~��Rf����ۚ�e<�`�B�g�lK��Ħ-[���|CkÓm�@�	���C$RYv�v���dehw0�8��1x?�[��i88_������Ζ�"#����ͩ���G�B3�@̒2�[��-2�p-6�{Iڷ�E���%�YH�:��Q��#d��H��KA(��Tv�W$��TǨ�.�d�$h��*���ͳ^Nqr��0-3$��Z+*5��ߙ���/�I[��G��^9#v l�
Sy��;2Pz�Y�>�K�g����'O�)�A&�?V]	1�a�N�|���8G&v�~ڒʊ�㖵g�А�۱�<�{u�fUpr!��p˹:��)5Hur7�B^h���եj�*ǂ*7 zL88g�x*\K��/����A�L�WV�#���6�i�k�]�Ax#��Q��Deny�]�m�n4�djR�'.���8x9'��~��7�=3O/����\��H�@r*aMF����g��a {%�2�qںY��x��0�'_:�S�T�x�0����M�A�4�Z�)��$��ۋm���=��I�Me�E.t��P�KHz9_���8Cp�"h6�ʚ-�6b3�[� VْP<�<��%�[)���*�ng@b��İt���|��^�K�,�j#���*�E�Y��V}�2Q�*o�ZzD��XT`�\�j�g{��3�A�O�a����K=K'X�|�G���M~m�
���q�㬏�b���ۅr\�2A�AY�@V��ס�@� R}�v�g���5�$��fjjRr6�M�+O�<A�VK4/4�����Єx�u�Vm-�j�hyyY��m��Y\�4X�6\Ncs���*#/�A��Ĕ[oe�4wƫ�t��2�`�nnq�Ǒ-Y*By��� �	-��B�h��B֊ru���k���G%�/N���Y�>V	p�b7�A�;j����	HG��"i��	�cg��N�"��K[��!�jP�IH�Y����ƚ���f۵$߆��Đ,:��ơ�d��5=Q�ڕ"ɕmÔ�)վF$�RR�Az����T(���t�J�4��zx�y��ϊR���e���֋�5f��������i��z"A}؉�T �1�c�tg ����p�&�졒�i�4���bib��<�x��y��$�֜%�.���x��Zy����Д��r��̏��F0[躽Α��qve{lsf�������$MOMP�V���%�n[ )�8蹤5A�uM�"m��^'�&/�i\(�G�J��\�L]w���8U�Ð�3ߋ�v��[�n���R���I����<I�L_;H[ln�̤��U�b�d�m�Ц8�R���y:����Б������@'QqK�[gu[�]��EhX��񀏙r�˾�Õ��1�W�ݎ�n�}:�@������!�4s�Dߚ�6��$�Ւ����ҩ�������� ��Hm�m��\PXh`�AhڐRr-q�`6���<A�"`-`�͍�w\�H|���[����A'���^�ˇe=K���5U��$�T����ѯ!8~��G����"k��|�'�vr�s�Z����`�fS�c�Y|?�W�}�1�����k{��n�� �z����i:����<xF�Q��2Q��v��Y#��Ĺ��9t�W��-L�Jg��_�A9f��W���X�r���Z��	;�|0_xr`GJ���\�r�D� 5���r��R;5b�THt+�M��� � <��<�۳�.ݵ���|�d"`��~�$�|�9q�5@E��Zh��f�ZRu.K���L��-M����KU�S9��K"�l�(��ulU�m����_0�?�2�`[����z��;;�Mӑ����2�J4�u!�>��1��Þm7���⁤�A�zJf ���K��gUK�W���>y�D�LA1�Q&��3g0+����|G���1P$p�tʹ�$���e$��jm۶���&��,�,�d���@%�Y��:��r����S����da�FK�옷��<jF�<`:�j L)X����.^Muá
�o�I0">�Hi3���K���sar��b�nE<�%7l���.��&�U�:����+���c'��zT�P���BP��0���7�^&�E�u��d�J�]�j�=�j�v���E7^}9��)����5t���=�4���I�,�aP$�GYf��x�M�&l+[2�;�&՘��ր�=R�B��NL_%o���@�ϼ�Z.SZ��~Ig���)5���h/���E�1SA޷����`E�L,�� R&CR�Rє�2:�D��%����u�� l/PA�?77�%��g�zO��ceZM�a���O{�u��A����|�o���s�@[�Y5۠�U��0L�
�2�H�Ce�S�Sl�So��M��,L%	nǝ�hA�κv���?(<�!��-�q}O��+MtyJgۗ��_�ؽt�5��2[%�;��+��=7҃����qj��xr_a`iV%����$v�2��ź���l!R��N����1u�ɇ�Y^����_��zݥl<��ى/X�U��S�[���z�}��vÏ_8��tE�(|�_���O�^75�ǐ3���n#�:E\,s��*5IG����昞� �ޚ����V��2K{�/�0M=[#��C,ې� E���8�)>�|��D�t�I &?�qz�<C �_�;_s�3���P˅�+WV����ct:S���ҒN�q|������A���&� >8e0�u�D]Xs�|�w���*��>\N�mFB��A�{�D	9F0��2,}����	֜w�=W����� e�Mi��OD���Y��/�E���J���vx��S�ƭ��GGh��R��D���|�=�����w���>�N4�6~֠S�tPe����w�g%�5�D7��K���I�Hv�t�O$�A�[��B	���G>�::3C��*��^�)�-��v���k�ŗQ7%鰽2O�w�r��U:r�5:~��ؕ|�Q��k3+ٱK4=��y|[|Y$��2C:�V�{y��S34xBI�k߹�h]�,��+h\�w�H��#�K���?�`�BCa"��v�3L+! >l0�$1�! �<��i9ޗ�Y�NL�~�)�gK�Q��<y�v��)���Ϟ��,�M��qԪu��1�<A�"�H��2Q�`
�E�Ӏ��S�8�n�J��
��=I��.�#G�е7_G�/��{�G2�_w���z���+�\j,�������i�a��Rc�e20}4�j�Ю��������׎�J���D+a����q��B+�#4#,2�d���Ve�v5�r����ao�����d3_�ƩD����F�L����Qry�SL�n������/�H~o�>���oF����{��P[�{v^B�y�A:y�C ve�;K�����7�E6�M�����_��,6��:�B��,��fgY<gW7ʃ�.���8ՓM�g�k�<�[��V����A��@��yn��xU�Y��+|�30��zM��@E��� ����	�0�/%^�Y5�hWx4��R�o�������D�kUd�_y�Utݍ7�iQ��2EǺ=��	�k�����ۮ�s���q���>L�>�Mn�����n��z��K��]�pM0~���4k��gf,����/�:����*1��O�%�N>�{�GW};�ґ���]���`D��J���oא�]g�c�_�n/�F���ma�����/Jf
�m1��*է.�_�1ߥ�ъ�v@
�ݻ�_F���Ͳ&�39N+'_�˯��n���C4Mz�;ү����mj��86��)IR���n!+��?T���{xBX��
UZMFV✁?[(�_�ɩm��m�-�I��P�u	�n/�V�Gn�N#�[hdr�8M�;qM�i��|z����Z�Dmh���r;L�rp����X;K�` �bl�S�^v���t�7�aAas�f��5��6M�g����s�
��PJ�*���Sb��J��U�$d��uf7]���<�D5Ϧ�{vҫ��DA�I۷]G#�*=��R?Y��������L[l���&�{��3$[9T�u�N�g�]�l��3��\gMZ�8G
Yɇdh��.Z�+c���+L�V�6�6�0� F+&�T`��j�z��Qk0�
A�^���]���}Օt�g�W^|�.��J:yzN�%�&��8Z\iH�� H�ȱ7�'i�%�t�tEe3.�]���혈�����)F��'b��D=	�#I�$�Lձ-46�Ե:!���Gh����&�r����-9����y@[�tP�S����J�:�S\_�۰=��"���  ��k@Y����b�.lG�>�ڹZޣ�u���xⰑR���'Lv���h�B�S�������ULg|�^y�E*1�.߻���7C�?�(����t��q����43{�>|�}ҥ��g���؂�鄤+��	K[�+%	��̮ʕ��$:E��!�Az�k�L7פ�%�H1W��LILFk$#���؉�t�U�R�Z�g �TM�Ypx���H�x/�yM]��*vُ�|�>ǔ2i7��@�8?���Z�62��t�~�W~�N�/�+��Z��|q��'��L]�p��)���F2{/Ϛ�d��Z=}�����E��V��}-/������Cg0��_��	�pl��Uf�j
�$���:�t5�}��uoK0X0�1ـ���b�|x@�S���`B^#@@�6˿�s�)"br۷o�����2X��� <���F%Y��Ύ���������}mz��Z
�ʗƵ�FF�����
Ę��z�ueSd׾K�뮥K�n�N�M�N���ôm�n:����1���Bq�؎(*v：#��Q#UO���nCrZ)6;L�+.�<����z�8gā��?��o`Ȁ���]�q4 ��f�j���׎��h�S��9�A����J�n��B �d08O���O�Q7��5腣3����hz�N�:� ��y��1������nݦ���U�ѩ��I嗅t)�z�e
�����uIZ2���,�|e�-L��J�;�CK���2�#�i1.�����=��hGe�^E��K���e�p%���Ά�
��DI΀�{"]�ď�}<��� x��P�ZEc� ��a��3�j����屦��Nm�Ӹ�ؔ `����66�~����y�V`g�&AI�˄�>���n�����|����bz��Gi���{������c�kϥ�̃��t�͒�2�����O>MG��^#3i�����Q���w�y�G'�W�1;:��:���[��d��?@%���%X?�\`F��Rtɍv��]�!�e�����K��Gj��J�	��Lx0,6��cU^���~����ߣ3�M��<���x{A�;A�!���Vap�Ȋ_lJ�\J����6/�gT�)f�$��}�N6�G4�B�5V���Mztݵ7�V5M�f���'���p�J�i���!P.-�L�~�v�ɗ�K�GF���|C���}�I��7� b�0\[�3(o�&2wt�Y0zЦ����'t(T3��0P��D0`����h%�/0 ���~���jw��,R}+���I ��q��ţ�l�t�nZ:�L�N�BέT�z�@M�b������Q�ɹE��ˬ]i���S�PutLF#=�mlhR$`�/�����>���F�wL�b�u��dט�w�a����!�*��%9_/UL�=��{/iC)����۲�,�3f�%i[g�}jD-z��?a�DtǍ�Ӗ�)���E��S���o=�|��p�R��:��Mi�f����C����-u�&%�[/�FD����:]{�^3���O
�n���n3��8�#�<B��_��y��I���@j�L�����|K��$���������;�Kc�u)�A+��)_����t��.�Y�xl3���s-�;TtH$/tM��K|�)�.Q߻�v���U��w��]���h���)o�?��uP=�\Zda.O��/�K���>�*u z�DJ{UQ�Ó���@Nm�$��k[�ȹ�hM8�v9�]h��XC
�% ���?��[���;&���C��4���ez���ӓ/f�ƶ.��V'\ct[����k�\.tF�Pl{�t����o#Y�Gd��"�����C�i��2��<�ใ�h�g6��H2�"��E������8wD(c��m*nb��/Wuv���K�i���#�73ף��|?�޲z�ڳ�2ih#)u�^Y��T�![f��A�8�3�'������Ę�ĵ� ��~�g���	�\��.�<�?����(�\x:�hb@�W�{��`��>���<�y!Z.��CF�|�>���f(qkl����L�W��,���/&����B`9�R��~w�fz�v��GV�1t�	�ْ?ɓ�?A_����3/���vҮ[)`0�]�^���OdN]��a�������t4}ߤ�`�R]�-0��ӳF!x[=�NI#����g__�72ѝ�R�DN�N��IA"��ԥ=(�ɼLR��}6d!����@��ЬP�C)����z�⳯��~�**�*fYhs:��/�s��S��e����|�����N�C$�k߲*�|M�n�-1���lj5W4}C����.½�e�I�|Nq﷧�����&0 8�K�IG�΁�g����fݺ����jۅOe~M������?vT�ˢ1f,c����o�`��D+�B��N�ѭ��F$nx�����I��QV�Hb�%ݱ:H�gJE�<�ʺ(V%��3�s(�$�~¿{��L�	߳kK�!�d���,5��T���!N;4POw�2Qry[��𔭓��N��v�g�*��G+��.��r�4�P�f#��B	.K�g����]�A�+ P�SW:�������.6E��A��!���b�Hĝc��cd6 t�G�F(��`���lWl����V�U�݂8H��P�z�&	}��������c��0�-M��r��8��$�HeM�6�R��i�<Ԑk��;���{�~�1� u�g��ΊY���8��9v�8��,�����hB#�1r�'}j�!��`[?�X�Q���!C�Ʉ�;�I�i*Xۨ��=֔6���B�5ͪ������0�q*��f�AH<7[���(Љr XF�7��(z��%�N�V��"���������wm?�?����B���#8D�mt���{�?!.@*��z�$�ڰ� ��vV%mD��9|re��d�LM]���uE�ܵ�>���J+�(ʝٌ��m7��0��L۩�ŝ4�����k|"+��$
H�r}q�XD�f^�����x��\w a��Yr2p&q������yh`���N��Jv�]��.�@ɓ�򁲙��\�4`8<�T*�!/ʦ�&�BS]	�_B�9���b�e����ŵG6��V'�����E���2�I��y��+�|�0S)Ñ�]ԑ�i�Gh���}�ƴU�Hi�A�v���QQf2=:I�g��(3�Vi�D�[�I!a7�#Za�3u���e���2�ݿ�j 8��&�\�*���b�y[�̪�#��hK�֛o���d^�o��$Q}M��Wco�t��$��du�����_\��Q�ё.�yӥ��z:��e���j����ox.�-Җ ��hWIDϊ/��K?u+��r ��` �$߯"gׁV���o+�<��/8BXV8��R��l)4e��v�!6v�ԎI�v<��o���]e�����I�i�����p��8����C��Q��$x��(�����Pe�#���5�!�#�t`F���K���{q���._�S:&i-O~y���yVD�
_�哄�Z{�G��}W�.PL}�N�-Q�S}|�V���!�l��9��?�٬�"�� U�X�ڞ-}V^�����.�.Ӌ2.<���=�����1u��c��yJL5���Ƒҵ��~��5W��}i%��ϒ�mp�6�m�V%�6փm}�z�)~�m�I{�'���I���t�n ��tƅ��kS(�^TE����$ؓy8�,! ���Ӛ��e���kf�Ia�k�(M�$xSj����2�Մ�Em�+ѥ9�I�72EK�%���T�w�PV�.��O&��"8Kk)F��L=��%�$�gH�H�Y z�$�-�XK�Dln�a�M�l�]w镴u˄8��ϝ����M.ۓ*q�@�7���}��n��k�V��2P-���Nr�^�`�SB�O~��t�uW�����1�G���ˇ����q��+uI@��=�R#sq�<{g�ϲ��h�*+I�L�謒Rv�P������ݤCS[���������:u���^L}ʚ��Fy�hO��j�<�:?H��g���-@k�u�{[�x H�8 &��4�-����3ŅZfݸ�$[f6���ry�_�-��|���4?'I
���kh�\����lf���5{|���6M�ԅ~G�O�ȥo
K�	���-�����85����֪�Z\����2�ZG�>����p{������뼮��/���9$� �(��$J�e�R+̸��^3�C��G�?�Z��=�m�$�DKI�b� AD"犨�r~w�>�=��*�dQ�.WU/�����}�	Hh��EQ�]|����?�sl�PT�Q�n.Vqiv�|����'�g'$c:�p^�*o����֣k�����7OC�M3���M������7�B���^����1�}0��^������9WQ.f��պR�kS��c�Q@K�Ly�!(�����B�+�q0gH�;��e#����{�|��� �*���0;=�_����g�igs�b�A,�`�uF��Cl�k�2������k�d	�4��D�aI�3[o�AWA4��̴�8T�B^O(?�B833��v�d}Va��������=������r�� �
_Cb\�G���ڰ����}[i��q\k���G�p}v		�!��NE���Vk�n�qE���H�eS4��k�dI粨�]���kj��s��o��X?,��.�j�_#{Q��HqD'<�9{��x�!�SO��no�eA��=s/Wh����s���{�#(��>r�[�$7�m&�-~��F\��8���{A��6Z�eD���"(ʥ��[rټx��V�X���ou��<V��Sz���1ij~6;�lѣ��,�7/��K������mf����˒#����m뼜d������2 <���q�F]���i��T�=���Z�c#�����DC�����7��J���;V
�ʃg��h�h,�Q!���E�3�w=,V�"@mp�QV����b�ϩ"��תb8�G/����X��kG�rv��"���V:h4C,o����E|��O���Q,ެ)���,`��D�:�j�ߴ�{�+�~�'X�_�Ǧ�[C�Q�\�]?V��|�#J(�0}�!q��|�~l�:?��h����z��b��!�8J����}x'�th 9�wmߊGy#������8��#/lTާ;�5�p��)lھo��6���c���G�d�d^�3*=����x��.3�0K���P������k�r��U�h��i�X��j(��\��A���p��5�U����3��.Z,kb5+�Y�^',j[�<J\�p��Z��:Ǚ��APu4�k�����u�|7��������o~\�'o\�GW��v�"Og
����<'��)1lQ��EU�����$~�ʿ���"�q�����:����J�������5���z�ѧ�w�LߜB&��:��������˪T�8�o�۳GKK:K��+�?�2p�:�IxR����G�ĨIĶ��X��woW��L���8|���$��:>�&�P��1.�И������X�fc��|�M�b�T�#m��(j��h_�x;w>�b6%B�Ş�[�v�VT����d�;������Y��0""�AMύG�֋�%���`���9�.{�L�Y����76ܔ�v��t �ՙ�QP�uŰ�v�=�C�Һ�m�73-���2
&(�|��a�G���;���v�Qm�%%½Ck'��)�?�
���(��2M�Q�l���~	fE���{vno��2�~�i��/�[�lƿ��ݸtA,S�����p��yǰMܫX�u�c���+!p�Y[�f\�Yzں5"�H~ֽ;w�ر�|�l)G������Z��FUOa������y�r���甗��7>_!�d�T]q#(�l�eb�Y"NZ�"$Q^��8p���l����9��Ŝ�M�J2Yrb\�p���,f���_+�_]'� ����$ω+â. �I�T�Q.0��v�{,��¤	������aT��t_D}�VL�ǂ��6>�Q����1p�,	:�}Az_�T]W`�ׄ�^"]z���H��a�n�ɚ�C��JKjm?<�w�
�t�4�rs����l�+�K)��1�xlE��IB�5�7�+���o���3�q����ʳ��=����SW��T��Y�"+�2�'1$.)�Fő!,�����

^.�B��9��zG�i�ZS'L���@Ga���Ǧ�������$(U�ܰ��iٷ�JCi��Ar_v���&�]�i^�Ù�ɏ��\������ �3��h���/��"�u2�T�߰o�����oazfIݎ�n��r��26��hL5��U���!4CC��`��,�f�[��Sy���N�&�_���f�n�&t��u{!��Gc�B���R�]֑��S���(���Ԕ�CDJpz�Z�y�Ifus��6�kذo�v��Z�8��F��I;����~���(�H�ؼy3������L��%��I���۽G���ܾ5��]��?�c
/\�/�(�%�6���2�<�T໲=μ�=;:��L�Ǒn^�ё(�>�h����g�����czC;��+�,7����]؋;�������7���U�z��;q��o�i�\��g�冱m���7/��'W���*5�>f�֬_��"`��NU�կ�����ܕ�t�6e�6�Y�'܇a���'�h~��Z�8i���ԗ��Q4������'+@�����e+QDS��
��n�0+��\E�]@����؛���޶�۷k�KEԠ �.$O�����˗��%b���.,��[����%q��E�_����Zr�d���k1��?��q�1T����}�0�%��7�ǭrCk��l�����%�l�*U��q����/`~����ỄS��h�覜gI�0�+�U�h7����c���0!��Ѫ� ֭�7іk���y"����9��pE�J�+!H��=$��[nޏ�����}!�R>�t��V[�8q�q=q��Ñ��D;/ꠎ5�D��#s�؆�87]���>�՛�H��kV��g�]��+��X�M��P�/~�k-���]����Dp€ʯ��Rɼc��oI ��'+b��!FbM�]���!�A*u�me7@<�;�\]�7�}�=gBg�X�a�Lʄ��k�֨�Z��1]M�MW�3��JZAg�z�b0�E��.>��(�z�vL���ҍ�BV��F�+s-�M���c��}�zC�le4fOJ(Бj�Tb�l[[���.�Ө���h���a��(kb-I���rsJ��
v���g��������� [Ƞ�4��*�"[>^|�\�rS�(N�[�WG����$Rb˘?������G���5Y����w�pO�/�n]�~ŴJ�sW�ߟ	�~t#��X"g<7
�Ң�K͎�U��m4��.1s=Nt���788����o<Ȗ]<{g'�K�P���q`�V���Q+���~l9gvt���
/^�ս�2��: r���!C�H�VpEl����X5�~����13Gύ�Y�N�7&�Q������D��v^&p6�'"ʄ	���q
�gT)�����&V]I�����	\�rE�"���Cwd2wch�V=t�$��F'���ÖD��3G����ISb�k�}Oa�L�qY8�&ϖ�^?���Hrx��G�n�xI_��x^�*��ko���>�J+�u�VgIc\�G2��ϲ�����|:��h��;�����i,��oq��Y�ٱM�K^C/^����?���:�te�������J$�E��WR!$�k�np�=��Q����^q���9�J]�H�%D���tV6�hz�p�EQ������Y�A����V�p=o�$�{�H�4n>sUy%� uo�tW�^^���,!�(-���xS��`��]Br"{���̐�\C��)�jk'V#x �k�{ʶ/�
�C��XL׿Wzt�`# ���x��ڂNW�U��^�<�/����&xJ����\O6)*��_��7x�����Ѽ��_ZĻGO��d�������BF /�R���{��)n��O�yD3E���Xi�Xq�2C�Qi��ob�ڋ���6�dA>Qܲp���~ �u \�A���ӎ�Oa}O��xG�-�%��<�$�[r9�'��7���<O-�B�d��SD�x��T_D%��!��Y�e�e<�V�x��g�� ���9��E[u���ԤNw9��,�	�<h�(,ti���(+'�lW�wQ��ҁ�%���U�a<��CM��}g�,�Jj/?�����&���}�P"�Z�:j�4��N�y�[�Aa�Ʉ�z��5#�kROg�{���.�[��q��<R>ף��Sjɿ�q�3E��)Rr��f���s�?��J�X�����}�1"	�^r��G\���bCL�Ccm6Wq�3M���ZGPD#��'�Hr�'5he,���m�Lߊ�Ӎ�G`Q�@xnE��h�B�u6�=.�ѭ%P�ˋ#�����	��l#2��������a����G���=���)'�(���>������� �"g]�j�z&������f�e2+�����	,>t%/lP�����;(|��(����^���}�j�:�H���㶵��Y��Q�+��Ik���ֺ}GR���A�]Rε���ĸj��n|�u�Ow\�o3���dFY�	�Φ���:1���t3��IZuc:C��ktmO�la�XN'�қ�3��sͶi�YhSY�\�駣��}���M�� M@`k���`4�c���nxl�h��21��s��:n�!�wF�9S�.C".��A2����Hw��ٱ��Bw���T��\#���۽����*w�s�<���y�ڂ�Ʌ��mĕ��AI$��m��a7)c&���2��I�"��q������N����c��nrl5Í�X��L�j��3�D�|1ה�j�]�R��xfUym</����0ƽ;~�j6��{87���]׷)����,�˷$ncg a}���P�Si�ؽ@�N��'��x>���]��n�LRyv�M��mB�R����g'-��}�v.nך��a�e6F�$^�u��2�cUB�Pkl�r;u`� ��3ͨ [N�ds�$�-�*:W��2;�{�(L�s!R�F��x*h�����]~\�ݔ�n�=���r0\�IM��ulٸ	���#'N���-�q��iW+�ݸ�X�kh]���5��4d �y)��ϥ���8�I>n�@��zŝ��x�j`&�]�Z>�4*|�L�K��-ڜ�c@4��c.�@GF�w��j�8
���T�rRj:�¶͛�a��cY4�CXJ��L��Fh�]"��r�S6Wp�7�=wN�d\C�L'>�(�S�H^��`��괈	�"˒F�����heSrOޓ�$4���T��N�:�?]P��D
��ym8n���h,Z�biZ�*RI�L�׊���#�Әi�5`�+nY��\4g��`>�N���x��u�0wj$ܴ�:N�%����O��cӎx���H��9"7}v�&��f0==��B�\���9�H1G��HL�qW4&TL���L
�+�׃�'����e�9�b���1�hʊ̱[��r��Mߡ��-ߛ/�&,W�w�s	�eVv���p3��1ϔB�u4)��c�RG��ou�e[ 
p���q�Ωy*l���ǚ�V�ܵ_��7E�������>^x�j5��!!PW�y*�X��D��;���J:>�od�b�����Ѫk���t�~���}b	�U/�X ���a?�l���(���GFQ���L�ͫ�>g��ө�~��g]~`t�"��s��D�gd!<����{vm�S�?���6ia�/Bsuj�9�c'>���l�!�j_5W[�MbDY$�
8�J51S��7�-�Y����#G�=#BE�H�P17������سnL��tJ��h5+.����mdI� �D���gf�h�_����;c� -���,
D���%ea�,�	��ǝ��
�ghG�˺,u���e�hQ����b��q�E�P�FV��O-L��dS�����*��r��B������e��(w�J��N)�q_�	1d7BmQ?'�iM�ID���Ǝ����;�o��IlN:���:�\��7����Ye��D��դ�Nf�xﰗ�E�WPJ ��&*�2
Ve,��C��S����[1�p]]�X�6m��mؿq~�o/kU*?*7��4:��@������#J�1$9Od�u��h�<�u���\$�����J���8u�x���l�<J��A3g4&���Gc�ґ[��n�X*KFpcr���L �):xC,:c����0~����ڎh����ve�
C�غ"�^4�2�������+b%��fJ�N`�/|(����tٔ��YiQ�%qO���ss�ʵH��B>C᪡ߨbH6W�4���YbHg<�e}��Z�c'��ܖ1Q��Z3+�t�$�f!�ElZ;��������(�$�'ҷ����"܄u������
&g�4;�p�t��=�^~
2��;V�{�/�ibC�]di9��,��Mk�����c`/Ӯ��P-e�b�� uhn-,��W�A�$�	6vl��Ky�,E�&����)������o���E⡖g�q?행,P#H�#�z������~�mD�"Z�7��Z�\欧�xlߵ2]o����k��4Ƅ�qñeV��NE���Ν�A�V"b��n��+���h,�oky�n�ϸ�s����o-��ʋ�!V���=Y�I\� 3��FE��\/���EyqJT:W��ɖd�^�ס�=u��H0���o�m|��mH�-��f��(�x�+K|�zj�(��ߟ=�{��C��#�ְw�H��c���~,���d��3wt�ɤT��cT6Γ�;���d�6���>)� �JP+n�zqӞ~��;z�5�њ(�;x��N<��Ӹv�*�y��ٻ{wm�嫗pczx�lř����[o9�N�i�0��W�%�M��s'bѢ4rF�s�c���Q
��࿖�0A�m���,'�m���aF�Đ Q�W4��{��_	��1�Y=�h�3��R�<���,_T��ߐ�(��?�N�&�0��RyP8;\�%)�۸�7�{6E
�
�l�"v�����1u�<���^x�wؿkؿ�$x��W�^��Ï?��/��7ߒXXV~�"tO<� ��݂�����;h�B?`ld�X[qI�cx��n���\w��p%�&��k���/��< ���y��,[c��ܲyN�iV�����[5xD��%�ө��7�cB,��P�ōK ��G��OD �k���~H�n^���7g�s�n�i\�vEyOH��دb&���x:���#عfH�]�ͪ�5a����r���?�on��L7��j#�lJ����,?��fD��a��������~�s�c(���)S��wBԨ���83J�g��f*�3�8n1��}vw���LZ� �a߭��T۶mC��É��h��Ts���׾��:�d=�&���b�Xs������"�~���!��_y�A\�yE�q;.]��d�yq����޺㜊%�^�]�M�B�U�$Z����"�m��;7���J�a�6ɠ*��f�{�^� �E�)�gb�9�An�X�������&gxsri�Y;��Hn��5(b��8�s3�6��ѯ-�ˏ���4N|�Z�%|�/�X���W��dhtT;���JyZNP~Ɏ�y�A΋�\��R��Ejn}��WpG6p߭�esܸ	I�㦘�����Fd�q,���Z0��g�>�3�)|��5E�ŀv�!�_^��%~8�8�[ìdp���B�aV3Z��X�,���<��Z�?.���<�6���<@!��Ȏ����hl?=wK�y�IܞϥuF���5\��T%~k�~���������g�xD���(ԟ��������g�ں�/�C*&��w�v(��-�����Vb��SZ�^���z�>F��̐4�Ў�ÿW1]T�u��S3z��R�����Lj�䚆��>�p,̜3��l����C�S���LJ3���}"��q6���>�����p��Y-��s���,�{A�C�D��[w�t��WO��. K��VS7��¸��=���Bi4u�n^�!P�0/se-˩��K�y� �l?@��񋷼���*E[���=D��l`#���-�.�c��-k7�a�o�
7E�?ʳ�t,�q&Fm�:�1ʕ:�#��!�cXlŐ�ǐ�Ɍ��;�C�Fnڼ�%�H�)(����������QÐ�(�o뛘�ÉO�:H�\^>���✬�Y��N��ҕX�\!�	A���]D\�U[/�l�=G�4&Gd��W�ū����{��'9��qX�3���Y��A��bV�~O�R�"���.jF�K9"�X?�k��8w�:�(��܋��!�۽���>9;��;��щ�J@�؀L�q���Ď�n]���ɛ8w�d=q9��tD��4Eo�jI&p*��lޝP�M$(ع��p�07���2,k��F���@��-���f��g��<~��-Ȃ�桃 o����de+��3yڟ75ƭ<7Z�;�1ݶ"υ��1��<f����$�'g�I��要�-����úv���;���/kFz���#Y��Y�{�b��-�_��ܥ�x�w/����/}o�<+�]�nR���w����{R�٭�ʏ�կ)��%��Ra����7ú��κ����'��Y���Z�~�Hiqñ�(B�ya��l�#",�ʂ.�����:V�X�X��K���g��7]a�FK�Ҙ6/�'��o^T�0�����%�V���(�꼫�4"[H6�Ү��"�r#S�e�1�u�!&<�F$�0�Z������8�Od?7��yD�Q��.�	I%��Xi�E,�Y�o�;MpC��~?�]tPdt�͆c��>Ǯ�@�|�nn���	�0����.*����v��2,�q�C��=�����ݠ"D._���v�W��ˈ5k���{�%��[\��~��ofz�ꝺt�W�F�S��J7�S"����ǧ��C�d��u_���XL�i4%$*����{���q�������y=:R�s��G,�S�ʱzK��V0�U��B�ku7����Y<��o �*vo��W��1ͭG�������o�8*�f]"ϵ�ƒQ>UԹ�,E�.����6抜���R ]�x����؝L���k�C&b/�b,�
V�ɾ��`$��M��MR0@���V�8�utmA�s�x(��s��(�s�@x������)�l||L_��qM��&����\H��[Ik�½�w�hBe���w��WZ:;Xlfm��G;FD���ry�4�{�P���\z<�=���B[�m��^#�s����"�i�����z�t�9Z4�(��V}?���HgSؿg��3S��-�����}��I����F�4��J\�#k�N�
P6��1��t��8���2P�m����ډ�z��X��+O<��;v"��kAojNb���������|��u�2͞�q�i���wV5$�XB��*�I�xn�ڏ�T4�Tڡb�#��}smMUS�g%^d�5��,��w�n6&�����W*˭P���znh�,W:�β�jxΰXȨ�s@�݂YH]���VƪV�l�9�U��v���_�i�L�-��)+��6����e���$~:�pXK�(䄦��͞f�[}7"�3��q*;v��� �-[A[O-��e��Q�L�.��gp��4��O����<x�^	u��Jl7W����Ŀ���*觇P�I����j�΁��6���^��`��FW,[ ����r]�乷�\��k�X;�Fܽ��j��~K⾶�����\{_CRY�"��ML������G�J��ϙ��Jh���t۶�B.�A.�Ҭ����+N���n𼵻���q�޵Rx�J�=����9jp�L�1�BbTy��r�	��H�ظ�I��5�⺩��abǒ3</��X��~�30�eZ"�N�i�:F�NTHJ?��n�Q~��ёq4�*�J�5*\�.���8[_Z9�ֵ=�9��3'8�@xqI˒�����
0	¹�}�Ɉ��˙*������g�c8��扵 3��B�Z],��,[$�]삸�:���S~�s`x���_��8V�^����nv�۶�'�G�|f�Ь�E�n�9ilR%�9?���	�
xa��,�q�0!�4�@؞#ޡ[�u�1��L�D�� DD&$���?��w��� �b�������Y�Z\�s���j���,�`1YԽ�a�dI�N�n{��u��kx�%��nB��F��j����~F�b���=tGGj�1�>���>���zD7C��W
�&�Ҍ!q��h�w�KH�ҭŇ0�����P��5�uk+���&!|�L浜@��R+�4}MJ�28[9.[FC���R����Sʌ�,��ĵy9�4<�le1�|F9z����h��8I�������^Y����R/-�1��%�M��~R�/~�X���a���sI�X�'��ν��阪~\�AJ���%nDZ��|�2qWWQ6)dy��ҕ���43��/X*�Q�Ɇ��5�빸%�et5v���i��o+��������Jf��00���u$1��Ab$�=�؊�l4o��l��q��;�dh�L�X�ZgW�w�,w���0&O��d�"@���y��õZq�+��3�{d/d�I.T�=E���ql�Z���+��:|��un�5�ﻹs�hu�5qB:�+m	I�:���9��)K�4��u���6�:jKq��*$!��EQ��{��o�֦چ�6�m���x�!ʚ�m\�������U���a��rYt4��Y`:R.���u��(�	v�%�*꿧�~��F]�����:~W�\:q��+3_��R��2i��.t
M]��M���|�����@u	�܀|�Ca_w�.Q�ܸMs�o�{��9�l��ʁ�e��N�Ng��h��@��*H�d%���i�`R��o�i�T��g�M���{����/&d�t�Z1���"���J,�\�MQ�s�X���)$���_�e�������/�K�WC60��T���U+��6z5�nn�aG��M�N���
c6Ӌ��)�Zl%�Ǭ��r�K�������a�������&�ܱ{1�G3)=���=�Z��,z^[�.~��c�,<_����9rR�&o�wY;Μ�{.� Su���kc�Y��\P�L������.*�	�%~L�.B�'b���8�	��7n�a����5�Q�@���N;������C���V0憦;�^O�"��0�ZNN���;�
�Үn�hO���\0��|78_gc^�����	�Sk����\Z�UQ�BS\6k��Vgb[�����XCT�v�oF�&�'ݰ�Ė�^������+K���~q�7�+s5C��O8^�f��}˺��vԝ���w�ɫ��F�-VETE!0Jg�kK������+_��r�H��h"�)Iqyf^����JՒ��,(J��E��Q�!Vm�V���C$�A�&R|W5te
���9���Oc�&#���#��{eA<�/ߜ��sWq��emB�X�,��%�4�R|'9*�F�,7}|ֻ�r�:GG�݃ے��[m��c�tr������,��W��,�s�g�H+F������T*�g	,������(/K��A������t~<\�c�Y��v��;�>f2Z7,�	���\?ş�[a�id��O��[�Q�X�~����%�	a{mq������_N䥐J��ih�V��6��QHڝNx�(�4�fL���6��Mz����i�/��}��ȡ���k3�x��)�8wM�gQ'@uu�A\�+��T�7��ޣ&�XYłL��Ǵ��UsSسe3����������t�)�:���\�����S�$�fP���9���`G�&�R[*(ZS�F�I6�����؀I�ʒ�/��
_V>b��lں>t��܃�X8�FA>p-�����gR���X*ګf�~��M��:�^�M�0�ΐ-<Vn�h�2���6p��-�u�i�d���"�͆�eV�t��-�̟uD=j�"�37<���Vp��jؿǯ,��bC��(���k��ڎp(���8CJ��X�a��IAa��X��snzC�����ɵI��K��������_�pN@��8QP���KG�/�������REλ��+�>:��覘�;�$��ҥ}�P�^0���l1�L!���s��c�ѭ�6��4N��uOe��a���-�OGO_�
X��.��x�tl��!�N]#� ��L��3�5R֩.,t&8�`dT|�2겑w�[�g?�l��1qoo5+�b#��wꪾ�#���L��=u�bJ�?����f#l!�p����V�21���J۲�_̷N��f։2���`�q�eW4Z>-a9=5��' �"����Eq��wD�&Q��:�@'Xwm��od{a���x��y\��s�=�+��3�TaI̵tkA��Ƨ���>��sc�*�Z�^1��9.���|���7�Ÿ�����і�������0��?<���«�j���Z<?�.p��=CJ��c��� {�hԘ�Ȓ�L�qF����=[��}(Oc�HQi�c�[�TmbǺx�у8~���S����7gw��1���t��ځ�QGNs��y�ڶ	��>�˗.ai~��߫٩Sg��<�T\6'�i��3�?D���4+�!�1�����2Kg�{l�԰��O�w+�P�@X�+Z���o�$bg���F
ktxэ���}v�y�"8�9�����&�𳢊�Z}o2��"��|��nM��?e+�5��0�%�b=vi׵����Q�{{��94�o��b�������j�S�,1ޮ��D��ڵk�����a׬߀�7n(����[�ar�&����E0ؽ��Ƴ��W�����B>�BN�j�z��m·��.^��+�.��rM�\���J�Ǫ,�=V��Ը�� 0������6P���رYf��K�]☾vQ��s�
b���Ø_����۱s�f|p�#�]�u����oS��_��J���k�8qZ��|�i��3vcj�&�o܄-;v㵷�����/0�~�����1�{��}���b�gǘ&/V�_����hv.:�����QBY�5e�s�SЩ�m�.t |�B>������/�(	����n�	�%_�s��F	�T�M�-���D�k'�Audk�A��,U��1B���M�w��yTZr��<�߄ܦ�ȮقY�<a"��+�����7����'X���ǿ�u<��38�F�ݳo�fH��|����XEN��#��!���8���2�ߚ�Q�X,����z,��o�(�oY��k�%j+~�K��U;�'��ʩ=�Uzn>1�Y�RD��9oLn�X1+��h9�t��[j��Ž��Q]��0�$r��qeM&Relb*s�:5�7?��X�1|��'�������a����E{������_�[��:��ԃx烣X��?��{^nRcIrg���Vkh���u��l�0�"Z��J릿��MТ��Y1
U������1s%s�Ϡ�Gd��
�z
��Ӆ�]�
�5k���GPQ)_L ��`���ϧ�)L�b�]S��VRA��~^�`eTt����=�T�Z��<BR�SIk	E\f�9u��t�R���d�S]S��]Q7/���%��e�����܇/?~�������'(���}حְ~������'.vJּ[C�2��o�lN�'4�s k2qbŋ��eL��x�܌{ILdx���j�a��D��L�B`rc�H@���<��FG�������A6�,��!2˅�9�P�����Iɭ�c�h����ƞ1=?�d��H>%.fC���C�w(����v�v[�f�.� ���oO\$B�+�,�A΍n�q�u-�$u�S�X��<(���&|l�'�E(@Ƙ+gd1 ך��̈́��ۊ���"ݹ�~9L|��劖(��}eM��	��wSK��0��NB��Y]�u��ΤեfS2nr�+^�>�~�W��ē=�nbD�����ћ���ؖ�hV\�|�s0�J٨7�ͥ�L���œ�(�E�M<+�fJ֣��!��k� ΋�w����d��e�x�©��NP�	�;+����iM��@�0��R5,�j��w���t�/����ǖ-[����Ӛ@�����ɩ�������nB�j���9+h=��:�[��v�¶m�5�Z^_�¹8J��	���=�ʁ?�ٖ��hH~cl�q{?�<�7ج��nnf㬧ι��0��ϡ`Ń�� f��	_˄
_cTZ���a}���&hF�|Ye�Q�fS��t���D �)�t��0]�=$���kٹg���|�%�cǎ�ȑ#�힞���˗u���Ç�L��i�^��իׁ�;�EӞ��(�X1�c��P_�87�s�U�9�jZ�{��~��U�t1?�%x�Bō���nN���'އ�k�P�wr|�R��94�5��=n�8yBgI�X������{G1���о�Ŋ�F��?�	��<�^����l�"�m�:J�ؾs�"� Ap[\�&���JO�Y����ĵ�~[�-z}�����`�GyC�	�	5��3ĈYC�xfm�i�6�[X]��uZ	��{i]�|7��)Z:siM�L@������(�:g�r�œ�nd��Έ?�p瞐0�\yWr"2)�JXZJ(���/�vk��h��_{Ǐ��OK�ƹ�7&�pmjε�g-�[�d���;�7ݏ]��C���ŭ_��J:qc�E||�N_���2ɴ�mT�w�!��wO:ǣ�A�9L�)&�.]W,۩�W��w?��� ֏��޸6�ф����w]�2�w�~�J�	?]ԛBA<E\
�i�K+a�\AM�5�)�2_�����#x��s��1�X���Z��_�u�܈��w�c���ĉr�]�̒���G,+�[�Md��@�a���ϱ,#ZX�Ӵ#l�I$C��eZ60���A
��)�}T!�M�nnCF���8��,/�#���wxMZJ��Q���Þ[	*������y}���i�Flٹ])�xeq��D�0-^����]΃��<5�kӳ
���Z�)���񜲌�,2��c�TF)���L�F09��_��6���������1����a^(�ޘǅ�^��<./T�e��ҕ��=�a���ah������ҽ$4���j�����(]���^|�(�*e|�ч�s��֡Ԩ�pTp������p��h�̈j\"�9-%�ʁ���и\<��L(4�w��HO^���zy��%����:q��6q���$E�o،gڃ��Cr�d�����X�����|�7�6��)h�Ԗ��a��	|��F�.Z�#Z��R��F�6�u)�4�,��9��`�`x���X0w�(���ː+����:�e�e���Yǝp���PBGX���0��g�h$
�����ӗP�p�C-d�>�^_�8tʮ����>+����)2E�V��jQ>��ζ`����T&��?:�D�_{��ٱA��nm�b���_�q�}rU��Dʴ�t����a(����t�����,S�)(�`d9���
}�k�5̿�1>�pF�0!?���U�.�gjI�5�6���8^<�K��)�
�NY!d}��;z,^��yv�Vf?!c��
f[�R��Mb�hC�t8�ެ�J��;����u���-�[ˎ�ܑ^����;5�������A6��b?ÄZ��v����ٌK,�@�^�G�Z�2��]y~��A�̱fGI�$
+��z[��ʵ�"O���u����y���YYy^,��U�P$�b|F�l��a��g�T�Պ�>�V:!��n�,`��	Ӿ�q��G�b��������h|w8Q�e��qwq(�c��qϝY���k��M�~�f��8Cw�ߏ/M�bbJ3VJR��Ě��&�h��Pi~���Z<�W��_��!�
SF)���6��C���>���e���5��5:�����ݵ�ŭ���D:�9(�i�O���q#�0Y��ì�k���h�h��fAV�:��(�2�D�C�0�~����%�rqk4ƌ&]���X�f���h�;P X������:s�øL������gq'��8~�.Ί ĳ
r��UE�$�e��,#b��`��k����J#�{�ΕQ`@;���lt�'p��<.M� ��
$��9�;��+̬'�l��<��uB�M�����j�. �{a���֞\���;�������գ���o�t��*my���V�5EuU�CW�Tj*���0��E�$Z]$�ӯ����5J���Tɔ,RS�jW1a��4�*�� �Q����ǂ���ܰܬ��i�@��3��DG��8K��b�����Fٗl�+���j�w3��h�ȱ���G&4Q��	�^Բժ˄.����. ����{��wF�7�*M�7q�6gr���4���ƍ��u$���fҫ;���7d3���1[.�1���3�)ػ�L%QO�¨��4��%���	��igK_�0'V6)��#8�����S ��Mk����ez!������� � �>3���%�u���9�]��8��7�4~��R���yts�}���m�5u����g�#_� �H~b�e-B�D��b���
m��`n��`���-�N� ������b��l�mnhKr�p��΄�h�(č`�$?��+If2��)B�5�/Jo��h�1J4��2
[0F�bNsy�w��Vs|��|?R^�/���<������츁������-^E���V�v��8�ƈ��]�}0:�V�rD�����)�]U$I�{���|nBb�J��?�Ԧg�2,0O�ݤ*�X�ۺ�)n[�c�����۬�,ǔ�\]"NR'f������'2z����1�r�y��A�Hߵ8�Vߥ�e����2�R�u6�g�q�iH��qv��x
��mA�5c�$v�8`/ս�,��`��\[��p��	�x�����dS�N�97f7I,�ZP��Y�M�K*p56�&��l(�޹���T�M��=�z�[���~����^�zv8w��q��]�^R�����T�h�O�é�ɴ��h�y���r�nGx�B�V�
��`RA��Ҳ�9KRqE)<r�n$�-ᓩ9�G~V�5s�p�L�W1��:�S�/)J\���R6���z�SZ�㜵���)����)�U7����2���%I�nU�n�Q��Rh4�:ƭ��+Ҳw�X%���\�A���`m1լ�SXڵ%��01��[ί*ϳ�����H �'U+(�݆��H��h����o^g�qXt�:� H��3{�_eCw/-n�ډ5�w��P�Q"�Z�q+
���K]-H�S�
�Dt
-M��Ŭ�u�|���2��D�m�!3�oC������t�J�0��}�YR�=���Y2C��9�S�T�r�e3�"�}��m�<�j��*k���a��<t?�O���ݜ��o�T^	��W�\A[�������U�U�k�d�5�ڲ��Fy�D�P0۵
�	�|tL��Ʌ
�NN�"
�^YRF�XW�uݍCv�òP����|�Z��A.:�-E�!n܆��x����.ܿk��╚�N�>:q�;���g$���T�L.8.�Z�j�ʢ�p{,�t�mM�M>���k���M��J���Fl|�tk�z�&J7�!ݭ#O��XC�Tݵ���?����h�L��e���iH�(/K��f�=�p"Lz�wF�a%=��O�N�1~�N�L�<�u��(���>5;�\� ��� �V	���3wħd�u(l���A.T�����ne�W�Y�c�Eʤ3(���(jX��Z��P�rTq\-����R6�\�:�H�rM%-��(��c��[����3OĮm���y泥�ݜ��N���O��<�MЗ�x/��8	7ft��ղ��l|Y�`���G!֎c�?����cX?���)!&���M)���ㇰ~|��_^��y�8e5�6::�ri^~��|��rURt
��眼�!�W��Z;v$�Ŀ�t�
Z�N�9�F����8�=	o�f7G tњ�
2��m׹��5�Ld�*X\gβ���K���i�͵G�a���W$#UfQY��8�,j�-bBc�����6 +X��Fb
�� �w>��˻���skw�s��u\o�'��0Y�q�?�b٤�"�v}�fJ�E��캱�L�s>�I�q�hV��/�u�N�VK�vpr^�sO<����l\+��)#�I�G�8^��u��n���1��c���8�@w����]<bJ�lN���hu��&�pߎ���ֶQ��7Q�2&��D���Cxd�v\~����o�Ԭ����i����MZ�r�֯�!�bB�� MR��kW�74��&����;)7w�P���d��Զ7��l���[�gҦQo��ot{�!���h�:�\LN����l�BK��a���<�H.�ZsYo��9$\�����p΍H���(���aw'N���cE�&zOc"$%/"������P�;�s���L���'����n��x,���Ȩ�_Ogc�S�S-뵬�q��6�J���,��ĵ��1�Kb��]���q��14<����^�Mk��ܱnDn/i�e�FFV\�ZY\����(޽��xW�;�T��\�6ޢ�����������n|BM �G��Ō�2�D���BC���n����%v+f�䣇�މS(Oψ��Q�e<u�ˢ�ֈ/��яO)(��?�Ν;�c�>��G�� ���p��Q����oLkccW�O�ժu��%9�s�(�\5���
�U#]NnF��1������u�X�`Sv��hnd2>�I��6������E�h&Q�v�E�5H�B��-Ǿ��6ZD~�a+Y��j��~�2�q�sg��;����oY`/���ZPm�|��˵�60�l�Z���.簸T�~ ��!<t����_������#-B[H%$���K_��}��I)�
|ΰ��p��^l�Kt*��axI�	�C�IP۬-���۰g�f?uF�_:5V��`+�Op�J�xZ��T�������l�5#��K*ti���h|2Kĵ������Qj�Q��12�Eb^.�1�|�����8��[رm7��ȣ���?�Z����������ޫ/��'����q,N_�����7ʈ���H����r~��g���2�&�YQW�3��lEp�31�T������}����抄�m@'0�Ii)6A��Fb�h��	��E�؏m	���/��)�T�� f7y �bO������)�� ��yV�NGL� �4�X����� g\V��H%�KSq���غu;6��峧q`�Z�g��Ͼ��&���g����>N����\Z����}a*��e�쇶ι닥(5ɽ�%O��e%�ـ��Fq�D[�|���1R{~8���p�{��tj �&���Ԯߖ�21kĴ--WBܮ��Y�o܎lZ\�{���h��~�&.��L�:�_��};�GuaK�fqk�:r�am����q<~�0�o^C�QÃ�fu�dA6[�ٰ8�F����z�6ғ|��5�^�?@]4sT[�%3f��Ec��f�n�h�,���q�]�.p������
佀Nb��t։VҮ��h�@�f�����ie* Z���������Oy����g7���Z�LL���2,/�Y�kif5�r��1�4fn^��������N�p���o\Q����gqsr�{\�ʅs�E��ѩ7Tu޽f���)L�P�XZ	����`Te��q��Q���*��n_{��=<,�e�lR$��C��h����[�.�ia�F��d�Z&H��n��&����x��x��A�N�8��l���O#gI��(�Kظm:�����Y���}�n<��Y�8���Iޟ��?)�zt�Yg��@�b\�`�������T0<o�(g���a��i�c�GK�X����{���Y��<}��3
cCZ(K�0�g4{�yXЧed�Œ/��9���XT��)e��Z��#��0e����/���{��}��sh$�"ty�~��o-"?4��q��0����kM�������Çq��qQ�cO<�M;v����r_�ߦ�eI��Y^ʥBP8�'�rI�\�ņyb�A�1��|97�ܔ��2��Hb��4��"���S��l���E
�z��Wb��8\T��f�:��V�+`F��$m2�Q����$>�ſo�N|��Y�<y	{����[������%|��ǲI�8yR�?s�\��`[b(q�R�7� qX�q��3�Z���^�P.�V�tz�L�B-B�@�L����o��N�;���DE,�����2��[�p�;���v��4���:��z˂ZK�N
�Ϟl�j�m�;Z?���YQ��h|�$�� ����?�ʫ;$�=�'DPB�v,�r���x8�7�H��Ǯ�w��� #.1�oɚg�����~Ͽ�
�*�;?4�^�-��7(��o^x7�ߐ���s늝<y�������l�K%4������4�-�(���_����y4��p#��E0�o9��|��8��XhBx�u�󦝽to=�g@aMN7N��6`ʩgs�<W�+�����*��Z�+`$7��E�.(�2#�O�3��m��)��rSmׯ�����S�E�D�=}���*����sطq�6mp������N
&�H1�ɒ,^����,�	�J�~BlyC�D�<f�9nnD��������b�R��|h)i�L)X���5/�]�B�/��[�h�P��Ւ~6�2�e��=Q0+�N����J
�	��Z�|m\�Eݗ0��������Ԓ��Ή2fO�_�O�7���F����ז����-\��o�eK���C%_{�#����8����֏�ѹ�rɡq̈�C���3
�'pP=&u8`�m?��M�<��z����ʱ��R��!L�/��/��7�о-HŻGW��s�.ޘů_y�N�G"?*~�/~�ڍ��HC��#c�=.����V)d�9/nȈ��ǒH粨��_��\�p*��ׇ��]���P�9��v���b.]��b��E�����yD�x��悚�5fWpGX W��}���k"�1&ׇ�ǃ}�|�P����~Q�IL!�>@;�h6U_�	����"۸>�J�ir�@,�j��5�����J��BI�NV�c򟒡��Ι�L-{d�n��b�8���u	�|��.h�E�XQ��.�y�<��C��/�U��<}c�+��R��c|�T��o�����|>G�l[��1��-S$���R��Y\.%B��!
��pnr�Ͽ��C����*��us5|p�<N]��~�J�[b�Z-_.:�^���k���;����>���γ�[,I��C��@\��Ęn$GlJ�$;4�l&��K�b49aqV���َ����`�C71��BŚ���+��c4��G<Uu�ĭfY,ia��,��>��P
����4�od+vӺ1����
?Ǭ�#4rJ�*B��L裟I���� b6����������NW[��79m��:zIW�Z��¨Xd&=�C
��\�8L�\*�(v1UD��E:�(�cHK��
��I5����/Ib�C�O��X�㵣'p����&D9�>!B��ۈ+�&�&��"�3��}fs �9����m��q���['��;GŜ��Ũ�9�]6Xq�m�����xFۢf#	�;�/�f�(���!	�7j:/Z[SX�m6B�E �5N����=�˹֗Jl0R�;��6��Tw
a,I�2�2yr�#�ZgUT~�����,B�*I	�Z�uZC.]@���A7�:�լ]PſJlW��0L�)�BK��`*����`M��ZV����0��ۃ��y�w<���z�Q��r�0d;nQ��T~=Z)����B���&[\./��5�;μ(�x7)oo���\BQb��S�퉵L�@H�����*�����r��2���U�t��)ee��U�
����grÊ��{y�
)m�g�>�Hi��L����W���5�к�32qǓ��K����iml���-�L(7D�%�}$p�5��c|������ڜX��b��E�gYǁ{y[lX(8�.	Jf"R�[)x~�_�����6;�C7����PZTg��/�z��2�X��%3�F��L%��<��i��@�x.�F%���
�D�L�����s�M���/"q���#�X�6,O�;���m�osI�\�VC���z�!M��G%P��Ck�����62����!.%A�I�p�)N��E.�F�ի�?j��D@c�C��1%d�ؕT����g�/� k�vw�u���9 c-�\ ��h_g��u2KI[.���A���@2�p��و(gPm�����^N�u���ß���5��BR
n:�D�K H��G�<�������p���<���h���Z��^�P.�c�W������)��u�c��_�(���3	���A:#nL��
D��B},g3���5�#����͘��|�q-M�K	�N�f`W����b���(�(yn\�vEa�\pD���Q��Ӿ��[�8}���"4�1Lu��M��1����v ��IX����R��N<3��:�yw]����)p��u��4��x�q���l��{��QZv]�7i2���� �m�(���ڼ|�@�:��.�ު'�B����h��b��N�c��v��C.rL�$7�'(��*-�Ih�8!��쭌u�)t�Tq�h�ɫ��S@*�<�5�U�9j�D\,]�V�Y웺v�,N��i���]�5�P`7�j� }A���m����D4�v�w5Y� G9)7��trJ/�s�U\���S�����:��W..��͎�q��~��LFҸ,6psb�^
7eyq�ѹ�ehU+���h�G�_r��D��+�+̌��4D
�ͪ���Xsk��c��6!2
�5s/kJ��:�/^<���/��H<ڕ!�����ψ���%���~L�$��Ύٻ3�ңzI\E��#�>�J���u�~/%���{�G%f&K�)�v����v୵e����
��a��t�_�y�����`�q`� ��Q���v�vE�b����4�xb���:�]*�iC�#_���i�p:��1��`�P�I���Z��L]r�k�2���
�1�_ΦF�z� OnJ��n��Z��h��9�j%� ;����՞�׻�u�F�9�ĉҞ�c#��i
�
Z9�����hlh�zF^kނ��%n�86��hTk�yN&qh��`��l&��U����C�jV���2���S��{JR���(�R$Di���;Lȉ�H�Y�F�����_���Q�=�1�뜡]�f�	�f�I��!MoC�gl�����\Ӗj�$%n���ת���5^$^83��Kw�X�{��Ǟ����(x�<٤\�����w�����uVA�K�%�I���ǧ�љXZ�%����k��pt�X�q�n�{L9��h2��ZՁ��\�~[]:�Ht\��7����)����e�)��
�QݴJ�_^�YH+�V_�tv��K�ԷvNm`mqԓh��Z���W���(ߊb��R��1��D����Ni�c�FK���u�p�9�Uז-CdV׌lYZؗ����u��� �C�y�^bPg�W�/�[�X0(4��mV��r��z���b����SB�]��&�j��f��SɄ�O�ڰ���rJd�y�f�>�SnG�o�����q���f;S:��r��^ě�K7f�K@&M��񠻙��Ě���$�`�M��|��b�/ϔ.������o����s�>�� '�'�!�I���	�ݲ��n��x��:�#��#F~�Z+�1�
V���$u6c�O�A�\Gw��D��v�����HP�����ltu�xC�0E�y�K���e���e�Zy����_-)D���<�;��kt�(tx�ˈ��A����,�Y5nFB�X>`|-�s�9��h������ �y��Fi�+9�rI�a-$x,��;�渞*/Gg�������{>�f���Z!A�X�%��.iE�+����J�W�r����7+Ðʏ�=k˾�61����7q��]:�)�y��׮Mc����i�&��Wq�ڴ6Ew"��v����Eߛ:]Rk�2 �u���'qՎ�����<���o@�J\�����z�T�]��#��F)�wo~ �h���\V�]iA�*A3*IU���W�Ep�ݹ�i
T���z������� w$N��.6�q��֊�sckv��Q��E�`�ޱU�kZ߂8�i��=�c�ˀ��-���ޔHk֐xOm��8Jr%����݀�baXDi*��f��
�X�^� x�w;��<	"�W�tx̜�6̥��9�Z\�G&x�יּ��F�V؆�Ѿo�fS9�#1{W�-U�
`)C����uU�Y9'򛔖naH�%����%�F*�v�;
��qz���$/����pd�v�[U�/�r���3�{�n����P�0��z�c�t$��Ȑ�sf;v/�t�K8G����b�Ţ�y��~���W���iWO�i\���:^Z��*��=�O��L��L�%<q�0�ۻK7�+���<��<�������g�v�={�7���)nio��JK(�2�KܲM^���V���n���*���JE�<��o��l�E}��������6݈G�nH�:��7�TQ����@���ڏ��se��{�"�΁�Z��Q�く��l���b�1p�W�V��x��31-�C˲q+i�e/��(yC�o�T�2�^7>�o}��n\�pKs���w��L1��}�i����V���7ޖ�+��x%��y�=q�}�i�by���عa�:(rX{�֌&��t���%J��v�����`�Tܩ�V�GQ,p�6��q/Z{\���ZW���v�cE�ٺQזX�2�%�Y�U_;%��"{nj	��������J�=�M�������x��>lY�]���o�˚丮�Nf�^����4b#A �M���YK#ylO8�Eo~�_p����Oh"�p������,98Z(��� ���F���]{Uf�|�ܛ�U����Q7DU�*++��=�l������������`��E���4Mߘ���� [���/�?���������Iݳ���Qʰ����
��W�\��z��Ҧ��X�ֹs���hݚY1c=�4���>s��^�ftpN���Yw ����,�Y��,iQ���A�`ZKcF��5� A���|,�t�B3�""�����+��,�#zt�9��dk������_�c��A��Rm����3*D��~�5��;�P*�Б}�w������9yhl�ǎ�իפ��4����>����#�_��G��@�Z%t�e���~`�о��e��Y4hlhP
�o^�H	��@�4�B�ꊶ��4�	��d�ʼ�Ng�U:�^Iqej�K�5Ԣ$���檼���S��_���B>K�\F�-Mޙ�,��/���U���w���̧ts�08ߜ�B���W����t���p�2}�$�AJfS�/�_^��ׯ��l���vk,���=�a���ҡ��<�p�v�3�?D%<�&]�<)�4w��6ri��Zf�p.��T�:峹�8�1^�n��V��s�U*[!�5-�c�
67�(6Qh����Y�KK�4SY�Kw�
�2�-5?{�~�ӟҟ����u4q�"?���ܠ�#C�?�1����L�}�������%��A�.��5���θ�PP 8#�7h��׷�Q���6�P�FI�U�,#r*6�C���������� � �I!�� j4_e�:�� I�V��I��Yx>H}���+r�`�9�B�<&��G�K�`?�я���gg�����LK�w3���9֮z��Z������qe������h8ǆ�m�cK�n�a/2w��Q��w��f-Zp���HЪy��Z[�G��
�6�;wf����MR�g�1����;
;F�	}9�|����Ʋ�<8��zdl���I���!�YC�sjsl@�_�t��+�k��/ ����>:�����i+�={v	ǧTM:r����������Q:s�,�_U۷�K�FQS\�$��E����B�%�`Y�-g�] 
�)�؆���@�=i:� $�����Kȣ����ybKҊ6�;9��;��"��I��4;� �<
��t���{Ḋ߲�~��'�A<x�N�<��m��|�m���d����ZX�c�<G�Μ���\���&�<.U*�@\�&�/Ipe��y3�9[c��Ռ��2N��,�yd�q�"D�F�L�v����|uk(�?�v~n��k@���D��A�"V*@��?�³C��k 	��{t?�:�9-����#�i`x�Fv����Cz��W��Z����/���:��Q*��U2�_�
�Y����Co=i�"3���� ����6\\.�� �JYK�
��(/J���>�R�X��&t���@Fk����d{��鳴o�:~x�t@-� �����+���%h����'?e�x�Y ��Ԩ��~r�>���A����_���*	��r�nN��8O3�7�$�����6�P��#�Ë�TO�Z]dD0��d��3�WIB�#j���u���'�*=8�^'�RNk�9Ko����\í$��������:>m��m��ޛ��"t 3��H&x���]�Fhe�NMO�
�ᅾ��J?���!��*P�y��o~NM�$YC"��ť�Gr�Rk��gg�����(D�b����/�'N�KON�V�|Fs}���,遗�gOх��p�z�Q�_����=�Ɩ�f�AKC�M�7 ]v��Neh|����S�/di�����A� ��J�hjf�N��J����vF:�����	��j�!��X���U�W���<^�t��%�Uص���la@������tht��v��(�Lx%ݤr�;f�ߔ�ڨ��w���P���kh�s�w���z~�}mm�)*Bg��[�v��� 4�j�s�L���h�}�k��t۔�NAnR�pd�a�ǁ��R�P�s7n�4���2��X���tg�&fw����.j9]�ͱ ��yI���0�f�$�t�*�z�2t��~J�:��
�)�,��>��<��ST���p�0l���<7����xR�$;��-D8��^B�2����
�X�|d���� #�qӗ&���	:}a������!No�F�\Q sh��&�.�ܚ�l6t�w�\�*��I�`z�l��Bfs��c�\�'^���e�.l!"�ޒ�
��3R,�k��D�l=9�&Y�s �fC�X�(@"t��7X�E(�X9�&��F`7_u�D2���|�����\�D�m_L����]uW�xH~��Z*�G#l�Գ	�23G�@{S�9����Rl�(�	@'�vg j�r�cK�O"�&eڴ#Ĵ�-�x)�rr�n���N�<�4���Q������M:wm�>:�&f˔eA+�S��/y�V��~8��H�	�F�EP@Z�jW�� �s�w�e�]:�:��w'�<�ڪЭ�9�����E��(�SI���ˁz�w*)�@�>0���S^⦳B�P?$2�[ZM�̲��/�WD�&�]��O~Iay�2^(�v�ς�	�;Ｃuk	�l.ŊVeؾ�ӊ�m��P�I��$u��L4������:v�
�J�Һ���t+�*�e�X?%"��ĸ�� '���� ;\�x�J�
5�U�ZIQ��&�I�#�ʗ��Rf���ͼ���#u����T��!����vS�[ +��@���zl:��)	>�d�(��z��8��<����%K�-Q���>%e
�;��v�W
?�(Wq�/9��sڧ_Xk�{j ��3�7/��!9��n貺0��Yc��sjs7�m6�uX�(ؙ���4��{I�;�hF��M_�ìEM��*�(��"�Yn3��,�g�>��vX_��AK{���_\���+�}��g�O2��D��ܽ�D$JkP,4�����2��B�m�RG����D�D/��Y��Ē
d:��Y��c�b�*<�h$h����k�=@�p�ͦ+�e�������x�BP� $Gɔ���D!�a�B��*w���;,��K֖J�K5l
i�%�[��R�-)�5�^}��Б�ߡ���i�h.0��[��l�UJUApׂ�8ӄI�I����8��1�H�Y�c�~���{����wQ��n6-�V �=v�\^��������uR��VY���%�Ӓ�
��g���� �9��*�֨�%�ms��@�ט'=�
�E'�/`q���P�mԮ���7:7�F�U'�6�<~���l%%��g��J��K7\�k���X�
�����9a�eey�r�$���-�j����s���-]�*e�G&�T؈S��+�ݨ�&A��_�F=HS�G�-O���[�d��4���x`hk�%�l&)�0���ܬ�pJ{x���B��H�w�	��`���_E�Yl�{)���Dր�d�'o����=����ƌ�ҡ%d3uq 2�<�@M4��)YX���������C��R�#�F-H�-M�NRn�5�}�.��$�����$���u8
ǻRk��19&=�4�S_�O�`%x���z>���&��̧�\�-�i���ܶ8V���DG�+>���j�s5����ԗ:C�r"�R$�1�I������S�h��Z��R��E_:�`�P�-G��W�y�H��Y��Ңr��F�ϕD0E��I�L\��[-v?X��R6�|q�*ͪ4���
���5�c٨\3on�A��2�l^�����g!ee�啝�n�4؎�7L��8H�\�Md�	���b�e1Č�����C�N�;vѝ�ɹ�C�|��ؼ�5�|�IN��-ixؒ3h
=Bݝ�x�Rk��JN<�����u}�y(kJ!kG`ړ%���{6bD�]mC[�cܱ���lԺ��H8\��I��&"���&��{�gj����Uд��w�����[F8���i�����\�.��	�h�շ���ҩWA�Hd�����ʫ���~�H@�4������L�~ �_87��	t������L�lphU����ڄќ�vpŒ��xl{ɻ(։��8�5�hUa�
فM���g�@O<����b?��5��o/��.��,�7Rbn�lU�D%u(�r��& O|=Lb�V]\Z�5"�E��,�0e���J)��-\��d��nDy��VQ5��(�8���Z����6�yc�	��|�5aEn���ȋBJ�lj�DcY����/��H�̞�u����7[?�j�z�]yۍ�(!�X�B/UG�Q�����f-���v�N�l�"6,҄�RZ4H���b�PJt��p\!*���S9a�J����YP�2����ך�)�fjX[�~�������H0|ͳ����q�2� �%�\�����$��2�kZ��l�(�	m�O�"ЂP�2�wA���:r`/���q:��a	�#�+� A/}�������9���lk�Ќ���l^i�bB�ာ��sPW��KA0x�Xq�e�����$燝�vR:z�+��6�I�:b>_|�k�6Λ����U)I�ϱ���m3����}�Ւ�캢Q ��T�Q���E��_��c��T~_��D�f�g��k��Bsr	]�5scy;�o� ځ�R�dLN>�!�堓��[��8��@h�Ō�yf�dB`�+#@�V(��V
W�}�@
6!w��o�J/=���#/h��l�����c���_�/?<%�fɶX9H@ρ���cyh�Ɛ:�rA�},n�W��=����"�t�I� Pޕ�)�R�Q�\*C����ܛTf������ħ��F]*���̤��W+-���V�Z�%���Ε$jY%	�> �};��DW%k$u'�m����Ys�*����T�l�q�n�$� ��K��>i�c�������:�(B��*�@Ϧ�E��`L@�{]?�(f�Z��\���[��ۍ|>��5��E�1=n��l����i�z*,�������W�o|f<��8��S#��,L����K���ו��x�$��锫���ty���/��r�Rl�4n�Ρ"U�*�����}�W�^i�o?9#���H�nl���#t����$/&��@������G����(V��2��|~���7��"��W����ܡŚ�^��K��=J���$z��u�1��v��ˉ��422L��G/^�����˿WX�	EdwR�Mݔgso���i���A&z��֩h������SHɱa;�n�R��B���oP0�1���g�^�,i���ф��|���0^H���� &pF[SP�Mt(��R��s�ũH+)S�����u��y��W�W�{W����kt�4�s'ݼ~]Z�-�/P3����iv3�4tbbB
�lY��
�3J�=���uieyC.�P�-��ÖSؠ�l�����|���]U�Q=4�!�ү� �v�c�'�؁}	uH��,=yp/�_���DH%���y*�����Eu'I��a{������6��d���WiLŅ>`�5��H��+t��Oȫ�/<+q�`�Ξ���C����7y�Z����i�A�!0�qN�#N���h'���Mb���]����i5����s-�|1��2����[e+���<��4��v�
�	�X�1Ў���K5[<�ѕ�f����F�P�:T{E�!P&�z.t���}��3��	0�l1=�f���ղ.}��ߡ��2��������6`P��U��9E�dZ�D�?@{wSm�A3 �~gi�����V���*�����Յ[�f�6�lf��Y��1��鰨�E�0�J�K����a��ǧ*�X?���%*/͑�/��5���Ɗ����f��ɏޣ�L��x��o������i����y���_�����? �ՠ��9���h��Np]Z��;:�Df��5^����K!R?H4�ێ�!�:���٨�(q�8��JZX��0!�����<i.-t�	��"�V!b�{;"�h���A����/�rh�U��=	h�C�D�FõE��k����ʀ:�x�8B��� �g,R�U]!�	�����ݰ�y#�5B�3�t�� F�&i׮]��d�45{��?�	���[t��ݼt^�ae��d��7�\6-�aK++��`e���s(�.�GK��߽�N��S�d�ɂZ���5R^�?���4�(�>�-z: ^�ة�B�o):/]����٦��t�\���f�9i�����Ta�U�0]��R�!�c�_XxQ���Aiu�>@�Ϝ�\_Ձ���z��b�=4���c`1�W5�D����h2�}?T�0�����=�y�tnR|#M�4��9z�w���;�.���4���R���aJ����/Α�BR9�����gT�����9H{wR��H��9ٕ��%�y��D�
l���B.^��ڠ)WH��i�l����3��V��k]73֘�]��Յ}�D��m����{������L��XK��e6���"�8r��g�f���K��7^���7$H74P�|6+��lb�����p �2)�[�Hs��C����D��Y���4�\YEI]&wI��ت�3U��p��%��Z曒2w~� �vA�>˚-+�ͳ�ej�,V�Y#�D@IZX^�7�z[��>=s�?�b��N��}ҷ��te��k�<���RP8 4�&p��	G�U���]8�j�	��}:��"�_ޏ��������2�7؇hұ����~�-���B��8I؎��!P�aax�=�<oL)����+wn#��"_�@U��衽�����N^�k�?'jԄ�(߈������t���J%�>u[���	���P}�̅�f�ܮܡ��n�N�a�#��@r��t��
�k���֬pa�~�%���1�90LWǯ���K�`�c�D����x�nݾ;�%I; ��d��qs��姴K^����tB��m;6[�R�����
��k�$ S����G������f���v��?
X��{�}�g�8H�Y���N�fJy;�Z���]'��la���~I���0+�����}�c�ru��Xǯݤ'?B��"qaa�����˄���	�����ifnN����d{���].��T�{�l��]�l�޿��v�eJ���ZU*zUz�Pa�De�%��X6'�~�R�oT+�L)�\�ϵ�م��k$�Y�E�z�v���3��c��B��6q��a3�0BC�-gxSĮ�B餑ViJ�G�\�1-/%EP(��t�wO�w���1뱴PI�����H�{�/�Ke���A�u��\ `���2�I�Ы5�;s�Į#"�`��4q�&o���{��Va[���L´�N����c}pn�Ƨf�,MIu��x���aѷW�0�.pŁ�N�4x/<0�I:���}���hx�^Z]^�����~�Y�����I�lB8"�@���|�M��X����k3�B���`� -�nT��M��,�1g�W�d��\N|91Od�$DҊC-dlu��c����5��Zv���iVX#�ȩ-S��DY�.kRϕ&��~G��+���[B!��俇HK,�����)�:5�M��B�F9Js�$�ا)��iаŞa������#�"O��+Jښ����zkv��-0�f����0����kAĝF�}�l]�1C7��$E4wg����W��S!��g�7h4)�H
�������_�����������R�.���t}z���oꂘr��]�H�r��n��=�{ <������j9���ES �y�-����׿A��(@�1��J��\�����3�~�}�� O��{���1����z�J���4�fk6��(/>a�?G3-�H�O|����B���E$�#��%L�gf��Z<m�y�X�q,O��5j*hW�[����EM���A�� ?�U!˕����/�|��G+Z�<�J ��~9��<)�{��Z ���MR��j����k����U�z!o�n'Kzi�,��*i9Js����J	~嘜��1U�&����7���jQ�2&ۧT�%����¦й�ĩh-�3�1�УΗ{���W���?�+���/ӓ����R���x����OЙ�"�o�5�az��psŦv��alM�4B�qH�!�{�.�=����%�=Z�ޘ��G���Jo��[4ug�*l7�a3��z6tA�;�p:k�I
�-������e����h��s"aZf���l��]��&$���;jS�wY��|��e���p�Ji�jR�3�4�)g%Д��>�^����T��N�Ӭ���r�"�q���x�ս-7XS��G`J�C���	�8��K�w�g����˷haj�7�������?�{Z�'i��$����G�Ǒ�$ $�p�4Ռ�)�5�G?�פ3�ճ�;2���Xsյ�>nYӡ��:�B�����^`��jBƄ�pa.�O�s�w޴S�X_`�9��3�gX��K���G^�ter���4S��g�Ӱs ���.E���Z�n\nYӱq�d��)��F��D&ǻm�w�eV�Eɗ]��a�}V6�*v�$�s��7�(�pa��  >{�#�sW٤�	�W���MNh�F --��E��WrNM�M���:���\�ɋyf���"f^-g���ȼD����4e������y}���6i�#�ͤ/�x�KvVv;�L* �BK����� jȢrst����4Ay�S�Y�dBM!�Q ��&�N�k�~*����ͱ%�6��`sճ��f:&�oZ�4KsVN�U˰b`����%�ՍA��·��Q4_*�6¬�/k��`�RU���L
�o����Ʉ���A��(!�o���Se�hr�6?�i����h"r�&&��F�F9
�\h'���JH�7h�ރ_nI�RI��sP�7���b	��b���� ]T�s#=��$�EYP(�I{9~�$�h�CO2�.�����_f��QlEuq�����旚Td�+�d�[��(����Eyp-C~��ozf;djDCn܌�4;3y<�;�g�&a���.�;�
jd��gG(?��b��7YUx�����Xe� %��Ҿ�\���q"�Ϧ��=�2p��� � k1_2�[(����i�`w�Α�ִ�i)��:%��vq�6��o�؞�x�G�<��j;�~��?R	� Z)�V��v5��t�4/|�M�b�cM�SD9NX��g. [HIm񌚱t*M��'t�T�����D}��ȳ��0w|L>�G����,�V�qK�ǖ�nG_����S��GF�ѶS	��?|�i:���>���n�w&^4 �EIH�$��y��l�8���M���Jb�>X��9�~�!sq����F�6O��~[�B�3!�^���P5�a� ,b�I�7� �6��܉ �A�<v�����o��#�9jGn-ȹ�m+��5?r�ȊXk�����~���Uk�w��z���#��}�E��� CIj�����вՕ,8�l��u�Iz�cKB7�W�ɤ�'n�X*Hb�_}�qz��	��k��	-�e:�JE��Ά�`3��z������Q�n���p}��`��e�C���׍u��p�nW �k�~�D����?�.v�~Ks���p����W2����`�X�B��쪤Q:6�&k;WS�et�)d�˫+���y���r��ɱ��pf|�����' ��`� ـz7ٰ�ӡ3��6�߈X�9�����U/��N�Ɵ�p����ھ�V���5Ts�tm����!m62w�p�b]��xa|�u^8���_�f��W�pp�h϶е�U��,\���S"��r�_I'�r����<�,t��v�\���[�+�f����zEkQ�PR�j��R
����LG��h �K`t����6�6;��b�M�Ưoz~���l_��f�V��n�������6�Z�e�{�X�����*?� �;:��]j�������Y<�Z��!z#��z���?�:�히�^x����������3���W|�?WɁb�^�J�t6��%�!*����|d�m�ω�q8
���+u�jq��e�G���q�5�����aA���jq[����u�붗���b�[r�Z���R&�FOʢ����MU����v$�s���n�1o��&f��㬹��1�-�
��{�U�9kwg���^'٘Ut�[e�1@��z�ox�!�0(p4>)iM�Rk��fj��\:��/?��I�k��0�����扽cNܾs����K�˫��	�HVM��~���_�S��O���I���Č-���F��F����2Q����Z�0W�	ǉΣO�かE��j�j\��k^�]w`|V�b��O�)���3�(W�����[p"G��������Q�
6T/��t��ʫ":"c��o�L�����b��Ub-F�9��4���f��T�,cǷ�넴��덮�B-�>��r��'���e�e�C 1�M?pU4	l��33T�~p����}�[�5�{:�T"Q{ll�I���j��6n�_C��v��>�?�n �]#~��	E���M�������|��{�{��l�����}	�F���N����Q���l���9��xX��5�*t���q�����m=���������m=���������m=���������m=���������m=���������m=���������m=���������m=���������m=���������m��$�Ժ�r�    IEND�B`�PK
     ��Z���y �  � /   images/483af35d-09f4-402a-a8a9-75c28eb4643f.png�PNG

   IHDR   �     ��   	pHYs  �  ��+  ��IDATx��w�$Wu/���Nw��LΚi���	� �D�/&0�,��D��3H$s1&^[`I(�<#��h49ϙ�S�X᭵v��:G2����}���OG=]]a��+�V� Nm��SN1©�ԆS�pj;��v�Nm�6�b�S۩M�S�pj;��#��Nm��������X,vX��hoo���vj��h{I�������\���f`E$��d�O�q�����97��������yɶD&`b�Fmd��g�4�<bsv�:hY�p:�
�jV'1B��i"R�7\:��Ct,�F�!���C�à?��L��~�}�m�!��8F(p�@ h�5,>�ϭ�kq�0L>6Xs��}_�z6�Ou<`�c��`��e4l#	���Sl�5��׶�1-W��,�~ðL������U��]�n!����q��+��`����a�>��I��㥉�;��r]��Ԣ�hrj|���yn���8�k��D�7y�|=ȳ���8����0o��Թn��,���:����l�k�u�{Y��<�$;�`0$���<u,��4�p#�h�*��`�Qjkk�x7�ct1/��$F�Iq��Rn�P�6V����E���2���{/���k�ɢ�(�JGoo����&'ݶ���ޟ����GG'���H��¸LyA[QO�˟�k�|Mޯ&N�^�j��5���3l�Bp���f�q�k荎�����w�i���oD����B�o�����o�O_G�W_����wZ-�Ҽ��;]��b���Y�^�:�>�Ͽ߻Q�#����\���x��__�7��)��=Gz���{�q$T�[��l�|������@8 u�"x��XV-�N�3�%���lvvz||�˽����l/�j+5�+��.kK��j�j�Ρ㊱h�j�H��r�Z�B�c��cӍ�*5{C�QR�VkЂTE�j��dY�exg�~�|�f���S/�^p���wM�r�Z��#�&�V�q=0o3��Fc��q
��$�-Z(Z3˦�[��b� }Zj�A�I�rq���_�>�M�|v��1��$Z!�ou}��@«y�&f3�Ʋ���q5C8�֫��i�Al�.��Þ�2<f�+,,%�Z��f�;����x̪��Ա<�ǐ�q�(��δ�ggg�t��'#��c|b�lV��%��v���;:}I��%����o�b�v�p4v�α+�	�J�@v.;{���\��?94�z�x^���4�J��VM&�/�Xh	,ߵ��'y��K3M�~���筂�ۃ`��7�X��kI�iZ������ٶ�r�,תT�1#���c������l���W[����Ӝs�\�CE�����Z�&c�k�ǭ�9�.3�-�ǟ~���T���4��������5��>����+D�1��M�������&��ݍr�*�����Qs>D�~���ӗ�$��C�p�n^+�]����B�ģ�
a$�IY2��]����l?9��x<�A����P0�XT-�V�JRM	 ���X/��P�B��B���JK���V��c��w=�yտCU��\tM �(�H�9f&.VF�hB~ӰI?o�y�Wi"�s���y�a��H~Z$)�������<�-f�ĥ kA��<.�������ӵꮂ(��¡�\Wω&P?LS�B�yԳ�5������95S��U��R�D�R���N��5LMM#�a|2�d:ðI����t�$�_|�y|I��h�i.�9�&$ְ;�U{�sX��bDԄ��t�|�m���;[(.��oظj�i+�.]��H��l�D���s$A�9�!�+Q�b4U�o2��V���K=uO�Hu�<��P6�Cf+߇G_WKX&}O�L&��l	��p#̗�M�gs$����zZzj��X���sX�c)���������u���<8���\3������5����g�c������fz�h�@���*�z{:q�]wbÆӱz�*���?���I{��z�����@�%H����h�Yv�7�=�B�LO�dx��p333����Y�o��O2>'^�z��6��Y"����$H��E��PM��[�r�Ak�<�� �"�	M�*�uL�zfs��/�[��x�^4&D}m^�Z-҄�u� �X��k�i����?6�h�m����3=&aL��w4�i���7�'&&ۂ-�i��|>�m_:�Ʈ��m��<��P��i;�mBD��rL����(�u��8���cn� P4���m/��ĉ����#�af:�u�6��Fv�f�֨'j5{�~ϳ��8�cd����$��u��ܽ{���m{�����w��?]�jkCgg'��
"AV�!�J�;:I���!����d{���e�fg�x�[\!�P��؊p�x;��Z�ʿY���LMl�W������Pڠ4%�|w�������� ;�!�5&���)f���Y��C��Aj��4JI_�cG��ָ|W���>NIJ5,�߼)�C��8y�k�d�Mk)ŠaW�PD<� ��#�jC�\��Wk�[�)��]%ٙ�z�5��J3�|G�|���ѯx�s�>f >��H�X�2�"r��9�b�E�i|�FNҳ�=V'o�x��.����K�F��MKv�M��b�S�g>���k������k������'_�_���?-�;Эz� �u��q�*�,إ����"�/`rr3"�&��u�@�I�s��1��S��I�J����C�����m|6K��`xD��E�Z���´P�t�A�B�D���H{�D���tN��n�X����f��}���gf���g���y�h�Kt/� "�~L�RQ����j�r����8~�6T���H�g����,i���Lcl�3�q����0CZ�O�Z;���^'��C������חǧ4U�j�	���x<J�WA4C�l�J��d"����ֳ6�<��o�b����G�b�R�6�}ct��x;_#��I[#>4t<�G�������믿~bpp�n�{����o��w�}%���D�Bx�E�f�rC��uwwav&'��vL��e2�Y��	����LZC�P�a8�c����}+|Nԃ@���i2�i<Gby*o�v��_���;���� Ē�%�	���pD3�05�����a�2#����HX	x��v�2C(��[X��ƞ#�f�oKܟ�x�3p�9��6z����0+�"�#e�/�����OZH�>-LX�ɜ0cx���m4Y����V�6���F1#E
�&�#��@0�ϠE0��Q%fh��K�-FtG&'����QSL���j�8��1�G�@��j4j1RI���i�OHj�`A�e���=g���L�/������5AFCaeȑ�+�K�H������Fc'��h��i��F ���v��P��5[��_k�̛��ބ�C*(�%U��iW��Wf�9���X�o��� {��+6�4�~|���JR���P�G�5.O3�~�C� �m[���=��r�9�.m��fP`���������7k3M�L4̸��<���}o?{������3���<HY-/��j|�P���a��"@�� o�Z���ڕO�V"�M�e�UEp2Cz���V�0N�n����U�N��z'2�?b�P8�Eo���MBCT���$��*";=g,ʋ0��Gǔ��1��pH
F��BDh�"�x�,eb�0jD(!�V��<6A�3^=�V�IU�1��{ h����~�TA�\���D�:M�1M�f���f m\�1�x�Ɉ��@�f�T�oM� �&IG4�����&�,��qkX�s�g���D��
R�渥�^M��S��ӛ��{����F���uRm����x�xc��qm{(�V�h�F&�A��q��1�LG���!��+�mDP��1o��h�%1�����B!�b)/���:�ce��TVvjR$G{{�TW�&���=��xBl�*��yƧ��Aꢾá�<`<�SI!5y�8Bh��d2���x���L�$�4	��-��C�y�K-���F��^��9?���c��ƚA/�b���s�O?���9?=B�U���,&�g��֨c����T }���q*�|C��7��4�j7�f*��B- cc�� -��{�K�3�Æ�?�6�h��)֜'�����g�C0��CU�C�u"��]]]��AC�pؾ3#�\N�>�?b�`Ш���ݝ���٫���a�������8��ޓ�Ɍ��{���C���(6n��իqrhT�S�� \k�>a���0��NM0D�:\b\����������cYc�n�%���?xq�A-Ʈ���2j�[����ox6��_e����C�М�G��I>�k�������H8^j���>?7�D�2.�*����B�4�Ӱ���$4F!&"	�A/O��F@��7��*�3<�.'4����u$���6�ک���-��|(�7ȟ�-R�a��R?�T��6�0�QUl�n�mČ���3$Ї�Y�*��T�}����Z	�x'1m��a�>/m�FYq��ař4��,�uarz�.q�N�1]�"�'+>�<���d�s�M�A1XS�O��p5�$Y��P��G	^�g\��M�5��֟����x���{'4�ϚZ�)����nIf ��r[ƣ
ұ���#!P��ݝ6G������ݟ�HL��F ;*֎����ۼ�+�1
�z��W�uf��F5Ķ�?��v��ӷ�����i���'%q�
�(� C�^�d�%��`
J̅ݐ�)���
������_�x��7����̘�Y��wH�s�[X��X<*ЖI ������Q����m�� ��=�I��>J���1�/���^s�5g�"�R)"BK M�+۰���0��R�&E��E���w�(�gہV\�f4@���B4�P�^���~n�[��:�G���6�m��C�%�o;軆�+��c�b����
+Bq\�QH2!�^�4��T2e���}{�R��T4K��G����(��z���0a2��E��͏PP�E�J-4?��Z��:c�_9B*Y�t[�p�Mp���r	���b�C,��i˧A��mbt:O�ff��@3����F���� ����O��XL�!x̜�H�-����h9kT� ѥbs��bV��(mDw�E[$,i1-xj�������3�\cE6�g2���'F���߿ehh�6����	d҄�"	���p�a˖-xꩧ�裏�-]�(�g�Ɓ�R������wq^��j���] �7���H���Y=�ju�`v[�����4m�;��Z9=,kndVѐ��]%���t1����=Z�c��I����h?�y�bZ�*IQ�!
(h��<�&-Gu\�����x�0*�9�='��������$q�Dᠫ�N�._ǐ�=4�MĨ��Y����g@>d���i�|��7
���	���;��_�ZI�*ө�`�5DS0�1��a(f��&td��y�%�t�o|=N�ґm�mrݨ�Y<�g���L�sp �aՐI��h�1��$V�J��e�@0`��$n�(Fص���/�+�-]A7(�Ò����T'��=�O~�Sؼ�L�^��S؜�dx��D*�42��<�N��%�0>>#��1�y�	˃4����"�,RE�f��^x��o�)fQx\�9R�좕�e"r�z;Z)���b��U�V2[L���13�^¹�~&͸B����u�M7�Z�PX�UZ��q����8F+�s��4�xD?ߛ��	�a��,�s��kHiC�^N����k�1����Dˈ	����n��`ۆ��iz�Խ��fгOC���lMª5
���șY��sn�Fv�*4� ~��l=�<���M���j����0B&�\���|�����O
����T�6$&.��2�����r���_K���'�@�--�ʊy8�<K�i��_�����4�.N��W�m4�%9��dh�n�V��Nؚ���'~��N��0ǋ�$7��]���I_W_s~bG��{����R3��K�c��/��������
[TD����kzLR��9���\��JJ�5[q	���ݭ��L�q�y��8�|ҡ�>z~x���n��I�R�����D���]�!�ʹ@vf>g`ft���6u�wHC>�Ł�H�H��p87��E3���'N��s�����sχM�-E��V*"Bk��ٝxr����e�1�߇e����C)�E*��]����F���E��i�w�~1�882���� �����$�GM�b+�Hzc��>n��=~B��V�n� ��F�j0k4�����DZ{n[ۓ�b�и��zQ7i%����?ٛ��O�����+�P��Wl}���q��q�����>N�"G�HAI�6Ļ#� ������⍓ySF4�s:L`�
Ni|&CF��Ő�]�|g�f5]֘c#�)U䣜�D͔���g���%8'F�_��u�Y�Zg	X�5K�*��::��q����c"�fu�x�2Tr����Z�/���
=��W&Ӂ����ghݺ�Ж��g���|�#�;�p��݋�G����W�{��A�TA �|� M����gf�k�H$Q��Q�k�)�|]��~�:O�
�(�Q���DU������$�@#�pV>L��"�����ؓ���61���ݷ�`��>m^p�=���؋�?�3��=ߏ	KQ��B�����JL�<���d�����L;��}�1!��㗔�������g���}��`�F�y?Eˮ��ul���y����=�&#h�Y�<F�A�'� z�*�C�=�1�X<����g3L�aɒ%81|v��e˖���AW��@m(u*I:=��avv�cccK6o܂�C#����'��a�_�ĈrH�k���dO�B6���cp�+�����S��s958����XB��
/h�Par�;�������r}��J�Gʥ��1D�j�O�$�J�������\@M�i
��dφ�#4>��\Wζ�
�5]>�ƌ���Ee8�s��:M�/�C�g,�b3Opp��n�'�1�R+4�wd���w'����GTsa��Hڄ��	��!lȧU�I�!��3~�x�]�5}��N�8��8����w�ms�w������B5Mmcy����L"�bQ�c�q�J{�mZ+��++rX00�Z�"i��t���z�r�/�fff�G���%�F9rL�𑃄���կ���������m�܌a��e�p֖3E��u�V��-o�w��=|�?����.	��I�D�0�45�Q�t2ĩ�pǚ�!�����J�c�2R.;�P^a���L�Z5�䳺�H�AЛ@�G0��܂ڝ�!N�3���jԚ��)��}�Y��7���h~f����ԜC%�C�ܶ����A+��ߕg�h��!���ǩ��|�t�]��b�x�U9�J��sz�?ݚ���s���y�	��<h�Z:w˜��<�;t�Fпk�d�ji{����N�ãY��B	�2A�A�ڮF�ua�J`�X�]]8y������$-r>��QF�V�s���z�[��i�tJP�o^/�BV�BFrA�;w������"��!�=����Utu�B�"	x���HT�~x�nYJ��1�v+WJH����%�;�s�5��:����uẖ�ĩ��y��ҒV�KM�M��W��i��&0]R��WD_��hEo�u9@ٍJ�T�Uތ>׏���~CٟL�\@�vd,��~v3��Cjl�8ʎ�OE���̉n��fW�N��Y�z>���L�p��7����u�hUй^��_��g�o�l�3Dk����*���c����qn}.���*5==}:|ScØ����݅�L�>��W����d's�T:�C��-#���{�=�)�K̀r|Cz]p�Eb+��m��n�5v�? ���5kp��1����u��z�:\y�k������ą$�{,Pހ@T�&WJ�J�D�u���\�D��pA>1Qq>��Ҳ[.QU�ɑ[��T� ���\��7�9�Oe-����(CrY�K��5��:7��	n�I��X����#B�@Ur�bM����M��{6�ϒU6<������G���!��������'���xSWnܠ���ꛃf3W�sɔ�Li_a[14�2��-$���gݑJ7�.��M2
vN�3��V쮭��qXwmK	۩��(M�1�T/	�Pp��ք�|	��$킑�?�1|��� hx�{q����g��7���=>��0��^�Q,�I���듭�E��"�v����bxǻ�-��^���}Hc��ߏ��i�"� }&ہ?Šr�hSІ7�C�q�&����b��b)_I�&U���3���{ß�_GR��b�iK��m2�����	_l�a�S����"|Hp�e�:S%�lK>>����x�\�60���^\,�ثRv��ݞ#���Ɯ��g��Y�s�Fs�s`�$��4�fL��j6���
��r{�Ze��Q�]#�u��L.ѭ�&*�9�~B��+Bvdm�v�a.��x��+�Ш+OS,�@�%�T�����`4�4M�~�`l��=w܊bvV�t<̉��L�,*��r3$d�$����v�E3B>;�'d��,� ��F��9�ozz���"�(I���nK.�#�ټH�%��I@M��l��"�1.���B�OB�/�2�;
���E�V�l_[Zx�e`<�33�b{�����^
�п��3�9���n������7J�����~<s�hٴ��q���K���q�X�����pp��D?�p�1R�Ѐ�Mb,/�
�����:��/���V��Bk�ϩ��(x���D(FЏ u��S�ǌ"-��L�
C#�t�ܺ��@���"��C���EѪ$D��8�U˖$����Y�w&�*"N�W�Ob��q���sLJ��3&|�]���������Uv{{���ѣ$��]�L�!�HFd�(6��=C$��o4;3#����KF��e���Nhk㜥�MJ
(o���sB�B�lXs[�`X�:��t��gcV:*Jͱ�Te�*��D���a�ƨ�3&d1f�槮SD��l~@����]+�\�8��K�g�tW<]�0�6!����d=m<k��^%�6��/�7S�Y���H8�@�Ag7��g/���+��:��I�jC��]E$A� NUJ�:A�^2h�hZr�0"n�V�6�`LRl*����/$�����������=��3����fI@�X�2�	��!N�T������=t�333��	�������&���)h���+���p�lFl��B>�܍�+.{Y���q���:͑*�!�����Uz��(�D�*�WI	GJ6�s�/�HR�UT�@��������
*AJA=��Zy!xf��ݳ��mF�%��l�kѭS�n! �Ū��F���[ƧOr�k L��(�̂E�0�kpI��4��;!��U=�:;��E�X�;�5�</��-zbg�pakD8���hn���t�|�.^��L�%,���t&U�����K�b畫�
�g�M)5���l'7�E�i��v]�TxF'}Ka�4���R��:�}����Ę	H�8aî������6CR�abb
Ufb�EP����}�c45��)k��ىR�Jq*�DOw����#�[`I�jQ�yp�� )��_c|�8+�5��u�U١�jL���^w����_�ݕ�8ǥ��Y��t��?u���wp<���z�u�"ټ��������K�Z�%)=��wf8�7����m)�ӕdry����RϟO#�G�=6�z3D�ᵒd�-�@�k$0E\��ż�1[L���$�M��ɀM�t
�]�O�#�ީ<���CD�1b `&7�R!(~~�-K��IFo,VU1n�`*[�Zq��ա{p��*3`"��)%���'/#���������kňΒ>q����t��2������|��z����y��4�<6n�(j��'�	���5��m�S���	�n�r����y;r;��&�Ժ�J:��y���/�㨌Mv�2��y:^�!�&T-�Il Լ���~���*"��g�R�Ѵ7I�g��Y*� ^�qԩ�"�`���f��[�2G���)q���ۘ�J5Tn0�C�������6��e��9-�Oxsr��VT�4$�D�'W*-�vnL��������@o���e�b�3nO�����EjrRփ#$�H�ۗ�L���i��d�q�vlK�%e�=�:n���`��	�H3\�����{��e$�!&؉b5ӝ4��4����ZwOO�N���[��d�%������b��T��-Q�lToL!8K%Iq�yg�B,Z<�P��מ��gw�Ӭhy:�ĩ%��V����_��w�b��jh��|���m���A�Y�KX�<�������շȝp�0����Noܥ�m ��3Zu�Z�h&��P�~-�t�?�)�B�9�tvc���6�^/#`���3i
-ԥk��N�KR���Ud��b&;����	z��%��KtnI��b��.١d�W�"���W+%�?�]̀�Uox�c�<쁫��+i ����q�e�4K���a��d�S3{p�	��t��ӡ�9�p���굫�8�=�M��z�Dj���$��X*�_"��9�*�Br*P�\��34%�,�����Ҩ�me�j/�^l}�?1k�������R�)�і7�:�Zo���y�G:I���y�Kh�&^��BLe��i�V��;�Y�A����-;��D�R]3�4_��;���cޤ5}8�j�]����b�T�;��ػ�k�ז6�A�S�D	�03S���)2�j(�|�]�b$����<K�ʢ��R�P��p�Y4�}�j��]G9K���tV��I΂�-�3�����#�N�����/ˠX��^���zUx=���.:7E�ab���G�m�)ds��$����aq}j��Z=)ŵ�eqLX��4SRX�kہ��zӝ�k���T�h0*u�\Y�����q����wq6}��1G���-�s�v�i2�_���4�K�O�6<�a;E���.�F��r��c�,.U��P� �<�Qu���W�ɐ��n�2�jS;H�'�u ��[A�5����1�{ԑ[�=0MFbc����]�[RCB�R�D,T�6�	����{�h'��� v������4�d��6-A�+�j�M�=��	��dN�<�QD�i�f�VT~[ݩ�{`)�|��%&^y�%����ĶǱ��1\r� �^��z=R��?���s�=��i"��DrU��<�֋WdB�m�&.���ԙV+�P?�TI���H|m&M0*b�Iq�Ǐ�^p�E��,�$�w�0��4_�"�?�r����̇%M�sU��|���+i
^Vf3�Xܥs;Yh2u0�K�����J��443t�1�v�[��>n+G����8ݴXK����>?��D'�'��*˫�0$M������=$���p�����q��P����%F-�%���b(d����`�H�s������e�p�La���+7151%�6�a�+�Du�t��~C�������{��w^��z#���tQ/}t���R\��{ѻ,���ؿg��#���9zP��Ϸ��sh�>�����S2T�hG8YM�o����O��|�F��ѐ��Kr.杯!�-��� �����3��8ßj<�f�c��(��js�A?o��́Ӕ���2��]�����iI�B�r�R��k��[$*���Z�-Ϟf��V�ڴ5d�׿���9@��Qsn�VO!i���)f$�p=	N�;�F\�ό�@����$
�CH�9�`���AvX(Us*`�7{!_"�@����KY�X,8�Ub�A+!���]?؃��^���1N߸�������|�#�чO||+��!Jx4^�F�DH�YuK���ͨ�ʏh�J3XWIqCuЄ,�ù�<�^M������kM��)�*e�nJ$!^CE@͠� s�
'�=_��5 s<�4��%����&���l�	u��7n~���V��2+^,�x��Ubˎ���+T��:�m����h��Y�j�at]=���6w�6=���[²_'�<�ő�b�f%�W�Ӱ��
v��3�*<��bL[u䓈��	ģ9��5���*�F�����:w��)���r��"��J�'�=��b+�g��Q`�PK�j��jt��X�2N?x�}�|F��q2�6o��M7ޏ��z>��m��ߥ������{���m��e���6�	���J��C�zQ��[������*�R���4U��61O
���@�Q/��[���VDz%�}4�@�����3K -ȣ�?4����ܗ`��?��%�Z��{s�El��E3��j�_WݬM���z��oC��γ	�{д���wh��s+k"v�ռ�D��q���s�ߓ��*Ub�R�G�=�n���`ܑ&^�. c7ًh�l�FCJn�B{� ���� [��1t�=�T�Bx��dRٕ�ؗH,P�c����\|9�_��u�A����3��#���u��O|�çcld7&�|��� z�:����s�P(���v�i��<̫&XIO�8���`z������t��ا([��!��J���Ҟ����JyA*^�0�g�>څh���;�)�D�M���< ����k*�d#Q������Um2\S�9��⹚Ik��Ʋ}mW�]��r0(���Q{ͮ�d=�2DHt�i޸�6$9��M���y^�:���v�3x#D8*j��}�n�f�ʁ����2a��Ot��1ۖ`w.3Ue�Gm�8�������V踲�v�pT�==?��]���5��%''�2dR�d`���ޡ�����eG*�BV�ޒ!F
s���ׁ��2:�ۑ�O��_��o���}dgǱp�b8�6z�A�;W�)�y^F�[2!�����E�z}rOR�v���|QM�8ҹ���$r��<��%�I�O��#�y�8-�7�z콏����.�A�������n�e�I��~{�����q/�H��g��S��T���8����D@zc�&ª@ͅ+���W�c:��̙�R��ƭ��>F��X\Өq
DAz#���[��ʷzC����jE'q��s�j�";G�t���F.�ڍ�ښ�roZ�cf$N��<�t�H
S3�R,�#B�l���0(k��_f� �=�{��+�Y�u�m��0�5�X�Ă)"�(ݣC}�IWg$��u	z�`�s�Fh�)l|���X�&1뱝����x�e"H��؁8>��귝���4ƎM�oz-�c7�Ǎ�Bg���T�����L:�f(/�!*�0[eu�Ú�)bYʝ89�檔�P4"	v��I��|TarB\8$F/C	���"��Q�O(*����D$\i��@"(O:��s9Ia0n���N�b�G��Z�(��)T�e)�f���H3������	c��x'��L���y9�����'>�$i���XuU^JvL��t_�g���4N�/��ӑ�h|���m+���{r�#�*٪K��k�MKJ&B�0���a$�]�.b�)���M�D���)�I�Di��G�!	�M��Ć	"ȵ��r�bE֕��������"ɛ��F%�õ�i"Ȝ����H|�[8�Č����|��G[�֒�w��"f�C7m�ǂ%.��O�w��])"ܧ�0�hD1�'��Pd49�;Js��u��gі�g	�qh�A,�A�<�'x�]��s��_���ތ�}�l>������89F�a|�vo��I�����h��^P#8S�C��j�F^TgD�]cd�8pe�J�/;�EհO��&)�砚�h��Mʎ2y�<'�Yd@u�~��\�%5�ڨ�$I!nE�HcZV�\���yt�L2! �������es�b�=:��&u�.I~����o���׽� B&�����B"�03�4�F�k8��#�%�U+���25����<yR��S�����6��w�mQy�`:B�$Y~�	��4�W�9��&� �`��b%�RA"�	"�NqO������a�J5'E5�T��{F��@:C��Τ�4SW1��ў��r#��%���Q�r�:ҹbrxRn�8;W�%�O���=�,4w�,_�R�ut����ⴵ�K����}]I��p&k��9��F�&'N���Rޓ��zi�*�t���.+4a�h���z3Bo��48y�D4Ɲ��Kp��W�mߦ��S�z~ǭ�;A�!N0*�����Ĕ����������4������,�c��S]�o���uf����'�s��3��t���$.�ŀ�D�5�]��� �	����z����TWB���4$�o���wr)(w�����m$���ZUސd*2�d�&8�D�L��0;3+���w�ٶL.��JRzH"&��f�9UA��l�X4���i�vwblhH��N�%>��Evz�}]򂏨���#����8��g&Ӊ��O�܎={��:Np.��KN����1�l�*���m����&%�)�ظy��>�����������7�go==�4$D�Y�c�����������Ё}� &����?�L�u�4�q�l�d15:�:i��Nn�[�v<����<��la��q����=�y֜�eb�8�� L�W��m���$�{�r$����pqp�Q|��Hu_���g�|�����x�;� D4��/2��ÊU����'n���?�Ǫ��0<9���u�!���C:�$�嚡qVh�{ӵ9k�*�����uc�������}|��:�@Dowww�X�2��t�6�b�rn��O�pjj��'��c��b�A�\�B���4B�8�͢7�M���$	"�όbf�0Nߋ����/_��V�����DEJ�j�H�2$U�(JD8J����.�d��L�������&��s��0���B�-�P�E��5�]�߆{�ǎ�@߲�������c�NH��Jsd=EZnfjZ4E�{��G�����A&Ek0[����寓��R�M���I�ep��7aۣ����5i	L���va˹���/M�/�2=;%�ϲ���[�Ç���gb˦��ȣHG������Ż��Nb�Ř�����6�g�#����}G�Ƣ��|i��:i���lî������ J�^3�Y.X$4�%(!��G��{��.��|.�H�M;i�^b�o�-FI�\��kq����Qq��k5�%���ўg��Fp8~�8V��õ�ہ�|t3��)�s�^�|�^|�C��uߺ[/ƽ?څ����x��g�@�篿Q����F�7@�[vpū�H��q<��c��/�Y\�����5+I �	�Gv��*��\B4�����,wwwW.)-Y��T�:�*��d+�|�$7���E)7��/�L�av��-#��Qz��8
�Y���R���Jvhv>��a~�#�{;r=��]:�c��₋�$��;��E�My�����|����a�wP%]�,y��/߿��q3�u���9��t�x�V.�+�fq�g?��G�����ƞ��?�\��7�S��V:vL�O`��%�8lq����<r���Adb����w�6��8�w���t�>L��z'��g�c���|�q�@J<)3�'�!�x������s'���XAa@v_ON̊�X�ظ����ı#��p�;�w����M���b�U���n��b%}�ط�W2����~T���t�:���o���ZҎ1t|^wg���/~�+8s�I����L�pز�tt�2���;q�%`݆���Γ��!P��;��>�5+������ũҝ|��{���=�UKC\��3���Ż�}�wᕗ�f�0�Fʳ�~����oD���m��[�#-�W�_Vc٪��͍���X�c��p��I�H8l�4�����\����l+���_�u���L�ܶq�ʕ��ق����~����ع��H'pښU�Jn�Ԯ�I2H�T�r	R����!��}����]���~�r=N&�"���ڷ�I��b��W"�#˂C�N�0(`wx�X3������&��B�Q�qrx��������ɑ	1��{��������D���f�6�Q��1�rf���o�.�k֭'�5�͒6��L���݂E��dc����ޜZq�V.�}�>�_������W{�K^�{��~�x�A;A���4��t���tG�*~M�u�i�. Gp��xf�i�p��nOπ��>t��r��� �S(��}a���V��$�-�lv�ر�� NdcOO��:������5�b�}#'����>�g���;�y	jr8v�֖�N�� �D�2&�]���܁͛7�"F�=�+S@Ħ{o���ا:{s0��"�Ր��7��x�{���_F����暤SW�	`ɲ~��>���������j�;��~|�_'"?�ի��s�M4�+���x�;_�];�Şg4-��w!���W"l���w'[��Ŏg�����4�����ů�����|3>�_cɢE�院�=r� :2mR]��Cø��-X�GF�[�Yo���@�9���%�X*�ŭƒ���d:��#��˕������d��s��X�t�vY�d:N�?���r#J�6�qIK�$�ȵr�r��m�?���(�.]�|)�g\��#a��a8禡^tR���|��u"G��O~�|�k�(��#pqҢE���7�A�[[������j,F�j�c��12v��83 Z!@v�f6�h��R������՝������0Wwq���8�e��cjf��~1��^%bm8z��K�!�dW?z�Z��Ix��5�,
�`-�<1�����3�16r�l���Y���fМ������3$��#�F�ܐ8�8=�U/���Ȇ(��捝	���	:�[�X�#�r�舥�(q�������/�=��a�P��eA�I"�M�ˏ�J�� !����� ?���c�N���ItwP����X�d>�q���A  �Lq���������?���>|!��͛��kށ37���W\��{�A���$�l�>�wA�*��n؄D�w������o�>"��b\��ޱ�)�1f㙥�b2���~��$I=�+��kR��w���2$)JY"���h� =;1�:q.gD;�1��B�8��g�'�~+Vwz/ڀdJ;vLp*K��I�(a�6�A��N FҶ�p���<��}�<~�	1�,A�6�;I����e�4���*�hT5'`������c�Q(�Po��wB���`箧q���0L�n'�
�yu��ɶ8N�Ģ��������8眥H`�㽶��4+dw�6����IafF&;Mp�:]#�UͶ�8��93�SO�D�P ?�;o�������°o�,\���c�,�<~W �ɉ#��cI���a�1JzΘ�v��h� � !fm#Z@���\���&!�˖���&#��X���A�4^ij2�gB���/Q�0���n�	��W�nD;Ǐ[Ĕ��=��+I��i�s��6ه���sH�O��K2�_6����_A���ec��/���O���.{+�Aҥ�%�&�,�U�V�R|�]	�������YӍj�	$���FO�a�8�N5����G^4r~�ß,$��23�h��~uC<���	�nb�v��/:$(�_�crlA��I��ս�K0IZ��C©0]ʥ�� UI�H�v���Y�t�:9#nX�v�$���[6l}���IN|��CPL:ʓv��}��8��#���=���%H8I�-ʳE��:ڻ�ZY����(�I����Y���x��M�WL��>��K~�yZ�H��БX�y��t����!�O6���a,��W/� "�@�.��+�"4f�UǦ�[į�0�a�!�]����w�H��3�[3�ޮ��ys7�L<YL��k��0+��:踳���'��-�2$�m	�E����4	��I�V����.�G�U;b�ի��G�$x8-�ͳ�IqQ3��t���&�Q'{�
!�b�,��_\���C¢�j@�ȜطdQ���8�!�7�e)�R	���%�XDh=I�^��p|#��V��m��9�D<��d�['�"�
)ձzI;~��Yt��B��~��]we�����q��::3�HPuuG@�o������������~�A�_�� 9'�xo�� ��?�h�U��h-�J�l0�����,��4�&�X!#�ZR����Y���w"���-Ӎc$�a���ea!n~�xo������'R�8�W��u��w�Ej|-F�M��D31���t}�}H���be/�	��ۿ@|��)9��T7-�������I���˪|d�D
��d|-��Z�]�8�F�W^BZ� �NT�~�D�}=��d�FL0CC�p�����05=BĴ��������p{�xHu�sLҢ�YLO5p>���xN��2'M��m���02|]��p}�(ݛl�ݎ�vc���x�y�w͑Z�
�5��^�񩝨��H���:� i�|I�^�T;���!��`t��}��W8�ɚ���$~�������?N�61�Ъ&Bg���dO�IB!,���8H�AԷ��É� �F>v����d>�$�L���U�6��J�苘�_Gϐ�cblm�(����ҽ�]iA�uX�Lc�E�"��4	�C��ׯ�[)�+_=MR�m��M����qt�� 1�/|y#���ڭ���E1��˟���t#Al�e����$)� ��������CpdT��zPFQr��n�PzҋH�,A^�b4- <;H�����~"�Ũ��f[aQ� ff9�H�=k�yd����(��1Ż���8�o?n��X�`1��<�{��78(Vn��N�hŊ��G#��.Ho�tG���_�/?�$�Rdde�qO�P̕��R-�?��w��I�	��Y���z�ۥH��.�� 3M"�
I���
λ蕒6�����1b�$6n�;w<�x?�Ug�Og�]z�iο����%���6CڭJZ���K��կ~��o��"�!C�$d���:�n2����?Ê5���UI�e��l 3F�B�����w�C_���8�!'Z'K�����$�q0G�m!6S���&�Ա"�O��%C>w\����!�^�o~ۻ��I�VM�1S��E�77�Z�amQ�`e�VK�.,";�̛���v�������8:4Ms���8F	22��8jm�mw��&mA���� O��ٳ���^b�*�O��#v�+N����H�Ƙ"�O����ĥ���^��se�X��b!����<��ɸ{V"��X����PeL�)�$�����2�1�A�)�
."�$zp��F'�D�CR��o$I��t�
"���Q'�H�H;u���CG��/ǯ��V&c�sO�zz��،��,Z���虂gـ�9a�����w�I)W=:A#-�����ob`�"UL��9�P-�t�cx�{އ�~�:�T��0M��6�W�����ʕg`2;E��&���ҙ^,[��4�,��G�JL==��ŗ^�K.�B���W�U�%�2E_2�"���챇$� ���W�W��h'M�o
�#h�!&�7�8{��Qs��W�Y�Gz�Bc�y�ϧ��_����B�-��@;��QbDv�v
�2�a��}�=�v>-�	֖_|1�>�\�6a�����`��pr��>���/@�T%�4�0�(��\�)�_�f~���$I��5i\�*�6��N�m�:~���%!y˪�NK��0i�d�.N�R�1K���$�^�xD�(q��ln�x睿��Y���\$�"�9���ޘ��3;:�,]���L�%�7�-������������}=x7,h�c;p�do~���������cC��UQ�A7OR(���ه���md�F��%_!����pp).��UD�dX�g�h�K^N��
�͒����7�����v<��c�1�I^�����sϕ���fs
��x�l�JUJ)������n��a۶mx��w���O��U�@n��hy���[6oŇ?r���6���$fݦ����$�f�h�Ę�!�T�N�<���Ex�;�-};9�6trg�ǜCdH{� 	g�]"�0Q(� f��K���[��'����~�x$��قdy�":�w9�]�Ԗ����:�2���21�9򮊩@�h�����Գ��LPbXr���K��Ȗ[�.��_�&�n��+i�86t��� i�	�Y,]���o#���(z�"�1�����{���Ύ���[r�,��`�"[j�`�'�D/�YzƔ�\p.V8��B��;v@l�
1;5�=D�k�\��=��]:���liX�j'	�nR���w� #�����W^)Ҕ7�@^P��rE�
oxÛp�W��� �8,�FF]�Ƌh ��c��&��
d3�!��Ax5O*0O�¹���א"B��=g��h�{�q�؈��-�#�Y���E3�?}�DZ��.!����Y��Pǁ����$��-�������k^�z����~@ܣ|m>�%?#?w�4�:@�>�(�U�!V�Z+�/>'��!)n��}��M8q�(A�^��#ҷh����1 ���mq��W`�GH��䚖�6��@ۡ�Dҥ	�,�1�)m�> ȅ�	Ҽ� "�f�i�����8]�Y�Ǭ��g�ǅ5N=�l3��G�@��;:�zd[��#�}�wc||��i�6m��e��i1|rBz�rw:N>�U���^:�Y�[����"v��<��'O��+.êe��Mu������Q�;p�d���=P+";=I�b�m���1>qB{q#�p�ƿ�t�H����>ch�jW��qm�L�$��؊Ik399���R����ݍǶ?�K^q��������a���?��g��Ĵ��|��8�/n�O��꣏>�����
/�U����"yA��u�cUo�L::3KD<HR��e�%�t��ja7k�$D�0h���)LΖ�12�4!�?r����1OvEZ�����C%�����dU0t�������[^�m*�iltX��I���+�T���XT^�Ό�F1�^�%HTޟ�a�%� BY�p����%(cccزq��{�� ��p��Č$���h�D����C{��N�٣�+p����$���g	��7�C�GI/�c�咮qͧ?�_��w���X�d!.��g��W^qff��UL
�V9��H퇉!7K�G?������7ѳ�fW��_�ܭ�<-";�tf���ƹ眉�=�����{�^�X�@��W7�� ��]��W�7p�Ȑ@�81t�6��^�x��q�=��k	>���~�I���p�?E�ف�ĉ�#���ߕA.;FҼ��q7n��}�w�伿���>����|����FYb�t�Ɯf�{i�#)���/�E!��l��¤�*��j.:��X�.���W� �Ds�=��d"
�׿����b���R��<�|j'���b�(WG�L��/���M� ��ߕ���3��ɇ	^��Q8Nֿx)6�}1�.�L��uB0H}u�zP���w��^��4\�����[o��^������_�^q�$��ķ��q��d%��&q'�bI����H���,9������T�4�bVr��㊤���;�/��6�ecp]����q�%��md|B4	�LÓ�N��H ���/}F�Fcd�������ٵx��*΂]�������Τ�$�Gq�U�&aS'�މ���)c��a�5=�];���?��O� �t��+��@�����5������Y��}ca�}ؽ{/�����O~�A��JI�%j�U4�����ށk>�!i�{�%	�u���4�=�<�G�ќ�� {�{�����'�N���7��w�E[�":��7"-��]����j����܏���=X�8��#]��8���<�xh9V.�����ҕ�$H�H��;��-FF�x��߀2i).Q�ˍ�A�f�~;��s�#����D�[�v��[���{+n��&LLqS1��N��m:�5;�z���6�J�X#x3N����߻�x��_�s�8[�>���\�Ti��-��0����؃�E���A�RX)SG����G�y�˱z��b�E������\�"�����ؿg7��p@���.������$�^!m"�0�g]G2GZ1Q3�IM8�Fsl���o�I��y�/� ��b0�$&��a-��o_�-��'?@"����@j��t�F���_����b�\n-DqfF�_ȍ����zЖ���܇��A҈'�ֹ��G��_��X��&ö���������I�����J���J����~#�x�����cc�`X�1�3�;;n��>��	Ff	V�2��$$�ڗ"@8���Ez�e��%8@���ӤEC�p�Y��ݞ@1[Bn�B/��,��	��'�/?�:>�����FG�K�,�5�����̞��_s*E��د�x���k��?�CG������ұ{3DCX�݇'nن(	-�����CX�h1���W�#{I(,$�\���Ȧ��]���^5!i���nU�2+�/	p�aN�����	�=Ӌ���H�-�h��O~d��Ё����;�p�����n���3���~O�x���8J8ҵ�6���
�>vz��K�4#Ud=$��� =����L���A��,��B=�II����,_v6l:���F)��w`��b�D�9)F!��3C���=^�ض��ؽ{�Hof��^eF�<���І�N�{������#ْ�i���+���� ��@��ޣ���A[Z�[�K߶���]�R�вI���c;��mI����s�씾�Sē��C�������\��&#��+W,� aXii)���h�������76��)d��lL��W���NC��z�ï9�L����ɾ��O���}_g+��%��7��%�$���rz?����tX�
�`��.S5n�a ,z�����(卶8:�ɭ�U��L�q�����y�RB��f2Ɵ$�?�z�vf�ʼ����-�#�aq��?���ށ��Ff^��6��x.�{�	,]0�h��eP� �D:aTy�ʊ|t�����p퍷c��Y8&�m<�	�޹M�����9h���'y�j*|{:{	q�PJx���T�T�Ƥ4�s	���J�9Ɏ���k�m�)�&�De*����c�h�z���c"�8�ȱ���t\PIp�Z��٨c�M�GZw��H!��$/���#$\C����Cp9K�B1:���@iqF�Z���QQϛ�<=��G��
űe�V��	��%��21���Ok��$��f��P?��l(��q)�m?�dW_��ʅ�_I�,)�0���P��C���s���.�hj~���H��ԉ*3��s�?�ˮ��gS"^P����۷��ƫUJ�y�I��?"�Y'5���0�|�6����ǟ�k���.E���B�bI]�$��F^RUcö�;�t�ͮ�1Z[c���$����q!�����%��GGQĬ�j�|���S�Qes�4�a^v1dhb��H�/�MQX-R�K�e�w�!M�8Մ����>�8�����&�B��g��"�9����~��n��Vb��_���}�q�lr��TC�5�-��!�\!�/��S^9��ؤ{$��	��H��l��^N��L=L�w���Qc9\���.��N�z!��ĬY�(+�E��S^Qh�1b�Tzh(ADC>�	�gT3�M,Z(ݪ��ȓo:+�rz0����y��<�����-��#a�߷�8���2�_VY��$̋vם�ĢE�c��S��Bf�X>�|�-[����o����TD����'oT�^�Ru���^x��E]�W�E(��^��� *U;k�g�d�����i�.O�洶�1���:<:HǶi����Z��طs7o�U�|��a�4��c�ɇ=��D.�ؔ؁��DbR��l! 3��X�ڻ�l�/ʙ�b��V�.-+ 	M"8ү�������yE(/�b�906��9Ss�2~:0ԯ��sEL�F��gK���8���z�z4�.]R���Q��N͘�n�y��p�Lڒ�������dPKε��k���w��k���e6��=:]�Y)&�|����'�-�RN��c��jJ��HS�:o�`t���JY����l���ǴB��C鎘�wVT�<��!���NF�0J��.�����A�_�V�-�m"���h����0���]�6�S��y9'��H''��`aQ?�b����}����dd/�������������]�]�o�;w���}��*r��҆%��yV�fI���y$s̟?_aЮ;�z#�ER.g� �5�Q.W>3PD+%��-�U�bxpXO-y�)��͛7��H���,~啍�U�K����+?�L�=9�('�����0@�#�k�(l��:��HΜ=s��a��&��-�&&�:� Mϩ�‟X]�\8���u+�l�����?���́��<0�dGƻP��_F�{� F,9i%B�2�A�wfG��Ձ�с��|��T eD�	�ڂ!��V�3�f`ߡ��'_*�( '�U�_�G��E&�����qrt#�1T���1�"j0��O��	ԖTj3����/6�?[�~5U�\2����Չ2	�94�B�r��4��eU����\HK�2�=%&�3%4}�:��"�+��<��d c����L���5�U�۷� #�(L9-�m~�]�4�3%&���N��aD���A��wx�b�ٌ:��=؅�]�ϲ����� �x��q;ⱌ�0�Ӎ��:��{��C�`.[����'zV!�_�eAB�����AA<^`���=����K��H&pH�H�DO�L��\ ��C#c�.��|�
a~^oa1�wt���R��� 0$DJa��uhy!���8���`%�{�ԖW�Ir7H��ꔙ�4�����	��ڽi�1��r��/�O}��c�.V���T���	O�|���>�]��qf@��dTʟ�}��Q�m�5$���c�g �5�A�A,]���:�S�A
	U�`�E��(FG�D�,��B��B�b-w���������@yu1��{ըƥ���]v������3�yF+�K�If�5�f4ј�-h72�g@w[]p �]u�.�����t�d��U��zݸ��K0g.�ڄ��3j�L&�r��J4xݥm��&U��r�)�9OT�]_���ɜ��/�ʃ�,���S��<�=�7$��E��#A�􍪶e,a��s�'|QI�IT���8Nb�3��-�W��0�o"�����J�af��8��(b��㩧��A1�2�իW��0�����h�̱~�:�b��e&���"twwb�w�2$@��xc���r�:�<�\(9@+�k�DQ[W��臸��ϡ �C���@H�rfPRQ�X<L���S׬S�3���T����]�={#|C#4�!:��3�h
ϐ�g��s/����p���{����\o��u��?��f9;_{|��~�Yр���8�<��nr,���Ui�B�H����HfzɅj*K`��u2��q��8y�y�"���|FzB�>�X�ׁ�b�����;o�o�í}��3q�g�V#���y�ȩ���<�,��b� Jj�1�|��:��*p#�$�J��k���է���׃N/�Q�h���JWae�h����c��f���!/����ť�(K��BO�-y�)h�UO0{&3Y'�T�D�RA�bf�i����4���@M�X�*�7�K�ı2L�m�nUm����G1J��k���/� F%̍y���):F�,%K'��ы�%�9�9g5l�H;��i`�9=�� �����n�%/ųϿ�;��L84�f�,Fue�	�	�E�肿U�d
#��ޑ,�a���hjjV\)?S[[�^BI���PQQA'��ݻ�uc�P(-�cc!̛ۄ�W�E}C3ľe�Ō�DQ�f�����=��z-��>�/��W_��������a��?�#�C${.\u�U��+Ǒc����B�R��W]���z��V̤�NԟekL����,�%�W"��ַ7
�38,\\���ۈB^����}�"8 ����e#�2Ҹ���b�9c��0y�.��"f��ȍ�&\�kf6�i6���"f���O{�n,����{z�\A���>��H�d���R�Շ�G��K���D8��u��P����c:�-�`��EZ���=�E�&[V9���֩�n*�{�Ԫ��5[ӺW\�l�2E6�i7��ܘH��WG󙒓پ��D�=�H���X��O+Y��W~���Ai��W�=��C4�<���@�֏�-�	�*7��S����N̚���8�6�"d��'L���_z�h�;O���q���D�V�%/�D�칁[#�NQf�u��ie�ȑ#zQ�����/�2�8���	�	3!�rj,����!l{o^{�-�ϐ��^�����L*��]��	�F�,F�^a�s�و%KV���<�����桪���1�$M�t�a�'Ɖ�s	c�P�-��3����n�g�!e@&����*����]\���K�=z�C��6"&4t�����N�VΓ"� �7���j�fi�f$��?b(�	q��qFf�k���eI�������,:� �l��9��"F��ѯ�m��2o�"d]�h����>>6��J����葉�HW�IO�6o��lj+V�����O/�>�hTJqƘ��X��Y�\Ô�yJyBv�CV nZ(Y� �L���,YgG��$�9M���E��QVZ��<ڥ�u�(�*e:?�+b����X>C?�ՙ�xx���¨b�4�xM0����%'��δdѭ��Ih������Њ�f�cb�'SQt�pZ'�V�:�F�����F����Cb*�P���fbrB��D2ݷE��d��o�.!5dy�2d$�B�F�����]$���vq��8g��I�א���
1��Cnb�Ȑ_!XYm%_w����� ]}z�t���:��
\x�e*E��!�i���e_u ���c4��HH�t�8��	ǎ���t�͘?UN3bZ�\]|��R�,.Ŝ���:1����5��K:fE�2���=V��{U����wqh�Am9��i��,f��!Ta��k���$鄢0(�K>Ӝ��x������� ����]��/��F�}�R����	�E�D�)��VWV!
��-o�HK�^{ ��ȥK�ˮ`=�r����V��Pd��3ߦ����0U5��aJ�_{���M�鞱魠�2�Ӛ�fY�hPB�ѺO�zzSC$2�ZË>�i�hg�����r�����售��2� ��\YQ��en��!�AF� �P����E�2~�K&��~U�����aG���h'��Eżİ;ۻ��y�
�����jSc�L�����
��۲�]�R�%��0���BA����C�Fj���d1۔w�;]V( Ѯ*�R��=��Ö�^EMM�ěz�r�Lθ�	?_+9��ʚ&����>�C��Hsp`����s���}�����f	!Sn��T�����?<��>�8�N;rMi]8(;�O9}.��F����(����hp\�Y�M8����~�!�x/e�籧�"�.ĝ��,.��Zfb���띒�1���͖��]�����Xx���`�ض�E<��C���~HnU_8�ڶRi���AV#�z��g��x�?V����"�M��c׎M�����~��hWY�p4��"��?��Aw7�BuôH����1�-UE���ͦ��Yqh�6ʟ�.��"�1����#A���W>��ͭ>L��hS��T:"ENĘȥ�����%B�.�^3��_ /�p4H�]:��䍑%�iQƶ�g�*he9�3���
J%ӹ:p��o�~��v�#��#�+���L���^o�zEE9#�1M{�%����4M���rQV�\yb�FH�{�`���fwK�;#�t�ʠ����QL���E[�^x�yؾ�-H6��6��8�K��G����y_o7r�����ձ�\�IGa�����F��/ۈ���(,[�aF��7"t�ǉ?��a<����	6���9�V�L�y�P>��1�;�<K�6�	�#aܧn��<O���2��(`v$w��4�u�\���^ӢB���7�K_�"�m}G��(�BY9|Q�	�q���/�=Orֆ@����3�\����5T��T�/41��Kj��� ��|�gDˑ�l�x<�*'���N�0�O8AV��8��¨�k��Z�%����T�nRϗ.�Ⲭ�����>RF`j>"C�˗.CYI)�U�T6BfH|E���w����b�~�s���M��N�;��e��t~:y�G���7	t�.��|>/ɐ4���|�+_ƽ_���K���z����s�p��uh�]gw��~�8�x�\̣GZ5*� ��K?(_/P`Ҝ9s��d:�0����>�E��*��2S�'8�aH�T����
���I2�V��Y�'���z�9�3�]qխZ�m=܆e����5z;��v���`��q�^c�6#��O�>�f*):Y�9�	G���߈��N��1v�Y�r̄#�C�u��2l��6��T��F�,�·���4>�� ������
#z���+b��~���v=
\Ez�"Y��t�X���u#���������M�Ä/� ��ߟ|��|;�2c��i�(�������IN�]��^��DlR�@��K��~�v������*��
)�M��F��]�P!�)�����ig�ڐ)�|��B8���L/>'O�1~o�9�͒���%V_���rz�i�=��.��;,�W�7.:���eF/�KԪ��z��"C2\7gR����X<����m��tQ���S�j�8��x��v����2BLj@�"e�U;�q��jQI�����!ƒ��b��]�tA�S	��իO@)�EL�>��{�+�ذ�Lť���3CĽ�8~l�:������	�R$pc��&�8���ct���5�*+f���/+l��b���6�Y	����P@e��w���#Z"��*#�!����������
\K�H��dGa�Ɋ��.�z�t�0���W^	%�V��]����f��_;Y�4��7q��W��� ۧ�̳�����햍��h�5S���|�L4x���$�J�J����dۇ1�	�ZZZ4xv3+֔�5���R
�M+\Ϊ�3n8w�@�ɮ�Jħ��Io�L ��8�/cP�}�1+���8�dAb�r~ 6!�@�9b	�鏶p<'�IJ�XoW'��H_���{�^L�}�i��P妡�th>D萤qL�&PU�q�$��t�V9W�Ф���x�6�$.Ri���&TeY��<��������{8�³���P��ё1T��a��m��\�J�����$)'���uTՐm����#��(��O3���I��!���E�@��������j��m�*J	�B��I�ЀIyQ�#i?�1�O�t�uw�����j�̷�"29���0P �d�D��ǣ!;چ�KW���H9�����1�~�����%�p�-���F	)6�Rx��a�<e��>r���v��&��*L)��J~�y�|����"Y����^-:�xfP�9��{�#'�h\�q�cCJ���`5��v�h���sY�.�2"g"2��kBg�I�s�4�̬�AH�&E94t���B&��#����--�d"��ܬtD�;���h�	]?��]�%ۆ��6+������{��	�TA�P*C��m�C�����F}C5lV�*MX�n��{�r�ujqG���n�p_�F�C^*��4������q-[�['hh�PI�3�t�J"�M�A�V�u�-�hn��}����K.$^ղe��d�7@�����Gu*���P�1[Zi*�6d���V�i�qo���5�k��qG���8�¿PZV��"wI˖�1o�"m�+�͈�H���z�f)�Kj㒱�}�$�I`�fF�}$��

<҈�pXMr�iǘN��u&Z��G"�LV9��!.�`�A#��[HZ��*u.�L�����q��c(N�91(s���[;t~YtL�dfCJ��ܴ*Q�ⵐ�>��**%,��V�DAC"���l��
֨�b�f'y���XE�A�����H����h�l�	��3#���PyZ�w����A�g���v�Ђ��,��Ѝ��n��Z��7c�.e֟p�sL;����/�8��I��˙�aP�~$G���I)l�޽h���$r'6^z��F�F�ڔV_�$�2��T̺`�Lެ�<$�!��͋%Q�M��^���Ct��8�$��GO[qaB���8���ٓa?V~���.��\��*:j-&Q:��ރ�i �8&
p�����LQ]]�'ֻv3���~�:m�k���IF���n������� O�-�˒g�!�w`ɒ5ho۫c�["�c���-*��&�ԇ�?���:Xɝ֟����OĤ��AÌ�jI"+伆(�ѭ�����L�}�L+�qoo~Q���"��{ND��k��'����suYJ�Y���E�U�*ǕW~|��t��x��UVT{��eH������A�#O;q��,_�7\s%vn{��_��h)������?&y���˼��hH�myf�F\}��x��H��2E���àfa��Eqe5f�^D�b��h�E|�*'�� ��,%�鍫�N ���OF8���$Y���9!s��z֢�k��*%{��i���PG�Y�pX��omڤX����a���2M3k�؀g��g��2�w�¼��?#>�eq��QP�Q�������),B��<z1�L��� ���x:���ATՔ�@�a�v�i�g�g��܁5u���� wf:q�p+�F:�����'�ӏ7^߬p��P��w,�[Wf5�Ж�'���[,.:�֜z��<�_O<+J�udSd�%�O�ɁX�ۅ��V=//�W��2©(�e9�1�'�kO]��?�k�튫�G��0�ݲFsT��<��Äy���0;q��7+���`���~șCMm->s������QX�yu��&%���
�pƆ�t�C:L���E&55hj��cm�ؾ�x��E^��*K����f�o�s�>K�K��$�{4����v���Am;�1Vi���ug�řl�0zr2��mt� �oժ՘�����֊Wec3�QB���(Uk֡y�VB��f�у��K�����.z��l�4��M��S�A: d�I ��bt��(�8p@�A�:�CC��ߏ�g��������������A�81�l�E�T;:��ۆ�:7�/��IB�t��j�o+f���3�b,<N:�	��A�8c)"�5�4�\��	�l����`���׌O/]��+V��o���Gn>��q=Xͯ?��'��֯2.�|;f͙�F�o��h����o��m2�j��Ԛeָ���v�Ǐ~�S45�GeUٌo~�� *@}�L|�_"�L�k��$V�U����q������@H��EB���2�w^�q]�1��v�T������Va����&��qU��(��~�h��H�Jm�,�1�y	E}�>���7/������mM.#�h�¥�䧾���2���CA%�"e/
���_��{Z00�gf��I���X�l>w�=Z���
Y�HWHw����A��g���^y{�Emu�`�Ã姜��g�ǌU�	��P��%��*a��e̦�O��rlPϑ��}��`)6n���ب�E�S2k���y�<.'|�^�Tv��ԖS]̮#�^���t�g���PB��q�s�ka@�s�
S���鎸�����A"Ų� c�0�;1�Bv���\��$�5e�hLMn�J=�'D*����T�+mJ���uu��HG��]�n��x��7�_dV�@1\t�X}�z4�Ƌ��,��n�Lh	�M�������X�v���<�s�Uʪ�k*�_�r�����rl_MH�ֺ	O?���~:�ѦNsֆs���~��á�92�����tW�ܘ\fY����䉦Nv�zKp�g� �/V�R'�oL@��8�=$��~���M�����
cْ�XN���ֿ�핑QJ�%n�� ?��|��;�N���	��1�f����ZL�IO�.\6���袒L����Cm�E�II}}5���=�G��G�M�X��Ю3���Ϙp�����s���&:���D\x�-� c��fz���,��L2���Ӏn��N!bG����"��u��,��3��Y�����IU�N2�	_�a�d*��}z��n��1���9�ä[��:�h�a��='�d˓�j�����I���BѦ�+NFc]#���X��.�He֋-Ds�ɧ3"��{�NcӒ_Cc������2�H�����X�X�ȍ�T�č�}'�9���^��5�*&N.Ifq莳�֪�jV9�(����뮻����F�|�t�M����ψU��z��55E�M"���Wj�">�s����봘h�JD.���OVX�2�%�2�g����=��c���o���H'f�3��
�Y�T0l��+%Du���^|�PE���=�"U����
=�!He3�n�d����.�̐��S� ���Jn�8�|_2C@��n��̦*�lf vW�����y���אʡ�Vk��-��5�5��Ņ^8����l�zڞ{¦�A�m`u��
1���׽�B�����B�)�BO	��u�J0��3�s-;�T=Ñ���/��]�!���Ǧ���s��a�4��,}��ӌ1��E+:�:UN��d�VD�C���^M,��8
	�$�������H!N��d�����H�p���h).0̛�5����9/zQ)�%�z#�����E,,mu���OӘ��0�%��ȃ�4DQHdd�A�(��I�U���P��Q�+���:�U��K�김��D3f4h$����~�h�H_<�;Ǵ��W�(�UR�%<�׋$(�(�4�����イ޴ a�l}��uFF��*�*9)N$��C�Yi����M��!I�r����߫��wﾩ�4F��ݰ#�Iz�e�����ݻW��d�s�9�Qѥ��rS�y��P���)Q�~����;�?4�x�5�a��T�x{����5y�"�Α���f��~�.�i�*آE���[���x��!mt��VL�%y����f��Ν[p`�6���'Ƹf��X�hf6��Ѯ>D��E6פ�A�c��MZh=�o���9D����`��'㺛nc���fO�ӗ�\�U�Y'�|`��d��������i�d�4���C������#:�3�5�W^}��z:/b��oI7�W�%9K���<^����s�G�VS+�jQ~��������7�\fm5f6. ?�bl<��HF�T�P�(���&�سm��A:�+W�������EK��4���Y�*C�̗et!:@��,�b�ۛ��2�,ItFinX�j!�r���!�
�{ڏc�ܙ�����B��ב���<��2r�U8��#���U�}Pr�������n�\�'?y^z�_|��-����q2o�i��%�0B1�Q�h,X���^�~p��;����#����q�=w㢋/�e�GdC��,�����Ƿ���G�n�q�-Z�y�7�ag�[���*OHV�$;-Vi[/P�������*\��T�Y�G�����i\w��򗾉ޞAԊD��m���r�e�֏~�Q�%z��	:�9�7^}���)�74����CZ��F�Y:��_�=�w�x%ńIQ?av����?������<���Q���T〈E�r��-G9�YQ(I�"��z��൑�]���J�uA����Gk�KF�����&��&�������7���m7߄Y��˗,g�GBW����0��BW�����߇'��("$A�E�����ݽ{���Wp�uw2K� ~;F���� �xH���
,h;���[�x�T��hy����ᚫo�g>�9��8�������5��Y��7��Sh�صk�}lݺ��:�����[u���L"���C:և��vo�+��7b����oJ�c�Nmo�Ѹ�o��äs�\o������o��>�����([�:�;����9?����ddTj�"_�}�n��_�yh䓌���y�4���s,8��s��-�qG��V����w��������(���W�g}])����w���~�z��L-k�Ԯ���z�)��ODeY��l���Lve��Yn<�K����s/��!�R,1�v�n��f~N���A3l��S�-��/��yP�Rm����R���3O��w^Cy�[O�k�*tN���4�^O���_⊫o`��?)L�M?x�,�S�u�9D�G�qI�\���Jv�L!��r�ş�'����&����l���3���M)+c�c��ϓx�ه���_�=[�KҨfDn&�={_��@s�'-_�l`DA~ZIn8�Ǧ�~���.��YT%�I|hw���:��G��(t'�k11مy�e�0VF� �ÏH�����08*C5�Y���t�����啛��ݥ���ݽJ�e�^~NNBO[{zV�El���6?�$�z���;�5$"2֙Aue���`�w��~�x�g�)�A8�9���v;��s�b۶��o �fT4O�NQQV���~������oR�y�H�?!�S�삦I-^nd%����(��/��"N=s=R�����r�݂7�}�]��<W���$��ω�y:��a�޹�VgU,��_vɕ�U�i�&�Ty��p2�,jP���x�y�W8��t���x�M���Ζ����tn5�|>�Y�C�͡p�� B�\��i֬?��΢�[v�^bv��sG�%�m6|jtv������2�a�(j�+����3�&+a�Mi0��� ��p9�U]Z�1�\�{��Z�&@���Ԛ�%~�4e���>�,C��Н����&���/��_�#�_�Ab;�ӊ�:��pKW�� ���}�0wV9�}�Ta���삐�L"�j�A�����{PH��u��.��S[�2��{�6]r�ZI޼�49A?^c����΃Ő�I�g'Tq���s���W^'hЋ1w�f���o�@k[�����ghz�ZuGW+�鈁�n�b]�!�K�q�"ě2���Qr$�x��+�c �{�3���h�B�#l��F !BL���)��
*7�|�q\u�ZM/�u��Zu8H���9U��D^g�1�s'�Gq�����B}}�rq�q�ڷ�zS���� ?_�{U���"�#�t��?����H�x�^_HC7���?��<̣�x���*�I�S{{?��&B�#m]�`#vI�(|��A�qh�n,\Ѐ����Ԉ��������rOj�F�hm9�5k70"5j[�&U�����j=��|f��= 3��k�/��+Tl;܂�O�@�ͤ�-an�r��]q��߆��\A��dY93pzJ�E�r:��0��?z�l�8�B������"�HI�i\��ecJ�X����ũ&!Mb�o1^y�Q��)I��]i:��#J�%���&�!���/ҥ���R?�;+#���eD2��E;��¹%X���x�OO��ͯ�K�F��.U��U��N�p�|,��i\�H9�b[�n��DO>�\x�������j�cv0�Tp6��C�%F�xZ�q>q�?��$6�{�
�����_��0�x�5�!Ҿm�ꠔ�͎�NM�$���0�|�1f�[�~'��Ɲ��K�#�
3�x�h��F^��$3J��.h�]��ɨ���Z?�^�I��2�j8u�V��;s���	�3���Z��BI��;��LU�QZ&������'!�Ǫ`�Q#r�m������'iF�3��>��zD���N?�s
�$!�R�j�؃?0�25� 2�#�~�Q-'9-(,���m���0�&ym��<(�exhH��������"�~-ۖ�̤�#@ W��lI�S<�<�y�V��?o���}�u�h�vttثjj�b�G		���{i,����aM�2�a�w8p�u���&�����M�N�#,�%v�%j��蠌�=�"SD�
����Q�2e5���$+#�B[��$��r���"���P�Vit '�i�Hxݝq�a�;�QH�<�+�9��hK���}�������v=��KU��ȏ��v+����!|��L�a���U�xR6ӧu��@�Szq�G���M08)���	FHh�tR��P� ���qm���ޔ�a���ӤSܠ����#Y�a�|�nv0�1.�e�1B��"�TZY���'E��3�7
i,cpe�q��zj޼yZZ�6�pX�q���4։�nq�3{�-v=yA0Q�;��:bp"����@�4I���
�l���fr\
i^���Q���B��a:FIU�v�� ������tH{Qje�ij_��rey$�F/�-�[����Л<�t_�j�zG�ۖ���#9_4�Ngb�H�Į۶�];iH�d"*��4c�.���K�B��<��碄���c����$f���V��N�%���	��B^<9��JGc�b�|NzzN.q�)Т7C��1F:F`q��@,&��y�s2#��pQ~"���,���Mc��猡�ح�lv2Z�O&�fJvx��f�p�J�~*G�Fi�v�^����'c�I�.)�j����:�����|J5Iz�t!:�pȇ��B�3���|τFr8y�'���/?#��4�X��(�,��Oh�``����a�\��9V�.:g#J;z�[�t9u�:�&m/f���穱�{��$��Y�TF���Ǉz��t��(�2GDf��I���ty�����e��|�
�c�*�|�ںF�s�
�zh��|�v$yu#48��H#�k��%��҅�m*�3��Ѐe���������Fy��P[/���qHԇ�t��s�Ĝy���U�Ř=Q���	a����zЖm:�<��t�B%�:.s�X�p�����=���I��{�e�d
��&� ��q��l9����G�����2WAjs��瓿�S���;����_�^s5R�v��&i�f;�ب{�Qoт��ػ�Ma�$�r��ԁ�-��� S��@mĪS�����ʊ�p��g��?��v����n�b�<U��%�zJ,;*�h�b�i��c�������98��]m�5��0�Ȗ����b�!��.'o�[U�Z��,������$����8�c�ò8X�r��'i���� �L*L8�u8z���uA�D�8	��>��"w1���_p���0�XO�eH��P+�	�c�_����;��a�\*9N��ߓ�����nĜ9�e�I�I�<�,_�p>V�X�-ｫ�
�u�B��,8<4�U+W�?�	"��v	����Á����}��p�?��m�"��NB�����u���7�!?�3��8!O�`j�����㷿���L9��7��^�NET�c�^��$墄g�E�2{�'Cb9�lg2f��r�$;��=}�r�L��džDB<'��U1�?�d,RRZ����a���F����ĀZF��GZ�n."R]t9��h�0�N��u���=>zsiR"�a�`!_��r4��דډ�J��Ã���fd�q�2f��)9���8F!CiJ��p�ɀ+��!�>i���LJ]U8yi���kw��i���19N��*��uX�t�.B��牌ic
���v+g��"2�'�-���>4̞�sϿ����~uu�n�Iq�M������������$���k֬�}��������"�p�F#1`����k�BoO�E.=��#��>�3y��zG��<��S���1�
���³�2j�Ta����h�9�_{֟}>�%!��bXhf�h�a��A��݋���b��AU�Xr����>�9>=0t�=
/�HJ+k��`���+n��ｅ�-�>)����Y8�|�!h2c�sf�(^�i}�l���8��eF	�P�!�����̊�s�Ÿ�3�UH�͠!]EZ���Nx&�_2�HK�W�!Д�Tw�^�Eތ��&Ԇ�V�����?\~l�>6�ϗ������������8�a�����M�ߊא��UXVv����Qמyz����^^�F�<Ѓ#�:@]�b�:�������F��^����V{1����d�o	&��+��+��j��h�3��ҧ��EZ���3�Ì<�8���p����Z��-hDU�2仪��˴4�$ͷ�u�)�ErgGyuz�0!P��&1�E�Ǚ.ìً���t|Q�$Iר@
��l��1m���_��
�qg�~��M����/<�����Q��7^t5�Z{_�GZ�j{H]c��ˑ��۴�t2k�U���ilr ���T鮣c�@ӬE:s�HWc�̙�L}��(	hvyHEy�������o��t���"�ᔈ�	�ommSX'�b`R�ҁ�~��aw⪫o��W\�`5?�s�-����K���Ȼ$���3�uuu���M?���w�����W�[�K	4K���#�mk L���Y9��eN�E{��^�wJ��yA6#�r��r��������UQiX0�vP:]6Xm&l߾F�ٳ��w܁��)M�a�E��/ة/��-;�L�
���s�N:�"���G��'¤0�!~͊�D��R��b�(,m a�8��:/N;�Q,Ǣm̢�c6@O����	K~��R�s/?�xz���~�����.LD@ȓ tqj�ns��`n:�ik/����c���:iVRT�Rw����3$��|�4/~�i[�#~?�
�_w���j%��u9������e���HYlR���F<$N�S�s�ԛ���"-G
.��bY�d��K&��,����]]�	�	�n݃�0�s�����L[6��J�k�J>e��x�ꌖ0��0��DH�h�̞�Q����\u�ā�ʳS�R�`#pV�9[���@H��?�:�@ʙ��d"�Е`%n�����*'��D(,]��r$"2�&�.�2�)=Z��i�x�ƛ4����TKv��7�:,WGpuf]�1+�f��Rf���Z�`h����ɋn�%�\���Pޔ�ٻ�)��������� ���7�u��$jfӠ���FȜ���r���S.��X.)�����O�&ٕ�� ���E��U��v��b&��^����� �f��i�t��V͢�Ԙ��!f<&;rI�mv#��#}#�$�.�f{I��p��:j���@1��^)\�ح9:X�s'�	����Ց��RE�E�a]2.*d�j�<��7oR��պ��ˮ�i�qh$��yj9�z��D���@?~z��u�{>��6/��"W������LN��[�����R����Cޏ�K�>k�z]כJ��}��+*�٤2'�6!��/��gx�՗QL�(ZOs��&t���,���b��Q���P��D���߰m�l{�nD�չMsএߦjv�x]��t�E�uE@iI9�NY5�X�J��Z�9z6e�:e��3C�D&�>L�������L�����T)��Lؿ�Ya�^d�
,� Өֺ�l�g�{x���x��X��I/�u$+W��Hl�*;�RJj��\@'1�cK��h;��o��狨J\(@ss3.��:��\�FiE^�\�>��)�7ӱX=��c��8��V9��f�[��Fr2�D��~:���١0&�"�AR�
b��]h��6�>�i����^u3����6���\L��PB��1��QQ[�w��{�=�;�����D�s�=�:!�Dr�8T[�Q^�����ڬ��{r}�~�<����=��2�7��*�2�,q���	�$�a���F��?�$��N|�_�e(�$�#%7\:eX�?�1}�Q��r��O��?�)~��س;+�,�5r�,�"�UU!j�����˵A���Q��2*:܏o|��8e���7�Cl��)ϬM���Z�{r�	<�ģx���Q�u���H˝�����WH���ڷQ?��}����[2�$x�E�)�Sj�G���%��?H�AG�&�z��U4���������u��l�2g[|á S��D������n�<�A��Aw�#���ԓ���ʗ�o;/�o���ߍ����O\�M`ɴ�W�Fg�Q�����_=�ǟ�;��+�bP\��z�R2�!<��s605���ՋH.͌fG�z| ����q�����E���՗q�^�|�L�xq��p�ބ<�8�yV�_�3ϿR7��u�]OO�BUE3J��+7�={���t�*_S���#;v��-��¨�I�z��j�r$[����?�c�m�L�x�l��x\8t�_��K��7��M��ߐ���|E~w�`fc�J�H�V�&�|�y3k��RZV�4�=�$�EP&��q5|�Mڒn�f1���!\IC����uA���hKF��ٟ��#b�	=9�z��ʬ�&�ж�?��	,Y�����,I8"�(�����x�0�B�/*v�^/��IT���~�k|�;?�}da�H��S�)=d̢���lD��۸M9ٲ�l�@��0���ߗ��bѴ,��H� �����\��T嫂��ϤQ�����.�p��?Vh��t�Z���7�W�����&����9��O��Ǟ�Ƭ����z��ϳ5��N���]x���o�2fw�q5 �æ�����ڲ+:;r�R�1�(j{�v�w�Nw��y�^㌬aUKK��$��x����M$��`��5��.2����t�<�C626�7u<bF�M��x�O����/��U���1��M ��>��Y�xYVQmj������\�5�
��3�sR����mێ��G�br�h�jUU��A���jk����5�}΂�[Z�ꮱ'{g�ߠ�1Ȍ$e҆�ܳϫCI&s��W�Lj_��r{
�ض}�Y7a���ҳ�r�9�xc3�v�6�O4PJ#N��D��x��gp�E�{=jlA�����=+�F�i&�xV�_���U�8�v���ìyU�U� ;!���)���א-�f�ӆ?%���l���S�_ӎ1�k�Jgr�w#�����r�L�@?�`3������?��9��SQ6����%�����o�M�
��MC�DOᤓNGEM�F���UQ]���z��:��w���2�}�E�e�z�z��֒��ʲ�u��^�䓏�ws��tyv���������x]�x�鿩���7^GMm	V.�ˎ�6?��Gmu��
�CϷq�7~��J�6��YaM}}���VT3�b<2��"F�!K�"̌BX����Mn?ގ�_~Yኴ#�a�<��9su�v�g��H��ug��C#|��T�C��́��֣�t`�n����!G�d��J��� >���u[��{�-�F$p����Ps��d\L��z���~���&\��cڡ)U"1!ƒŴuyr\��Duܱ[Mhll������N'>B�ə�[�B8�AQ3����	:	3�!c&!���4k���ڙͺ�g:r'%p��#����I���"�Y4� �{>�3�I����e��'n�#C{�fg��O�Ta���{�q�?c-2�v��S�E�ͥz�Q60�$1����p��e��c�r'�h��Dyy��B�P�n;�wc��9���!�a�&��۷��֪!�WK	o�7��_�0V:�(�x�Ǧ7Aڌ��QP^�'Żv�EQq6��H.���Q^�U�3I�e+�~[/�"�3��������q;�x����|��"���p�W �RR
��y�0���*q����n��§�V�w�yK�>�J��ɢA�vGv4Qn���<d���J�U�&=���x_*L2�,��dV* �n����	���~�|�:���;���T�H��dǒ��)gӈ+��r� PJ����H�' �����$���&�e�Ӑ�"̬\ZR�+��^��S?(��3�%�	�QMt9�����ڽ:�$-�-�Fcvِ�֪R2��-M�1zp��-��;�830��pM����q�GryT�W�z�-}"i�m�9C���@��cGT[_$XD�jtx 3ʲjČ��v}~�^{��J��?9�(V��㝽8�rT'��BBM68\&f� o�}*�0��,7-g*��1Ih��=oQ!�	+�I�W���AR��n����qȒ�*:(o`�Bܧ"a�}+bc��Y�� y�U5��iږ�ko��I��=�����{���A�R�j��bR�F?��%O�]��E����Vo�!����?/?�r�j�9��T/.d�X�D�[8���L��HD��"	b��.��+V��3�x�DO�Dw9�l���a��'�D��C?!��jh�� �Q�-Q�K��"��g6�"�kB�3���Y�Q�~�M���̘5{wo!��sB/o�����1#7�ys���s��ժa8�qjׁ8@:����F��).��3�8r�ȧN��݁j���OC���_�u�P�������[{��,�R�0�S`�ڵğO����ܮ=ⓡQ]"�1;!�a�BCc��Ki-F�,�=��%�>���V�D8*��eF{� on���H�{���CJ���ܢ4�93g5���L **$��Ew�}��b"��ܤ#���l^�.����������aIf�� ��4�:q��m��'���ጵ'���8B�l_M(Ǣ�k���714:��"O#]�2^8��`֔f6�B��!'�rͤ�A���D{q� �p'?���@l�V���W1�\s�UZ�9D"�o2W�)�J�wuw��|�ޯ�3���d��ܧC�;�<��j�Җ  }FRM��I���={�:�\kY����CX<_����/~����Y~��Bk�A��hЙ��9��ݤ�T��FG�-.��/��?�����
�D�� ��P
��Y�`���h��R)ɾ���M�(6Jg��/�R!v�'����?���S6����B������p�ͷ<�m۶n��,PEQ���x饗�RN������$�}���%�Ξ�e˗dS�x�)~��'����?��������4ZXT�}E��HΧ1o�|UE`ԑGE1x�Q���t�� 
LL�l�A��rLy�麛U� 7'��oJ�kPY��с���i��%$�MZ�FM��]�3�ȦM���8�z4�-\����n��'?P5�P4�¾Rm�,�%K7nܨeS�Tt�Vi�޾sǉ�r�)�l�n��̘1C����~`1H٥�~�z=x��n��,ߗ�p$ϲ�_��V��5%��sNGAY��a����?��aͮY��b<g�}6��V�"V�"�	����yș$࿭��;�H�3�D���D��"�\{.���)�S2r;���n�h��I'��ǟ|T�t��ƞGB����4�7c��s�X0��6�Y��:�{'
#���Fu �kV>����-��"`��X|`����S��ó����͛7�+�#����\���jo�������1�� #;�bPŷ�3f�������Bڝ6F�*��H{��3��O����Q#F�j��x{��F���p�ɫ�����8��b�\,X��y�_��+��31<�Ǜ�A��>��4���/� ��XM�#��G���+��"��p6����o�ͫ��b�6��2��D�)TW�����������eE���l4���y7�4X�O���{��耍���.m�W]q�
�n}�߁E��\s�Z��|4\��2�A[��1#.��F��oڴI��d%.��VkdZd%�O��EAQ��Z_r�%Ȟ|�)%���3p�g�Sw}��6}6
�#�/�g�:!���^z-�`۶wa���9g��@��ٽ�FO^��)mV[��)�SO?1bz�R��4��v;E��*l�p�jI�g5�s �f��Rz�HA@`���u�y���@�/�>3����1=��AG��!��9��Y��6QM�H,�u�Zn��I�U�^}:��z�$,���X��u�b�p��P�,�h&zDzKyE�z�}��1��ؓ��� �@���n�g�;��L#��uS}�0Ad@��D��]w}�g�#��ȐGC�� �1w�r\p����}��#�~�{SUY�� �=w%��"l{�u�6B��n��uX�&~��W�X�\NIf:�u�ܼ~������7������$o���n�L �M����6������O}J���۟��wgo�h��C&Ru��-�UʘaD��ݎO��)5N�~���z5!�ݔ�
�z�"��9|n�r_$+l`��L!� �.�]p��i����e%�3mQ(*�v&q���s�?�c�2m'ﻫ��o�+�K���P	��!�<����睿�����H��i��'Բ��vѮ��w��$�D�������-��Sd�`�Ȩ�<=�&��͚әq��ZUʶc4h����_��`L��Z���z�� e���VfGC�X��T�~���I�)ӓ`9�������%2�!��I��$�v*���o��P@��=$��s�!^���T��:PY#�]R�-ߦ3Q=��c���7ߊ��.M�Uu3Ո��<������C(.t�����׭���G�w�IVVۮ
]]]��:�4ݓs �(ATD��"�>*z�WT��^�  %���LN�s�����뭽O��^�I��Ǆ�:�����^;��V�J44/�g�=�D��4����̦��ʍa��Q��3�J�8���/���+����\۶y�t`^����K�c�h'_"9����m�\M���������#�js!��6^|a,N�����=τ�}1b��B@G�����_�~�c��\XG4e{���n�PDa��8d���i��09���:���2t�g�z�5�������Mx�H��޳{;�{J[��*�BN��J�`�w����r����"��i�z�?�c��z�)�N
˖���3�YT�mƑZ�0U��5K`�aR,_�v��v�����Og5��#���h�V�}��g��M:�W��}R���M�ޑ�\ӳI����n�ŷ����t��7�Q��3z��h�Yd�9�LL"����w��K"@26���V�W����1���XԥJ�c�J$q�5No�\t�>%Y��{��г��s;���V�=m_ԍr:��܃���,jH:��8ǣ�T�!˜�����ġ}�	4�_�1o�ǫe�v�!	iw2!�թB�@��\u�N8���R����/3='�Y7 K�jJˠ�t�>�\~�庢J�F���{��4�u3���s.y�ź���L#���{�B�	O��I�IW(��Ɣ	|KC3��<����կ�<G*F��.<�|\z�e��	�u{=ᲨhK���?��`(r?e���dnŋO_u-N;�|UIϕ�T�RJ��5H�6T_^z�Y�{��x�-z��C�v�Y5��׾qz���f�T�%u)oc~c�r}M�@���a\��w��h4��oC������(�UUi5aǮ=�3#�z��U�q�d
����P�\�[�NZ6NF�����=���v5�L!�#�XJ�o�%]��K�C��(aK��/+es:��\���蠶[���e��Շ�ԒyV2�|�?>��=K	o<���1�t.Z��Y[���0�|}~�Ûb����uM�X�|9֮?
'�p.	Z�z�O[P�c�ӰM��p/F_Epl��8��C8V�Ѡ��hn�BcS��!��&E�A絴h)��[��^�^���[~IXi!��_���qp�A�H��L���av��K�Qn`}Y#����n�}�߫r/:C��j�I���ˉ_��k|��o��:�vu���m ��#���\�/�ˆp��Fz�{�1�����ǖ����J__�1�%n��v<��꠲'M�[dd>�����ŏp�o���FB�r-��~������?î�{��/}�3q�.;�&8�AN�����15xK��	�͘&�n�c���՟�7}�'h%�6k��F��[�A�iK�P$x;i^��b޶K&���?GH��E�G��M���-[�
I�T�r�u�����
�B�56>��<���7?�7,�h�����ꈞp�ػo7���~/�f�~��	��Z�A�U�'�-ajl����?a����X�N(�Ui�#	�w��?Xܵ���������n���[_}_���E+Ioc��XZ6��x�al~�>db	�{�u�"����.WR&sԓ��*�3�(�C�O��!%��c[����އ�wvv�@��P�8q��7��_���lA"�@-�V:~�ӟ3�e�ɏ�h*O'�+����
�l�0錎wJ�N�D��Q�������M�}� JD��
�t}υҶ��A��2�"�T�ٓO>Yy���l�����q�t�XSS�� ����V�j��_�*��n=Qn U	GG����.�GBN��<��b�uͨtW��m[��c�`��'�RyM�"FL�������@/���r+h@`�,g��ud�W��)n���tH~~�F�g�]kf���R�W[�	7���C#��g�%/?أ�̢����t���'I�͒��7_�-8'�t*����ox/�ڪ���v��&����ĥ2xn�#8�U�{v����n��A��#J*�����1>�,2$o%���x��%	���̧��_�{T��F���0>r�}�ϱby;Ȉ6x�����_����ah��"�_������I��fb��8Z#*}Uڣo�Órg��r/
3n��q���H�j*Y������cd}��Dr2�^=�ǅ��i��g�8��l��ͭ���t]R�é�@yȹ|RZ��s���h�Sj�3�Y�[3����a-yz<�{u���c��5�6J��!t���?����)�j�2K-��w�u��U�f�X.G^��B�(
&fw9�xa�sX�v�!�BÓ(�<�����v�r�0h/�uɼ�t�z�MD�����S��t(��zyf�t҂�|H��$��r$��4a�>�6��r4≱ADK��W��r�.>���r遪pb	N�Bf^J�t>ʬ���, 	�b��wAz��Gr%ā|���),�
�epNg�H��{��*���L`zb�V-%޶�׶c��ON�H� -�m�R����k�V�P�]o���R[��nG�XJ�O~�n&\����03�����I�}�ȥ�L�fu=��xG�l�"T�|(���,�4;��6?�74��a��)	�"�&gTdJ�Dc�!um�|�A%��*?ڃm$,꠸h��.��{uH\�H�%*�si�u˳��9l}�U�w�9*��E�(1mJ,+��\J�ɬ�2U����d�_��8Ú5k�����y&���~Z�		g���1�浍Z �~AY¾>'�2|��}��{��1��*]HX��Y�:$��n�:t� �9��$�
�V�׻�Ƚ����k=�@��)J�3�Q��R2���B�X�%K���3j�쒬W�� $P��f�Ɩv��r�"� p1�)�W~L�+s�U4��*Elo'���������̴�>!Z�w��
�|�r����yxf��7����L3<�nT:�01�G����9��O�`6)SY�VL���?�uG���W��LJ�g�f�����I;�03|��u����;�q�4�>�]w,�)���ͥ�C9ٯ���	Է��!lۘN,���b&���$�JR��B�U��n��g�"���,;�IȉA����&��Ҽ����L=�$���編`���C�!��N����et��7��v����"6�Axn���D�C�k�F�ee�<�ݼA��g��t�9���m�+Vuaˋ��iu�'U/�k#]:%J2X�L>9>��^�D)9a��L/�q\��תl�N��s\����@�\S?���C��)F0$|��!���*�E?���Ja�ӏ��V��m!g�x0���Ҟe#�*�(3**�ƛt.?9X��U8}�{$2�q�*n:ߟ%2?z2/�@��|��`T�*�������<�6/8�;���?��%y��rs%���8���J�����i~D�����"���� )�	��ٰJK�� -�)F]�Q�UE��X�zuy��� �,nf�~7^{s/Rѐ�^ĈI%���D	�����9�3m�0Fx��w`���:����_k9ȩ-��\^��L�)�������f�Y_�W���=��F�єFg���c��'U�t�:�2���}*�F4���!o�C��.2C�S�u�r��hyxe��&Aq���"����T����|&L�(���"����M����3������@���+��Jص��]�S24#��4��;��� I6)2O4f�P	aH'Ss"�#P��ԎU� �O2���c�B���E�B1��K������A,Y�VK�R�=UmC�A/�Y��7K�����9Ec)�.����eG�W��.j����́IE������e'�=H�R�a��?O��r�|Q*Mo�	^���K�@��6diT��rm�a�b<B��F��,�&��!��V��rW�����x~ۙ��}*�"�9�	�����3ڤ�b�-���""�v�t?X P�fF�t.�xZ�\�t����|�"�B�^[c��aD$.���zFё��nOBsqTU{�W0�ut.g�zA���sq��F�K.��O�gu7�fhi�E:�0 ��y\��q��$��bQO�+�
zB��Qf�E�������i�jh�Í_�:��� ���C���?��|���Я�@eҴW��8c2��IǞ�3�<#3�!��KYZ7���lB!W�B���w�ӄ\�r��	�͢�����W����v����S|�ir�F�g�lQ���#NЌ`�ѷ4�����n�����-����Ui�D/��@um=z{G�)���'>��SSr�Y�٦�{1�����~	l%�5F�����?;2F�Qf��g����>��hN�~�y��c9c�e�j�Z*�4����-�*���Sg��韎,��#��T��&T�X����r�|�QǠ���˖h�T:'Ńe�N�שk��~&&G�K��L�"[*�ڵG�[,��<�XH�gs�H��o�+ZNtJ�Yl%�^���t�E�^�D��e��h�Zں:��+>J��38�$�����'U�I�a���u�tVoZM|��G>�肓�/��B��e&�o:�쳱�#v�lop��rUtHɐ���=�9���Ç0��7�����E]����$�I/���M$�������h�B�(��Q�ུ�+d�c$���a-���hRN\e�ˬ�vlt�Po
N�U3t�U�As�V/	umg'V,وh0ol�t�#�fp�g�	�a۶�(�Q3�$���$5�Ё<X�d��oH+�`r9���
�YԹ+WnT��^�D4'��}h�\���D%#[4�@�pV�IdXK��W�Y�G�zK�vcd�#���Ho�Ϯ�x$!�f�ǧ[t�y��B�[E)\�P(�9X8S��Q�y����XB}GG(+��0Eֆ�ݻ�l�`�ZM
)�j�I�na%3��L{.&���O�q�AϒF�ɿr����U-hj�!��"B���!#k�fcsI����!89���0z�`�����Y
]1�4l%C�3�Mh�i����G<���6�Iډ�,�;�с�c��zZ-��r�#�"v���AF�jTF�̚��yQU�A��գ�z)��j�>�k�y�Ỷ�4#�9a!���ᇞ���q�ZY`��#�4b9j[jTN'�!:_�_�|`o�N�{`�q�9dsV�m���W��è<��@>�%�.��,V�|��uh���)�բ��5t��\�D��&~m"�މ���,b�dfݳ��صMK֖�#�J��	T6��S�#!�±���WU���	ttu�3W]��O=�������C�Ʋ�+�Yy���EmC�{g�͛��q�>r�e8��#���c��:u���`ͪը�o֒ym��X�[(��d}��yi��4�YM�����2ʧ�ڹj6�[���B�pA�Y�U@H�t#F�AmҘ&	޸n��M����ػk/�8�L��zF��go��А��C�0�|���v^�!eR�'��2"������FzY2;3�����o-Z��yk�vñ�O�@T����'$�d�R�ku������To'�N��UC#�{�`�G�F8T���	�e��AIz`Kenb��h�uܯr2�d9��pW�jb4읧�"�s&x��eFSc'>���}��W��j�j�bm�)s鮕�Q'�������JeX��x�\����н`Vk����(
gFE�Z���f��T(���5�T/A���%Ǒv���e
+���2�G� ��ʴSV�S�h���{�ٶ�]Gj�V���I�����<�kwvR$�S>��?H��W�4���Q�E�@�dǃ���WQ�#ԓ黁�^���L�\s�L��~�ʏk?���Z�ɪ�b9B��1/1�2��Rϖ�x��w���Ӆ.Tm�0�5��NE�wt�p8b������\t�E�b!M�X���ZI`��fnvz�4ԅI���Q�V�\�+�1��t�S��J*�H�����:�_D6�3�K�Ih&�s-m+�t�&{�z�'���5E�l�a����f4�ifH�n	[X�s�t�#�=9�L����d(��;'����%�VfT/m�äP0�r�\8��ƕ|�e�9�|��%��5P���s�<1:
	��A�ٞ���8�jF�M�֖r����JDu�M�C��H�8��@a��1�i<#g\�Ý:�P��Q����I։2�c2<�hJNS��3X	w�Ji�yd
P~�T��}���PF2OD�紋)�ɩ�ͭ$�M���B��9��c��)� |m�iȌ���f�x��Am�۾��|#�9��6۵���A'�mE2���ֽ��׮]��?��j+̉'�e˖����	D�/M
�,��]����:���?5�R�B��ؑ���w�z:N[���%dya6៝*�KG ��b��pD�$�^&J�BRd���ؘF����
+�H�2s��Ĵ�("�(Z���SQ�p>�,��E�@���oO��,�� ֓s�ٽ�:f�9��,���QX��IӘ�B��i��݃��R=ď�-�kDeM��4
�Hr�-�6��C���ߩ�c���߃Gy Ys
����T������rL�B�l�D��d:F�!�L���9�dz�$?I�17"�� �1�!"a��XА+U��D���[t =eP(�H�GQ[����,d�'N�1�I����Ǉap������hi���,����8�j�e�Y��	�j�
<�$���Sy>&�,�ncpzͭ"(A���Ώ*_	�"B�.Ͳ"�S"��HG�{$#ػ��%p���B=����g�u.8�C�v��K2�XU�����"�%��}�r�&�շB�}�1�G����G�|A��'P[͟M��x��cv6��7�.� �F*�P�$�¢��К��W�v������F�׮~��g6�+�T��tD`�ǡ)]<�ྜྷ8�w̌"-M~[
�q��ލ��g�гp{���9��D�	W�	��B�ݘ�!��i=�f�x�o�p��ꆍ'3�U�Qj�ŜH��#1|��1:D��4Ԉ}_|f��"��ע��0���s+)�D��s�׋C;^���ݍ��v�م�����j����=��λ�������;jwZUO)������/#z�)-Rf��V`d��e-܎VH�����g	�����������w֪�����P�وJB�R��*�L�v`��S��[��\��� ��2�}�Ń:!r��h��E*'�9�eb�I����ZT�4G�z|����볨�1Z���*ub0�,�1��|{���,��*�!W|
����£��??�'{���A]�m�V��ٶS"7�����t�C��j���T?�$y�gq���o��3�cvVR�B�,oa~��5�L�M�f1o���ny��-�
��¿0������z�B���u���1�ԍ� C��r�(%'~�S�I��w`'V.9��K���14��(��/���	C*��z��k̒ ���!�ұ쨩�D)�ȋ��N`_"G�lA��O����ʤG��uၭ[P��+�u9Q��Ѓ�b����6���5��Q��$��r��
3��6���Ew{36m�$��_���L#K��{~�K>�Y]b�;i����ov�AF�VIa�J�p�O���k�KX��M��g�=KS*�/�@���^�:Q�b
�;If���܀��$��Q��g��^:�YC#���1�kXx���,F�w���0���,*�DM��c�AT�f����'1��7o�c��-X�ҧK��G��^!WyB����	�3\IwG�cz���݄��I���[p��_ACC�,�%�:[_yu~�¤ӌ��!=��j4S�2�_�������K�_w-��'h�Nf��W�h8��X�r��3��^�6U}ַ�b�}F��H��f�p8���O*Ohmk���ob��ᦆjD��W�2�nVUO��4?a���c��#�Qq
E^(��=��~�8�Ĝf���%F�Q`Do�,�I��~c/�:�t�����d���k[_��t�H�I��R�%��W"ھ�o��/��[M�jl��R[4Cg�'���p�(��n�43��D�n����/�C��RQ^��ld�fB��L��([�2��.f��}�κ��[�2C�P�Jr��e��HP�����"A��Y2���SYi"�H���T*���j���壱��� ��dUN��lhv���7�כ�����:.�Q�B!;�2��^"+#�l�!Գ��"3��\l�0�;�������� �;��I����}:������_���i����L���n]|"j�`���N��� Qȯd���g��G>�!����G�v�?%�Az�4��"��.��
��ҽM�Θ_�B�0g�o�>U�T0��l�/a|d�[Ҋl[�~���Fm�*���U�ᅦ���@l،ddZ��d/��D/��1�[n9C��6-l�3����Ԕ�Q�QJ�@��.�8��f��ɉ��!q�i�Y�A�J��f����̈́$T�bt)���C:eU2&�$�C�hm߀U�M���Vw�~+Ih몗�hn$�Y��@ st�,aJ�� ����2]|mD��IJ�R-�!N'V�}�>B�"=4��F��J��h,�u�R㖽ϲy�L�y�\��N~��1�ɐ�No��M��Gve�Fp����	�G� ��RG/�E����.�5{�M#�HB���D�H<�3��S7H��h�A�������aA�D\� d�!Z��Uq.�����������F���f��h2ZJT��Y,[�3�c�ͅ016�k�ʓ������H�@%}R9f�htN�X�@6��j�՞�
�,=�3!To��,�D���f�����j��Ywhy��&.�H�?:�=;�RYtQ_�����k�]~ �s9l8��7b�(˛]��X	��3����;*�շm�H�|)$BA>H/��8fiF3+�[�@�e3a�n��@�R�0DĆ'��c1V�Z�$�2�"ID7�Ic4cǛ�g����T˔�����#�
720���&���ͤe�p0��� Bl�lBV"9�>���m�ѹ����r�8.�`8�'�n�I�
�Ba�MqZi!@��L�#��n�� ?����s��9r�*�z(�?�PXUn�������@������LT!�K)w��t�vaJ����L6���IxVC��0k�CTVi{Ce���0#�Ք ,��q��tY��FQ�6@�&��N�j3Ety��/� *s̵u5��-A�.��L�BF�]Dt�¼�����-7�l]�k�� �1[t�K~�8� ���o��a)��<%�م�|�߇F���[���Y!�u���(*���ۉ]ݺ��Xȡ�azdjy�u���e�L-e�b��J�2U��Ȗ�6-�ׯ%lF]m�JF��x���0�;�d�X(F$�I2�@~���V@�]{{q�l7��t�^��XM$��v�����8�����W`���d�6#N�*+�~|U�V��@�W�qV¢L)Ig�j밵����ڟ6�𽬺���:�w���f�y%u>B���(|�6�L�DV���B������C��Th�3� N+����DDwXK�N&�|e��/ٙ���B��/ɂ=)c�Q�+kI�3
�B���W��P����BRK�V��8�F�yj������1�*�%�G4I>��}3�"Kǁ&��u9���If���%Ku���aáC�� �NNo #|��8�sUC�-hG.rBi�*�W�P ��)���=�7ٽ�J�ftO��U2���}h���= ��EsrlTu4dc��R���5�7?k΍��	�>��t.�)Qd�t����"V-*I��}
1-[�C�v#I,�+R�)�z*��M��EhH-�ڐ�'�5ƈG;�0�{�~�	t�ib�$�zfIc1A'M�q�%�k���oAmS���P���zZ�l]��Z�UȈ�Z��#O3��y#����i��ñ1r���g��5�����J8���g���xwNF
	Q|�5�ѩ�1���ϱ��B&螡�3�:Q��"��$�M��j�V
�BIɲ�`�mr�P�\Y��o�l��BdK��y:���m�jBL?���i�x]��:�m��=J�(c�S![�k�T2�	������	��5��\�,'=>�(�A�Z֒�\vFaO!��1G����Qd�ݪ�r
}�	'�����?�O4���׬�wtp\�.��b�Z��0�%D��*�Ì'#4j����)4��� � ��D·{9�����3�A�g�A����s�uO��#L�G<s!Fֆz�����&���p��7�猨f���0v�ُEK�i�e�}!�l�&:K�� �S�@K��V��Ҋ��@,����Ť�9F�$�o����Of
�h�I��U�:�\��x�6�ԋ1b��A�hR��G�@�R�
mS3U�h*D��/�֗��� ye��"7�`� 2�
��t:���!�2�I$cX&���� 9����j⃢�H��D���0�����/�{Y��i`j��i}���@"�d%�������m��C3�\��4v"�4{����͕*0a�.SI�Ks��<�h�Y^����v�)X�E�9+^~��;�4v������ ��ȝ��k��L��l>�^"��ӡ98�6��9:-3G>L�ֹx�%��_g�h6'�RE,��W��[T�H�,D%�&�\u����㢋/VU�ҕs���5D�������R�).�Si��1�']�o?G(�j�;�s��d^�a��;;®={��<�c��CG`d��`J��xk_�������U�)P�Ŷ}����W|K��7Y�p�0�H"����q8p�ƣ�\<�}3�*���Ɖg���4�rw�$��O�D�r��Ha�_��8�� �L �(�?,�.^�q�{/A}C3I��녍�Z�!������L��`/��r:�Wa��Ո�O:�L�fb���8�	�N㘔5���9Tav:$[u����W���Xܵ���.�"��d	�� K0������9�7��h�V�GO[ʽ�;D�ĭ�|��E�jђ2j�N9�È�����H�py�����A�
��A*�{���^�d$�k�i[J�����f7���ӛ��(D�._t�̒��[7��9��ix*h򴢶���d>'��A���sq�U=h��Sռ9>_i��^���`�с;�o�ܩCI;v�@��EX�n�*�<��(í�<�J�;N���* KAʅ؛�K���1[��&-Ʋ���-�]��¿ϫ_�Uӝ?P�E;��yVuZv���N.��L�cX�v��(�Ā�4d�ڛ��QA&���TЊ��P�2�R>����n��I�>~�-�QD��TVk_�]���.��"�"*s������߈��LLM��A$Wk�.	F%��BKr��&e�*-Y�H�'>~5��&{wo���t�k�\�Ab�X�s�t�a��(m��'Lo��ǝCC���>d�ZΊZ-#5��.Z�r�e�7(ɞ�9>ga��~?��,V�i���z���G��7�t�5���Kf�LK����Yַ6��z����	Չ�V�Dt�(�� ��C�@�I��k=L�6�=+�CU ��b%�ҵ]N�T�"z.�=��"cCC�Z��:�^nn	�ޮ
:��W�RrѠU�u�վ��>�Y�5u���YO!	�z^y�h)�5�mm�>�2�!D��.Y*��9H:w��,�;)]�܎t-K� ��Y��Gm���0o`�ȿ���L:SR����c��j�H
ĈF"���Bg{��Z���rI,[},�I�V8�CEjrznBu/pI:������X�v�*Z��sH��Qm�����zms� z}$u��g�^�ll_�jB0����Y�*���JYUR�`���4�$oIZ�Ě�[p�q'�yG��L�$�qXk+Q�"��ϔ�9\�Dcg;�C1����-5X��4��1�'�f�xԨ��lrd�Ҟ�X<����\�;��Ӣ�Z�3����N~�M�C"7L�����d��ƿT�d�ܯ03���F#h"G>!'���If�Af�I�r|�f���i�k:&�7vZ�Rs>R~����1��	鐎���i�5��XL�m��ҩ���ͪn-����*�cSx�ɿ��W^�,��<o)U_q�'��o`6�@�dCh6��;M�m|^Mz�����,a��}��Y�s�QYѩ�6���J�1hSR���
�:�y�����B�s�K+I&˿�CM%��'�b�����1��/_܃��zC�.����|�1I]e���0���c��x쑿�?���}C� 	<��#q�I'k�l��W�	��Ѥd�DU����cýx��q�=w ����Dy�*|C}m#�I�����w�O�
1Z>��c���3��g��-�K{�┓���������Ųr�����nMR<������?�ǖ��^��30K�V�c��%��F�������@SYS��t�>Y^ߴ�Tu8�������@�x[�8��c�&��&ly��c�� Ο�Cj�����*�t9*H��ѱPY��p�00���^f�8�άb�9���p��3�4�r$CQf{�f#�5��\/��.f��Q�!�J��4�*����!B �A:9��vӺ5xc�����0CL�@�dv�}	��݉ǟx_��w�b���I0��c	����-�|�<p?z�~ {vm׳����w�7�����������Di<�3���}�C�ba���-M����[:�R��^�[�,��׎����b!����c�����{���d���N���сuG��*)T�ѹl��\x�H2BG��������b߾=x�'pݵ_b�܀��}�j��\���##�<�׻���~�������1z��ߎ����w���E��-Y�V^�M��=�k>�9���\эO�ț��^:���0��ߏ�^}j�pܐ��j���Ww��o��7wण�����q~͢,��U���=G�%���YB�r�-��E���a�k�s��W�ÚE"=���
� �]�H���7`tNZ�|�}8Ի�d� ��zPWf!sL3Nbtvqf��V:�l���B��u6�kp��~C�Q�Tҙ!a&M�f��YU�EwU�IB��nFphkH�T���-�����x�Z2m1�h.1��Z�IQ�3�u ��I������8���Zĸ	M�d�(��צ��~y�O��Oζ�cA嗲�W�6#����������=sX��UyA$8�j�[�nǷ��5|��_�
*,f�K6J�&�}�`l�\(��FFfX(�ʟ�����;g�eJzCv��/�b�ڕx�-:k\]�ǣ{@�K7ވSN?[�*=�U�������|Az}L�EOgzv����8�{��V�Z�����t�u���w��[����:q��ݜ/������/�]=����Ҙk��R��/n��*��޳03���4sY:�$��Y,]����9f��rr,���^}	w���8���1;��Lr2�2�bԯl�Sņ���p���`&Ql[Y��e� �AUmm�O���]8$Q�Èі����:�,���|�)	�ӄ���;Tv�H㰖�+�&a�-Δ�Ps��v��KBJǐ3��:=�3k��m%�·����+0��rr�Ɔ&U�hj"��9'�u���Xl��3�Cãhm��Y��	*�]��wv���9g�b�!�{(<#�V<QNH96�_�_��:#-�"���Ӊ�}�F~^w@�+���됓i;��C*�����W\����y��I�V��o�$b^o�������&�a�����8BCc��I>��>� 6l\�=��"S�ޑ�i��#�x����6�<��\���~%�������ߟ����̇P�ʀ�u<�䣺g�c��2ch&��fhb��H�m:�a��������aͲ�ط}/���� >�>�#����Ք!�l$�\��N�Ԝ�l�/����F{�����{p�I2�[-� |/�}�>��܄ #���x<2a�������YM{�Ӵ���)���8_7�7�|�����]�bjte�q~6��]V�;��`�I���Q���"�{c��=DZ)����xRU�#c-��L�[��ϻ�p�HÐ}Y���g��f�5�g�CXD���2=X��`3~��?�6iC�_U+�'r��'�NË��B:�&[�d}m�pLW��u�1~��X�����T!�3}��8�ԍ�7VC�v��9�����*��%=�����s���Nd��ȉ��=x������y�!��ɬzkS-�FK��m}��}�Ft�lU-XєjR�ذ#�/ꀪl1?�vx]����q����lVk�/����t.[v	�ۃ�E���xm�5����nƣ�<��n:Q�Yd\�~�:;�t��L���LjK���Z����El�PN;��ԐI��������TWT�����j052M�Q�)-ؼy3�{�����8V��N�T\�,�|y���ʍ��D"1)�Ms$��q42��W�Ӊ����=�>>G�j���kc��/��z
U$���:k����l$�H���7�߹O=��VQ�Vŭ"aBN��Y�$����p���(չ_��g�`M�������GÌ��Fըg��zF�H�>��g�����	��H����YU�3:/K�R���U���Xu���\�jNf�i>��Z>��Z"g�F(�����ڶ�q��'{ژ�]�r�&����T~bd�uMz�^�͚t�T"�{��	I%�H3��R�p��{t���E)���9dQ�p�3Zg���úe�LW��I�����/�h~8�T��.ԅC�����;:��%�J��H����,:�)o��"Y������Y*���mzZ���%�]��5������Q�'g�[��	ޖ�Ņ�&�?C�#���?0����>YRQ[U�C("]27��+]�ɤ,I�}&��t�>ɗ����LN����H?�D��w�0���o���#spT6Ȇ)���u�!F���Rط����EL�4���;LL�h���o|:2���4����J�p�tp�L���f��61 �׬*e�\&�a.g�J�˦�B�N���$�g���[�LXPْ�����`9��\�L�Vj�RZl�X�畦�8u�OJ�R�\�������VA�f�Y`+8�RF�o��a#�\J� 8�D2k���$|N/�6B���(�jk�\��g��Y*����Yk56*��u#4��F?��ȿ�^��S��S6�־#73�����,W�w1��p\�DX'�D�h�WvJ��-5��;�߽#dS)W6�׵�r\����L�Y]y�����Œ�k��H*e�����e��$!�js��^�><d������&B>l@�Ǯ��M-���6��32�H�S�v�t�*���4�g�%t�T��2�,�&/���f��jm'�EMU�~6�h������[[t�H�D�DT������h MN1=6�����w->���G-+u�Qmc3��8�NN=�Tr�)�Zݦ���I>����b*mV\)�C'O~"Z�7~���r?��!m"p�h)��"��G>$� $��y44��	��{���}�r���H��2��c���(_���htb��LH�ׅ�^s�g𝛮�4���ʊ�t��&m"���DoqW'R̠".&��Z�:q��p�A��qxe��R�hE��Txt���3W_�s�f��lxN�1�І�G6݇
B���$��t���M�wtc��0�,_�JO�ә��.�q����^��0b���>5��%G(w8%����k�W02<������=l%.#�`K�n����a*��#�����s��y��%$�E�_�U._���=��#�zFI�r�Fg�}�.*��7��gd0�XPZ�GHv��c3A|���4��ڵGG5e@\��n��{��7����1b}�Z�0B�u�4���'>s����3�I˨����U�1�Zp����6�gi������o�����g��M ]�=!�#��jԆ��h������S�(��G!K���`�����sAG�Xۢ'��/��_��^{-
4�F�z��b`�M���o��$���$�2a� �e���c��C�.�RPQ�xD[��x��p�����Y!Ѽ	Y5�X����'q����J�F�D*�+�F	�6n8��q&I���	+;a��d�j�oތ�>w�E����*������}Twgê{e��������p�����%�$O���Oᥭ۱r�:|���I��i=ܳ�L�C8F�,3A��k'�[#���x���wt{�'K�d[F����v56YHWȦ�t�J��b����]�����(qksF��u%Љ���?��o�f�푉1���`���z�j|��ִ���]r�b�`8����9�T�X���_�i��`8ECu̅2|�k_���C}��]*e?���Ez�w�n�������f�;��eJ���/�����/����i{dv:L�����Q�+[wa��otn�=�л�U����uW�ɛ]�LR��LCn����0J&

������8S�l_�?��Zf�g�� ie#_�s^z�L��dH~���Z�W_�ic�l\5�*�n�:)�~�ySg��3)��~�����eU�����|f�d���:j﹜��҄p�ի6����ؽ�u�P��I���)���c�;u�|?�wyJHu�DfF>�l$�I��|�a�VU�v�ֶ%�~s�E��=��HlNO�E�H�^��Z�'���>�({nnjřg^�MG��KV0�T�LG쌯��"��^8�����m'�_��A��p�/!�M����&F��������!�`����Ќ~��t���}���M��E�H�Pv.Z�N~v�xS[�[�\��c�ڕ���W1������W鎱ޱ!ř��L�ڷo�K/o����'������k����>�����es�:�%[\|����Gpه/��O��aF�A����T����P�D�I��ѳD����C�ON��܁���8�w;�a�^�����r6�YW)�����8��K���ERW�2����clݾ�����f�0�/_��9�B�E���Y�o��1Y�>::B���M߻Yw�f����O�"�KZ�Fg+��*i|��<�:6#x9��e�~��r�}i�W����\\%�zbwXT#��c�ɼ¥��e��7o!,T�'����z����t�`4�s��c��<p��G��$�+��?����/d ����3�d��-��#���`�t�󋸘,~��w2���-��)��U���T���H�i�&�}ݬ��F�m(��o��� ��9ļ�r�x4Rol�4��Þ�{�c��լʨ�\�X55�#ݥ{p�]O"Q�&f����.���y�F7��v��1"Jӕ�N�p�&���\L���.��t�����!�?M#8����TbͫP ���ժ��@)KJ����pک���QW�>-c��YOT��7:Ї��������(s���^x����t���0&Qp��cvh��ǉʪ:F����d��aQ:�ҥ���ܤ;�d��[��ո�����rȥ�tF��DW(�ѽoق�g*{�D��X�ي)m��9Hc���f��u1S���G��8�@%!�&�pb�e"&S\��/�v9�p{��y)_kA:g��_�X]�Z�ٽ�2S�R� j��#���눓�e��:��;w�Ѳ��\�*�ȭpV1�;�:XFh��֤��RȐq[�,�w�0F�<)�7�7NSSgU�}��VT��Z����k)yn��b�֑J��JʘI���N�.�#�m�����1j���Gnđ��kӛ�@�é��A^x9v������9@'�����+�`�7ѫk�D�fכ��kQ�;'��2d���=wh�OV�nX�^��?3Đ����ؤ�A/I��b�,��֗1E�.����W�ԝ�c� Һ��Ub����4u��iU�����v���W��aN���c�Q����x�sߛ��V���e��tq��1;���x��^���E�ty��Y��˗�T(����H�*,�>���3��% |������^�g���6m؈/~�Z4��u;L9�΄UF�4��$d�����nՔ�"���'w<���T��)�����ɠv������B�'�x���*�%��R�;��Sp�5�'9BF��D��{�H#���F��/�<���ƂC�_�Gq��G謓3��MfD
��!��\�MX����q߽w <3�������)|��H�����)DW�2r�!�Q36����%��X�,��J+��Ė_�:�f62��q��e�꺺C&�)�/d]"�;M��y��rr�)���`$����"��S��������%K����^�|��LF���篻{v�s�G����Y���t:��qh��јD3j���qtb�0�_���?�RW��C�Q���	?��&�/,�D��[�l+Z�ʥMX����ڹ�v[a����گ���RҪ�T{�A454������⿾�]��j�8s�~����%8��p���Ȓ�N}5t���A\��s�����ܠzώ}�/�-����g��1�"�qy�^��m�8��3t�K N��R�$�����/��S�駞R�'U"���&il]�{�?�7�x�*Z� ��4>��ؼ�9���_�ZY2.��2e6;;M�i't�����8֭Y�ٙ�A��E����a����ˮ���3#����!;�d���;���n�)�[j�YQ�짃F�o��H�E�Aޓ�zn w�\\vKK�N`��C�a������T�Q�r��Y�px&_r��}�% +^�6������a2�yL^Xҙ��ɬ��,����7���R������q�o�Ӈ��r+2�9] a�k����}���P(G�jV�'%B��}uc�����������M�8V�}�C�b�C�k�#tY�:16�O|���w���N9Y+T��iB|��:[��k�A��]��No�JY8H&ۏY�[��&�ۏ��;��-:�)��S�Bϼ�Q��%����`�Ms�P����^��} ]?삙� ������k����
��-�Bf93�F����g8�ēh���N���%L�֡��}�K��AFf�Q��1��cU�=��7��e����<��p��4�!>3n���
O��i�^9GH���_7��)��7|�������D��df���Ď��u=|kkk!�R�;�c����N���Ӫ�z�{/��L����`Yr2B��#�b�nf�jO�l�9|�N~�~��9�U�ב,[��Df!h�U���%ϼ��S�_�B�U������#��Ҏa��8�ZX)U,��]�H�ҩt��kĐ�rb+�$��������2�<����Ie�����'_��߁��{���v�2B���@���woA���ǔ/����KJ�C�\�n~����߬"]�����ࡇ�st�٢)Qj�r���\"�If��7��#�:�Xn�O��%�������l\FB>�����m�(֐����߰��3����tI�Jd�y�����!�E�L�T��}d�`�`w�T<��{�ť�X��!�������Ҭ�V���L�6j���Y�"¿����/~MN0�;���,f&G��c���1�ߧM�jm�Z�@wtu4b��jۋ����2;��4�?���JT5k#��Q�k�ז�T2�v>����\�яc8V�ho%�݁�}�|���5��"*N��+A/�2hi�����I���dW�<��AF._}��r�ܝ&���체�ˠ�d'mg�к��K���}6"~Q�?��-�Y0l�(���4��~مH/_j��=E����X�#��w��us�|I���a�X���e�J�����IF�aM[������Ri��]et�������O}F�.9]��i,���/�>9�H�S��#P��Pi����.�X% U�T�j��E�Y�9���=�QOR�j|�Ձ v��*$@H�o� ��au#� HD�gĪ 	�|�=8v�jjX+R`��
����0�����.�$�Vvw�����| I��λp�'>�I}m���ЏS�YE�5�3ж?I�d���N�  ��IDAT�E(��s�PUPe^f�'T2G�.I�g���Q�I(8	�ۥBY�H��ބ<�?��bú�&f����d�&��)'�]��G�ӹ�8����A{���[N���=;eT��p�ܹ�N<d�j��M��B��ك�k����)�HP�I8�Ղ�o�#�� �<��,_c��n��N��B!��^}K��թ����	QB&o�I܋.jA�
&�Q_�rޮ}�Ѐ��|��Xpa�᝾��#��KA��6Uڗ�I[����C��6��BJW�J�/CR,Q�UيC���fJ��dk��Q��]��H�i�I�[����@ʬ�(ODbIF�Q4�6�I%��PH.H������Z�U�%��H$�{�t��J~��pXU8d�]��:��1Ի�54�ꪅL��{� ���c����aTz|�=�ePY_����6�j�zE���%ዧT�H��ʺZ����_��ITh�V�C�̈́����Z���*����
�3�&1L~QS�#7�C%ў%g!���UYFn�RQ�+���f�ۗ�-eL�g�����I��.�I�iLm��d#N�NTc���|(�?�C1���m��!����'"��c��ڬ"�B/j���2���e���I�V����GN�����z�/�:�p/H@T�E�IJ�%�E3�[�a2-^��������3ƻ�F�!^kYy�hQV딙1�&{Ĥ	L0���=2�V#����	�Cz`#Xʤ2
(v��u���$�4\i ��|���B*"�#S��[Y�Ѡ�7��0z�.��7�#OV�m�FCV��%-o%�,�C�r)+D"��T3�i��I�%���m^%w���hk�T\��j1E��o]�#�5#:�+8�kHͶ4�.3ߗ��ZT�r�r��ߧ��D"�����a6)�G�f	K�t|3����aAMkF�֬Z3���]B4�QyM�46�Z�W^ކj�	�b	�v'���D��(�[�'�_����S�6l:���K�=6f�Q$x�.�VE-����(��O=E#�p�����V�hn����{P�̕+�k�r��IS�"şgPW�.9ߐ����d�ݳ��g+�C�p�=*̜���et���v'tu�H�(�m�Щ4�B��QKD�,X�oI9��#�ۗ��������^�7-V��b@2�')K��$u����<���.��r�S��:�m^��P&)�7K2��x
.�M�X�l9�<��v2�~d�oO$2�b!���c�jLr���Ä��֤��٬��KC��4���Z4v��EG4i/�\<����55��~�F��*%�^B2�z���(�FzH���##S8�F��3��+� [/_ڍ�����+ϣe�ZU� ��f�!I���uGi�rfl��ag�s!^?�ŏ�gJf�]�*����'�ܵk�~�/����"�B~!Q��S���Y���fdlH��~��������\x�{�N�:2�gu*��x�8���h�����FKK�:�4�y�~�73�d���O�L-�y6f1,Y�w���n��1}��"'�m�vO��gW�_�@Y�S{"�#�Œ6��3߃��a�a݀d��-./aR��e��+�@u֭ۨs沓:��D���� ����Ə��F�H��%Kr�w�16�f��%B d�@6�n��MY��!�B !� �����ݖ�޻f$�h4��ɰ�|�>��c��̼�{�9���l�fEz�#QD�J�ZQؑbƞOJ�_��-S¿�Ɉ��a�z��b��	��P0L�"m���!+	W\u��[i��)�&�Eh�A��K��f�|���UV�[�\�`�ړ-���wx�3l�����}~��^>���X#�����*�hG�Ԣ��ny��a�`���i��ǟ��Bye�)���h��Q��aK��W��7��<���\�\e�;[ }���=g�;��T	մW7�h����t�zt���v]pN� 3�2��X�to1���J�Ųh�	�`��`�ࡽ�C�p��x��N����E�Y��oN�ލ���^3",��_��+���܋��r�T���hJ�����5�Cc�l��I��w�6!o��w�{�y��;5�� �ij��Z·������C�;�F^��q���U�O�����?�Ey�<����3���5'��k��6��n5:�g��BNA!���z����Q����7�3vb�ٛ�NFaq�m�Q�HB�.�
�1^�L�&'�$O�P$�cN.T;��ӧVds:u���s�D����'�_�����;[T%nT3��e��y���/��o��F�8�y3<��7o!�`��F}��˱�ep�R�h�1ހ"��'U�����^���~��L�l��h�2�r�����E̸,Z����y<<�a�5v�~�0�w�����U��yE�O;m#���&z�"+CШ�u�ހo�v'|>F;�,Y���xrLj}����j6^y�ct���F��P+��0֬Z�}�;�c�;|� \�T��7�� ��� ��J"�)y�����Mp���X��"��WKJJ�K�M�o#��(��ŏ���}g�Y�A�����/<��-B��0_;f2�2^;P��w�z����w�û�k������p;֯_O���Ϣ�����ͦ�����m<�<�����{62�Y�\���=U��Mj�p�ZG�D�}��,Z��ЉO��=zB��\�r�>�b,Z���3������X�GaB	%t�'	��@H]��2�0&����N��u��<��~���@l����?�]LWר]�>@��D��,=�65C3̪�PV\ER[��]���.���E��!������1����X���J46�Y6J�^^�l�}!U�h�<��8nLm����u��s���C�M�Іo��pme�4#�z���%� =���^Sm׬�/�r�����i �H��ƒ5kQ���~��EH)`��1�0!�	^��ׯ;�]�������	g�B̘U��V3ʑ��v�2�U�\���w��a4Ŝ��P<s.�Htld�ȯ�ԕ}�кآ|h�i�H�:?q�N�|�L~���x��C��UCikoBG׀��;*$� �@ﭵY=}��e�97��[�ƗOw���ާo�\��N�J�W@�{���:D.�|���y���;��d�T��Oyh�H�JDy�z���X֝�����*�j��ͥ���z޺c�&� -\�\i.#���b���zh�$&4#&`��<��5�s��.Q3��I�i�2�h��<4�b��R�m��m��a(,.����M�Q�#Is��t��V�~�q>�,�Jb��~_�`��iҍ�C!,�T��F#G�kFuq|�H�3e�E%��V�K�g�u�~���$40�`08�eb�$��QF�І���J�[�G�R˖��V�(q�/�H h^h<B��Dɢ��D� ��H��=X<o1�����ߍ�Kgb��}��������eSWE����Tn^〩��kg�@74�1r��>0�)�,	9u���TUWۊ���D�,������GO��_@���2���f���{�o!'*Ʋ�kH��*����4��h"�,��zh8�䐭 �쀔U��G����=�O�d�;lh(�r9���݄��n��6�����ϟf�J�����y�,ϭ�n�#8zd�u�j���Y3��}�L�?����?2���>7~�y�4�~��Zi�D�o����hdO��ˇZ[[��ϖ�E�!�j�j�	�2A��[j�@��A���1��R�Wi�L_�ɫW!����}���nK�U��$IN7ɒQL��}��/��W^0}�Z�I]�,��P(b�J**+�C�6���!�9����O���$����A������V�[����6m�$�c4Z'L�:ep�G���_���?��L�;Ń�7^`=�*�|���:�\%8��M>Z�:��m� /?�
v��І�G����+p��� �(m-�<�QƤ��v=��������;$l��v�v�����N�=ej�P�j��p��0	���^}���R��Z���+&c����=r�,���D
�C~>�,����{��P����4������٤�2h����o�4�^��f[>_NE�T��];���/>���z^[&r��,+u�a�g��� ��J-ݭ�q8c��gx�ߺ�?�����3� �5.[�W]}=�=�|�ٽ�>�B�h�6 �`�_�8.�2�-G?S\�B<�k���:R�c
�"��Ħ���O<�ݸ��+��Yl>���&b�d��%�M���ކ��}�b]�noF]�ean��1�<<��CX�z�LR7���Ⱦ� =�ÿ�%^~�V�_�hox'_�NB&X�p�rSJ�N�c/V��a<8���w�}��m��<���h;���m���C��W�BkZ���,^kn���} �k���������;͛S�ѡ B|�I<���ŗ������-�����"�������Q<�����SO�8{0k�\tu�㞻��#��>�(j��-c���N�����yVv��sq&=8������%���-����7���Q+:3��m��?���yy�Q��(���Ռ���N|�������5��	�Ծ��Ӎ���8|�0V�w�u������0���݌���lܸ��FQm����8i^�OO>��{�Y8e���Q:??Ǐ7_������&S��㩞>�T�;��PZ�����طg�x����1����w�����gl�
|H�4"�)rl�)�Y��ԟMA����w%��!�rs��G��W��<�tt�ܼ�H�1��/���]gz�>��ɲhwXVf��ɇ���D~�!�"+�UUT�0��5W_�g���I�ŉ7�P�Ij"o8�oƵØ00?;��{��+�������5�R�K�2��P�c�6������z�N���53�N�5@����O�2���R�4�� ��G�����E��H�E5y�6�����m��c)��+w`�7��?`5�Bz�S������9f��:��fF9/2���C8e�J9t�FD������2<���h�Qe���`��$vQ$��m[���V�]ec�J�l:KCG�ly�	sr2x0�7��i��>�>������o���Ɍ���81�+/���?x�F����cv*K�h�4�B��?�鏱h�+����V�W�������1#����e Z���))5�����r�:̘������k-�5�j��������ڈ��D��̠��Yjz���u�M�E��� ��Z-��@,)b~�&��S�2�V=�t��FP�TR,����� SD�>���εF�ݻw��A,˛�p����f���>�-��0���\8R�h���8�^��uux���q�ٗ�j���
�)����'����?d�o�É��>5���l����n�����n���>��#�ک��c$���A�%i�>s.��=��ϱ��s�p�R� �C$����|�R]|z����>�9o��׶o{g�u
=�l��CYuz�A�w�fֺ��J��Ɓ�{QX��J���0̣�=�;n�:�7�J�_��+�=���V/���X0��I�L��f��8�\u�5��=�4���--M|�hik$�JGuu6
K�ɓP��P+	{>��X��$60��1n�u˖-�;{�}�H�4I=^�]����LoO>��V���?	Q4��ʫ��H?��CS�a���z??��R�ҳ���70k�B��|�<,#�c��7w�H���ح^c�)rJɱ�[������ʖ+����M���I�ǩ��T��o����k�j'�4���/�_K�x���,��H��b���ՂtO:>�_��>�u׿�@��=x�-c!�����QBl\������D��K�r��/��u�]Dx����mM8|`�C�F4Ӳ������j�e3R�8Z׀�W]m�>T��d�L�={QR��O�����z�zg��md�/�݉��yN^9	����i�.���g�������b/�t;��QHo��PA���q"7)�0C#$�i0��CG�����SbZ7C�����.��3�����[�t�e���6�(ΕX��fh�����4�#���v��n8�f�����;0<2̧�a�*�1Bvw��ܾ�{�z��tu��P���J�FCQ��w��4��Qk��QƸ��N�$1��=�6��U�mc��F�3U�ӻ ���IcUu;� ��3`Җ�O�����x���t�'B#�����6Ao���ǥ�M���MGQf%�Rǽ������7Ă�f�d�T�9"��_j��
�X��9�Rfa-c�A�F&�|ĵ�BY�AT��{�z~��e�����1��q���J��Fx1��e$K-|�q-wPPm2s����-E6��EIe)>��$��[IҪ��N��F3z�Q���t1���b(���oi�;3τ��˴`�td�Gx�K`�	����"ț�7U;�+�Į��<D�1b�qL�.�uK�"��������!�JvVY��#dtrY9^����VQo}�53���چLߔ�K=|m�9N�FR�;t��^����`��3���I���E��^)���o�-�d���k��˨D.33=��J���%z&R�6�|�FJq}�Ȫ�pOS�jˎ�T��/L���[�I�����X�'�ו$���P��v��:��ɶ�/�51��Rwpp�gT������ċ��7��`g����#�٧�J�֪�2���^��*�Tm!9�s��)'8��7M{����dU�>���ظ��Q*�PH7إ�J9�����Ǒ��_I����
�"-9Y�6#<�ؘcv!�Ӑ�zMy.[e� ��rެ�HM�3��RI?�� <���1�&�TVV�=��V�)�(�D��Y��L���[Q�kLb��.�<9�����h}!L!���֪�~������:?�I���U��Ԣ<�ˤ�x\&A��7U�'$�����)���G��#X1Ml�Ԋ*�Khٞ2BU5�6Ю�-A�;��:n��W0��"����t�҉���4Z[[�l�r��\Pѭ�v��[�;?2(�&t� �А�"������9{�M����ä�إ�^���}ʞodbКÌ��ZE�SVJ�G�Nr�j����B6��e�]�{��nӻ�P�Slپ1�ʨ��������ދ��	�c⹉�IL�����O��m2�x�R�m�$j�д��O���X�d��q���
MI�+"Dc�}}B��U�??�|\�"v�a��I����N1p��c|�(:��m�ZC�a^|��@7I�I�fق�C{�l�ɥ�`i�~Ls����;���'�)�2|Jү��+O��w�������<r*ᆋ7A���a��5<���$Z2f�1N/��/}	�>tj�+i�](�w�OO��s�I�-�+j0�ظ��'���z�t���ݯ�b��}4�ie�18H~���*��3֟m;����M�y����c���ы�r��6&��H�L:Q}Z��9��17ٓQ��y�����~��C�-�fB�s����}��k6o�l�9*4�_ł&�/��>�x��4ސE�'T��n^N����Ɏ�.�P�йI�`��K1<6���}�8��>	���@J�_u�fkk���&J��������w�1#��ed�b��L;��5GZ&����:���(��>!F�K.�̈=�	���1�ozy�62���ƚ���/���g��'�������ҭ2���QtR[�25�<5��X\?1CG�˟��r�iؾsJƅG�/�ìYs�L�cfa�%�,o^����څ�����݇��#<�ڝ���:�W>�'	�]��K�ACk�m�Ԑy�+�d֝u�n�x�=pe��+�#D���Z�3��"Z{U������i.z r���_��^}�9��������$���#���+����ѓʚ:e۵!'�W^s��Ã��¥i�y�
����r�|�X��d��I�l6z���p�����nśolA��v�,����9��ё .��R�:|���m5Hb|)�G;v�C�R��VT8��C�p8q����H��U��h:�`��53�������(�'�x��[J=O�B�ګ��o}�0skG��qbk-lt.��<W�Z��[+�x4���z+B�r�-������2:�@5����j�@k����Zl߾�E��1Sپ};|>n������a�0"���	6ۤ��=���LY���Ut^���!پ|�5�|�Ֆ���Ti�ƣf�2j�5�K�Ǧ�p��<��ӧ�s}�ݧ*�������CsƌYغc�ɡ��[�䗾�Ư�"s0(E�4t���&δ�\$���ʉ����n-����)�e�^��Yk0�Ћd�p8i%S��6����u`�ϐ|���~T?�w�p�����'�c�a)dҫN�;�zRM/���l��g���]�Ġ��L/�|Xt�\s�M��3�~E�(�s���ߩ|�sQʈ�H��������1Ђ�sO��|�xEɠ �x�f��
��]:0c�t|�o♿>e�þ~�	�*I*����Н�&r=�)v��y-�����7��}�6�n� Z�%ޠ.Z
i�y���:d�Wչ���Ν;q��!�R�㌙�f��R;���8�2.��yX�z��C������d��4k�k��;|ȌB��ľ�!��[G����oB�r�#��A^7�r;N=�t���!�(3#ˢ`���j':�'-_�;�[?|�G����g��o����S�M��.WbC�~"#6���/g�;��)�4�6��>�IJ�?w��o!�������-7Dӱ#�3{���a����kѶHr6q*�&�dR�kN݈�T.��^�]�&�Tzl�X6�F�7
x ���Nq�r�U�A��0N�pf�[�yQo��f�CrG�#�����&S�JV-"���|�����w����x`�qg��ꁷ����0♝E2拢�W�S#�TA�ן|cC�8�� #���g���*8l	W�Ĵ��34���Z2�t��\��^�<S�k%<�@��#5��ե�')�l��1�ԍ�t�2̙>� ��|BQ�رF8餓��A���/$fo2ܭ�OM�b�ZI/z��:zբ �R�J֙:n;�J�B�Cs�)����k�L{=Y�^q��A�����Y^�"��J�j�<�/9�3q�e��,�d�1�y�����Hk����x�ZD�,4;];c��L7#�u�_I�Q
��<����%��d���q�=̶{6f;������br��e��5k��<�-�'���߸i���p��g}�E��<�AzT�j���2&<>J�����$8<HV�F `Jqy�L��NR��N�����_�X��8>H��������Eh�i���#�$�*-/C��X����A����׾��vD(/1�sE����aP'k5�Ӻi���©�b�<�m�皨�����c2�rg����ԙ3i�5e�xx{�푧R�AGP�ݟ�2��[RRn2�J�ڵO>�m;l�b�
�u��v�iZWW���&��'F�Ki؇~�h����,-3Y��s�YVI�M�_?�>�gW�_r-o���A�Ox}��6:�ґR󡼭Z�u�D��~:�2������K-��6��/�����.�5���jI����m{�Ӵ_]|�R�PT+�uK ,v�Yy�j,���G�8ߴaS������kg�xݤ�iJb��`r���v&���9����!͕k��*��J�˴����hG��~F�ޏ��8�.���
�7�3g2
�P	�C�H;�<y���#��`��?��;_Ę��Pʉ[�_�+N��ų�GI��ťF@g�0<�yh�:�??�(����Ó��#��sp���a��087�5wF�e���|��R��z��o�e{�I�%z��W��6a�i���0��t	ځw���xEٙx�՗�����0z�@�Ǔ���e��&Q�kiW���;�a4�����M���}�M���+����12U/`����ҽj���p��O?�g����rtv���?"�r�����_n�~��j�ٖ�L|��%#�6
��ƃ�U�:�Ͽ�
�<�L�t����[��Iɘh_��3����?��7�z�Zi�f'y�Z/�T��N����L�JE��������V\S��F:�:s�i�p�y�x�̘

K��� �6���{����ű��B����%��g�7��v!�Y$�ҚSO��FN駼��_E��VZ��~8�m7HP�'š�����X8g9qx#J�>z���ҺhF1"H5l���$'�d�9��(�"5�M�����4����i��k��jQ�2'%%e8r��-���_�#ݍ�rV�+Acc+�^6��j�q��1c�)�b6��p8yH�Z���_��x3���M���<��㣿�Qb싯�����Ӯa� d&K�<�s4;�%�X3Y���1���|ؤh���oD=���5�ǃ�~���yCy`�9�]��6��z�W��(ŪbZx<dT��2��|�{�j�ض��8�<�Kءt��A���K7c���ܴ�U�A��?��E��y�D�S,�f$Ϸ����r477Q��'�F�}�����cs�v�H�K��5���ÿ�N��V�Dy��$][��J�Jp��Z:計�&=�>�-����v�n��n[�դ�#�l�4��b�R�s75�y\��s-�S���7ʦZ-9^e�?'.�200���a����[�7�o������_R�^�Ҏ�Nd;BX�|6��:z߀��57c0�/84g�e�>Z}���OQUG_O!z�� �C�����q��;H���BE�a�䗡��Sl�O8e=����Jxh�F�(;�~�m��'A	�/��#��	���S=�̚���ubC��t�q���SX�zr����NzX���<س�]4݅����4���)}�`n51�'�������oŞ�G�YK��~��K*m�d��Ox_9|�)Q���н��P��YۅDՑ+5J��i����HOs[jZ3�?�N;�B���uQcdܕn|b׮]ֱZG<�ޕ(^���DQQ��u�?ڜ�7�$����um9�y����4<��d-U�*+5�u�$�KͰ::�li�
]{��1m���\�礣���r���0���L���OɁ�QY3Ӷ�ʷODbV��K�ǎ/L4�!�wjY�D��[*qb���!E���5�%#��+���)�)�9sfم�k_AF��׿&2��� 48���<�V��y��f�\HҴ�Ш.G�yn�~�#�%�1�ׇ�Drܚ�$ ��#��~�]���$�=C���̰mC8�x�;�hPj�q�ީ�mb�x�,]~�U�����3ܖ�#�4i�;lݫoD��!	uR��O���{��� �w���)���HԈ`�j		�#�|'j*��޻[���s����Pc`�>;|m�8^�^�������C�6�`�v�dO�^Y#�%l��!=j&��*���MP2��V(��� ss
M�E�DQ[pKC|A2�k��W�#�����)ǖG������z���/��2<����g̚n�Dc���.���񉈣t�����W�:��9mֹ�y�(����.g	fͨ���k��T��Q��>:�F�M��3T3U ����Td��)�{����.���z%k�7Y�=��
k8DX�����3k��#2��>۾�r�Z�H�K
f��̵�s�c�h�ً��TK^��e����[�`�_������(J��`h|��!�J�-؂d�=U��Agz�y>�p���Ψ����]8��s08�O.�Gza:vm���cVq<���++������1�!EC>!F��L�!��b��J4�FIa��C���b�޾a����F�D��_5Y��;ڽTF��w��uk`�OCC=��?��d$�ԯ"��3��»�q����@o�M
jrOݻ��|�3thf@���caӆ	mQF��.8�"�A�E$��F���WO:T�-|�%K�`3�P�w�u�-{�q�3r+��[c��X���&X,�4I����2�C����R���u� �Ȗôv�a�BnJ�z�RRR�W�u�_�����D���T5@�$�6pd]���5��d��F�<r0
Mh���Y��{y�s�U_O���p�ϩ�7#���0�,�FZR�Z������,ۨ���G49��F{1Aҩ�Xg��l,6�3�7#C�
E�ɛX)���re!=Ǎ���j�����L�?I����g5�	�x�z���"������~F�d{SM�14�k�_�&6?�ԁ��2D����x�])�y��FJ4��xL�������=e˶6�22Jܬ�Ș�|F�xR*��#fO�	k.����<p��	+��YtM#�6U����A�Q=�ji�э���Y��(]K��Lޠ� r���Hi���R(Ԇ���B�EȻ���&�F�EFB�%4ܻg���9��8ő�	R�ț�����y���n��SE��RD7#�TM�iӼ���%Ȩ�29H�V�碹�.�	�|C��ɰȡA!s�D,2t%���-5��<����(��a�4��jS�`jٸ����g���6����C�
�J�/0��8o�̙�q�)k�9[�AϞ��MS�QQ̐炷0^`��Pc�R������â>�����,d��at� ���^�46��Hf�,B]s
��}v����/�COUX<i�.�u��,Oz��L`ޢ4d���������/B;=��Y��o�Af���U3���Q�X4�0d?�K[O�IFV�@r
�jg[�<��IE8�'��a���M�������#&Hl��,dpF�i�D:��Z�|1����a/�l	��{ɊR���;w�E�ʲJ�E���2�V��T,T$ҿ�sТm!�3�[��oR�v���6�+�����'�p�B����-�'!W�� H~a�e��[-���m�MC5��VR�v�؁�l�-w���v�?�`)j����̝?G�lъ���~��d�j&J��"v�����5W���V�p9���qF4w�E9���d�g�BqK�Z(1 ^����罿�`j���3a�'����j��'��M�����gR���ZܷG���?	�2�eá0Cp�zdGF�L���ц�H(%��m��EuI&:Z�M�H_2���ȄiYe(.����
��0�C�9�����N-B8��!�%L�"���IH��X�'��Ƈݎ��
ݸ�.��?�_��<�HfH�%Lz��Q6}�ym��M���.�E���4��˷?��h�DphU�4�.8c�7I��`�SPYU����jj��4�֭[ͫ����f�%7���٨�x�_DM�P�����*�m�N�VuhuXB� C�4TZ�{��v�i�7ir���Ɉ�����G�"�W�PA3�J|� �}Zw�:��H�䥹�ֱ�����W]�ė�|�5>��M ����.F�k=WǬj-:���ڼ�r<��/mf=F���sZ���k�;'�\�������c6o������6���oL	v!���$�/.��P�KH�$�3-u��O�$��=Yd;qC�o����X����lz�t��q���ӗ��7;v¦ӧf$ӣ�A�tN�tb�|z�n��JNE�| )������ɕx+� 6d��7
o�,�/[�do::{l�ީ��\x�+q��'�_�u��n��g��Ϝ�k���� ;����4��^]�az���*�>����_�������*g`�?B�X�Ј��-C�G��C��H�H�q�X;��_��n�Gxx�:�=Ry��b$T[���'��\��Q�]���0!^6�{^�u�����V0�K�X�
�-2Վ(�";�s<�������#>?�rM@AY�4z�U�O�-_�͊�jԏ���2��=���o8���w�܅�������bղ��ƐE�v9,�@ap�<B��������>8z�H���n�^$k#�tY��4�<vp4�LF�V�Ak{+^��o�u�Z��[���眇^���F;�B���$<8�o�.��ɳ+K�*)�DL�"6�~�*���:g5d�/�#��!���2Cd������W�W$T$���m�u�ҕp��=��Q�������KO��Y+�H��IG��ic���!��9��Q�|=��;�����~de�(�yJk�ѫ��E�u�Z?ш Ġ9�娝���ek�Ar�.�Mq�a�9p���H�+q�H3�5o�Dؚ�D��),~�_DE�,l۱w�u7֭?�P-y�<̞=״�vr0���Jd����Y^�&Ժ�g��ѣ��{;�B�b�
̜>Q��c-�ġ �(�d�b̟;��A{{�VIό�E�J�E�0�HM[$�� �2;?����8���s�5|�F6��<�`I�Yڧ����b�%���}{M"EY���}ՕU�n�bTȱ��>���=�JX�0&���Kqq�|ӟBPUZ�lj��a̰���h��22���Ʀ/��g�I��j�����a񢓈6|�;��s�dƧ�ri�J{�}��p����NL�NaEm.9��L�"Y,1���L�"���qVR��bXm��	B�˕qM�8�����d,=�5U֑�`�X�l�d�I�oڊI�Q'���C�8��JE�E;�R�)�ҩ���P�n�'"����0q�OAyI���ҳ)E10B_�Y�"5��q�雭�DDP[42Ȑ$�LP�W;�SH���WMj�0�>3�{=�)�^���*����/q��'�B(�($�>���>,[�uG�ȴ�X�p*�J��=a8^�+N��Z��4����*�,-GIY.m�Q�CoW�hK����p��*��N,N�0O���ô�%�� +�-ݦ���8!b�=͞��ɦU�ơ�����Z�c�Avn��|+eK�E;F�G�t'�:�����-��8s�]���E��\"�qF3�<�ԍF�ĕFx?=�r�h\��T;�R���G�H%�(�|�h��ee7��ktRqp|b�P�й�MUF)>%�8'�AHlδy!$M �s�\�/�k��!/GHT�� �FU�e�!���R�!>�����*��M��Qk�tp�x��>t�C�Z-$'����f�?��xV/����͑��ۑ�LF�H��ɏ��~zM5�EPX���a�vӓxx�L�D
_+m�b�l����6X�̧��6���砨X��
}�|_�뜜,b��xj�.���s�z[i����N��\s�&�Fh˨X0:JL��C����=sXu���D����b�G���H������������]gj��R�[�~h�_�*:0��S���a�(��5_�c�[ob۶m&�(���gBQ�?�B��&�O��=j�;f�b��D҄�c�F��dۻ���`���fp1KM¦���Z,�9�S[�mVY��l�;�$fUJK�MqPݥ�����E(ܗ�2��i}TJ���a��X���X�2yMW\qf�]��c�ƥ�yt��:���[9�$�5�W�'�FxbbrcN�G��ܑ��#w���x䑇g/Y���̛�<��@4� ÿpz�'� \�����������Q���<���$de�b�_1J��0Ҵ�M������k��D#��n�����j�d����4��x		x`5O�����ڀ�%D�P^U���l�9�.'�L�r~<%�^�^�{���P^y�|��!�vgf���~��k��M_�ͭ]����y�mԼ�fzc�t|���������_eL	�v�z��n�n	��{��E&��>����^K��h>|� ~���h�}����;6�?�j9�!a+����b~G͌�oF��-�Ev�57~p�>�\z�fS��g)T�h���m������q�:keѲ�ΞNC *���؜0����F����!P��^��*�)r��;ɵ`߾�i��M��^��15ۏ�������������6�j�`�?�ѿ`)��%�^i+�Ba�j�]�^r t6F�c�I6t� �e5���R	K����ѱ�,ӂ;��m����Á{	�+�m����۰|�2l��9�e�Hu$�l�]���&�%�4��B�y y���&���V0����ni���}��>̃Rw�!���9�`��q8�z紤B���,~	�N���� J����� yn̞Y2�� �F'�k�扖.[���P@j� ���Q��?���(�/CQN-�\���B��N��/��u:��'E�5�v�9�'�E��}�*K����W�x;v|����mipd�"��Ou���w�6���C��?>i��~mSb��V��pќ��-����G3J{���Iǵp�t[�����Xu��K.�D�����R�ݽ���[�`�R�42q��3-*H���'��5���/~>�:�֮ HU[[���C���<������
�T�"�s�<M�4��h:{9yr7y^6>޹���1�乐�N��%��m$���wY�x�g�;̣�p��$
�� %z��>��~=��a��D�����)>��ZZ���iތd��H^bΏ>݁+#)݃��X�h]���J����PV���ɱz��g��������JF��<�uğ���	�n~�q2ze�=V�w�1'����S���(��s����3�e5)>B�B���g7@�4��!bŷ^|9eį�Ҥk_x�P����cx�ݦǩ<��d+�ky���믽��.���	�7w��ւ��~���t��a}�Qk����
��ꫯbÙ��{�lz��?���ڼ�I�F��'�DD5l��]����,*�6*=���^������0�˄�+Gh^�����ƽg��a9kn�-B�aZ���K/c����$������j�[J2n�����K�5��\ځ������[�f�r������OIV�-��B�s�����o�V�M���Y��9�7�f�מ�ý������d�gϨFg���˟�x�*�{
�Tcp���S�xUR�^LBJ�J"�VN�����v'$R��Mw��$=M^������74����XJO��[�~�����!��*\�Ԕ 2\��u��z�H��B�ԟ�`p� <���I��5.Fp>�p����Y�ę�B:��?�e�T��t'"������Ƶta���h"��6�=�0<a����1�A�\�3xC'x홅���C�1�հw�!\/��E*�{= �M*qm08�W_~�&�2�ҭ1OU޼���d�L#�%�:����q�.�p��z�_z�%�v�?���1Lm#R�WdN��Ё�;e4�*6c����+�`ӦM�UQ�PB��g�+*�EP����99^>|���f�6���oiUɡ�Ϧ���(%��Ov}����0Ւ�476!Y����]s�β���Do}m+jg�$�)YAG�K��NO�g���Kʅ*ک�"���aSI����{����f{"F���R��Z����F�U�z��לe��	O?�[d%����?#��% 1=��/�����Ie;�Y0�<�.B���I�&���ʫ$e��&R�1�UO�B~vR��ۚ�� m_��O!��dOH�� ���m��o"�g�����u�C���JRJN��dB�8�v<%�F B����J��F�f�碳� J�$ٚ���&���{lB��jDŴy�.iE��<4".DSq�p�	պ�J�U��wiI*Љ��R�5VP�liН;��@Y$�ϰiE?=�����pzcS�qߨ���i^R��^��V���D_m���`zB����ڶ�r���j�&�$���NeZ��G^Yj�1�d2���+:�¬� �����Ri�����'#1,�(N�X�2�~�<I���bX��D�ڵ=4�g�8����h��(���@O�#�Qia��%YYƈ��aKWix�g�2<a��:`��t
�~b�Z���D�M
���(Yd�E�9�'����OU�52���;�y��p8K�^�}��iU%���f�a�T�Q���2#­|@�1� �Ӻ�m�Y%���r����9�&1$J
=fY�IrZj���uy���n��aN*Ն��#�]�֎�-�˟^��?	���LCw�����W�_[���ܗ�y������E����64��1����;x�ڍ�hC:�V�qYPGg���Ղ��)O�,1PTRe^��3!^�q�䤈�,��f�أ�ʔ��{����USڔ��y�����WPqK� �=Tн���H<4�� <��E|]�Z�u0<YnK���i�ڋ��x�zd@���܌s�q���k�����4NE�N����R��L�F�KL�1��	��4�,��Fg�}��y�m%�Z3�mi���(,������J��MJ2)>f$:B�҄^����!�����N��sؖ��dw)��I?�E������S��Պn�oa��&&2����)�l	��������<��3����x��*fX=��فOv<��l�nGyp�,��P{`6���̞�9ӗ���гx��?�����}d?=��
7V������^�<�����Ə���"D/{�g����j���CIG4��\B:r���f���H�*�y�2L��N�9A��t�x�W$�>	�����6�C�1����k��O9�C>�����h��x��4�T�T��Xn������-�Zܷj��2� I�s������yIq	zyM*0��mje��Y�{ZYQAs"e�<��߸?�������0"#:&�Ȇ�����7�|����Β����:{��5!�I$M�����|"�S�]F�1]�6�ϒ|����K.��7_�[�.`F�(��ek{֜���[�9蝥}��r��W���������}rl���$>��F�'��.Kx{�{�L�^�2@!�]NN��%��Y"�[�dS��2�D�K �A�zt䩺�����(��HJ������/�
�cO��u�(cƢs��78�BO����!ۄ��ӋO��`��K�~�:A�D��k3�!%-sg������?} 3j���X�0:�i�7�z!1z��D�[�<��_�b9�?����y�rH��Y�ԧt�全�����NaYȓ��`O���f<���G��T��-EM;q������OFSS�y=AuI
����{���܋���(�/�p���RnFE7�`�����)���./�6�=�|��>"DH��!�BeQ֝v����㝕����W�EUO�5	�ǟxºF����#����r�Whl��9:&�_�l^��^n��6'������Gݫ7�|��0�*z�Y����sχ���ǎ �塳J6M"�6�q���M8��-M��4�i k(A�5�x��7��O<B�ic�#��\`<���l�^������dJ�	��AR�r��(v�35�xT��E�ڮ���M�c���!ģ�T��civ��.;=��KR�D�����r;f�_���#=������+�i�O�3O��k�y3���������x�fb�\b�vx���P�(ʲ����v�����PIR눢�)�M�\�ko���{�^y�2IR�v�S�M= ᮨ�������(IX.�6q^�t%ν�2r��k�],wJ�&���m��ΥW�ì����O��at�^.���PQQ���`ͪ��$�%�v�yѮ�l��0��WY����"	���;h��gL/�g<�Ľ�N���r�6��Y���[�b� [��i�^�:TO���8k�R�H��#�|�W���g?�!��ѣ���bن�X��\��)������y�b�ר*��|ʔ��{�=k��t�E�η�\�lmo3���-E���OF��g]�W�E4[�H���5-Ʋ���ۧ�R�I�d��6L� %(�jg�С}�eG�w,0��+�ш�EiY�ـE!����fFTDY���#�d�&��:ty��G�'9���~MJJ�!��g���3��&��55ڃ���˰�;g�JSPC�T+<B�1f2�m<Ϧ���
e 2�s1}�\���Z���c"����.e<�j��a|�?E'����~���x	����{!�Ph�އ��C��Ko6�Nĝ�閻b;��ӏ���EqI�io:��㪶o5әHč��6S���[q�闢������x���8��z���R-ߎn;t�nt#w�`媓�f��&��NR\�_b�+V�2�������3�0. G�tѦ�ɻ�,�)C'R����<��s_�0֝~��B*�d;x�Z[�ͰD��{�2�!Q���ݖ-�X�럿�m�y�!��NF(���ȴ<���4��;�X$?�g��-�W��n�kX�},`�G!�S�T�4�M��4��4�@V��~Dg؀��x"}�L��
��v$������0?#�f&	���8ܱ��폋M�M���7	��E�S��{����Su����j�q�4�f뷷�h�u�:Ɂ��L)�n�����8�����N�����a
2r�Kx�?>��"13��h
�z0g�b|��cT��IH�f���p�TW"22J�Յ�8�?���7*N��é���6,^��9�&7�6��$t�v��-%�i Icd����4y�d�eų,�?��$�^�����r����2ܻ3�`iI�9]B<L��0w�b��1�'㫥����6��C�$��Y�1�V�X&Ԋb���v(U�UE:M�?��H�U+C~^B���X����ԡ��d<��5���g��{VQU�9�fc��Eh�1+âyf5��(&��e�����ub���A��Qb�����E�O�י���h��m"h==��I�N���Ǜm���"TUV�ȡ#&�����6�hT�[{�z�fL4����gJB�8jSz��2�Q��m�3�!JS����r&"�4��6����vUlu3���'���	#�E�K�H����2�bf�gl8��V� �k�XR }$Z��$�S�x2���W_Bݱ�<�Gy0�p��Xw��<�v�㑄�YVV�y>�̌�ք�ч��Ȧv�%^]t�զ�Zɰ������5`��إN��T�v4��Q�X��wԙ��(���ճ'������>M2yF�T�)�	��o /��t��z�<�w����a��P2�⃼�T��/� ]{ݕ4�!o��G�t�b[����'����b�L9�'�����3���	�����ߒ�.µ��@5�Fhuo"������I6�&���/ei[��F�����hk��CYF(���Q��O*#A��	�Lv��V��/��\\y��6�0����W>�V�q��n�G���
^�3�Z\}-�)at���/Y�o�c�G��x`�F9�c-�e�ؒ�������f	.��>I�]�z2� g ���+��j~[KvN�
��۹u��«�2����N"�=xt�G��_����l�dN�8��Ӂ�|[^߆K����"����?+�7��Y�/~x�z�z�����ol�Eմ���?�ͷ^����{�MĲ=�FxS��6ޘ�o������=ĸ����ZA_w���g��o���=�4t�t��@�k�c��W9'^|�14=@�ы��5Vm>�>��D���_|b�1���M��E��ô�b<��_��[�9�����H��ۯ����}�s*�q�7�C��[�k:P�����w��W�I(���d�[����k�>���{�_=��r:�6#��#>�ނ<|�����;�HR��Usx�q`�^�{�=���_��g�@���� U��J��3��Z'��jp�X�
�̘z�Q� ��n�����(��P��?}���R����0z0ov�x?؈+���ϩ�)i��,��(ǚ���+x�O�b��i()t5!�{���=س�^|������g��j�KJ��V�]u��ԙjT�����/H
'�W�:���{�2��X&�����N�2�3�H}M?��=ن+�U�UW��7�0���sk��N�4J�NbXUV�������f/[�(�*�jXo��/=�׹����cZe1�`�S�#������oY/�B�
,jK�Jw�'?��x���?l䭄���hj�?��Ω!QNE�1q!�67;/=�$���G�7�d�-|r�t4�a����� �j&����h"��e�����x����[:�`(���m>�-:ۛ�Ir1�W]��3�� �*J��/Hl����\s:���>�L2�����~���S���ɳR�
�����o�k�4ّj߭�
�CeQf�(����￉����g<�G�M�_Ww/>�.�c����M4�5�2�2��9_8�3���;�0o���F���\HN�F�g���L&�q�W�ž=;p�iy�1B���[L(XGn���/ҨSm�ԑ���x���!4*Dc� ��'?Ư~�#F�<��*�ظe�<��v�e�vЕa��5"�vN�B��ɡ��SŶ�MΙ���b�r:���:aC ��W�Om��j�1Qχ
>�J
����`e�&o�7�^X���o��15�ɑ$d�sN���ن�"/&�L����ư�#Ņ�����v;| �j���S1�?l�L����lz��0֮\E���n��i�;ﾁ�.��!?hZ�%�n#�Y���K�ܣ�0f��ۈ}_oz������2����\��۷~h]����k���v
F'T�B��(v���/��͗\`0ғ�� �k���̬\���m(-��@�y���y��|�/]{��0�HpxKJK��/V�p�)�Z,)�e%!I��!h��Ҍ�#G1�I�� nt���[ǥE�Jժ����!D��6��������'�vX;�'���˯��¼�.f׽9n��I��<(%�w��;�\B�Q��#yzA#��z�֔�NM ��&����Ä��;:�֖7q�Wn1���t&D�4�,��<u�Ö��ۘ=vL*XL�cq�)񃩢����x֖��T~��555�;w&� ֬YeJp: o��VbI5�l0�G6ayI����&4����b��Zh��zV�_D^�
F�I���H����R''�A�LF�ښr�ۮ=�<k��d�Xh�����0=g�v'��:�Ju(\�+M�f������a�����J�Xf��̨%e>*MB�
�ʓ]i���M�ڑ���Ho_?V,�M����� ('-�^mxCqy:w��ܲt,�|���ۈ��^z�v��WTR֨��������m���H``���FFR���.�=��Y�b^��,/) ��@J%)K#���=��G���ٳgы�ޏB�`-���6���U2����=q y���Y���$-��'޻��e��ٜpQa��8�	��H�σ¢L���;F�G�~~f�� \4�@0Q؂C)]'�����=�����1)r��HVR<����M�E���R&G5��9��l���H��6X6>nI�ى�Oi��|�$��NuD�ZEb�)�-?�!��#��. �� =�ǶTj!x�7/$jM�aKA���σOIH�K*��hh�|����ɋ��T��U<�p"�Xd�H�gM���{0���\�۽Ϟޥ�Q��,ے-�mܰ�Ml8�NN �ܛ�Óܜ�=i$�%��Bq�E6.�-�꽎F�{������_kK&�	���<��Z������SgX����i��S�*���N���LSKu&�,$�ABR�"�PB��Ī�l68�ϐbD�p&k
�*ӱ��X������e����q�#���Fqy���^�k�B��Tc}�$z4RUU��]##L��R;Zdi�Rj �ʂ)�<@�� �|��j�"z�z$�#J�!X�h�JI"m���U����(!�Χ�c�$��j
š$�s2���[T�67�6���,���n��˓� n�&�U�Y33��G��h~լ�MF� ��va='��"U�+*����#�kW��Tք���N$�tG�g6�th�zs�.�`��5��'ׅd��o[3��){���7�h�4�.��B�t1a� M�#����9b����6�F����[W���	�cƦR驐X�Q���<2=H6T"Q44�)˖.� t�x&Tʧ3*C�$.�I�&Yǩ2n_D/I�E�x]��*�������Q%9:>D�W����K��U�z��?�8������PD�����f��J2�j�9�ͽ�%J�06ɢ���3�0>>�~P���R)�ɼ̹�RT'��Pҍ�Mʲ�wѩ�V�[�`1;��v���̛������JR�\��454HT	���EF�L�O��=�����3�Ѡ�G�7e�1�9xP��mmk㡻T���U�!{���-�m��əs�Jݦ�`l:�!.[���:<ud[��,�푖�z%�Z�7@{(�J������R��Q"���ֽS�795M��f�%���X�ae*��pTl)���h&C@������m}��YЏ���/Y�&�캈9z�	�� ���C�$�x��ߤ��tC�fH�isC!���ѽ�裏*��I(���2G)��RV�&HHZ����5W��5A�s,؛�����)o�xE	�)-�+t,\ ��ƃ'�,GX�d�:}!��U���pLU\���E258���D
�DÌ!'�%ɌLI@?3�u��I��drT
�Mj�l��z٥�P�P&<2<IF��|202���#�^�!=�0J	u9��П�,������bjeLͬ��(�Q����U�4�e��E;{���w�u����}K�k*��͛eh��,���Q�}�n�I�<$��pB���<�B�E�>HG1�>LA��Wm])�u�4q�l�w���5J%���/<�Y�պ�ɹ�jo3+ �RI�G�/jv��|W�]1����A~�A�1F�}��)�6� ��j h���6� W�Y~􄃠A+�x��f����w�W�h���T*��U��|�3*��OO��HP[���{��I2�42?�rVy�U�]*��S��h�N:+���;;;��Ӈ9TYU�7+�T��>��r���R�,\�I�Jy���*y:�Mת�ꐡ�	¶�y|L���e+V�m�9�BZz�3{���+�(��GZU�C*�KA�Q�N�ǧ>���/[�\#��엧����P� ,�޺�rY��2Y�v5zc� p�cJl�_]}�:"�TI��{����,�4X� ���ʵk�$�\�ֶ���Ò�K��w= ?����^3�s$��J��/]��K��%���EZ���O-R���+(Y�A�ܼI�~�Ie�n�2����u��U�M�ġEbD�F͘>��;n��?�N&I�E���GN�����Mf!t���ibOy<��=,�5�D�	���Vٳ�+Eׯ�(�����oPϳ^�~{����*�7��G�Q����-��aZO6?%{R��"{�r�w���8�%'�
|^�*t�*0��ӽ�z�����_P�ʨ���9�����I�H��E%�=CJ4�D_����덊���u�^!�9 \(�0|��$ܥ�,+g0��[na��MJj���4���.���ݧdnzN�,�"{�����	�(�������m����v�N��)��T.���H�o�*�P3bq5	�V[g������%�:dy�*��q�d��e��ﾇ�״�Z�Jl`���heD�SM�+��Ns99t`�:�SRS��_m��^�N6nڪڠRטP��"�
jz0j&����7��`��W$��Sͭ�2ܽw~H~�OȂ�&Ր=�Db6�Ax���k䲕��w��ġ��B��M��ֆz���6���|n:��7#G�f�(�V�Y%�7nb}~T 9���g���0+�}���m�߭f�<!0�e��-��ʙe��C��e��[ rIp���'�����{�[ϵJ�v�vۍ�/j֌�\Q�W�3���ɧ�R5F����-����ɣ�q�e,C_�f����[Ș�ش�_��Y��7�Mi� �4���0��2�oALӍ�"m`�M'&��� ��g�/W���e�b1���jJ  `�����S��p�ͦ+�06=6:I`�\V���}DJ��ՙ�MRIX��9�:$7�_֮٬Ri�ݔ�]'U-m�2�����a�E5�\R�r�����KK�����(�Չ��K�ՊY]C�J�>����ʉ�g ҕ����;／&���Pƙ�`4�0"d�ơ�u@(A]c(�w�M�ɕW�S�E��QILԊ ��S�֎V�=?�&�W}��8�=h��^�\V.],���t A�dVd{U���8�Jh�G3=�#~��mٲ��2JB�0�i��fi��&V,
� U!8�T��d���r�>�:�����yZ��IKcC���ˬ�;Y5_���.gt.��L�z�<��22����ʈ����������ɢ���{8x<�-� ����g)�э#�C�}�xP��ti�0J�e�@;��7�a&_�XC2i��,���%3�ިf������� hL�lHZlN%�=���cL���R7@L	��=��jF�,�f���26�g�U����w$y*����"{:3�-.�������A�c���%��i5_<2	�͆9z줙L8e����E�a�����bT��'䡣��&O�T���B�����0JWM1��8�PҌ���I%���F>Si1�/S�V;t��E�&�qG_w1������s a�����545�	a�0[�𡣲��W��cK�Gԉ�&�0wQCЁ�^3҉MDL�Ç��fޭL�+A���v��Y'��Jo����9��C �%r��7-mif �<#G7�t=+e]�Z�|>|�>W(X!����\��x=�׍�IW�aj�5��S[đ�%�P��~��:�f3�:*qf����� 4`eD�����/2��a��˚��b�K��w� -`�f��&ª]1sT�T^2#�b�6]KI��R�������M���+#��8%��Si���^y��%�:�������{jU�b` AN�AU("N`��<��S�'�H*��z9r +�yr��[a��+�DL�P�ׇZ��]^{�Yy{��J�%ּ ��aӕ��oP��w(�:s�(�˩�Gާ��ɋϿ(�g�2���l��Fٰ�j59<D�ce��Z�74���ex�G����G�S����JOhM �]�e3˨Q<��O���~����'�`d��`3C*��_�O�@���͋�%���ꄶ��|���O}�TV�D������r����=w? 纆Xڍ�xu�@�C����=�3�9	!P؉�{�k�QG�.ֳ���e�V%��#Q]gL��N���_�z���FD=�ʮwv*sn0���'Acz��bN�?�D_�<�[z�w2`�d<�q��%ұl�:��!�=�b�Z�鶣��)�ij�6llh��e:q�K.�4қU���.��lܴAFa��F��_��|����^�<k�Ϟ?%�,ӳ����wd��eAs������0X�/5�z;�)�/�P�b�u��֩�ܧ�3+u��t�; �=G���!�*��=�TQ��uJ~�O'�,�C�M�*u��g*�u#J�66���ʏ����ׄɌbgVU4ɨj�o<��rǝ�˒��T�^���{���T:qP��ͯKk�<5���QuB'�;��gGdR%�ͷ��BD8���Ѣ�qd�O������Vb�I���;XK��'�����������c�u=* � G��/Y���&�K1��!У��z�A��_~E�,_$'O�UӢ��@~�G^z�yy��g��	s�fuo��NN	W���9�'�E5W�|���1�<77�kp�Uwg'q�jnݼ���U�gCC#�³O���=�}D����TWp2���Ӳdi����vy��(-Q�*VF�U�業`ƣ��sOȽ����kX5�A����
EQ^��M�O)�bAZ��A���5��L#�]�Ϙ��Ob�)��������-�S��s錠RkNl-p2�@[�h�|�O��*�k_�m��CT-��.�������\�RRb񩭯�-n�^�;{�]uN#25�pe�L�M�[�=�nd|rD���+�I���)%�0ofh�L����wr�=�H�ج44/"���؀�(1y{ǋ�PdRqm4��Qj%]9x`�Wę�H��J;@����e	z�W�L0�U��5�!�����/��ˤ��͔�)����SO��ħGU�;)���쏩�<�5(�ʇ�j:�z�Ⲁk�o��[o�cR ˜"rh6*j��ᐼ���j�4� �Ӫ:�,����Nd�+y�E�J����P󵶒�(�_�$�l-E4}
����}!���j�'�2��&�V˾=��_QW�� rH����8佽;�\��S)�V�n����VQ5�����*�p�6�M>�۳K����$�Sl��,fQ %����zkW1�K8�J'�,bo��0��&�i���L���a"It�]?p��?@���E�j# �m:<0.}=���m^�mNUܤ���+��\)I=H����~A���R\�"?)����-�R�JB������RɂA���z���V�,Ɇ��Ɏ�vɶ�*�[/�)�d�5���/=-M�a�8��(���%��P��HMeP��#7o��KWI\���PN="ݧ�l�\p��*-=e���9����ޕ?4O�p�Q�4hp�����U��	J��tR!��e�V�_y�M���[e6��D;t��I�!�N[�i�[����gN��"
�o��o�g���c#��7_U�>LL�&����R��_�/=�g�{(����Ԡf�w��8��31�nql��A�,�������Ï|BM�!�f�#G�ʹ3�Uۇ�����5� ��2�CVF}r��Qi[�X�x��yq�7bP�7������V���B�ݐ�����s����s�Y����BT�,��]n��j�������� &��
B{����ۂ�A�6�/����@o~��vݧ�<�C7?*�z(�u-���d��wd�:Ic#3�TWI��p\�~j�����f�!�^�@N�t�{��!gϝ����&���3AgaZ \��x�U��j��$70L�3j&,,�٩��㌫@ K@
t��Orj:�1����'��$�����)��0;�'�E!_D)"��]��%TQ!�Ϟ��a>��P���M/0)��!��~O8 ��jUf>%�Y����`w/�M5ڱw���f |�~�i�5Rp|z�ɯs��ōp�:�+Fe�L���5��G^?}������2p�p�`O���
cmQf�gl.���O��X�-V�%���x����Jk�g�f8[�=��&Tc�6��D�r� /�&�̌�kxF�&&�:Z���-Wo�HF���B��� �;"o0�1"�K���$9�ΰV�@�
���ϰ�À�yO�B �d�|>pɌ����Tjvx�?�~����HH�ޮ�9;4J�fP�nZ�� �t�H���[m̚���%�R���@��ͧS20��J*��:b�E�j�D�JLJ��c�J0��v�����C�uFeb�>-�s%�g�k�#>�O�A9t|P�%�
�L&��?1�z�bM3Nu�fd��i�Y �*A�[Q�� .uP���X�!n��;��l&�v�S��u�|��A�K&�dEn\ttdB��ODp������&����M����`?�s i./0ΏqO��������0��C��U�P�@�i�������YSF�(���(�d$Kr0	� 3�@����6lk��Z�2�
�cu��Դ��Iʯ�������Va0VQnг��0�d��b0E�ʌ�/�cy��o���9o#���U35 ;w���M�l3��e0J0�h��1C�0��of%�ds�����`��t��D�е�.NGTq�\:�r�K��҉H$����8p���sg��5�l�kL�DS����v��*��\%7�x�����r��W�94,]tD�����,��._�x�J��G��)�1�YU��9H�<��
@�v�E26�Z�XM�Rt{զ�Q:!�;�2y��?RS`L�'��7�%5G���70'd!��|�JW��5�͓��	�)!E	A}����2?"~%֣'O�#�e���F\l�Qb(G,1���V�w��N�PJ��wzbJ�����$ e!����>(���g�)Q2�b0�p������z h2����r�-�~H�����D�6G5��X��	���j�^���l�F���M�qD�j��]�l�l�YՀbA���	�1�{Эu֫=��sAV�{8>6���[�T����:�L*z���M��߶@ͻ�f\��J�>˱�d��:�Gl�K3D�
WhN6�c2��!���NR}��<QE،cU��e,9���I���tS�yMMN��dI0�'��Qd*;d�ڵ�Z�R�������J��/ɪ�R]k��H�LM�u�*��n'��e�����R�#<D574�H�[��I�H$�*%*i^���OJL�����#ʖ��[���q�����ڲ��tƽF�Ɗ*�J�9���d�שI���>u�����m�|�s�+����R�DՊ\�2�f�_����t��;>�l���� a�"��~���/�>K"7{l1�&�*��*$�}��_?�(M�7((_���,_���#�<"��z�{�����6��|��e���j
M��1r��(a=��9����k�(s�\E�1����� �&�ԩG|��n��M��>����K"PFs�x���s�**�ifU��SK��5���o_���ٟ��t��Y]� �T����浩�S�Sg���џ��;�0wTCg�Y'o�f�j�)5������G�U�t�d/:��޾@�	 	4��G�,@dش�>d_4j!� |%0L=JV��~�VM}Pekk�o����[�|�)��U%��,������c�=Fb@���(�Us�[>���)n$�?�<��n��n�U���V۳�2J)Ƃ��F_w�M��K�ʱc�U�֑�**�UDu7Ȃ�K���!L���cSҺ��~��nd?��3�T:����0l$��}�A���;�O5�#)р0u�5��l�<��y���	U[��8���n����HT��j�V�j�C��B4��}���~I��տ �v,]̈$1�0�qyt����v�����qj|L�������f)|��1�DʠH�XA6_�En����g�=����G��~��!!LLN��J @u�TM�G?!���w���H�2ΐ�C��d��7]�(VZM#�24� v`Z2���������Y]��E*YԽR�k�<��do��L�� �cFDP�WI��k�ɫ��̞��I���1>1#m��>	~����;��V�����Tfh�窩��犬q��' ��,�zn
�~VF�'�B�4�9p`���]^�����~���;�"�"��]NG�@:O�.]v���W�����=�tV���eA�fRc�"�)'C�)uX�%�~U��]3�0+��[�f�t,Yav�Mq���wI7�3��1��^YۻVN�>�C\�j����.�VI1�0m�aw��N.�X(��r�6�-��������ÌouM-mz0�8ly$}Pǃa#K�������d���W�������a�@�9G}��p�y6o���BP�j���5@������Q!����(�����|��Y�%�0W�p�6��I�ɘLA�9iz���_�[>�a�u��o��m������q��jeD�R�JG( <�
�]���cB0�`v-X����`��>�N��(���o��D��p�G~�>�I@�(�Y���)�N5={{�3�"��dMQ&�h¹�Jc���$8�3��B��FeK�Y�5?�F��O7͋��-7�&��{�`oy��La%>,��(�&�m�jv.�I�����%@�/H�7 [LN'uC��HUs�C
�>75��%ϥ�)���A6^q�;��(�k�	�s��6�~���!�R�%��%˥}�B,"�3<6.��@]t����Q��8����y�a�fY�t�� �i�v�
��	*�j(��{|��:��V�\#+V��-X������`,z3p0(�CB,ɥڂ-�J�����@�VOҘ����3�{|�?s_��GG[cC3�����W�
��${�yO"��g��2�<5�,�y�G��[[�h��2��+��p����n��֊g��� �_D$.�#x��PtI�D����<<�;��_(�u�0qhvր ��FÄO34dN%FG��f����;�Y��J2��0h����nw�I!���M��Y��]	�{�yx5~]hҨԝ��kU	<@�l.W�`HmC=��\�R�����H\�8
�����Q�sv����H�|fv� ��0#�2�XH�AJ�3�,����x����$Q��UՈ>�Ԭ�� >w&����G�%G� �B@(ky`B$Ri��q���[FGk�� &�`M]�Aϗ�u�'N��}���Fh�4Q�3�-�RD�@��5 �~M��x�s��f2���c6��� �Y]?�
�� $�������aqN��bE/���9j��"B��aL���!(�#�n��p��4�yP皰+%>�{�07�]1%	Ql�������`Ϻ{��oU�5|��̽t��Ē!��.BàtJ&���w����e�x�Q#�%1BN����&��jd���@��2�U�A���aJ�z�kP������ǒ씩S���e<�Jqp@m��$'��؞?6"8�FU�����	 ��N����q�0��qe<Ē����"T��Q{�v���֚�`�BPm�@� ;��z ��,5Nq���#0�]#��0�� ���IxE�h�8AX�
�^��81>N�ճI+�@�E����w���'�P�T����I&`a��>�a7�÷������Y�Y��T�lG��(�Ĺ��4���v�z����\��
*����(s�b�:�,�@�D},"N�,��S��`��Du3�����&�(Z�+OU��Ŕ^�8>Eg���)$�2��7V�f3�R]�a(\z�&�RM�w�D���j���ly,���pF��!��z�w�� �A��nR�i���� ���u5�ah9D`6 ��`�*�VC���1�gP�%:UsCA:[��#���@���K�Z2g͞��đHb?��^`^������G�'����٭����}=�I��~H|j-���b8L0Ըj&�m=j�є�AtX�'����IJ���r�/	�"�sb��4!�1��E�'?�vú�c!=��Q����U� �kT�>_�S�'2�^]����ա��?�*���dg2��ܥd�
���G�Q,h=��bt,�EȜ1��E�	��`�4���.���$Ϡݝ���|�R�L��p6ikTB�h4�[@q�@�)���}`����$�n�gU�aca�D����0KZ�Ŭ2��C/Y!.���*����p��Y�2\�`w�qO���u��T�T�bVh�e*1���Ą�K&��qgɪI/��>oI"Օd.�}�
�LRL�d�e���=�cw���B��LZ,Kg�<�)�L:�wD#⽠�P���rjd,��67y��*��m�k#��L��6{p�6[�bUfڵ�0�\Vd�6p^"�C�3R��ϲE�5�>bVD�i�tY�� f���4
~g��Zё��Q�a`	2��9�y��nC�Ng�8�%�ȟ����/Xg���s��>{,���g3��}�)��Q&�3-t�vD"VU��ً��
H�$R칸9�]AL��u[^R�ͦ
e´7�\?b��a�SB��فg�6��\d��񫜟��e�Y�fڟ�8L��j"�����8h�������@��ɂ���h�����ʇ�h0G`������#@c�0����s���(��S��5�a��X~w�ALr�EԊr;c�&$���0>�*j�|�AM����#h�y�g�c�߸��C��4�_@�� ���ɸ)�3�NT��,��_iaG1y\0����"�k1�.EC8W��M�����pr�#pߩa�l+JKk5#�B<�t�K��}�����5�Q�Sp؄b�nہBi@I��0��B�q�^�ep���a5^C��*�d6��>D ^e7l�m,�@N2`s @3(��GD��Ļ[�æ:X�nKA�l�)Z�\ �y\���5C'���S�b���벉�F����I��2��3�?d�/�x�p{�Ņe����S�~c�����]��4���/��6c�1`��߂�Ρ�!�{�)�J�w+c�k���6ҸdȤ\*��ۃ�Y�K�i�(DV�q��O�~k4{\dO�P�0`h4F�j�N���&����X���iZ��jN%�b$q��A()5�� { f�Q�8xζ��Qi���q=yH�,����k[b	���0v]t` ���D�CL��{@��3�A�b�[B��删"�j�NKes�"ui��)8O�:p�A�������:4 ��RF%Kڬ���|҄)�6J<�@��sZ��%�ctcT0M&o���A@��ܮ������[�""�؆&�Y�YY˴��`k��iz�Mm�A|�}����>³��� ��`��9�2����<�#Hw>�4N�0�b�G�8�bm�y�*����n�c��s��0��h1����}���3-�{��O'-	��?v	x�v��5IeeÒN?##�C�9]�n���Z�i��:���.��fX\ɘk�e��%6��Q���
�J$�~�uH���$�e��LSr�	�����h�2����"���{��=:�a5gɲ�/lb*�����bN�%��ږ"��^
�f z��.Ʌ���Y�\�����$N��F��m�_Wbc������x��0�ՠ��nXO!W�L4G�0����i��b�B�^K���D��辶�q�/Xʚ�໸��I��{�$/��Ͱ�ri���[Ʉ���D�L�t���l�x���s�fg4Hڅ����(Cǽ;;���r�J�	\Y��8d��O]�.#�}�v:<�A�4���I�:��/5S7���a��a�Z8,��n8$��Q�¢N`�9���|�Q0�M��a�rem�ʤs��&�>�4��gҍ�FR3�b�N8L���Lq�-y, �������bC��o=b�5@ =�[	s�6y�����ht.IQo���oi��r�3s�;c���!�Q0���d� hPZ�N�˄cK�d��o3eQ��zʄg4��{C��/�aU���00>�=��4��qm���tY��<]ֽ��r]t`�|���:�a2��/�H��B�A�h��Sr 8�����
�G0��`@��^b�H	,�+�*]�v� ;����Gl�x2�Y�����h֨M4�;MU��Z+Y��F.Ƽw�9�I;�S@���3@��av9-�c�n��d��&����G�� ��h1��G@�����刌�F�>´���vN�����߼!^��Ȯ�h
f]���Qފ6��.���~��8�a�21!�kEz�Y3�
���&��%���8���#�Rն�m;��\.���mk6?c�%���-�7�d�Z�:]8��y��h$��P��Hۣ��H��lʙg[M��[�IjaV�r�KW�g ���)q�r:���n �h������P[[�UG��X-�F~�#�)Ý��7Gυ�eԶ�bq��'^oy>���Y���� ��D��J�yT}E�p�~S���r�T�s���Q�!�p���HN*�b�L�{��~��yӷ�&�[�	��<��WF^�!��8����L�}�vӌhl�,�Z�s����!!��P)i���D�\��h���:;�&KN��Ŋp���g9�H���"���I�*GFl=���l9|� ?�t"��4��Ĝ���U{"����	0X���f,Jqs�!2��ꔤ>�����$�B�SC��$ijED�ް����{pc���M;����Ԅ��F8�=@�I d��I֥�.���gߞ�޻w��	���Bʲ)�������p�O� SL��I|�`���o���fc3�W&��b����h��S&!Z���4qt�dvz��;�
�E��W�\Vy��,;	!0Y�J�����!����*I���w�ҁm��u��c�DcC\�o��2k��r6�&���$�<d��E(F"�9]��/DD�U��41Q8f��ơ-4OM�#`�{�^�;�2Y>�MĎ�s���$1`0��0fM��̸�2"���� 2h �L��D�`]�M�h�>
8��mɘ�^"oX����nO#��y�`���~$�^��������*�f �j�_uEm�;��qp��2%���3{U���n��=|�k����̳�|*O���PM9�����%��03�@@���%�jUU��i]$^ ���K�ԧ��"\<\�ryс��ì�J�V	��.J�,	،�-Z!Nض��(K<X,V@�"D�7��<���5��,���(W6�T���E��M�p��s��΄�p1D�-G�p�=.k����~���<m|��|~� ��3���ޘ<����U"�A���B�pҤj��.+�b�A�`���4!qH�T2U�@�0Z�*�@�KK�Bh� �R[Žu!jXppx	��LL��v�a�PzC#)�@�A���|~	� �,�ߦ`i�$�(���k��Z3*#ސ(5JF��RY�,�`C�ң�5�!�*dP��|�����PwP˗��V�X��;v<�H$�a�����)yr���V+�AJrHH�,[��p�+��&T%f�	�R�vX�u����&�__nas3u.��,��)��9���`�$	��}��
F��IF�=@�F'pWY��LQZU����2Q��e��M��0Ȣ�P����(.;z���(���XOP*C @&a��ɆJR����P��v�!��)Y���@{U�V��`��N~-��h0��\̊��Lx��D��@B/��dh��`ޠw�ծ(�@"ѰuQR�J5*�Y\���
h�l���Jscn3�����Ř�VH��}q�\:�jX�'�` ����H(����$M�R�O{|j��|���̙N�AmS#��)��	y��=�.Q}�h�+C8���I�#���h�韦�:::�:t�x,��鉉(�Aq���\���<�a � �㝝��[��ZZI��;P�f��ܹJmi[��B�)640��c��S��7�si+��a���#G���(i@X/OX�
%	lY���@��!� �2�N0��MiA�3���Aj�9�
HU@�� ��
'��17�=X�)y0v4P,v!�R�����x�ɚ!�|�jjb� ��F�+�A�V���Y�fd��&�`�r
�ה]8�2EtxUA��Ω=�``��F Q���8x� ~x�W��a�"�c��AVς����r�F"�'�s
LBy�2���*�9f�"�Q�g����655F�Č�8�W�W����(9�Gs��*�U���F����sD	���90����Kf\�֭{�董ߞ����]�Ci_�@֬_#Y5���8��g$�t�Y��$��W�����t��%�䵗ˑ#�T�(A�j�V�~�� h����Y� (��j���"R[&�"�F� ��ۧY%�Ϟ�����\�t�[�;�\�i���Ijbz�*DII��č���A(��f�+ޛ	E5�9�ݍ"���Y�	��?O�5&������3$���&b�ɖ�H������|�4��B�$|/0$�dHW����ѹ��mbB���.�8"S4�l�{`� ���<q[[��ņ���	���t�"�n�{�]oI}C	���@��ei�p@�f�2L�����m���%f�����kxU�n�b9�M��	�_�XEs���yik_�^X�eù� y�p B����.�쮭�U��O=n6o�<*J��_?�F(��>���GX�a�`L�<�\�L#5�uR1:B,|l���/ɧ?�iv��r�n�<9|�4�կ��ɏ�ú�Ͳd�R?|�uŬ_��A�b��]n��&�ĂF!�OŔ��0q8�p`�o ���je�	�y�w������lK��f��r) ˸�	N�q2DU2gi�$sh�5���r<I�L� ����V_�<�'�,/i��Al�ʥ��$�c���Z�t�3Q��ć��	p�7`6��C/�a}(�%���#f�4����K �W�>?
x���K ? -�/د���E�����Q?;�BD�� �;�	@^F�� m�<�����>��5<D!oY�^���6�/�_ AeldH��G�
D�+(u��ֳR�/��l���&l)]���1B�Q
@ Z�z.©�O��'�廬c_ޱTv��MG��ϣ�oϞ}��s��C}@|ʡ Lr���ԜA;C#�+Uh�>�Ŧ�����PPc4H������^#�o����9³$p�B4R��(1�j8G�C%�9���(qO;�I'�T��q�#S��a�ä@�����λCR3�f���Xd��kl13�����g��!�ѫ�`�'7�	8)vk!��"��$�&@�Cw LS�(uV3��`0���u�<�F܍�z������G����6��I��lij�gN�>�}�{�u�q���^�%tZ�o�ۄ>��Jet��ggdtx\�5d�0�"��k�J��,�.�c]����{�I8��E%�f�/\-<�	Y�d{�zfx� ��|��x*(9{U8DU��ͨ@)��Bͫg�s�M���e���9R��j�ɰ�_�M���V�tN��|3�n�ܮ�{}��X�r9�%dS���jc��H��>���I�������Ɵ�<�J�e�tT�!�j��I�S��o��SM�#������%��)���׬]-�l���WX۱c�h�G��5^q�4�`������H[M�� �3s�+�k�o��U�s���
B|#�@�/�X&G�e2��,����$"�5j�2�A5,�gߞ�,�^�~=�`F1M,�A`J@kA�y�TA�&��k��4X�P(4+*�9ZI͋���L�^�N���ֆMB��D�~ۼV�3��-Xܘ��!E�9�k�V��ٹ��\�XjTc,X�P��v��z&��3c�n��N"�|'ɹ���j4OQ�| *��u_#z�,��I5�Q�hU)���2��׬S!������0AR3��K�4K� �>n���?�~fF@�����Ib�'M�@WW��_V"��XL���=����P�>�,SS齽{�����Y��N��xρ��'���L/�Jȝwޥ���8D���8N���Ɯ ��0�\�~B6_�E6n�H\Q8z�̧���ke��MR�(Ϙn�c�y��wI|���s��:�Z���Mc<ʯ�~D�<�,F�����w��a�a�@�n�z'�W_	�_���(���#��~���v�Ю��Q�`t�CP� f�]�u+��3���e�d9��
��<�L�ƍ���U�Y�{�I�m1�B��硁a��o��nذQ^Q�	9 �]�T�~Z	}VR9�S���]���+����E�4�k�g�>��1Yu�R���JP�d	n�x��P�(0���8C��<�Y8�!#*LjZ$���� �=������\�r�7�)��Z������<
��0�V._![�\i�R�dH�7�x���:TR�o�G� �@���MG���Z9����{1��A�@tسg��|�e�	��L҉�QaBY�CK���?K��	L���P�8`͜޼��{���ٱ�D���H�:���0����iU��vw�=��O���w�T��.0�0�����/���@X�Bs�&�4�#fО��s�l�|�;���Z���Q	������U�_��|3�֡��կ�A�|�?���yFͼ%RS]G_=!/��25N�h�?0_<��[W_�&Z�,h��	; �����^jȅ3ҳt�j�5S�1�p�J�^R�o�=�g�T�A{��~�5�r�-S��'/�FG��-I,��:���$��s�].���o����7e�[o���po��G{#��6�&Y,��X�wȡ�����3'�mP�p��w�ɽ��8�u��!���ۃ������7��2��zp��C�����]�vɻ�w������5K +o١��٢&ǜ��l���Z)��5=����l��������>��0��6mb�s��l�Y9y�#��6l"�<u�<�ρV 3B�A����$Г'O�`�<��7~oW~���O�-��N��ň��\��Ѭ �B�P�>?��S��]4�p��2����!����r���*]1���A� &vù�Ȏ�%t���{d�޽ A��;Ьb�?��z��v��ۮ�^�\��	p2`Z�Ͱ �߫Z���O ]C��߿W���3Ǐ�y��۷o'b��`~�&� ��U�Mf%�F���(��w_���埾�-��3� ��x�|`������O��u��I�ɳ`b({�P~������{�e��,`���d�]��Q��Q��"ygכ�z�Je�&��C�����8cj{4 ?�i�K	�v}M�n���DC� ���>��m����)�}�~9q�$���p�����քJ"�T�@�0&\եz��t����ٳJhQ���d|d��F���ˊ�Ketd������k�:�D�� TP�
�����<LdF�����㍷����˗ɧ�q��;���LR̫	�������˖�qzb�N3��P�Tg/����x�@�7�x#qQ���E�+� S��2���+/�Ë����:��De�WH�n�x�~`0h$�@���#��t�"�� ����hb�V�ZM�	{G�4s�U�7_��*�{��ɷ��M2¤�u�|�Y=7���`$.����8��ڽH6�ō�΢A�����0�:T�]��C\���ƨ�������*3�*����x\�b��%?�R"�3P4�,q�~��E�p�~]@�8�=*ж��T�N�ا�]��(M<��� Ã��L�Cў�����i%�Ԥ�d�zp�v,����c���0v���z�
�|�F6�#���#_%;T:���<$�pį�bL��nrX�!K鉃��ȜUO
�TL�L(s��C=$_��_���GeJ&w��� Ni[�R�Q� �Z�j�|�Pg�5&��m`ZAZa~ ��]w��P��>+�}�$z$瀅��|�E}X�}�H����s�<��(Q����A�,^��C����W��o��'y@�'0܏R7n��0�����$x${�32�?���[�r)%?��˕`���%8�Q� ��Z�'z�AQ%�~�"(�y���W��[Y���`�Wo-q�N��$�RB;�������0�$����o��
���n��N�Ǐ�	ݛf5i�*�'�{d�l��nY�Rf�)Y�q����
�R��t��"#s>_D^u��8z� q��R�|�T�@w��{:9�n��g����k�[����h��!Zݩ7����)7��g��_��&�Tw�����6o��%|�R1�Ü~a; W ��][[���Jr��?�j�=�&��-|�y�8�o��LT��={XJ��������L���� i�>w�<�����a�����'��	Y��U֨m���x�BS��5 �:ϝa���]]ݬÇ��4�^`���!�BF��Y��׾�U���+�F��e"(#�H6�3���uݺ��7�4A�(����"� s��d`����h��p��ٟ��Ҧq����X�K�Z�x�w�/x�sʸ�-�~��B0=#���C{��A6�]'��Z�����V	�����d��v%�S�� ��xl�K���.4��JM�ljFz��3�ߓ�5!�:$�JK:1Ǯ�Z=��T��x�;�R-���2I��!._-�%��m�L�fU�2�����T�L�����p�ѡW_Y/�_������*�L�U�iR�ת��
�&m_#�}���wߛQӨ������#��a�}��r����|aͳI�4cϐ�M�4�*J�1i�9�Ub*}W�X�6�:��|�A|��a6��ɡ#�eD��i����_�n��;��ww�~L�UV3�ٔ'$9�ddt����F��7����A�x�G���Ѷ��@�
�� ;���Laf��qk�\FBZ�z��ۿ�lCB��'��8>�O�ɨ�[:�Rmr�},�FT���<�d�}{ޓ���4�~�]mu$��z�M���w�D�y8<2F?����1�P-R$�ü��K/��>�"�P�bt�A��WS��]��B���|���舃i8>1�*V�C�`��ĕh�U�ի�Գ�c��*���M21��;'�j߇���U�{��ȫ��>!��O}�q���X����]H�����rG�4o!� @FGGh�Q?��nf���_�T�����F&��+١��1�ׯ�c=	 ��/�ڤ^�Yƽ{�����e s�덑L(��� Ke��J6���*��W�#)΢K�:F.�����|�����!�V���/��A�6�7�*d��Ң>�;ＣN�jT;��!����9B1�ؘ~T;7H��s��]g��>P$m�-�Q3����y�,��=���:r�0c���*�!�Y��Ε� �Y�&õ�^���η�R�e�?|�L
��)�����@��z���9Y���d�QJM`�hP�O�1��t��1"�+�B��X�̹NN�?����KF��R��c�	��[x}N�n�U�^����lN�BQ�N����h�i���bN}�ʒD*��s�y)�U74I��f!���g3R�Gw���3$�y�T���� =��j���y3��/�e`{KqP쉵��>G��Ynw���kbο�����=����b@X������au#���x��EB f�~f�"��(�*��&�H��f{��E�ٲ֥�Z��G����
�ϐ2ޠJ��J�Q���aUI���mAU�M(F�6��@;!˜PIsl߁�dd|�0,�0ӯ�&Î?e����I�t2Ni�IH�믿��&�� P�#�L���$Fh���7��!��i�)ͦ��l Q���'%d��DyY%7�FϢ�e�J2�j�_ �����\ ۹쵁�qR#�<E�54Jlf�IK���<�ك����)gՉF��YM104���"�}
�7��̪���D�º3���Qm�)��W�\	8�8�*��jħ������52���ϟ���C�9���tL�����,kB�j
�~QF2k��M�N�Ȑ���������0;QVtxC�FXض���/O{R�s�P.׍`�{��ZLh���U��&jQm�dT���H�T
e�G'�ȡ��4|��]4��h4-�*�0ѓ�Q�W.�`4䊫������Ij�-�g������~k���1�0�C�i�,�D�~�m�����q �[n��U�ӂ�� 0��Ĕ:f^�'PW��$��C Q���2��T��!SG}�ˤ��:j�'IX�i)���]~�ꫯH,�d��	+�'۶m#�!6��'��%=��U��y�X�`�N=���,�j�V �l5X��z�*� L侘j,�0��r���w��#N�n��A��FrqI*S8|N�~N���j�n��J��G�&��ő���\n.;�ɧS�P(77;�KgJ�@�V]S�Y�~��ٌ�X(8��K5*`ԟCPX����3���A9��a���kٚ�?�������6��&���LZ2�9&I��U&;���yD����dE^�
W��=�I'p���o�#=�'��Hbv�v""4(h�gb\����O%��J�0����Q*؃ J��N�,�Y�p�"������C���ݻg?5�+@�@�\�*�3k�DQ�j��E"L B��VU�{I���P�F�馛�x����b���y�Z(�X����f��MK�,���&o�x��e�{D�uv�43i�� �60�
�ȮN���~a3h�HHF�"��D��.�׽��v�4����Z�a�.��N.�hY�2�8}5�S����R�ڳ�",ѺΝ�ܴjB��U�)FR���[��������������YhR���֭[c������IL'���������y�-��L��5��]ۮ��;ǎ����ٙ�}}�~�ף���&��U	g@u�8���h�v�RE��r0�*�����IO&��o�B��yN�uGA´lݪΜ6��=r��0��@����{��'�$�|b�w�I![��0�׭g湧��q}�p��M��ݻ�����n����ij�Gm�%ł�[�=0��#˩�� ��y�����e.A	�]ڨ�u��1J���-��C&ӑcG媭WRӢ�&
����y�>�駟�M�6��U�Y��߃����s&O8D-U]e�wb���Γ�^�N���2_jk�� zD��@�0�H��ɞ@�:(&��N��s�Q/��pQ��U`.��rπ�a@�5o|aI��klRB�s�/4J$Z��:�1�=?+��o5G�����O~��{zz��}�)��LY�/��]~���׻'N��v�r��t:�u8�c���B�:�HV�b�L.*fKn咂�盫{ᡀ�鬯������w�+����w���,: �>'�M�Jd�x�l�$��J9�c.�L]�0�gϽ�cF�n��C4�Po�I��m���uN���N�A��{ͪ�Xk� M�1��*	q<}�u*��'�ƍT�#�u�0�@��-���W�����I8$�<��SҬ�5mLSH�N�GvYƂ�6�Qm����#�����[(_�7%%Jl0ˮT3qP}\�#h2���'b�����\�m����!!1��h����O}�SԊ �-����)�9�5�6��m�1��]�T�q\N���V���̥ٸO��C*`�~(.�$s��}��j�:�-mGd_��"���t�	!�����9��ѥN۔���'~8S[�Ⱦ^\P��j%�wX�|�,loU����`ä�ͥHd�}��g�ii�ǑO ַwA3\��;ir�\?�±1Ge�~�&����������M7ʙ3g�0�6�;�DJ ����+V�`�*{@D���)�Hl!����zo7�S��G����&��%d�1�ɷ��6m�@߁&U�Ù�	�w�z��Q���}��ש)����'�R_j��8s@������}��O<-��}�}���gR�d�_|��U=f�A��Ƙm��D��E�O�p���ep޼�Ͼ���2�{lq�ҳ�B�������u �(�����\�l�8�K�T�e�5���-��wp�L<Q;���m��E�j��U�Uݥto������3�/㚝K6`�NZ%-:��j9�Y����QU簐�^|E-n3Hj�:r�U��M��b�r2ώ�ޖ7w�m�p����m��Ч&	����L�v �
��Q�M�
I�Z�38̈��K�s�� �D�+;w��߃Хe_0S���-��ǽ1����U�0%���4u����(ߞf6� Ͽ�,����7�l��� ?0����	���>K)�Yl̝��i�Y��7	~��	��^{�uٶu�`<"hp����Z]�	v�А0ˠ�.XLm��J>������}�����3޷�L����?hv	�pJ]�Y\U�D����ߕtV��q��/LW5�Ճ��j}6N���d\��c�2������b?�J �p˭�J,�2ǆ%�*��j�d�D�!S"�޵[�z��>W*��V@�L�)���p����P�
����} a�=|�w�y���a����ah���"����hU�/�LbCb��[;wH�:� BHlV�",�|9k����s�ބ^���wr
hC]�C2���<y��
��!l��7��E^ 6<4��v��I��eòc�p��Ԫy��s8�7�|�<��3���oP�$3�r���;d��5��D���o��ZȆ����zX~��%˖un��x(�qX&4�7��m�O���/�reX���TLN�:�:��Y@�����J�
(���Ff�a.q���,{м^�n""�ڿ�(/ ���c�
h�v�=� �-�!lrSF��id�R��*爑��������JX~����{Ӭ������:-�g89T� �h�A��#�L
GĊx9H\�S_��f���7#�T+bM�[8�x? h��/Qm�	������C�OX4(�-=~�����kL�K����3�+t�Z{�ܓ6����a��+��Og���@�n(�y��[���w��aƭ1D9",�@�7�c` �	!`���-���	7%2�F����["k"u�kX����'��D��n��ǝ�&sM��`���]	
�y�Ȧ$�`2@Z�-��#�2��T�446S�y���
����H�( s3��8��!�|W4�@jcmP5Pu]��$��x¬̬��߁�m;�D�S��c0��&j�h���$�p1���k?�`Zp0��C�GG�j�ʯеz���_{��I��O�p|�_�#~����!����h���jl<��$k��Uvي�u�e�6Us	�����, �v�c�@��p�H(l��Z��ք����D��A���a��UBMG�ib�v�q�lJ�����U�h$�lTd���t���86�z>̗�5�
� fD�8��2@��4Ӳh��/{�oJ1����&��cna�6|����Q�v>�n�KC0S-%j0��
��7G��Ϧ.^@�&>Q.*C�#���p(�7ɯ����ܓH&��]�Vy�[}�K�>��㪮�΢�5A7_NB�W���HO�9o������	y�ٗ�O����Ɩff"�U���i�T@xh�'Pm._Fy�Q�p�!�&��Bv #T�d�&w0~g�c�|V�Β�B��GM��� 62L��?\�:4 ���;?�S>�`�fs�=�R��>xC��_�.kf;Z�f@�vk+����/�cW��ݦ�,�	��t��q�L!3T� ����ژ��I}~E�~Ů��.u�av�e?EN&�5P�?�n�����}PU���G��#l�l2�a���i���'3���S��=��b_�ς>4�4\V6Ղ?���8l�u���`���u����A`�������e#`�'ؖ���x�x�2=��h9k8"|83^�]�4B�3�Tf� �����?"� ���e���(�ڎ"�b2��Y�)S�7~{�;6,����F�����O���9��;�W�jln>u�왼��m�`�>¿�@�Og�G{���:��٫Ծ�*^d���8G1��ћ`�8�U�*�9"�a���jxGQ""E�Dɐl�A���(3�]�?�C�9bUM Dq�J�u<(����mj�����QF��������#�e�[,��?o�6���*�E�f�E�H��3d�:��m���FD���2`d	3>�� $�UJb���yHb�B�>H��>6��p�!��=���(��NMN��}�)aWH��I�U��Z���{L�����������:#�R��Ў{�髾����q:�lI$g�ZS]W�{C�T�������T���1F�JH$��L(D�%��|=L�ڵ6�4�_	��eM����ٓ��/�Ϣ������)q�����/X&�2ٜ�"������e��e3���_���3��6���أZ��n��2C��'RI�����+��������b���H��xZ��A��#`h����X�v6�52�kpa�m@Ò����z�;��W�R�Щ�0�묷!=�9U������J0�m�6ca�/���[��ZXХ�^F_�W,:�z�(ttg��`��?p�B�����˥����A��[
�;_>�J�\1_T�_t!��0/����τr�bD��W�WfPZ�{�9%6�~'�1�LΩ�q��Ig.�se�i��`�����Q��T��J�N�[פ�,8�(qb>��W����50��qu�A�o@�{�oP�!��_��J��H{%67+�x�jc��N�8�����ئ!��%!������{C���t���;�ݴ� �����i�P���@ą���o��,�z�	z�{�^�z��Z�V$�
)-��ڝ1v&=Fq���HV����.�3�A��b	�fN&���Wq��9�c�����H�@d�7���x�#��o a��!��h���(��m��]��m�Z�*0�R�n	�F���D����{��<GY�)ڢ�����:	Q n�2
��vJ���R`_��D=�cȈ�|��H��3tV,�����6�~�`�`c��KAw��+�p��X�ڲ�-x=G����rŲ9!�h%\�(�Zk)MK,AИ�|;jZ*�i��w�m�;��.��ֺ�SL��"Q�����<?;K"�a�1�(d�k�a��	�1��MϵI���S��[��0z��V.��n���d2��[����b��,�Ӎ*��)<��H�-�cs����ǆ���x4Ƣ��z��Žz|�V�E�J�P���a����Y�N!f� �N�W*��^ r?���~�J��WW�f0]ܶ�uDD���A���'M�
鰝� ֘��1�N��Hy��H��>�Z�������Dw-�#�t'<4�l��^�jB�a!A����� �WAwTX,/�6B�ؓ�g?�~�R�u�ܳ{&� �=�=����N���=��GQXg:�^�r9}{���Ų��`,��� ���ppxBA{���m��᫪��p��8(�!� 8
���;�0^b�SY&9�\Zn5E:a~    IEND�B`�PK
     ��Z�9M/�  /�  /   images/0a03a94b-1490-4d51-a356-eaee23e4f5f0.png�PNG

   IHDR   d   �   ��<   	pHYs  �  ��+  ��IDATx��}�{�ו�{���,KF�Ifv��B�i�t�N�v:m����t
3�R�)e�&i��q��$[��������}G��p���'��{/|ߵ��2���?��������PȾ}a0 �@v�yy9��hh��W^~�W$`wؑ��	���k��1c�� l6+��L&���F#����W���x�����kL��"�;u��J$L�h�Ǥ�_>QO���yN���WB�Db�.��3���a	�u��?Q�������?qmN���M�uq�.���d�<��<>aĵh��a�a��f��j��k�������aq7n\��מ�r��m;n��)u������?!##n���0Gb�	*�����јܧ�g0�D�EJi*-���8y�&�d,	��A��|L)��R�k�7]S���~���E$]R�}4��BI����+���x��bA8BC�%`�Y(섌��1Y�M2'趢Ơ�6o�#5iRc3&d�fJ.++Y���N���`xx��Y��B<�	5������?ٽ?u����P�����_���ͯ��_�����6���{>k�X/�����.WjGi��b4�jL��Q����Ѡ�D!�M&���W��&Tc\���&6o�� kD����/�'��8��F�d��DҜ�Je ���D�*4j�W���=#���G��k5��T���U����$��x�Ƹ���AiN��r�^����C�w6+#��5N��P�
�\���_�kr��W9�a�Y$����P(4�31��U��#%�&�?���eQF�Yƕ3�ei"��hn�>UTrW�F��S�G�q]H2�7��G��=h��A�&�_��͚I/G2�)/���I+���,FW�ѼQ�:\w�v}rd}ݻ��*�4�"��:�4|~�钢��g�����=��LQ�O�'C�`(���+����hok�c!�é^���U0���é����kԅ��Q���1ݭ���LZhRyFM�b�@�ԵД4��Jr�bIf�5�h�LL�0�3�1lJq�Y�O�A~�2�+�����4�C*��1�ͦL�m�;bq]�q1�^�2DQ,CD,*��l2�<)Iy��a����p�fN�GC^	G���J����;h�͹�`�47/�����<���{v�v����i{OW׿�c	k������b(��ADU��j�a4��a=@��Q-	����Y��T��z���p#N*F����(*7�`���{S^$�ǵ����+!��I��x�R�2���4���n&��(@.jNZN�٭ؿ�?����?<�`8<��o����]!
]1dى�f����^��?:]��VW׾t钛�:;�T��e�紺\��h�z��qB�UC\�$}P=<�a!)�$K�%#4�)+TsU�P�(C0Q)��!D))���E|_R�IOS���c�"����QB��6�M���C������<5&���8,L�I�S
��G#2W���k^��X� ���d��(+p��wM���ϱ������B�%$��|����Vc(��j5������ʽ��2�jPa*#�,��&i�!����`��D]%^S��9��&�\}��ܓ�B�����8z�JBGKɰ���We2i�4�y��_ݧA�ؔb�|��^=/D��H85����>'P��M�	������│�ؔR#��r�;(7ih`� &}�p�R=���X$:�?��K/�!j�����<��������X�ਖ਼�#�鉰`!$�����LFw�%���u(�ǌ���Z,���PN�d0^V4(*�1�4�s�I�����/-$�X5���J1�@���3���_T�k�%�P�b0|�)��L�W'���W�sC�^�y����R�ۨ8��k��Lz����N���Y��݉���7��W��U拌���.G(�G����J+�plN;����)�	{��R���Z��x�!9�"����ĪO�hK����H$� Hrq}�r��s�K����@4�Jh������d_=�j���k�3��T.��dV�r=�2�ə'Fc��L(#��TH�TJ��@]���F��T���	��x'`,4dx��iK�Õ�_��?�	~��c�����j��!>2�U�ף��[���0���t�t��gZ�0Z5 1�2SlM8���$G�P
��V����iV�}�u�A�s�d]B��܄�xM��JH�9׼ͨ�x���5�j$�zƬ�M��j��(�e
J''�=�(S�ِdG�BԠ�Aa��bCh|��`0�"�q",T�+'?�B���y_z���/��ņ��+* #-=y�d��
/�����}�V�@?�Ucd��x����5mV�Xq�)�ay��Q4f�� �N���+7u��td��T�����B�I��ߛd�k�8Hz�ɤ�%m|����&�3��5Mq�xB�.�dhK�_%���Е�(o$i� rD�2������3��b&a��`P����#���vσ��_VRRV����\��vwubl��9y�,.@�ӊ��a�e!�
�x�p]�/��j!Ȣ!%�]��4�	o��j��6�$Η�ğU�M�)D]h�����Q��+qGєm���E4�jaҬ���6?����N),�<\�;����@���`L�!���X�dg���ʛ��FG'A΁3r��<khjjFWg;2R��k�x�8���xI^~!���p0���B��M�R��z�(���a�N���1]9�����)�/V
3%$�)G�qݳ�E��T	�4�&��L����=�pT��~��w��¢�5���1!����c"n/5�M����[*���W`G�����<a����Q "�YzzjN4��$
��r���N|�Fb��!
Q�|������ d�Ϝ%aKA[�نܼ>,Y92Q�^�3���+�W��tT$�ArIb�S$)&b�+�h4��B/2��D�Lh�)OL�y"��ŌU�G����eH�k����a������<Y�&�sL�eѪ%{7�x��P<��.�!q8�尘B������6�83{v����Ob���F}�@�MZ�)DU.�}��\��~�g¦be}]���x<�{���&��	�́��2q�Դt��NZO�PPH��h\�])l
�J��L�@u%����hR3k�Ob��F�aM�4?W�R%�x"*�'Y�����5��y��aɐ$�n�g�*��������¨�א�"D��&8�|�NL�3f
�֨D	@��P "��b��&>��O
Qf��mF��!���u{	��s�ph�!�_�����s{(�˕�a�HP��3����N�������'<0r�^NjbbB$�!����I=K�iu�A_��^0�Xj�'�{b��Г}��dΉ�ϾVԒ}2�$c�Z��I8ѐOL��RC3H�T����i��ٹ�Izy�JsF��!4��46�!���3B6�s
�T��gb87�4h>�å���q�jI�w�0(d��O�	�����g�t87fg��"��>!���&!%Q�nJ��^Ґ���_�:�D��u����/�/��F�I�҉TV5Щ�Ӊ]2<����	�TNJ򔘮�����
���Z�|#���� e�4 �N:��	O��[1�e�
�G9Sh�!��X"�VJ3�'fW�;�g$d�ȮJ/��i�p�m�jE� r3�#�2�N���4�}�A��9�@�U�SE<���&��Zu\+(�R�!�,G���Jh�E���8%<f$,<��Р'����UL=+Y�P!M=_}��h�֠������$��+W0:Y�L�P[��J��g�٦�¨/�)�$HMGpF����/V��%9~@��5�a�`��	:��(d��T<�^�J��2�����Q'��|j
���C������Q[^L��b\JJ����E_�0Ȥ�%JbJ�+��	�t�STm�U˺&�i��*�Qgʚ�'�
�dW��X�Z�UbzD}r�!6Ǔ��a뫅j�Pe[��J��w���8�)���J�I_ZԔ�Mlj]�  @y�Q���C�&�Sj����C�{�!�	�i4��f�6F�{�1üSG}�b��47yH}���:��|\�4�\����t����^�*"�V�'O��S?=16�R�EwK�x���k��y�T�Y�
#I�$��E��Z�|&��ص2� ��p�����|e �'���paQ�V�,@y��P��%#A"��Z_W$R:o�J���*�âx�ũ�u�`��L�e��Nz]ħ� "q�\�jKjj����c(/MG^nP����^�fb���28f��j�� �\s�z���������e1�I����(��\�-��pZ�z�H�AS�ɠ5$�ܡ�z�F�����}�Ѡ��ԓ"^�.A�`4	�<!!����~���-��}��c�b��(�8���HL�P
q��gr�&���C6Z�8|�򛄏�Y�<�+j�&�0a��bHwXq��~�]z�.�G�����B�Ӏ���x�,�2�����2����2Ջ��J���h�B��ĵɩ�HT��p.�dX��P�#�Ԡ,\ج��+�1��"5�D$&��-ZyjD-F��$jkJP"CL���E��Vς1D%h���⠁�Х��y���`�f����D�ʒ����hAr�<=%�@@�Ȭ*k��q����H̜�ݘ���[pYRd�T�E����=����Q&�+f�o���|����k6Wj�o�~%�W�!THB	*��E�yU}�ts�.c��T�0 ���,"�p����K-Q
$�Ŧ8lD���@HdL-��v�Ec�VF�|OH ����1�Fie6+Q����O��x,���NZ��D���E����1�?uii����Ay0o�jV>74���-�\�˧1$�%?I���w���J��V�/�=�;�2I���fʦ�Ǝ��ҳ���ee��
)F;��*���?�MKɄ�m�g,GZ�	�_%%Y��Be$v��"�Z8]���O�J+���4]����c��T�΄�>z�Z4��z/���#��fΚ���x�&�L�Ӏ��?ľO�����x�(���8��ۯ���������;1�a����	-�8�w7گ^��pp���ͫ�<c#r���j��ᱨb6�l��D-!�P�M�����Gg�El�҈u�7S��b�����? �'���:3��b��p82��8��{��s���`�
؋���7��͢�S�LȪPh��g%p�)����RR���C�a@iAN��@eE&�e&�,�ϋ���:�����Bzf��c�^f!g)̙��(++S����WZ�����@oO~��_�i�$�
]�>V�f�K�t^�ţo#�/���KX����ꥴ�N����i�D���<ݍG�
�5N
����K/<Gk�J(������OPZZ�gƱ��wq��G�t�Z�烗�v�(*�ǩ�0�����j"�CG� j����7 �s3���"���TN�g�`���Bd�9�ɉ~d1$�A�^�@ސ��o��a2��{��?>��lc}�C��ݷq�C��r��cX� ARǜ�F���˩�a�0rL����� RR�G~)Ce�I%����A[�f�ˣG���ӼEO�+p���҉��EFf��jK+'a�E8w�$<�p�gq@q���66�<���i��V�$nq�1As��Q��/��p��1qA��l�.�O��w��o=&��:s���$ɘ>�0-ﾽ���
�;G��ˬxB\/�|YGW
���r�:Ê��q���g�váǎ�ƹӧp��$-5�B�+��Wq<��G'$�hH&&�Bv�LѰT��f�g#5�A�l0�7��qX� #����Rk6F�p����"!�H��CZ&�Te�n;B�T&�z��4 81�:�5Q�����aT�ɉm� �	���;�>��O0TM(+;W��b�~��q�9��2a������nу�9C���I+𥳐��J�;q���t�r"�� ��%��������艃�?y�
��T&u�J���]-��2�%���ԥf�� �-\������ �z^~6���pBẲ���C�֎��4D�A�͆EK���7��6�^�7^=	�W	�spfcå��ߌX�f^{��C]³���t�F&���������Z﹣��D%DR[�(�cEI�C	�xeM�71���Q؝F�1<�B~I�tUST��B.�"Q���DUM��J·r�Z%�A_���L���7g#C�����n1��=���>df��v�̝�A��B<��o��}'��֋�|'s�,]�B����n���������ػu�fl���z��rÍ����d��Ø�d=�͢{QZ^�96��a�B�r�Z�Ϛ-$Q����3o�ŋ�-[�s�/e�"�p��V��ʵw���*T��%kQR� esB"8RS�bÝ8}����07���F}O�4���ʷ�رq4_R�HZ
=�b/3Y��#���8��[VL�"��qNY�.�ĸ~�"Wo!�֥)���*��`�<��pPeeσ�z��H�P�W���
����Hۑ�=N�t��0�򋑙�GHL.C4����:ڻi��()*8��<r���~CÃ�x\YQɤ�"�[眶2����0<4Ȑ`F���J��C�5+7o���HMe�L4��Dn%%�X�z��%Զ��hz��x���3�b�mX�$��zl�B��S�Q̙=Ki ���V+)�qw/�?A�eź�%�,@~U.
�Q�T���ZZ�2t[PS� %������� ���.�"���s����e78\�K��h
q�C�v{���~����������i��>�����v��dtU������5�/�N�z��E���.&� 6mބ���b��,}���Ge���hinAnvr�
�k������!+#k�Q ��J�@"��'���X��%+WcZ�,���C~|����@_'�I�+kp�=_�02U�F�'���h����q,�?�տg^r�z�x_~�p�de�p�d)��Zo��t�� ��{O!09
�g�^�����)"���}��Cx�g08:��!UZ:�/<��a��P>.�<��w(8�s�m�i���/��̃�V2a�|�<�TSH�9�Hb�0��]o�����ݛW�Ǣ�7%���/0d$�7�;��ҊHl����w��s���$�'���e��+r���R��>���;غy���ؘD��ދ_���P��7ɐ��΋(*��a5�#�����w��"�>!��7��%����^��S�PU��<��s��
��==Id�<�[���3����C�ً���k�����p� �өG�Fo�;�����u�%�r�W�BQz��$�����=�n���玟��ߍL��,�[�8��� ���"�J(j)W��
�Oxm������tUg��V
���0��g�G/�8�����,f�-��H3�+����������p25L�s�Y�0�2p������pv�s'��y;��]֛ǔ���S�h!!<xP+I(��J0��f.��{�[�J����cشi.���]��ɰ���9�I�?w����\b|���.F��A"/ȋ�/�ޡa��0
��k�!7݆�g��),9�;9A�G�������l}�s���>"�A�T��	I��`�u^�y�A�"Z-��'�P�0¦Z�\Zw�2N�>#�{f��EmUnҗp�6R��Hpҝ�����ƽn=��k	
k�:)��	M� �~
�DD��}��Z�q`��a|�[�D�+֭�r����~�mQι�琙�M�:���
�����ҥ�P�!�>�� +��U[*(e��!�dEz��a�L*����[o%�8F�y�����p�R�X~덛���o`7�i�*�����8��j ���|�1�QTex{:f�[B�IXl�`�����u�-,���0�B�j��u��Bo=�GP�N!���Է�gd�B��t�\22ҵ�P$bP+�*ϩM7����an�\Þ�Chmo��*�_�;�h��^Y�L4���=yN������D1�H +���޽iA����;��r"URI��0��]o�2"Zg0(���+�wێۉ����JR&,��+Wn��BL���[160��wZߒ�[�~���.\8>���p �T�ZBԹ�����q#f�ŝ[v�j�	F�(��ނچ.��\	T/�ʍ���K�D@K7��
�8lR?�6s<�����cĀ�s�b�L�#�D�������i��͚=��.�a�Q�3,4&��c���k�k(��C(��FU��C&Iv|����� t���0Yf:��^���2)�Q1}=��v�aO)`�1�;8��}�����E%��!�e��ta��B�ԠRS�d��V��"=-����i��ٙ�C>��䲗a�}�Ы��3�(/�Fww�UUU5���{p��7�J�2�IN#h�m����X�~V���08��@ϚDk�yļq̨�K/��.��y�H����Ο�8�v.�X�Y��Ĩ�TԠ�� 𣖂]�x�-h��v���&�ڞ�0h6���S�O*TedeI�BJ�+a��E]D!fU�1��z��s�Ϸ�X2����Bv�WL��A�[������5�!F
1�0uC=g��r%X�d҉R��N��-��b�Z����!����CQd��2WeA�`���`}�_R�Z��>�1.\:@���e��R
&+��������%�Ԏv/��||�{�o��!B��_���m��̨�����,M4��%��Ï�m��t��}�0x~��r,)b<����q�H�P��x�{���<�7$F�ҟ~�p`������<�$\ٕtm�_uE��m)[_VKjy�����$��Zߘ)����s�~��Kre�/�E(0��^y�d��`��)@K/����A��r�m"�A&�l���W04�֛71�'�p�X���A3y��ȐV-b�|A*���A~��	���`�ʵ1������
[q��i<���1�~���}4��GTbA>���˧��s�ǧ�2b� >x�5\a�Ia޳�������l3���e)�α^9GR���j\h����<����+��K$����3�ɧ���z��:v��i����[����iT3�b���ػ��N�	h�]��&�S����e�ج�K��ե�������á�N~��k��jT/-��!��U 0�v����LCԚ���s0x܌{|�#B�������WK���`/*�U�,f �詣�==�(�˓Ҋ�q����R��?z��Ê��I����	�%06�;�&�s^ڮ��ڮ� dMK1�G�����{)����f�����"D���K-4��)���+Dq1Zk �#D���ΞV������������n�ݙ�Zzƈ{�H\u�`xl\[oW�i��n�3�O�yA�MV��bx��d��4���-�	Y�p̣ҍc�H~Q�U�!j�m,��y=�P���R[����P}(/4��H`2aA�d�x����48H�NԔ��d[��v�Ot�wލ��3�L�r��eBh���`h9�q��t���sX�d��U�**����ḇV�y��Б�	�ՅȺ�4�)�1���QA���Җ�ge)W�� ����Q��T�w݆[��܆h��GqW
�m� ۧ����;w@4^�v�"?X�h����F�-�7��f2oQ(����a�
��ɏ��R5��"K����;�>��l6�U5���6F�h�C��D������Åŵ0��$��pv]w/6�����k��JG��Ay�"vt��C�S��Ӧ�[71�nN���7I��{�Y�"���t�2�H�m����"|��M[oi�����㮇gXL��b��hk�&L$�	b΂UX�d5�o�%UX�~;N;(Ž��q-�A�I���Y�5[&p��	i�X�l5s�v��F��J�7���;u����m1���&]*q�����Yz�A+��Ō�	��RAs�,B����t3y��PQ3��@��x�l\�g�UՄ��O����JVۮ�ҍ��7Q��B�R0]�a^1|���W��K�v1�����bu�f�p7҈�
Kʩ�(��=����sg��ee�
+�I�g��Nl�%�O�AvK�I�g�0��-#CY9֬�Ƽ��kj��:d�� Š*�X�=7���{�
4. ���SdER��7c	=A�����ើ>Y�/-.��oŪ���]���Ö�&i�5����o�F�ZPm<�N��0w>�n�Q�J�^�Z=ۚ�]PU>khV���U6����+�q��V�9MVP��'T�j�6I?�	j�mS�%�y�j[BX-R�BT�)�(�~wthh ��	>̋Eӗ���AC��`7�[/����I�@E�J�����L��Xڏ�ǚ��q;�0�����	
̑f������@*��Q\�����S����2��B!��QY�Tu�3����w�w�a�▛oƢE�$�(̟��8u�4nO����~�kp���JK�'񽧾C�֤�R�f���r���t�N����6.5�"y��������9��RP}�=��/�����a,�����S_�+�H������~�ޮ&��a{�O���dO��QtĬm�SZ���I�Q�O�W�^�D'1�������{q����#Nb��WB�=���_Bb���4t�:Cp�Ӷ"�X����w��D�c���SLƝ����Aq���fB�}���q��x����m�&�,���Gp���	U��[o1��j!L63v�~�˟	jR��?��e|��O1����/���O�8l;��Kg��_^�ß�M3�]ｇg��3����K/�G#���7^��g`U%�gϜ����;B�o�f��8��6r���8����+����~��d}���}T�9���������g��'���R'4���6�C�򃴩��d�ќ��z�׊���}0�#�$n�fGUYƇ{Q�U���f0�f:���ɏ���,Z		�@�q�h*��P]��es���መ�{�����Fme���"#8z�lݺ��h��f%<���T1��0�:�1��g Bv��{�`�[��e�ؽ�#�iX�$h1H#������sZ��H��T����*u��$ÏA�[.�3�:v^ma�+/6"4�v"�v�	����H�i��-�͆�l�����}i��KԶ?��B7���' jRJ�KK���/mR�5�G(�PK �\M!�ɠ4��Ox�1"���N�y�h� ��CE�����ǧ1^-rR�#i�1d��Ts��̣P����C^�bʊ��lwv�^���B��*�6������aue��Ȧ�Mr�&���`딆�)RTT��'��{�H��`��颸��砷{?�o��'+��%˗�V]��[�m���0:x���߆���P@V�z����q��aY�6� +W��Tb�5�Ås'�W[���%Kf5H��BM�-a�<J�@k7���Ƶ��k���L	�.��S��-i4�
�Xj��PW�`<lB�@3 /����v/R�҈�i5��p�Ӄ�?�iy�,^��[������<֋Qϐl�:������aJ�+��[zZN�"������Ӫ��������
�����J��+��o�e�z�]wݏ��Q� �r̆M����{b\h���c~�=��dш9��+	@��*j+z��у�)*ذ~Q�MF N�BI��/o�z[jK7�t6nܨ5q���K����I� TW��ƍ��x�,���	�_�����|$���5k�~�A�r؉D#>+�m��fP��X����l$�&=$��bJ�ʲ�M�����#~l�if�\I���L��[�?}Bq?�A�[]��&�!�IX����Y���u((ʧ�&�4�>2�G����.�_PO�]J�;��SK�|�=4�ˈ���f�X�22��OO=��)_ϛ;]��}��2��lX�AB�Z�Tm��#�'���X�f/�(h'5-a��>�Ie�u5Ӱ��;p�M�I�t
ў��������fϜ��o��6n�(�b`��j�(=j�e���曰v�����?��0P=�z���J6����Bi�3�MQ���� l-7]nz���#�d�Ͽ�k�-���%ziĴ鄹�X�=���+8r�(�tEŅX�d#j�)��4?4�9��+ǥ�0����m3�s��)Or�־���-��nD�=��l*3��=N{/��>"��BU��W`���R-����!>��}��=k}�P[)���<��_���CPp����>�?O���q�?�яp��aI�s���S��gY95Y���7��$��E٨���|��o�K8��gIrI�Ik/(��C��Ŕ���8,�]���֌�9)���v�͢����?]!ݴ����^ߤ�;8Џ��lL��������sH���CG�Qx�<�ch�I7��͏10<�lZ�ko>O��o$42�O��4��"/ہ7~�>�7^�s��L���ￌ=��q>��v�f�t\!��2���;�^~g.M��3�����֭]�=��rR,Z5��9x��L|��<߿� �:�u"��8v�/��������7^Á���n�rt��Y���g���.�7^G�AIA62R�h8�ګ�������M!3�Hou 0ڃ�����xP�N ���PښN���6<u��}?Jr3�(�豣�Htv�K��]_����^d��"L��꫻�~�������A�a�"^����X�|)�K�+�f��DmRj?~�	�68������%<��~���/z�F0���_�u��0-8.���A?=�lܴW�/K�����N�s8�F�R��1������L!T�ɖi����ޡu�3�vttɩG�V��JF���$^kGkK������I�S������$���n�˭DGv��n-�����5A'��ndk�u�HǾ��(���THYI	���/����q�w��Ҡ��ˢ�>�1\��c��/C���":�k�������p8.Jq0�}~8��#d���X��+�� ]�@�y"�M�8��"��՝1c"�@g�q3CC�JuIar���x�7�@�W��f͜�T���/[�G�alxT6�i0�-� _��h�{�'�arR��3Ż�Nݍ�����Cz��2`b_��=a�gf�b�\=� 	�1�d*�cv�,B�4���v��A���Ȩ���/��̍�Q"���]ʚB**�.����W�W�6SU]��v܁SG�a�	��w݆b�
U���Y�ūV������vd���l���(��%K�x�r�������/�|��e�v��3W���	��=�S_�y�Q;����~�V�8�����e�����¤w3gN�}�݋w�}O��,Z��;v��Z�_���߆7_C,qݺ����[��D5U,k\��?�0�!�Q���nټQ�#J+_��_|�o��5=͎��7c��m������Ř�{p��Q�ek�W�VF�k�l�m�P�à�Q���$���C�Ό�����
p��ں���|�{R$f��E��ˇ{�MT���B���}�����{����ZuY1�.�+*0K_z�oq��U�����BYi%y��p4�3���S�i� �H�,g�Ȕ%UN	Nr��>�$��wpr&L�3��8��wbӆMQv�5)�2��'�RTT�m$��׬�%۔�t��������0�N*�v�"C	T:;;��V]��w܎[n�Yv�:�V���sD��ѕոᆛ�/o��	�3=ˏ�d�jcgyE����7"y"��t��'p�S�#��j/c�Kg�bnuB�{�+�XWW���Z"�|x�0H~�ή���ۉ���i��X<��!,��~~�	Z����a��0�a(.	.��Ǐ��W_��&�|�"�M���C�;H�72z#݇�`¶z,j܌�yy-C�裏����&�uk�Ѫo��槒������%��mh`�֝!�ٱD?��ϱk�;����[�$�LKːNG�g?���1������o�����w��1&���}�9����x�3_#+274և?��'hm:+b��+�#_��u�?m_�v�Ţѩ�ͤ�B<��M&
��Ǉo���te���Y��(kɢ9���[a*3�k���{�[��⢑$����O�-]���_��KC.7�a�������_d�`��	?���&�j�����6�@Ϛ��v�D?ښ#���������	ܺu;����O�o����3':v��<�7���w��)�=�A�;|���'�|B�����c���kWV)��ٻ��y�OJG�{~HR�����f滎��<#�w*�����8{�$j�R`�ĺ�^®���;��lx���wp��1�ӓ�!���x��	���u�D�
B�Ԛ�Q�
`h�%q�������o������>211�A����DZ�x�����}�t}?�Ә��mȪΆ�
��axtyY�0��W�oF^��8{�$�c���e���N�S�0%y��u3fo�&9�L���X�wM0h����p�֝D2Q�ݳOZ��S��G��ўh0[p��(
�Oe�Ҿ�jm��<T�m/��`gB�d��D�F����_(��TW{GG3&<����{sL�Jmқ~ޮ��2��� F'b�LN"�JIs����MC��f�V\���������K��uI=����#�L���.�
g>Z�7J��7"ӑ	'9�ي��u����hЄ�	?r2�O��k3aU�G�n�]9�jO�ڽ��GX�d��0Mg>ʐ�!X�v�l����=@��@Ii�A(UrXA��m!�#�w���X�aY�tz�1zi��&!�y�l#S@k��]�ҫ�>�Iw3*����P�۷mFa��g��	d2'2IǬ�u��,����#SmV�$�\X?���%;�V���I2}�!LL�eU�q�B�uR��A�Gk�[�K)'����dH�wث���RLV�ġ�i�+"�^�r���P����`�)H����z&�3)܀E�(�n�P�%��֮Y��y�ar�Y{s��߄�X��kf/\�6�pR	�ť�."�Vd�����P���Pe�7��NՎ�p�8�������,�Ƨ�4z��1�Pii��V�NK*����#��q�4\�u�.jD,LC ��>���i����b}(ș�����L�+o�5�S��Ѹ"X�i6n�Cr���bV�<���`�����u�fl�v+�A�-K?q<�:tSP�D(��P��99����a��/��"jk�a۶�ƴ��L���1�l(����L��i���+a��)|0ڭ��`r
��j�斡�r!����-zņ�1��JÍ#���5vzNH�b�����D�Wŉb��G�����1���|aA��tza�f΂�YJo�!�$��"����Z�2��1S�XSyDE]�ƓH�ԡbŨ)Y���E�aY�S���#zO-n���_w��#�C�I;�PwV�ϫ*�p�NB�nP[>9VC�Az�ԑ����h��zr�Z�3�	�oo�.��b���	��3\AHظ\Y�_�B>y�/�a��|�BT̘���:*(��H���a��rQVۈڙ��RT�iFg�i� �֢J�W�@Y�\*�(]M-8��;p15̩Gu�Ԧ/c>pp�!���$�W��e/GfZ5Ҝ9t� z�1avQp��#��x�7�dR{]"�����pv�"^9(+�B�d�����F�0���5n�����Jx[���pD#�xi�؆�������_�.rs
eW�ۃ�쟱w�i^�5���&QYV��Qm�H�;��s\�S���r���&��vb[R!+W�*ߤ�����/΅���ݷw���ԕ[��b�dh����v^\9���6�5<��2İ`�vy��ԉ���h�@#Yo;�1�y�6Q�>�C�DZ@�3's����d�0m�N�+�\E����0F�Ֆ�[�����j�h�(��ڰ�`X�!H�]Y��&#�ng,?;�#�3V���ׂڒO�!Lx�6�C��BBjݞ�T��ey��.�5��=��4��q��	y�x����L�=�v�䉣4���q��I����'�xB;38���e2ŧk��!ّf�eeU�0���M����|�2Nu�>�#���c��s)� ��	����e��~e2��r�B�j=���¨N$%�7��BU�*�U���38~�8C[�ɐD�ɯ��M��	։��3�x1}^9�1
m2���~��E���N6sp����O�����W���GhS9�����fh�F��B=�1�tF"�؄Ω:A�l�	Ǚ#�**˩v��I?�9f��kƉ�,00�v����$���twu�a2A5>J[ջZ�\�c����U�I� [���Mq9dS��DB;��s���.`��t�M���I�U���B|�� 7�E(b�z��@j��ɷ͗.�� Yr�|�䈈����
��}Q"���4u�>�Ak��z�}(�d�&�R+��HL�R��أQ�����]�jװZ�Wv��*�Dz������EE�F½x*t'�
s��q"F���M�0>�l~_�1��W,��*�����8�	�;2��RAD��gΕ,UZQ�r�ޏ�OZ�ʺ*�/_�TJ��$W��HT�)'��R61h(�MIz-~�hBQH"&����`��	JUR3�sp�����?��C�H���¥+Q\\�c�����t1�.vP8��Q&�e�N�Ɖ�kk��=Љ+�Ȟ�
ͤa��u�;�P����12҉����n������n�?ŋ�����{�UjYNG	
�������h<#s��^!�]����r8��)��vWJ:Cvv=J˖p�Y�4���+W��e���hrJ�VH���Ӑ�5�cW��3��y�2l"�JČr���Kpӭwb����,�u��}��j{=�M?�ʨ������B�Z���Ȩb)�G��@��ǐ������o(S��F�E,qn�B�~����]i�U3KZ'#����v�f�j���d碴�^unK�*��\q#J��?$R)�

I�)G���ض�^Ri����V^c��������W��e��X��^���|ZY��y�P��9u��X�f��9�Z��Ɏ�����M~�*�x��V�͖����ɡ�3�\)fB� ��x;|���;�0;���@t���*��%ex�����e�KU ��mm�҄^Y^!�!":S	�Q��R���L]�ቲ���i����)�T&9����#|7��Ee�L䪐A��v���a;uI�r��[0g�B���)��x���9y���y���>KVS�!M���� ��*V�ЭEy�t�H?.^8��^zsf�0g��d-FV�*9�*�c�}�a�:@��ir3� �H���c"t��;@�_����p��
F�>��d�4g�盦�,�fιT�s�b C}���0�Qq�CE�}p��D�@���G���L�FT�}�3O0��]�r �/~��߿���b�%x�_FfV� ��U��j�����J=F�e]�!���!�n�}=�]8x�0�z�qy�̝� ���'�g���{���q�r?�.���~�=0��:��ݿ�.��σ��������7 k$���Ʒ�E��M4������{���?���@G;���3K}AZ|����P�����K����Ig�x@[g�U�QQ�c�Mh��KK����s��cA��̃E��k�٦c$q�-r"����;�&��<tt������'�r*��� z{�Ǌe��$	|�{Nۃ�<��-��_����?�5Ż����q`�.�JSF�;u �{Ƃ�}�;���"�������a���b�������Ʊ`�|&5s���F0�����;�p��a,Z���(�Z0cz)�m��J�p��Ҋ�+V�ҕ38��<LX�$�=y�$:;���Z�x}��L1!J6�6)�8q;�����2|s ���h��[Č���[J:��˻��db5�K�r����n|�{�Ѿx�/�H"M��jǿ��1�g�1<���'����?��Pag������vZ|o����Q9!H�[&	T�ư|�Ҥ�?܇��LzbXN�N!��G8���f#J=�4{�Q�h��`	�G{�T=L�i���z����)�����%��u�,C��3	�/��Q`Jkj_`\�
�F3�3%V��{����(x�C�r,f�`���|�m�+yGNN�4���S�����q����,��Ǒ�OE�F<���.~�c ��y((��P���
/)���x�Ř�ήV�_�r{q^1��Js`ɢ�x�M��F$�{&�a�B*+��+�U�����7�M�	��kܰ������\9y��8	���	a���OmĘ�q��I�F��G�-����P!�h֎2��m�������*k
�3�Z	��QE�YW#����kK���+� V�[n���W��c�a��}�3��D0�NW(��O=�_��_12:�����gPDh#qk�5�q�a�����i~~1n��a�	��.XK,?��_E4m �ӧ���1�%�fˆ�.��C�9�=}>z�!
���7?�i���_�K�\������bH80k�<|�s����ŬF��{>Cnb�������G,G�,\�k6l�s�q��_M#�!���,[��7�H2��`q��t��ǲj��a>n��N
߬\;�\-^i�q��h���7�����KFuM-����c��X��Ș���̨�5���Yr3r)��sg"&���9�y˭��>���ue�D5�EI�e���w��҅�

QTV�I��&,��;�n	�χ�e(J#7a0Y"p�j?��/a���L�F���{G�z����ؾ��߸I��r�8h��u�sn^���v�NlٸE��)鲲���*��Up����OO�&����L���"�ʕ�b��۱�q��<e��#̨��ܤBP���[oǺ[D���1��L�v0�~ҵVl��	�I�kL$�9ԖpZ�rR(��+Վ{��	������!o�
�Q?�%�D($sv��Ԇ��4z�Q_�*��´�*����|SK{��w�EC�ܙ3���>c.=J�\>w{�y���5���ؾ����=m��_? �p���Ý�oĬ�yLSv���_���_���(j˫����#���D!��0~��ë��F�J��������+��5O������7�x�V$����|�)9�C"e}��?�}�V^__ۀ���<R�IhU+�����r�䔊������S"5�	�O�4�O����?���N\�Er�nB?TT������i��o�t���FT���y�n��)A`b8�Ǟ�G��?�&�9���Ձ��v&~7��Ʒ��x9Y�?�>._�����h�0����Jl�����{pD'��I_��"��>��	�R/~{�<N��HXq�gϪs������x��	gjyiNZ�U<��_�{���le8}�8>x��J!�=u���K/�����A�H���|��뜧j�����<�����_zB6�~��n9�i�H#�:�b�ǯa�ݟ�Hq��] �J���A\�z��}�m�ܭ���ܘvX@,�(UzӚ�d�V�����C\W�U�jQJ�z��	T�ʭ�dW�o{�eWy��~7��o�(U.e�$$!!��$@�Ɉ`�����M�ƹ���~=3~=���=��׶1`r���"HH(�R���Vݜ���>�d��֬5�Z�o�9P��:�������N�>{�d����.@�� }<ee4VA���*Y�	�C	�"I�`jsz.vS�Zxb��4H.;�c<<2���r\��AIEa	/��BG
�G"2�G��Nu�\'����<�y���������01zmS��'�a��}=��c*����͗/+)�^Kp�:xr|��x14Ї��Je�F���t�=�51"�S�h����C�w��[z9b��nإ3�5f&���5�qp]��Fl��M�+��M�10�Nf��SW���r�͇h*���X��� u�7?O�¾�k)�I�:�F�mT���Y+�T4a�J����;���	Re�
�<	z!��$�n��(V��q�onzS]5bN�"�\8`낳̅���{R�N��i����Sz�c(-��D<���F8h�"\��Y��x����oa�r�O�*�)!��9����$z���A.n����2��͝�o��ߏ�"U=-�"Bv����>ltԆ$2�qf��}TEIŰN>Hk�����f��Tz�iY�����V�:P��f���L�����J
�;o�KO?�b��Y��ij����O�_z�63���e+��j�������;�|��Ӟ�ukn�'ϣ�3g��z�m/�߰����$��W�t�Ln�(v��D��Hi*�����4C�կ|�<�b� V���|<V����o~[_yNOͲk�b�[���9�M��p��_�K/����K��7߬V	 .X�<�=��:mP:���Wb9Q�Q�������<n��+(��~غ�o�"=I�I��clFK���I�?˃�宿�0m�#��J+��/)��-'�@U�W�� !� �
JPI��Υ}��kf͝C��Cu@~^1=�Z�t�DF�A��(M�~���E�X���*q�7SZ!������\�{e&��1.?�{%nY2f-��(�_aN�hc�X�v=�-^����[��lWO/���M-^��K��s��V���~�A�u�n͍Xz��Q�r Q�=��:ej����\{�j���e�3����m+!{I7��_|�&�
<������I5�Byeev��'&ep�Lv�j�����,�g�dC��H�h�,^�siij@�:�HI�"�	9�6�u䗵��{�Ĵ����53�KT���J�<ƅ����6���
޲r8�6�>y{v������b����Ь��0_���x��xbƱh�5�~ӭ�1��P�Z��pd�>���s��/X�[7�A�٪�������/�e���ɏ��S��k�3O�G�B�pj���w�jZa��uԯ�+���Ƙ�,�G?��
Q,�V����-Ξ����鞋�7~v�WmJ4>�g�|�~�.n�ͼ��_��;���`�,�66�re����y�~�O#���)'Ǔ8p�C:�!N�<�Eڵ;v�M[��w���W��u��p��\<}���_�����~;w����b�߉�����7�
fW������[��PbϞ9��g/�'�����O=�>���/Ө&q���5��?���G��>:����|_mӷ��߿ϼ����e�pN�9��%���?�e���x덭pȳ�9�x�8�����O��.��ݻ�ګ��96Ӧ8	w�_��_��?�	�%�}{?�����Z_B;��ON6l��ڋ=�v�����#��?�#~^5n�r�g���YR�+-	��>CY�?�!n�vL�����w�A�S�'�#Wp�\�㈍�a��jU L�x���-���O��~�cC�	��\��7������h�`&iQ�fA]�(��ũ�w�6�8:C��D~a�@t�8����>�OIІG�P�b��w����I�C�BeY��		��˗�*ǩΤ2�}��R�������K�(�r�Ϟ7f,r1�*�"t^���(����*<�"�i̻��T�Z����2�hZV�x�c�=�hl3W�ax�:\̤�;�%`��FVdr�П6D��\�hn��.H�$�K(������뵹�0g��{'�I	YE
!����4l!��^8w���t\�ЗG��
=N�����X2����i�qS�|q����X�=yJ��Mp�z����6JAMD/.OU���_юȖtFI�p��ِz�HH��\Ģ>̦���=�~�m�Lx�K�z|J�,^����`�X0|�7 H�-�9J�4C��$J�Np���7�s[&��o��dk��g�����LZ��+���'����zZ�;$��_dg�_G������*L�d�������
W!�wvj��8��G_�N��s֢�j���pݥ�m�/u#�`aٚ-p7�O�R\]�5�n����Cő�_�e��F'DUS��܄��{��WI5�m��/#/��/���þ��SR��b>��w�ܦ�f*�����i��F�y��:N#E4���{��W_ۆ|��r�_�!
��46Oŝw܁�w�G����˰�5p(HhZk+��~|r��ڐf:�+V������Μ=7l�����D���[��o�m�e�1EHĤ�#�ٱN��h�"���u�Sq�}_�1��3����X`���T���>�Qv���f��w��v�P5m����`)��S^��9{��ݔ@ۢ�(�m�JDqI	��B�M�%��%r�����ҭ���ڕ�[X�CR(��{/n�a-�Omm��?8��G����*��,\b�#��ϟ��4A�]��o\�%�,�*yi��������`%]Z��Lz	���_A���+���28�E:#$��6F5.�r�����y��#%�J�o2��֘�+=�,�2L��A0vC$`��J!�$����y��ǐ��3�+@���)���+�'1_7.{��p�Uc�;��3a)����N���O�@Ay�����u��;w�\�����i1�`��[PP=Mg��R	t�8>��4�uS�7��z�&�����s/h�`�M���}M!�ب`0�Ǟ|�ą�g�T_��|��<I���8�W
���踀�Nb���x��ā������?���WX|U�\��}�!j2�xtJ��8���u�A+����<ETS�j�|=&��L��eg�f����xiA��t�����6Y���3�R�����ر�e�޷��P�4�+2n+�v�zoE��Xt,ԅ^�U7�������}�W����@��%��tw���kyO4�?��(/��K��q��{ 7��CU��n����RgM�~����m��^�:Ձ��|��Ҍ����,&����UB(S�� ^y�.Jn�qa�����_�o��ńC�����=[K'�;�-6�X�A,�>>سG�2���	�em��ͷ�fgΜ�;;�0dh�<8s2'���Mw�ʓmͩ'�lۮL;4
�h���Y��,]s6�>Y-w億�@V�%��ݙ����45��cJ��T8��F���!�{u�)i]�f}��s-�FG�_�F��4LkC��M5wFKN\N�o<��X��i�9'Ν���9�L/l¹�'�x����(��ȥ3T�T}4�&��Ǐ~�Uko�����86y3���@�u�B�)��jcccX�f���*(��%��~:�>���R�
[��m޼Y>Bǯ�[�<�K�~��_��!�������b��==�}�Nkv)Y���&�t2��B��-q<S�)�*K�)����4"�8>�Ҧ���/?w1�H����4{�L�]AEA�����#��Vs��_�6�i)�KH��B��bz�|�G�"zi1�����sst8�,H._<��q�B]]=|QJ%�j���'�s��Q�����S�"h�V���3��¥�.����'Գ|	�N�R�]���/!�n��sڝ��c��y8��Ǩ���W%Fh+��)_�y��b'�f���w�ԊL� a�۵j������V1�����R�%�N!LNKp�^��>c��ܩs3hJ�������Q���V�kل�nݍ���3���.cx"����U�h	��U
���9�;3���9�W6]	���~I�z�$F�"�u�!e%St�{qY���-:d���{~��ip��Q8y��!T�M��E���S�k��.�>O2aCA�o�A;k/����{�.M������D_B  ��/�|3B���
l��%!����jnUB}��ru]�}���*��n%������l�̙&���o!�H᪫�ƍ_���T`��,=�6%�����O�MJ�ղ��V�iM��~jCr�r��ZZ��v"!��˛����(u��&cg�i���F~�f��@xJ�*�"�t�|Z%��iF�̻Q۴	y\�j�=~iA�c���P�8M�DgO�B�R*��˗�E[C;��G"�yN��͠���^w�V 
���@I��t�]�����I�5��֨��W�ꅋ0s��D��6'B��07"յ��x���y�{�GH����H(���؋e�V�}���/.,����� �vD�>��0�4��؄�:[]����a�źGÑAV�3Er��z*2�?���ö΋0w�L��4�]1M�A�'�KX{iQ!+��V"�kʂ��Pp;aq�����ϛ�p!G.��c�5q4:>H����T�L����S�qfާ/�����+oFIE�MHFC8zx�N�	s�[����5D}���v\��$j��Q����޲	-MMJ�J,�	|��>%�,+��}�5��Rt�;{�"�^����� J�h�_��"o}�8rh�z��|ǽ��ʴ:1M`�KO���������0{3��"��2�8��*�1��R�l�P�ELi
@"��ѹ�!��^y�``(��3�چ��7��GdՍ7�/���)6�&QSJ�H��dw�[vV+Ppx`���&t��ਲ਼�v�����Obb�C�����ǎ"��G`�)���e����I&4��q��>|�/�G)��G=��S�*�f�*���D ����m�����GU��z{��م U���ϔ������h�{�u(4|=���3O��Li�|r�>�ZZ[襇��}�����x=��!�}�-��|��r�'x������D�h��w���g�P��IgN� :��ƻ��gt��T�@F}��0����Qfreg'~fC�bq3q�Ip��1"� o~�3gcjyҡN�J"	���E��4�G�Vʑ����"bOL�t���W��rCcㄉ6��"��釟�ic��;5���F��jG|��Te���n>O�ȍX�`Lؿ?n�r�0:6��b�\���Ta!�Q�?��M�1�V�x���̹s��Sq��\�=��F��J���Ӣs+=�K�Բ�V���6�l���k���K�;�w1�3o��ph�W9���=���>��6�FS�� O�ҟGY��s�2.:.6��ʌ��a83v�k�P���f��	OB�0�c9h,���?㰖!+���c4&-D's�\X�@x&�Μ|D�#4da�|8U�3�6"���.g>�c�J� �ʡJ�:���,�+u��L�
���44����p�2����|�X�C�%���܌��z惆c�M_r�"z�.�U�j�U�K?�S�����ra����0Qe]��~��'t|^����ؠ���͝�҄Ӈ�K���T�i�S%ڋ%L:k^z��%A*���&�F=Z2�2g$Q��"�F���[\d�Aaݗ���1k�2T׷!m�A��;p�c ��>h5m��s����� 5���#ڜcra͗VÔ;U9�XNd��'i��T�׬��h�M�3���Zڌ;���#@#^1�w�~�x�|�ܰa3���*7C����w��ˌ2G1���Cx���1A��GX�F���:��ȫ���^����3g>nڰ�P6��?��G�,_B#�,]BT��B�@���&\�~3�F̝5��V��{`�i�����������Y-X�j�2	k:;�QYM2FZW���-��3S�?���D�����_��w���A/��3P�������~Ӄ�q���+-^B>L#�WE3������-��P��(���X�� w>0M��x����)֒�pdVW�Z���?^�1z�U^�Q�S������kW���9�j	:��o���ćD\S��Ԃ��kpO��|w�'���R;M�3��i�%!u�d:�7���e%hji�/���A�a��q�����(,.��9K��ڮ�/���2�$��>V#U�+V݀�W]Mw!N��Qo<�J�s��Sڠ�6��u^"�A���i�����͕�A�����`ks[�B� ����5|=�P�oG��ܠUp���8v�#|���s��f�&,X0�ŕJ�}�8���5�-��	{�k*���'����Hxen/֮��к��:��	;v/�}���9�|��5((�Uj׭�l��2�MU��o=�e�C��f{�	�����f��������)Su*� �yZ�@`�~H)}��~WF�U+���A?��Ǳo�.����l��n��TC9�R���p��A���������5�N���	#b�bM�j�CL��
ӓi�s:r�a�)svx�B'ATUU]ڽk�o��չŅy���{�pl�+��%�O����-���|����uuŔJ7���*�쨨n�f��ﾊ��3��������{��9y���8v��"AA����������� ��< ��'�c�6\u;q��x�;����W_��x����x3�K�����x�����+�T"�A:�O�o=B���3��no���h�bg'^|�9�����?|���"ʽ���� F0����qa���Ϝ=���wq���󔜿�ڛ�z�!��&�2�~$?b�r.J[�d�]��R��3���!�B�+JR�`0-a��<�>s�G?A��ҳ.@�4D5q���Òr�=�o��$z2iUF���J�:<ԥ�(20K>řC��ax����c>�z͹��[۩���:J~��wbX����edܭp�/�#1֏��8�*�t�����*�JI�F#QUE~
�W@@2��t�,S�����B�������/(��2����=DWiU7=�}:ݡ��@+⣑	��ABҗR�s�I�r(�&ʴ������$hJ���M��Bff1���h���d���G��͓�Om��a'�4�����:.��V"�c�S�NЃ��杚��KQ�6���a���<�:r�Dԣ�N4�����ik��v� �/��"�h�s��*#,���Q��9�_��9u�t�P{m�'�������u:PU^��קO���J�����DBR5�B{��M8s�KgJ	������"��M�8y�L�I��0=�a�Z�9�B���mhl�$�"�$"�F�TG�DmRGiy�n�i<��Y��@]bW&�=u %3�6x�R�"9�0�8J��d���蘚���g7D�;42\�c�*.)����k�cd�]]��a�����Юܤx�u(����ƕ��z6`+,bX�P��'��Ξ��{����$��QPT�e+nĎ׶b"���K�_���"-C�W`ٵ���{� ?8w����f��(=Ʋ�K�����	���^�j�n�O)�y�:��g��`��mX=�S[Jʋ�b��x���av�b7kӭ��7���"h����w���=b֜��r���m�h�ӊ�7p��܌Sho_�{��������k��du�4}��[���w�\|�OT�3-mr���H�<o�|��),��r�W�Q)�=�Z�vK
�܋-�>�B����������d�o���w��	U`���c� �H՟�j�����G`��t�hZ^ !��1k�"L�Z�Qy�ب$�h��k�Xs���؜.��j@/��a��|��Z].RF����Օuh�>�u��Ε�)m����E�'���TK��[�kP^n����*������f���'��� �TY�F3B���0���M�Kg����\[�5k�H�n��"��=c���}	,
y���g�A'��2Lx:�D��
a��D;3��~�
:���n\����yT�Pװe3��́�R26Ѕ=�^��B��e�Q^�H����|��i|�λ��XR^�u�o�BwJZb8r� v�z��S�����V(?��پ�<xD3�/�[}-�ϧ�KP�x��w�[ZX��[�-[@��iZ�i����Ocǎ�uzB+7sӦ/�(e��&���..��P�2**�1�}�T�����8q�0N�<�Q���Z��_���R8'����5�����������DҚJ����T*�v�S�kKJK���n��w�W�<��լ�h�y�JUm���^d�΂#��x�ᏹ�J� N}�E�N�]LI�)ڻ�yG.j}<<�7�x�n��0׋�?�/>�Xx�G��3x-�Ö�����c���aJ��4��{5i��w��ήNe�/,S�8�����t:l2W���i���KJ�l�$���嗞�w�)a�'��G��D��B��Dϥ��w������:���_��]<�����8{���"�|4�"����t�|��:���a��_Rf>m��9"P�m��B�Y2��d�d����"h�U|[_z9��p� /�H�W��=y��¹��GIN	�ʌ!�8���Vf;Ν�#�Ok�2KB��}�ݨ+jU)���z�a��Oc:��|
�8�Ǘ���͏��u!@�U�� �j�'Ǜ'�'L4�%tܺ49
�U'�o��@��x ���"�F��_I����RK+��
�+�U6V"^j
�V��I4�����=\���"�� �8>6�q3�����B��@��-�ڪёa�A�X�3P"�C��e��1�M��F�X$fSTٕ�	o��=���~�x4����:�A8��6�y�����1��),�Y�A7�����X�N�.�D܁kn�����
���a�ݙR�v���~C#�6^��@���><ooqë��b��Pҁ�>��,a��uz��OmFSC3:.^T�1a7Z�z5�{��?ZZ��-����;�EA�s��<=�
���`u壟�'�)���RY'�E*q��q����h��%^�R�"mA9Q��[��C���ryPRV����.y'��('�6�1)!�Ni���~���fΜe?|�c���h����]A�1����@?L�~QZ������m>���T4��+��~�����N,�-J��� }��}�R�u����[�h�$���ʼ��{�ڶ�2C�bo��&%�����W`��_�˯<�(�}�t�vǽFP�P���ݏ���?�g=�~�Zl��dL�����k|�������ƍ_���p6V���|O>��&�͙���7@Щ��R][���m��w괃��z̹�����Uj�&��W�c�����޾��a��(�J��.��ҿ(�rf�g2e���bY��䨽���������bH'/�ˀ�H\�/�p��z��#�Z-nu(��D���Zq՚��H!E�4�bP��L*���~/_4���݃�pHI[d�eu�<�͇�j$�6K�n���%1��s���I�Y�IY���;�'H���L�r��J�P��q�R���
��?�6�@cP�	,uR�P�DT���Y�/Y=):��LH��}��\��is5Q&S��T{~:�2�Bhs��jGc�L�F����"���P�Y}��w2��d�Z�83�/�3ڟ�x<n�'l,"|��0퀄��bI���j�#G�E%F#�H��h����l�٣��P$n��r3�hLXO�2KVS�2r��-+�J���3��[�� �n��K�N�y+U�H0N�K�
���#�\�d=�9KϪ�~���Ji��d /�ɳ��g�qKi]��	�1f��RZ%�C8ҙ�F�%%Bbw:u�����}���
ad�;Hk�1�Ŭi]���f�;�S�ϩ,�ذ�lyq�i|Ѯ��I{9R���ňb�g�H'���h&�����>�I��f����t�,G2.!{��.�FU8�L|�j�Z����d��%干�R���ް^��M���+���j,ͪ)����Jd,a�_���1V��6��hѱ��
D$۩�"<�c���R�r(j~CR���Y��[�7�T�H���j��s�Wnd�ۓ4h)I+JѤ}YV]u_��K\��YG��?s6���d0� �5g?Hk��FpM�Gz��H�D�ɂ2)��D�ȶK&!���X1��!hu,�����T�/������$73���iլ�H��SpX�W�����r�ZרF*�'�Ѧ��,����y:�E(3$�n6��*�t�$�U0�!Le�Dx~���?����3�a\�=�R<R)9R"fj)��YF�Q;L�yM�H�?�����2�S�ZG�6�%�*/��,�$ӳɐ�TF���xVɤ%#z�eC�&��h��B�F�)i�8a��LT��p�dO�xq�t5e�Y�4��� �HkL)�-�9�\]��疚�%k��Q
��b$a4��}LFC�n�P�%���2�;mnJ+��S[ė l2FQA)���!��	J@\�WZ,�m.��1�d	�e�}R�U�hlL��Y4a��ɞ͖���JT��f4��P��V��V�~�%�͓��eyB���@CM����0*ge&�,��nS
V�=!�6�(��V��&+�M%\N����m�c�){r���V=�Z2!M:@�)㽍�g���<��h��l���SFH^�'>M�Lk ��"���ͯ�˗-�H����ƥdI$�f1e��E	Z'G"�v��4�9	}:n07��z,���0���D6�������(�:��0g	�-��[�ƔL�~fU��o�Ȓ�g�g1�\����L]D.��#o��n��!�ae�
XR՝���	rK~��52�C�C���ڕ�W�UfL.�*YAB"x�OArH�PB
�~�n� �gx{��Љ�7nC�C��J�Xm"*�&՟�cF'!pL)}6w؞�FW��I�Sԉ���J�T��q��oS�#��()�=1\��g �� -q�LƘ ���;�j8[&e�6ibIة��«�1�Y���QR�f�`ƽՆ��OSv�	��k�Ôְ��%���%7g�^UE�L\l���M���d�yB�UB��%�/SH��@ea�H�G	��섷�ݐY�f���� ?}�'�jkk��{1�;���H���~K�=~k֮Ess#.w_V�������*נ���DB�TJ˚��Α���`1bf���J\�c[6C#��,�aQ| ����&i�������,�tTE�|��,n�U��*LQu*VIc���K-�ɪQ���VIb�<u���
�L��^�ΞM�%4BW�+��^��XZ�RY����r~���O��,S���dl�_D]�#f�+�6��[��}zC.X�C�)�e^A�����Qz̕-�-���Ve7)���o�[��������R���v.BW�]Q]Eg2�q@O��c+�����BJ�UՖ�1<b��i��U$&�H���
X�����0�6����\�.r<{"���A{R���r���0S`d
����ƷR�����ԯ���D�'
@��dLI�w�*xoA>b��z���[R�A:�DN�d��WR�57n�#GJ`'���W0��?�C�D�*eڶ��ɐ�OwPA{�>,�0R�eI���+�ܱ���ֹ�?<��Kt��D�G���@�C'N��w]����1b�8]�K�-�/����]h���>K-�G���e�/s��AKK+^zy+���:�,�P懵kVkX���cZW&��N�6p�|�ZD���,[~�Ny>{����S�j���C��$�z�i����6��y���;5v&�&x@Ǝ�/���jk�t�VoW'��JU���D8�@҄�XFa��ֹhjm�fG�6a`Qν�<�K���S�+��Ŝk�Q��>�!W p"n�CY�%�gi4���H��.-.����Ȱ�T���
}����Q�p�C�TU�D���;:/jΜ�ص{�Qyaq���ݶm���Ŧv��G���v\��j����D̆�;g�,�����
Y'�R��X���2���vC�SҚ��PL���^�����]v,Z�ˮY�g�}A7R�nޢ,�߮ �:�i������^���<��!t��,�t����
�?���2@�����0g�t���3�S-�P���A�X���1���s�ry��l}Y�tҢ-m��9���jA�%[
)�3)=2����y��|����(/�R~�KbZɠ�vӰ�yJZS_۠����cZ?��ܦ(IYp����S�z�Jx<n��cǏ��R�,�r��@�W�	��M��z�|��|ٵ��B����)k�������M:�UF}��6���x��T����Ʃ�sAw�������J�dȽ�^z��8H�"�Q����#���8���%����jq��)c̻����nô���Nj�}��q���$�+���Zf����ȇ�uG����\ a���)ʬ#�m�g�!�5�שm[���*�)4�g�Kq��v�j��m:�j�P?�	'O�5�qʘȐJa֌���J=T���,?���Os3�Z�)��K�0�vJN=\�j.�8��D32<��ׂ��J�𡃔�B�&ȼ�?Klұ�'yj�)Z3��9� ?7Z�U����0�ՠ��^ͯdL6)��}}�1���E�H���&q�<��� �>S�C`��|�?����v�bj���f�Gy<�Dy�8�:���>w��c
��*�����1]�S!L^�V���4��+4f��j�yq�W���K�mz�N�i�%�>>6��J�湉����Dw�yC�#��.^��E��8?W�gk�SKg��sq���_C�D���խ�\���U�E*�P�tڡ��n�P������؈��M�=� �OYI�xi���]�gQ�S$�l�QXI�	���������b��X$��{��8nps=&bi�����.��,��Գm{u�:�fLB�l6ۍ���?ߐW]E��*���k�@`����1�
���	������:ih�E"�uq���p�CD2��oQI�n@k[N�9�c���C��)��6f��gR�r?���'N�U
V���H�J^~��[�abC���ǅx��Oԡ�g��k�'���c_G�0m�Ltv��/ �����Ι7�Z<���>�&�	FF1w��.%��j�LJyLZ`!h/�s��{� 0:�MD����@|&���T(@}K��K�-<6	�6Я[WS]c�FS.����S���������>E�U��Ӆ�5Y�y6��csp7�D�&�HaIE�������nqX����MI�y3��ݘ� ����.9yW��/8`�R�R����k�e-Oű�G9=r\f�@؈S����b���H
��ix[��x���×z^#�gĖ�1s�L��q��a�R�!h�
��|��$�:62�a�Ɔ&r��4�K_`<�51�!?m�@]kơc�����0O��N;x2��5�D���;���r����*�~{��o��v��E�i��Y�j~���¹ �o�/�ǅ�N�?4�ڳs�sxx�Z����i��A@��;ﺽ���)h���{�k�C���F=<AG(A�_����f�c��aG|ia��������'�L$m�� ma���!�OTTTp#k0AH,(F6���@�d��Iw�Ph��Yhi��v� ����rt�sM�6�`�e�,��L��܈)y��Ր]�NiIծ�ղ;���ŒՁ� 1<]h�Y
=�@<�g6Oy9�*���z9��٣�'���ۑW�����&U�#z�on�\_{�A�<y�.��M�᾽�1�pxtd4�皡#�}��J5�q��HQ�Q������p�8%BB�.JR�V �O�P�Te�Kuȱc�5�"�'O���8q�O�d�)�,�c'�H��H/u�2v��'En$F�C���f�8y���oI�P�$��F�@M�q|�(�58}��r#��\9r���QGwr�pR�\8w���n:�|n���fx(�v9�f�:�"d���fȵ��8ymۺn������/9\��:���h2��on�\ӧO���ZHL��i`��6,�%S�d%�����uZ����#�o%'�0�K��eq%���k��RIY�ƙ�<!��]Ւ@N�<Fc�y�y�F�j� �Pd�OI^��O�D?���T�{D�ķ,f�ե���Ӛ����c��&�g���i��<�V��%�}A|�G?�M�gW!j|Ҏ����\3n���3�����XU77�-�V��_�l�p؇Ϟ?����IrIa)��\J�8R���d�cF���&љ%���NB~�t�ٜm.tخ�~]����C��R"��"�]6�E�Al���e�5bm6~^ǇkZ7�o���R�'�AX��y��J�����႒Bu~�{��Ǐ���g�,+Є\�"�!(�m��8�~���]=]�S:ׄ����X����G��1���_2�f�PL�āub�DX\�y$��T�$��F^B�^�����,甑�#�L)#�*FXT��y�b�w3z��Ň�d�o���P.�gI��l�>�I��J�fB���%�(Er �*J����s���͚5���4N&C�eϑ0�\_hC�������O�:y������Ο^����1��f��jOfbvq�bј�)��x,f�B��Qw8�R�	�I3�i[ p��d��&c�F�VɆ����R�&z�����f��ĸ3)���D��pZ�����6\I{�G��$M3f�%�d��CC��ϟ;�"�.F*٪��t ݽdɲߨ�O_�"˦s�/�����yb���'eWrr�Іl߱���.� ~��8���q��҉WO�b�h?��4��B�d	�'��|�>�h��S.}�v��W6ac�ܗ�Ņ���	3����g������i���	[,�S��ۤ�B��h$b�j��{�" ��j�rS6K^41Q]�0�og�e%�p�\ΎC�����_~������/r��MAaa!MSd�'����ĉ3:��m��3�$�k�p��t��5�W.%�R�#�vAD~�H��D�DmIY2k��I�)������:}F'4,�EL��'��o�O%C��ҭ��c�R��$eˁҸ2{]�''�85Q�\�1�i�O?�z����/�����K�l��clb_�Z�`֮�n������S����{n�w���6d�����uen9/	������4�B�(���a:��&� =���
�1#�����q-X0�>�X���4�Z~9�|���ِ�/\�)�U�ڋp8�g4�����' ��7����u��!�9�?'�q���!�/�Xs:������kC�']�]C}���}�����?3���y6    IEND�B`�PK 
     ��Z���BF BF                  cirkitFile.jsonPK 
     ��Z                        oF jsons/PK 
     ��Z����� ��              �F jsons/user_defined.jsonPK 
     ��Z                        U� images/PK 
     ��Z
�8b  8b  /             z� images/a7e3301e-fb46-458d-916f-a05c0bde95f4.pngPK 
     ��Z'�Y��  �  /             �V	 images/4bf63cb1-3675-4452-8ab6-1403298522d5.pngPK 
     ��Zgm=� � /             [	 images/793ea4e6-6f4c-45cd-8a04-0920ddad3581.pngPK 
     ��ZĊ���4  �4  /             �o
 images/627c2b90-5d53-4228-8b10-5ea0a126027c.pngPK 
     ��Z���  �  /             ?�
 images/7260fbed-8271-43c5-b1e8-f8e9900a221b.pngPK 
     ��Z�wp�&
  &
  /             D�
 images/e3aa425b-adcd-4ef1-9309-97e806748a2c.pngPK 
     ��Zpg��>� >� /             ��
 images/1c06f444-5387-4cb2-91f2-17a999ad4bd8.pngPK 
     ��Z�V]{[� [� /             B� images/995ec925-f4ba-4c8d-81fb-fe52a7fea57f.pngPK 
     ��ZVX��<,  <,  /             �n images/6bfc6843-1883-4a57-a768-11efac5c5eb3.pngPK 
     ��Z��s��  �  /             s� images/9d204b9c-624e-42df-9128-467635275a1c.pngPK 
     ��ZP�x&�  �  /             y� images/9296751d-4d5d-4f26-bb1b-b9b3216c4bc5.pngPK 
     ��Ẓ;�  �  /             �� images/f39c2bb7-8598-4025-b62d-e677fac223ba.pngPK 
     ��ZFI��  �  /             �� images/3d3e563e-9ba6-48b4-a3f8-79399330dfef.pngPK 
     ��Z��C��  �  /             �� images/89208456-78cc-4fe1-a1e6-da24e243623e.pngPK 
     ��ZP��/ǽ  ǽ  /             �� images/0b351edc-7875-4477-b820-546ce15be531.pngPK 
     ��Z$7h�!  �!  /             �� images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.pngPK 
     ��Z�U ��  ��  /             �� images/ae1d0bb1-db79-4eca-b526-eb1d648f9ad0.pngPK 
     ��ZJ��F�  �  /             � images/1348d1eb-e6ae-43d4-937f-d455f2ad4bcd.pngPK 
     ��Z���y �  � /             p� images/483af35d-09f4-402a-a8a9-75c28eb4643f.pngPK 
     ��Z�9M/�  /�  /             �h images/0a03a94b-1490-4d51-a356-eaee23e4f5f0.pngPK      /  Y�   