PK
     ��Z�l����  ��     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_0":[],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27"],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_2":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_20"],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_3":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_21"],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_4":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_22"],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_5":[],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_6":[],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_7":[],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_8":[],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_9":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23"],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_10":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24"],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28"],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_12":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_29"],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_13":[],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_14":[],"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_15":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_0":["pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_0"],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1":["pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_1"],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_2":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_3":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_4":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_5":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_6":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_7":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_8":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_9":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_10":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_11":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_12":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_13":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_14":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_15":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_16":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17":["pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_0"],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18":["pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0"],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_19":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_20":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_2"],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_21":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_3"],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_22":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_4"],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_9","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_0"],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_10","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_1"],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_25":[],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_26":["pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_1"],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1"],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11"],"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_29":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_12"],"pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_0":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23"],"pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_1":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24"],"pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_2":[],"pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_3":[],"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_0":[],"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_1":["pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_2"],"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_2":[],"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3":["pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_2"],"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4":["pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_2"],"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_5":["pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_3"],"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_6":[],"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_7":[],"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_8":[],"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_9":[],"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_10":[],"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_11":[],"pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_0":["pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_0"],"pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_1":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1"],"pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_0":["pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_0"],"pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_1":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_26"],"pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_0":["pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3"],"pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_1":["pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4"],"pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_2":["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_1"],"pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_3":["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_5"],"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_0":[],"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_1":[],"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_2":[],"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_0"],"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4":["pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_2","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_1"],"pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_0":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_0"],"pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_1":[],"pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_2":["pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4"],"pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18"],"pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_1":[],"pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_2":["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4"],"pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_0":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17"],"pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_1":[],"pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_2":["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3"]},"pin_to_color":{"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_0":"#000000","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1":"#e8176b","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_2":"#0E4CA1","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_3":"#9E008E","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_4":"#010067","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_5":"#000000","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_6":"#000000","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_7":"#000000","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_8":"#000000","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_9":"#FF937E","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_10":"#005F39","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11":"#774D00","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_12":"#91D0CB","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_13":"#000000","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_14":"#000000","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_15":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_0":"#C28C9F","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1":"#008F9C","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_2":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_3":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_4":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_5":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_6":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_7":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_8":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_9":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_10":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_11":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_12":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_13":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_14":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_15":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_16":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17":"#FE8900","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18":"#A75740","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_19":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_20":"#0E4CA1","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_21":"#9E008E","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_22":"#010067","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23":"#FF937E","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24":"#005F39","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_25":"#000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_26":"#BDC6FF","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27":"#e8176b","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28":"#774D00","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_29":"#91D0CB","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_0":"#FF937E","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_1":"#005F39","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_2":"#000000","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_3":"#000000","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_0":"#000000","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_1":"#5FAD4E","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_2":"#000000","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3":"#01FFFE","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4":"#968AE8","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_5":"#FF029D","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_6":"#000000","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_7":"#000000","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_8":"#000000","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_9":"#000000","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_10":"#000000","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_11":"#000000","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_0":"#BB8800","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_1":"#008F9C","pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_0":"#BB8800","pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_1":"#BDC6FF","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_0":"#008F9C","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_1":"#00AE7E","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_2":"#5FAD4E","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_3":"#FF029D","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_0":"#000000","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_1":"#000000","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_2":"#000000","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3":"#008F9C","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4":"#00AE7E","pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_0":"#C28C9F","pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_1":"#000000","pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_2":"#00AE7E","pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0":"#A75740","pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_1":"#000000","pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_2":"#968AE8","pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_0":"#FE8900","pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_1":"#000000","pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_2":"#01FFFE"},"pin_to_state":{"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_0":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_2":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_3":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_4":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_5":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_6":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_7":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_8":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_9":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_10":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_12":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_13":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_14":"neutral","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_15":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_0":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_2":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_3":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_4":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_5":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_6":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_7":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_8":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_9":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_10":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_11":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_12":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_13":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_14":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_15":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_16":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_19":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_20":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_21":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_22":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_25":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_26":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28":"neutral","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_29":"neutral","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_0":"neutral","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_1":"neutral","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_2":"neutral","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_3":"neutral","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_0":"neutral","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_1":"neutral","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_2":"neutral","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3":"neutral","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4":"neutral","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_5":"neutral","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_6":"neutral","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_7":"neutral","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_8":"neutral","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_9":"neutral","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_10":"neutral","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_11":"neutral","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_0":"neutral","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_1":"neutral","pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_0":"neutral","pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_1":"neutral","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_0":"neutral","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_1":"neutral","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_2":"neutral","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_3":"neutral","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_0":"neutral","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_1":"neutral","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_2":"neutral","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3":"neutral","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4":"neutral","pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_0":"neutral","pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_1":"neutral","pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_2":"neutral","pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0":"neutral","pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_1":"neutral","pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_2":"neutral","pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_0":"neutral","pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_1":"neutral","pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_2":"neutral"},"next_color_idx":29,"wires_placed_in_order":[["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_4","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_22"],["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_3","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_21"],["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_2","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_20"],["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_19"],["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_10"],["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_8"],["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_9","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23"],["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_25"],["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_12","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_29"],["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_0"],["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_1"],["pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_2","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28"],["pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_3","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27"],["pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_2","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4"],["pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_0"],["pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1"],["pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_1"],["pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_0"],["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_1","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_2"],["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_5","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_3"],["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18"],["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17"],["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4","pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_2"],["pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17"],["pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18"],["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3","pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_2"],["pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17"],["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_26","pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_1"],["pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_0","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_0"],["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_1"],["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28"],["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27"],["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27"],["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_4","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_22"]]],[[],[["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_3","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_21"]]],[[],[["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_2","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_20"]]],[[],[["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_19"]]],[[],[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_10"]]],[[],[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_8"]]],[[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_8"]],[]],[[],[["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_9","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23"]]],[[],[["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_25"]]],[[],[["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_12","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_29"]]],[[],[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_0"]]],[[],[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_1"]]],[[],[["pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_2","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28"]]],[[],[["pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_3","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27"]]],[[],[["pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_2","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4"]]],[[],[["pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_0"]]],[[],[["pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1"]]],[[],[["pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_1"]]],[[],[["pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_0"]]],[[],[["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_1","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_2"]]],[[],[["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_5","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_3"]]],[[],[["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18"]]],[[],[["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17"]]],[[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3"]],[]],[[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4"]],[]],[[],[["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4","pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_2"]]],[[],[["pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17"]]],[[["pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17"]],[]],[[],[["pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18"]]],[[],[["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3","pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_2"]]],[[],[["pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17"]]],[[],[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_26","pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_1"]]],[[],[["pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_0","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_0"]]],[[],[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_1"]]],[[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_3"]],[]],[[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_2"]],[]],[[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_19","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1"]],[]],[[],[["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28"]]],[[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_25","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11"]],[]],[[],[["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27"]]],[[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11"]],[]],[[["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1"]],[]],[[],[["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27"]]],[[],[["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_0":"_","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1":"0000000000000003","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_2":"0000000000000002","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_3":"0000000000000001","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_4":"0000000000000000","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_5":"_","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_6":"_","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_7":"_","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_8":"_","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_9":"0000000000000005","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_10":"0000000000000004","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11":"0000000000000006","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_12":"0000000000000007","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_13":"_","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_14":"_","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_15":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_0":"0000000000000011","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1":"0000000000000012","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_2":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_3":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_4":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_5":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_6":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_7":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_8":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_9":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_10":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_11":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_12":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_13":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_14":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_15":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_16":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17":"0000000000000018","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18":"0000000000000016","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_19":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_20":"0000000000000002","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_21":"0000000000000001","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_22":"0000000000000000","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23":"0000000000000005","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24":"0000000000000004","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_25":"_","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_26":"0000000000000019","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27":"0000000000000003","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28":"0000000000000006","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_29":"0000000000000007","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_0":"0000000000000005","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_1":"0000000000000004","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_2":"_","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_3":"_","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_0":"_","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_1":"0000000000000013","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_2":"_","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3":"0000000000000017","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4":"0000000000000015","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_5":"0000000000000014","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_6":"_","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_7":"_","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_8":"_","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_9":"_","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_10":"_","pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_11":"_","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_0":"0000000000000020","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_1":"0000000000000012","pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_0":"0000000000000020","pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_1":"0000000000000019","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_0":"0000000000000012","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_1":"0000000000000010","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_2":"0000000000000013","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_3":"0000000000000014","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_0":"_","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_1":"_","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_2":"_","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3":"0000000000000012","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4":"0000000000000010","pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_0":"0000000000000011","pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_1":"_","pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_2":"0000000000000010","pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0":"0000000000000016","pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_1":"_","pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_2":"0000000000000015","pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_0":"0000000000000018","pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_1":"_","pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_2":"0000000000000017"},"component_id_to_pins":{"c22d4b25-2814-4177-aa63-9deb5a414cad":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15"],"a3fee46c-a59d-48f1-92de-07521e484019":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29"],"bda6b162-0205-4660-bfa2-67789d801a22":["0","1","2","3"],"f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14":["0","1","2","3","4","5","6","7","8","9","10","11"],"f69d84f3-86e0-4ae5-b3df-45f565ec0def":["0","1"],"40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0":["0","1"],"834400c7-6892-4443-abed-984a8d61dc5a":["0","1","2","3"],"e7dce2a0-b706-44b4-a0b4-b091b9fc73cb":["0","1","2","3","4"],"a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5":["0","1","2"],"9009a5c3-2860-4512-9fb9-18d8067446e4":["0","1","2"],"575981ea-87a6-452f-b72c-c25c47ad5693":["0","1","2"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_4","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_22"],"0000000000000001":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_3","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_21"],"0000000000000002":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_2","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_20"],"0000000000000004":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_10","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_1"],"0000000000000005":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23","pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_9","pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_0"],"0000000000000007":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_12","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_29"],"0000000000000010":["pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_2","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_1"],"0000000000000011":["pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_0"],"0000000000000012":["pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1","pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_1"],"0000000000000013":["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_1","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_2"],"0000000000000014":["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_5","pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_3"],"0000000000000015":["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4","pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_2"],"0000000000000016":["pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18"],"0000000000000017":["pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3","pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_2"],"0000000000000018":["pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_0","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17"],"0000000000000019":["pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_26","pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_1"],"0000000000000020":["pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_0","pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_0"],"0000000000000003":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27"],"0000000000000006":["pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11","pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000007":"Net 7","0000000000000010":"Net 10","0000000000000011":"Net 11","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000014":"Net 14","0000000000000015":"Net 15","0000000000000016":"Net 16","0000000000000017":"Net 17","0000000000000018":"Net 18","0000000000000019":"Net 19","0000000000000020":"Net 20","0000000000000003":"Net 3","0000000000000006":"Net 6"},"all_breadboard_info_list":[],"breadboard_info_list":[],"componentsData":[{"compProperties":{},"position":[74.31793149999986,440.08338049999986],"typeId":"ea67bc39-2543-48d1-915c-5686eed5bac4","componentVersion":1,"instanceId":"c22d4b25-2814-4177-aa63-9deb5a414cad","orientation":"up","circleData":[[122.5,440],[122.64999999999998,450.5],[122.5,460.4],[122.94999999999993,471.04999999999995],[122.94999999999993,481.40000000000003],[122.79999999999995,492.19999999999993],[122.04999999999995,512.8999999999996],[122.34999999999991,501.64999999999986],[19.449999999999832,440.29999999999995],[19.449999999999832,450.35],[19.449999999999832,460.4],[19.449999999999832,470.9],[19.449999999999832,481.7],[19.449999999999832,491.6],[19.449999999999832,502.39999999999986],[19.449999999999832,513.0499999999995]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[294.1861825,665.8400614999999],"typeId":"26347ed3-a6fe-40ba-bac1-eb0320e06540","componentVersion":1,"instanceId":"a3fee46c-a59d-48f1-92de-07521e484019","orientation":"left","circleData":[[362.5,560],[362.5,574.9999999999999],[362.5,589.9999999999999],[362.5,604.9999999999999],[362.5,619.9999999999999],[362.5,634.9999999999999],[362.5,649.9999999999999],[362.5,664.9999999999999],[362.5,679.9999999999999],[362.5,694.9999999999999],[362.5,709.9999999999999],[362.5,724.9999999999999],[362.5,739.9999999999999],[362.5,754.9999999999999],[362.5,769.9999999999999],[227.5,560],[227.5,574.9999999999999],[227.5,589.9999999999999],[227.5,604.9999999999999],[227.5,619.9999999999999],[227.5,634.9999999999999],[227.5,649.9999999999999],[227.5,664.9999999999999],[227.5,679.9999999999999],[227.5,694.9999999999999],[227.5,709.9999999999999],[227.5,724.9999999999999],[227.5,739.9999999999999],[227.5,754.9999999999999],[227.5,769.9999999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[55.48029399999997,916.2790489999998],"typeId":"092faa81-5159-4edd-9101-4b5e9190799a","componentVersion":1,"instanceId":"bda6b162-0205-4660-bfa2-67789d801a22","orientation":"up","circleData":[[32.500000000000014,845],[47.500000000000014,845],[62.500000000000014,844.85],[77.50000000000001,844.85]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[746.9887495000004,909.1916015000005],"typeId":"57a52ffb-0cf9-41cf-991c-9b8593978531","componentVersion":1,"instanceId":"f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14","orientation":"right","circleData":[[781.1803510000004,854.7028520000001],[768.4873510000004,854.7028520000003],[755.7943510000005,853.6138520000004],[742.7383510000002,853.9768520000002],[730.4083510000002,854.3398520000005],[717.850351,854.3398520000005],[767.3893510000005,960.9613520000003],[754.6963510000005,960.9613520000003],[743.0908510000003,960.2368520000005],[730.034851,960.5998520000003],[717.3898509999999,960.5998520000003],[704.6953509999997,960.5998520000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[311.20404699999995,921.7023425000004],"typeId":"bef26dfc-4265-9461-6fdb-ad28abcdc659","componentVersion":1,"instanceId":"f69d84f3-86e0-4ae5-b3df-45f565ec0def","orientation":"up","circleData":[[287.5,965.0000000000003],[332.44937349999987,965.0000570000005]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"HLMP-3762","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Broadcom","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[219.16975000000002,853.2927500000005],"typeId":"82d731d1-c75f-e131-c68f-ff0e81dc6210","componentVersion":1,"instanceId":"40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0","orientation":"up","circleData":[[212.5,935],[227.5045,935]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[727.5000340000006,614.9999615000006],"typeId":"da65b43a-b07b-4269-9c87-2ed695c925da","componentVersion":1,"instanceId":"834400c7-6892-4443-abed-984a8d61dc5a","orientation":"right","circleData":[[782.5,470],[670.0000000000005,470],[670.0000000000006,762.5000000000007],[782.5,755.0000000000007]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[548.4687384999995,284.3815789999999],"typeId":"646c8823-36b2-4192-89ce-6ec44eb47b6e","componentVersion":1,"instanceId":"e7dce2a0-b706-44b4-a0b4-b091b9fc73cb","orientation":"up","circleData":[[497.5,395],[520,395],[542.5,395],[565,395],[587.4999999999994,395]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[455.0457745,492.29286349999984],"typeId":"bbb07cdc-963b-4f77-8585-9aff4347bf37","componentVersion":2,"instanceId":"a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5","orientation":"up","circleData":[[437.5,514.9999999999998],[467.5,514.9999999999998],[452.5,514.9999999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[455.0457745,747.2928634999998],"typeId":"bbb07cdc-963b-4f77-8585-9aff4347bf37","componentVersion":2,"instanceId":"9009a5c3-2860-4512-9fb9-18d8067446e4","orientation":"up","circleData":[[437.5,769.9999999999999],[467.5,769.9999999999999],[452.5,769.9999999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[455.0457745,867.2928634999998],"typeId":"bbb07cdc-963b-4f77-8585-9aff4347bf37","componentVersion":2,"instanceId":"575981ea-87a6-452f-b72c-c25c47ad5693","orientation":"up","circleData":[[437.5,889.9999999999999],[467.4999999999999,889.9999999999999],[452.5,889.9999999999999]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"132.78623","left":"-36.84623","width":"853.25223","height":"876.20049","x":"-36.84623","y":"132.78623"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_22\",\"endPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_4\",\"rawStartPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_22\",\"rawEndPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5000000000_665.0000000000\\\",\\\"160.0000000000_665.0000000000\\\",\\\"160.0000000000_481.4000000000\\\",\\\"122.9500000000_481.4000000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_21\",\"endPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_3\",\"rawStartPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_21\",\"rawEndPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5000000000_650.0000000000\\\",\\\"167.5000000000_650.0000000000\\\",\\\"167.5000000000_471.0500000000\\\",\\\"122.9500000000_471.0500000000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_20\",\"endPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_2\",\"rawStartPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_20\",\"rawEndPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5000000000_635.0000000000\\\",\\\"175.0000000000_635.0000000000\\\",\\\"175.0000000000_460.4000000000\\\",\\\"122.5000000000_460.4000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24\",\"endPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_10\",\"rawStartPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24\",\"rawEndPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_10\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5000000000_695.0000000000\\\",\\\"-42.5000000000_695.0000000000\\\",\\\"-42.5000000000_460.4000000000\\\",\\\"19.4500000000_460.4000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24\",\"endPinId\":\"pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_1\",\"rawStartPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_24\",\"rawEndPinId\":\"pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5000000000_695.0000000000\\\",\\\"47.5000000000_695.0000000000\\\",\\\"47.5000000000_845.0000000000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23\",\"endPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_9\",\"rawStartPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23\",\"rawEndPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5000000000_680.0000000000\\\",\\\"-50.0000000000_680.0000000000\\\",\\\"-50.0000000000_450.3500000000\\\",\\\"19.4500000000_450.3500000000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23\",\"endPinId\":\"pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_0\",\"rawStartPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_23\",\"rawEndPinId\":\"pin-type-component_bda6b162-0205-4660-bfa2-67789d801a22_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5000000000_680.0000000000\\\",\\\"32.5000000000_680.0000000000\\\",\\\"32.5000000000_845.0000000000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_29\",\"endPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_12\",\"rawStartPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_29\",\"rawEndPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_12\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5000000000_770.0000000000\\\",\\\"-27.5000000000_770.0000000000\\\",\\\"-27.5000000000_481.7000000000\\\",\\\"19.4500000000_481.7000000000\\\"]}\"}","{\"color\":\"#00AE7E\",\"startPinId\":\"pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_2\",\"endPinId\":\"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4\",\"rawStartPinId\":\"pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_2\",\"rawEndPinId\":\"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"452.5000000000_515.0000000000\\\",\\\"452.5000000000_545.0000000000\\\",\\\"587.5000000000_545.0000000000\\\",\\\"587.5000000000_395.0000000000\\\"]}\"}","{\"color\":\"#00AE7E\",\"startPinId\":\"pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_1\",\"endPinId\":\"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4\",\"rawStartPinId\":\"pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_1\",\"rawEndPinId\":\"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"670.0000000000_470.0000000000\\\",\\\"587.5000000000_470.0000000000\\\",\\\"587.5000000000_395.0000000000\\\"]}\"}","{\"color\":\"#C28C9F\",\"startPinId\":\"pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_0\",\"endPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_0\",\"rawStartPinId\":\"pin-type-component_a3b8ab88-13f5-48e0-9a75-f72ccc0a5cb5_0\",\"rawEndPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"437.5000000000_515.0000000000\\\",\\\"437.5000000000_560.0000000000\\\",\\\"362.5000000000_560.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1\",\"endPinId\":\"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3\",\"rawStartPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1\",\"rawEndPinId\":\"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"362.5000000000_575.0000000000\\\",\\\"565.0000000000_575.0000000000\\\",\\\"565.0000000000_395.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_0\",\"endPinId\":\"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3\",\"rawStartPinId\":\"pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_0\",\"rawEndPinId\":\"pin-type-component_e7dce2a0-b706-44b4-a0b4-b091b9fc73cb_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"782.5000000000_470.0000000000\\\",\\\"782.5000000000_440.0000000000\\\",\\\"565.0000000000_440.0000000000\\\",\\\"565.0000000000_395.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1\",\"endPinId\":\"pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_1\",\"rawStartPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_1\",\"rawEndPinId\":\"pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"362.5000000000_575.0000000000\\\",\\\"415.0000000000_575.0000000000\\\",\\\"415.0000000000_980.0000000000\\\",\\\"332.4493735000_980.0000000000\\\",\\\"332.4493735000_965.0000570000\\\"]}\"}","{\"color\":\"#5FAD4E\",\"startPinId\":\"pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_2\",\"endPinId\":\"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_1\",\"rawStartPinId\":\"pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_2\",\"rawEndPinId\":\"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"670.0000000000_762.5000000000\\\",\\\"647.5000000000_762.5000000000\\\",\\\"647.5000000000_815.0000000000\\\",\\\"768.4873510000_815.0000000000\\\",\\\"768.4873510000_854.7028520000\\\"]}\"}","{\"color\":\"#FF029D\",\"startPinId\":\"pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_3\",\"endPinId\":\"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_5\",\"rawStartPinId\":\"pin-type-component_834400c7-6892-4443-abed-984a8d61dc5a_3\",\"rawEndPinId\":\"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"782.5000000000_755.0000000000\\\",\\\"812.5000000000_755.0000000000\\\",\\\"812.5000000000_800.0000000000\\\",\\\"715.0000000000_800.0000000000\\\",\\\"715.0000000000_854.3398520000\\\",\\\"717.8503510000_854.3398520000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_2\",\"endPinId\":\"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4\",\"rawStartPinId\":\"pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_2\",\"rawEndPinId\":\"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"452.5000000000_770.0000000000\\\",\\\"452.5000000000_830.0000000000\\\",\\\"730.4083510000_830.0000000000\\\",\\\"730.4083510000_854.3398520000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0\",\"endPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18\",\"rawStartPinId\":\"pin-type-component_9009a5c3-2860-4512-9fb9-18d8067446e4_0\",\"rawEndPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_18\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"437.5000000000_770.0000000000\\\",\\\"392.5000000000_770.0000000000\\\",\\\"392.5000000000_507.5000000000\\\",\\\"205.0000000000_507.5000000000\\\",\\\"205.0000000000_605.0000000000\\\",\\\"227.5000000000_605.0000000000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_2\",\"endPinId\":\"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3\",\"rawStartPinId\":\"pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_2\",\"rawEndPinId\":\"pin-type-component_f3a4d962-4b38-4c9f-8e2e-685a8c3e7f14_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"452.5000000000_890.0000000000\\\",\\\"452.5000000000_920.0000000000\\\",\\\"602.5000000000_920.0000000000\\\",\\\"602.5000000000_837.5000000000\\\",\\\"742.7383510000_837.5000000000\\\",\\\"742.7383510000_853.9768520000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_0\",\"endPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17\",\"rawStartPinId\":\"pin-type-component_575981ea-87a6-452f-b72c-c25c47ad5693_0\",\"rawEndPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_17\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"437.5000000000_890.0000000000\\\",\\\"377.5000000000_890.0000000000\\\",\\\"377.5000000000_492.5000000000\\\",\\\"197.5000000000_492.5000000000\\\",\\\"197.5000000000_590.0000000000\\\",\\\"227.5000000000_590.0000000000\\\"]}\"}","{\"color\":\"#BDC6FF\",\"startPinId\":\"pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_1\",\"endPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_26\",\"rawStartPinId\":\"pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_1\",\"rawEndPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_26\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5045000000_935.0000000000\\\",\\\"227.5045000000_950.0000000000\\\",\\\"182.5000000000_950.0000000000\\\",\\\"182.5000000000_725.0000000000\\\",\\\"227.5000000000_725.0000000000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_0\",\"endPinId\":\"pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_0\",\"rawStartPinId\":\"pin-type-component_40badbb5-58f7-41cf-a0db-2f1fbd8aa7e0_0\",\"rawEndPinId\":\"pin-type-component_f69d84f3-86e0-4ae5-b3df-45f565ec0def_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"212.5000000000_935.0000000000\\\",\\\"212.5000000000_980.0000000000\\\",\\\"287.5000000000_980.0000000000\\\",\\\"287.5000000000_965.0000000000\\\"]}\"}","{\"color\":\"#e8176b\",\"startPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27\",\"endPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1\",\"rawStartPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_27\",\"rawEndPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5000000000_740.0000000000\\\",\\\"182.5000000000_740.0000000000\\\",\\\"182.5000000000_450.5000000000\\\",\\\"122.6500000000_450.5000000000\\\"]}\"}","{\"color\":\"#774D00\",\"startPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28\",\"endPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11\",\"rawStartPinId\":\"pin-type-component_a3fee46c-a59d-48f1-92de-07521e484019_28\",\"rawEndPinId\":\"pin-type-component_c22d4b25-2814-4177-aa63-9deb5a414cad_11\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5000000000_755.0000000000\\\",\\\"-12.5000000000_755.0000000000\\\",\\\"-12.5000000000_470.9000000000\\\",\\\"19.4500000000_470.9000000000\\\"]}\"}"],"projectDescription":""}PK
     ��Z               jsons/PK
     ��Z|�%3  %3     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"LoRa Ra-02 SX1278","category":["User Defined"],"id":"ea67bc39-2543-48d1-915c-5686eed5bac4","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"ae1d0bb1-db79-4eca-b526-eb1d648f9ad0.png","iconPic":"1348d1eb-e6ae-43d4-937f-d455f2ad4bcd.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.31437","numDisplayRows":"12.64394","pins":[{"uniquePinIdString":"0","positionMil":"786.93229,632.75287","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"787.93229,562.75287","isAnchorPin":false,"label":"NSS"},{"uniquePinIdString":"2","positionMil":"786.93229,496.75287","isAnchorPin":false,"label":"MOSI"},{"uniquePinIdString":"3","positionMil":"789.93229,425.75287","isAnchorPin":false,"label":"MISO"},{"uniquePinIdString":"4","positionMil":"789.93229,356.75287","isAnchorPin":false,"label":"SCK"},{"uniquePinIdString":"5","positionMil":"788.93229,284.75287","isAnchorPin":false,"label":"D105"},{"uniquePinIdString":"6","positionMil":"783.93229,146.75287","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"785.93229,221.75287","isAnchorPin":false,"label":"DI04"},{"uniquePinIdString":"8","positionMil":"99.93229,630.75287","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"9","positionMil":"99.93229,563.75287","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"10","positionMil":"99.93229,496.75287","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"11","positionMil":"99.93229,426.75287","isAnchorPin":false,"label":"RST"},{"uniquePinIdString":"12","positionMil":"99.93229,354.75287","isAnchorPin":false,"label":"DI00"},{"uniquePinIdString":"13","positionMil":"99.93229,288.75287","isAnchorPin":false,"label":"DI01"},{"uniquePinIdString":"14","positionMil":"99.93229,216.75287","isAnchorPin":false,"label":"D102"},{"uniquePinIdString":"15","positionMil":"99.93229,145.75287","isAnchorPin":false,"label":"DI03"}],"pinType":"wired"},"properties":[]},{"subtypeName":"NodeMCU","category":["User Defined"],"id":"26347ed3-a6fe-40ba-bac1-eb0320e06540","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"0795b188-35ce-4b4d-8dd5-08667f88bf32.png","iconPic":"28e7f2ff-99bf-41f5-8f78-c92be5544a69.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"18.89764","numDisplayRows":"9.84252","pins":[{"uniquePinIdString":"0","positionMil":"1650.48241,36.70055","isAnchorPin":true,"label":"Vin"},{"uniquePinIdString":"1","positionMil":"1550.48241,36.70055","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"1450.48241,36.70055","isAnchorPin":false,"label":"RST"},{"uniquePinIdString":"3","positionMil":"1350.48241,36.70055","isAnchorPin":false,"label":"EN"},{"uniquePinIdString":"4","positionMil":"1250.48241,36.70055","isAnchorPin":false,"label":"3V§"},{"uniquePinIdString":"5","positionMil":"1150.48241,36.70055","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1050.48241,36.70055","isAnchorPin":false,"label":"CLK"},{"uniquePinIdString":"7","positionMil":"950.48241,36.70055","isAnchorPin":false,"label":"SDO"},{"uniquePinIdString":"8","positionMil":"850.48241,36.70055","isAnchorPin":false,"label":"CWD"},{"uniquePinIdString":"9","positionMil":"750.48241,36.70055","isAnchorPin":false,"label":"SD1"},{"uniquePinIdString":"10","positionMil":"650.48241,36.70055","isAnchorPin":false,"label":"SD2"},{"uniquePinIdString":"11","positionMil":"550.48241,36.70055","isAnchorPin":false,"label":"SD3"},{"uniquePinIdString":"12","positionMil":"450.48241,36.70055","isAnchorPin":false,"label":"RSU"},{"uniquePinIdString":"13","positionMil":"350.48241,36.70055","isAnchorPin":false,"label":"RSV"},{"uniquePinIdString":"14","positionMil":"250.48241,36.70055","isAnchorPin":false,"label":"AO"},{"uniquePinIdString":"15","positionMil":"1650.48241,936.70055","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"16","positionMil":"1550.48241,936.70055","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"17","positionMil":"1450.48241,936.70055","isAnchorPin":false,"label":"TX"},{"uniquePinIdString":"18","positionMil":"1350.48241,936.70055","isAnchorPin":false,"label":"RX"},{"uniquePinIdString":"19","positionMil":"1250.48241,936.70055","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"20","positionMil":"1150.48241,936.70055","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"21","positionMil":"1050.48241,936.70055","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"22","positionMil":"950.48241,936.70055","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"23","positionMil":"850.48241,936.70055","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"24","positionMil":"750.48241,936.70055","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"25","positionMil":"650.48241,936.70055","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"26","positionMil":"550.48241,936.70055","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"27","positionMil":"450.48241,936.70055","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"28","positionMil":"350.48241,936.70055","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"29","positionMil":"250.48241,936.70055","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"properties":[]},{"subtypeName":"0.96\" OLED","category":["User Defined"],"id":"092faa81-5159-4edd-9101-4b5e9190799a","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"8d902f4e-ab09-4493-932a-1f1db25b6d7d.png","iconPic":"4c416a15-58ad-47dc-949c-f0bec13a5bfd.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.97687","numDisplayRows":"11.02769","pins":[{"uniquePinIdString":"0","positionMil":"395.64154,1026.57816","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"495.64154,1026.57816","isAnchorPin":false,"label":"VDD"},{"uniquePinIdString":"2","positionMil":"595.64154,1027.57816","isAnchorPin":false,"label":"SCK"},{"uniquePinIdString":"3","positionMil":"695.64154,1027.57816","isAnchorPin":false,"label":"SDA"}],"pinType":"wired"},"properties":[]},{"subtypeName":"SIM800L","category":["User Defined"],"id":"57a52ffb-0cf9-41cf-991c-9b8593978531","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"b5c34fc0-5882-471e-a80e-5adb517f5654.png","iconPic":"5f4f8fc5-f884-4b46-b794-7d87214b037b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.90730","numDisplayRows":"7.92230","pins":[{"uniquePinIdString":"0","positionMil":"132.10667,624.05901","isAnchorPin":true,"label":"NET"},{"uniquePinIdString":"1","positionMil":"132.10667,539.43901","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"124.84667,454.81901","isAnchorPin":false,"label":"RST"},{"uniquePinIdString":"3","positionMil":"127.26667,367.77901","isAnchorPin":false,"label":"RXD"},{"uniquePinIdString":"4","positionMil":"129.68667,285.57901","isAnchorPin":false,"label":"TXD"},{"uniquePinIdString":"5","positionMil":"129.68667,201.85901","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"840.49667,532.11901","isAnchorPin":false,"label":"RING"},{"uniquePinIdString":"7","positionMil":"840.49667,447.49901","isAnchorPin":false,"label":"DTR"},{"uniquePinIdString":"8","positionMil":"835.66667,370.12901","isAnchorPin":false,"label":"MIC+"},{"uniquePinIdString":"9","positionMil":"838.08667,283.08901","isAnchorPin":false,"label":"MIC-"},{"uniquePinIdString":"10","positionMil":"838.08667,198.78901","isAnchorPin":false,"label":"SPK+"},{"uniquePinIdString":"11","positionMil":"838.08667,114.15901","isAnchorPin":false,"label":"SPK-"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Piezo Buzzer","category":["Output"],"userDefined":true,"id":"bef26dfc-4265-9461-6fdb-ad28abcdc659","subtypeDescription":"","subtypePic":"36e83e0e-fd9a-4553-9782-762f273f5010.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"5.16729","numDisplayRows":"5.97302","pins":[{"uniquePinIdString":"0","positionMil":"100.33752,9.99995","isAnchorPin":true,"label":"pin 1"},{"uniquePinIdString":"1","positionMil":"400.00001,9.99957","isAnchorPin":false,"label":"pin 2"}],"pinType":"wired"},"properties":[],"iconPic":"edd00682-873b-4230-8bb4-282089490c70.png","componentVersion":1},{"subtypeName":"LED: Two Pin (red)","subtypeDescription":"","id":"82d731d1-c75f-e131-c68f-ff0e81dc6210","category":["Output"],"userDefined":false,"subtypePic":"da48ab5c-24bb-4ba8-ab59-39208c7b2ba2.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"62.87000,0.00000","endPositionMil":"62.87000,-341.89000","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"162.90000,0.00000","endPositionMil":"162.90000,-341.89000","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"2.14670","numDisplayRows":"4.05650","pinType":"movable"},"properties":[{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"b96c8ad8-7845-422d-b49f-326b2968fdb8.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"DC-DC Buck XL4015 5A","category":["User Defined"],"id":"da65b43a-b07b-4269-9c87-2ed695c925da","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"14f4e0bc-85be-4a63-979f-9a3c78ebf9d5.png","iconPic":"78e6be4d-468b-4075-9957-5b4cf1a5366b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"21.25984","numDisplayRows":"9.05512","pins":[{"uniquePinIdString":"0","positionMil":"96.32559,819.42244","isAnchorPin":true,"label":"OUT -"},{"uniquePinIdString":"1","positionMil":"96.32559,69.42244","isAnchorPin":false,"label":"OUT +"},{"uniquePinIdString":"2","positionMil":"2046.32559,69.42244","isAnchorPin":false,"label":"IN +"},{"uniquePinIdString":"3","positionMil":"1996.32559,819.42244","isAnchorPin":false,"label":"IN -"}],"pinType":"wired"},"properties":[]},{"subtypeName":"POWER SUPPLY 5V 5AMP","category":["User Defined"],"id":"646c8823-36b2-4192-89ce-6ec44eb47b6e","userDefined":true,"subtypeDescription":"","subtypePic":"483af35d-09f4-402a-a8a9-75c28eb4643f.png","pinInfo":{"numDisplayCols":"13.51513","numDisplayRows":"18.87938","pins":[{"uniquePinIdString":"0","positionMil":"335.96491,206.51286","isAnchorPin":true,"label":"220V Positive Pole (AC)"},{"uniquePinIdString":"1","positionMil":"485.96491,206.51286","isAnchorPin":false,"label":"220V Negative Pole (AC)"},{"uniquePinIdString":"2","positionMil":"635.96491,206.51286","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"3","positionMil":"785.96491,206.51286","isAnchorPin":false,"label":"GND (DC)"},{"uniquePinIdString":"4","positionMil":"935.96491,206.51286","isAnchorPin":false,"label":"12V-24V Output (DC)"}],"pinType":"wired"},"properties":[],"iconPic":"0a03a94b-1490-4d51-a356-eaee23e4f5f0.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Potentiometer","category":["User Defined"],"id":"bbb07cdc-963b-4f77-8585-9aff4347bf37","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"0c8b7e0a-6698-412e-96f2-fdf086dc4925.png","iconPic":"457643d0-fb24-4111-9541-c1c501ab524b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"5.00000","pins":[{"uniquePinIdString":"0","positionMil":"33.02817,98.61909","isAnchorPin":true,"label":"5V"},{"uniquePinIdString":"1","positionMil":"233.02817,98.61909","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"133.02817,98.61909","isAnchorPin":false,"label":"SIG"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Potentiometer","category":["User Defined"],"id":"bbb07cdc-963b-4f77-8585-9aff4347bf37","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"0c8b7e0a-6698-412e-96f2-fdf086dc4925.png","iconPic":"457643d0-fb24-4111-9541-c1c501ab524b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"5.00000","pins":[{"uniquePinIdString":"0","positionMil":"33.02817,98.61909","isAnchorPin":true,"label":"5V"},{"uniquePinIdString":"1","positionMil":"233.02817,98.61909","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"133.02817,98.61909","isAnchorPin":false,"label":"SIG"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Potentiometer","category":["User Defined"],"id":"bbb07cdc-963b-4f77-8585-9aff4347bf37","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"0c8b7e0a-6698-412e-96f2-fdf086dc4925.png","iconPic":"457643d0-fb24-4111-9541-c1c501ab524b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.00000","numDisplayRows":"5.00000","pins":[{"uniquePinIdString":"0","positionMil":"33.02817,98.61909","isAnchorPin":true,"label":"5V"},{"uniquePinIdString":"1","positionMil":"233.02817,98.61909","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"133.02817,98.61909","isAnchorPin":false,"label":"SIG"}],"pinType":"wired"},"properties":[]}]}PK
     ��Z               images/PK
     ��Z�U ��  ��  /   images/ae1d0bb1-db79-4eca-b526-eb1d648f9ad0.png�PNG

   IHDR   �  ,   G}�   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  �VIDATx^����yލ���[���+Q	� ���R)�jVq��/����|v�=�K9�c�D�-KV�%Q�DR,b�������~�g�C$!	.�>/0w�����μ�[�m��lZ�:ԡ�[�u�C? ꀮC�St���:��P�~��]�:���:ԡ0u@ס���3N7��R�'��f��h���F��lFM�BF#5uR��H(T��C�D$R����D�M�T��c�O6�٬�Y�n�yD��:�e��`u](�XT�������������ޡ��:���T�Vs�J�w4r]�&�l�����H�	a��($ �_���
�ڬ���Ԅ�d�lX�?7P��^&vuhZSt���z|��ԇ�]]��
���WT�Q�W�ba�h#j�:�k��<�|�h���M�g!�<P3���f�?H�\�M[�t�\ *�G���U�Y�m�,Y�X����Z$!c2��IY̒:OF�;�D,b�$!j=�KH��J=6��~�^1�l^�J�CӘ:���j<��d�?we��zF(���5�V�؞����		l��\�i���5e_���.\�|�%cqK������R}_#~fy����������r���]	�M_:|����MY�+k�������V(��0�w�d���)��t��׋ѝٴw�����Q���[=�c��`!f{���o�D��.�MK��P�R�>�~q �:V�Y*�ᓃ�����/~����K27!kԛt�ȻY3�]�zz�w~�?���|�U�!���#a;8P�o�E����4��Ow��hD�uKqY<&-V+[$���Y$�_��\�R��%�	K�Jƭ+���D�rф�jf������E�4��.�X����th�Rt�����Z�^��w��tlX:��;�u����W����%�T*2E�VmT�)��j��gՊ��[�˷X]�fR��4k����5�A.���� Y��PȤ�8oZ��x�p&q�^��#φ]��LO�tM��(�Mc����BqŢ�S����������A�T �#�-��W��{�g��b��tr6��N�Ns�4Ѕ��87�����.
�K�k<�� E��WŅ� N��CӒ:��@4j��E"������3D8:(����~�m޼ٙ��d�ݗ�lv7���@^�A��k�v����k5l>��&bzf�M�9u��`^B�Hԁ�V���ؘ������8q���Ƀ��������O:-Y.���t��4��.	p�f�U>Z*�H8�tww;`$�q�@�H\�a^f2K�ӧz.�d]�n�St�b��U��A�j��͛go}�[mѢEX #��^z3��[o��7Z�Zq�!�R��9u@waȩ&��5@q ��D�q��C���9Z,�}Һ��^tӜ:�� $ 5+�F3
;�E�qv~ڑ#G�<�ځ�zօ��߾��o[<wi����uh�Rt��ѐ4S�M��ܸ�ܹs]�\ �����q֬Y��f�5�#י�������.5��P�J��&��1�O����4 �l���ݶm�lÆn���L�!v@7ݩ�@�z�� � ��xৡ���Ld�X>�w�P�:�� B��-u@w��$��OW,,�YA`c�%�)h�z���)�NH�����{��-�JN#v�\��"���
E�-�q�� �\`��E&y)*�z��LV���4c��u@w!(j�Z�� V�Vl``���]wْ%K� ��Q�9�0�a�9۴i��v�mڴ)����kJ#���l�ҡiM�]8r�\P�\��{�����)M�z��~g�b~�D���Q�Mw���*��NLJ:Q>��O�q:��&?V��:O �_�j0N��Y)�B�̜��݅��Sr�� $�\�֭[g����oD+W��I:�Ι�	@�40w�Cә:��@�ղ�j ���;�í��f��#�B��^q�v�%�8-��g�8��������.�[��hjj�v���|:���ٳǆ��`���i�uh�St��P�ѴT,����b�X~�_tGz$�ȧ{��쥗^r�.�b����uT�4��.	7!z1!#",���H����MK��òe�l����x�`�A��;u@w��%�p0N�*�R�h���ΧHL	�@����-���:^ �b>���K����$ Cw2�r[�}��_�C��!��Q;��~�W^q u+DhN�ӦӜ:t��Vo���~���� ���?j�	���f����z����wj@��F�ceNs��BP�Bl�P�W-��8�����9�"g%��˗������$E	�X��5u�Q�ѰD$f�f��X����]w�e�ׯw=�gj6�� �_{�v�嗻�]�.w�=�t��4�N]0
P�l�L6����}�M�TD�����v��14�嫬HP�N�Ns�4��h�O\U�i٨T�y���ϸ�Rb�h06W?=>�Ǒ��/�����L��o���)��i�iN��@T�0/��K��.�x����w�t *P���+�_���[�x����T�`x�MvhZRt�2�p�����R,Zwwή��Ɔ�ui>��t���o�XK��K?�N�u�t�S��.��L�T�FGǝO��'lVۧ���o���=>� �y��tӜ:��@�0m+�z*!4~�1�Z{�����] �������F�3�r�St�����H�k
dl�w�u׹-�j��)sӱ=xS�)`.t $|�	+�ˠCӖ:��@���]G
.$pe2)�r�V�10�i�v�y������S{����Ҙ,}��;R�;u@w�h�Xv*	sQ*͎=n������K��<Ӝl\c���>��c{���Y�3��D�3OMn�#d��]nYLE�35���&F�y`�ST ;������J=  B��{��.�=9���6�yr���5�\�U�<{*^rӞ:�� �4b�Lt���)�˯8�(�͜[{���y�"V�ON&&����fXq;4���D�N��l���,��<���n+>z#=2�Ax���7�z:mɵ���;�崧�.5����?v��`�X��/�`i->��p��O�k=��f�0$Zm���|*���.ET���f�	a��;��}π���"�믿�MìdءP,�!A�5C�Cӕ:��@$�LbƟ���Nz!�$h��Z�͆99g�T�x^����:������f��o�w�u�)�;�*��l�z�!{��_�Ҝ�etӜ:�� $T�Ba����8��10��E4���E�� j(��G���8���
���Cng�Mc��B�L�r���S�����8��oD"15L�"!����LP��RS��/a�1ɛo���mXo�rŒ��
�e��:4���ER`�hB����~+���<��6�;�h:�#��ŋ,��c�D�T�F�nu4�4��. 5��� %��ڑ��Y���~�}�����Ӂ�w��ჿ����'�x­2Ǵ��ɔxtӜ:���ڄ���HG
�����611�yy���G߃Y,]R���J͸�h�Ms��ک.G,.�^�Z6�ex��mάY�S����X{�7��� x)a��Mo�����v��"�S)��JfNM�j��'��Zڏ��И�"�P���ج���� ��9��vQ0��!��c��(Q[˃�54��'?�){�ɧ��*����pf(�b��5u@w����9���˱?J!?ٺ$_��<Ei�v>����c�[��ʀG]���� �FF�|:�s�j���v��w;����ͭ1n|?� q��� �Oe�]�n��KF@vhZSt��:1C21陌FB���T��H`c�ߍs ��R��-���:�n�St���j�}�`�b	�r���/|��t�\�����u7���b��~�a�= �h��ŕ\���iO��@�L�CE���F�U�5���_�%�QK��IiB�4��i�=�b�l4�1Z�0\������h8\.խT,�,�H:_��.���F��q>"��g?�`A��,���	��M�
a���\/	w�Ph�E�д%7Vԡ,����Ή�ǖ�w�����Mf,$q���-?9n_��g�gV,�,�X���k���~�����̹mΜ>��
���S1n6�"�⵳3�AN����t���X^�z�\)��dl��W׭]gWm��m&�)��c4Ӿؖ��6^v���ң#F�\a|��B&9\��t��.t�r�����H�kj�b�b�j���F�&�o�T�j�� ��>�5>5n�RѪ��Œf5.)-װ�r�s��h+�MS�������D⿾rb�+u����"����E#qkʅc�"�*���,��	l!�����̪�f�p�y����?�Օ{��|��1u@wi����r���>>�;5����'��+�Ɇ���ӏB�&�l�a��O�ʊ��_�㱩 r��3u@w��7��_,��Jdu)"��pC@�hwkX��ćE#V:+u;��;�O��D���"��.0u�Ӄ�[��z�T��dZ7���8.����)���b4f��Ǎ��:tQPt���P=	UÑH�\�ZE�� n�p�c�AS�R�fa9vRv�H8�z�Cu@w�I&d=� �+�ݴ/,���Y��N5[S�P�c�ݘ��v�"��.0�B�F�Q��&�%S���\۲��3����ζ{u@w�I���F����7�@�L�)C�h@	�� �ա��:��$ �YW���
4��T
��F�i�@����ښz��~�"��	b��tV�qjT�B���ON����M���,hU�p�ˢé�:tPtӁZ�Z!w&�|�9���,�a�
���J���;��"��9�%K��Oz)#��k<h;�܏J�%I��D�Ӊr�QtӀ|��𚎭������c�0��u����S��]��4������\t�իWۿ�w�Ζ.]j�b��}�{���s�{"Ѱ[$��`�=ۡ��:��$���� t�-^��~�g~�/^�Zp��ngf
q.:Q�5�Ltu@7��p܉?6W�ʄ�/�\U��ղ۪/���-䦃E=*׮�T�.�nP���F=T��R*Z�\�F*�FC�h�-Z�[L��9
u���4+���V�h���:���D�5��P�H��yn	�����YHI�p�b�HhHW:�����i@�ӟ>r��'v>��T�&0	F�����@�X���ʊNOj;�M�e_���.Z�.�nЬl��y�������D�x�u�4��F�O�k~�re��}mq&��h下ԡ��:��&4��g����gB��p�\E��B�)-�t�k���t�fs*�H�ҝJuv����iD�d�X=*F�1i9T[í�}��C�j2�r�X"6�,�(��iDukF+�P.$��)a!4���l� '���b6S��EI�M+
1�$̚�ӽ�>"bn���.�P�:�t`�.&�n�@�fa��ϛ�u�Z��s�X\Qq�L&�t�"��5��Tـ�]�3-uEAw�g��EJ���N�l��%�vjo��"��EH�M#oA�	�hZD���w�ʋ�:��F�ر�a�421��Y7^qew�Rtӈ��`��§�ηs�Vઑ`]�C#u@7�H�b%��պ�8���j��bԤ� ]gT����QG��ܜyy��k ��C��K�M'jZ("��m`[&?�C1׫�=>��5`�.>�n�P�}d��N�	Z�՚�%�Ȭ�ts�N;t�Qtӄ [�وDB�HH~�����eX�	�:{5$;t1Qtӈ���Z�ɗV�o�zsCg�g-w�Rtӈda�J(����tt���1�2�h���D�F�R�V��1�r�N�ß;�:���KН#��f3,\Dk�F�Ro$*�z�\��J�z�X�e�j-[l���Z���~MM-(U��H���;h����� .�+����~��$*���fך�J���z$�'&�~�x����;Gp����Qpp��o���D�7��ը7�`�j��NG"��&bk�j,�Z*���O��>�1�����o��&*+$�c���wcw���4;tQtg�4Wr�RY;�}(��l�zju˥#�XѠמ%mT QG) ����Z�k�5�iւs\�'�N�وgj�pTw�kɜ������/|Ѿ���mӕW�P�l�Lfd|����2Bz����6�W�];���̦~8g����L"�r�l�*>O\+W,�"���q>s%u�c��BXל�s����B��C]�fq�CBP�V�V��,�JX�X�w��N;t�}��_��kך�M�b'KS�j]w��H�C��!i�Z�b�#�l�C�ʅB�h!oYk ���X�rBM�L��x�RI�ī��q�A�x�T�k�^=���<f�1��{#Q��y.��T<)�����r�j����k�>���z�-6g�\˗
&_���|:dZE��EFMע���['����7Z�W��U�	;v�];vؑ#G�\,H��mjr<��ǫ���}e@f�!U����n[1��lU���5��rJ�)[�Z+ۃ|���Cvզ�������a�&�+��p�6ش�f
��s�t袢�D�r��?L���
�C��5�i���������m�e�FM�e8f�h�}��l�G���3��9�� �[�6�JB��՝g'��3$W1�XTx�5��n��Z����v��+�T/[Ut�i#C�㿿2����Xl��:tqQt�o��5��7S���x�dIi����'�������3gڝw�iK-p�@h9����_(Ш3�M�,���X�/C�Q@) B=��ɘ]�f��[}���]V+U���J˙�xtf8��Y��.�P�.:�g�J��|nx��fv��o �F�1yѮ��Mv��I��?�#{�[�*�W���P޼D}�� �xgV-qØ��F�t�q�.UdbƢ1k�S�! �=��*��ʁ�?�G�gW�����t#�������^՟����X6�����}����ŏ����o���iF3Pj��,�w��z-=�K��Ѐ�<� 0���<=5�;bZ��M��ev&Vг��[�zd|셩���\10�Tz��;tqRK,��j��ND1�����a;4x��tղ��,�N����H\�'c�TZ��XCGB���D��҂�D�Bɸ�4"��^��cHǨҊ��IuY<�m�d�oc���J'ku����r�'-"�)V>{�ȧ����_2g�t w��?{Mwtl|�x8�����V+W-��������/���۟���iz���"`�RP{N�Xx<���k�f$\>�5i���Kyj�F���Ӫ0��'|ȱ���{!��H�6���z��/�b�����'����@.w��h�.r�n||�x$�����U���H.f���~������??��������ͤ��G�>y�f��<��q5�p($�K@i4#�f�}a�M�+�Z� �Cu> ��J�a��JF ��UR��������ݡ��!'����������|� n/M�7�B���?5-nͿ��ǛUE�W�'�ͱ��ƿ�oph��itB'|7៽O�J�	G��烋���}�PU7'���,���Z3܌F#�h�<١}o��t2�j,�~���|��9b(�hT�6VuOd�Q�`�:�=Rt�p5������b��ꍈ��Ռ�(l��7)>�Q�E��sv�C�;����jn���W$�&����`�@&d�p8����ס}��=�^�sW��ӵf3�dĭM��B�w�n:�1'�t�'ϑ���n��>)���TH����+��ի�|��M��F+4�ءѱ۳�3~ef<��:Q�t&a����e?��?o�W���m�T�f"6v�X~9R����L�ayw��]Z��wk+�w��HO���NmeUD�mt��z���A���O�����ǂ{��p���48����\�*C��C����_u��9�pJ���=�NN�<3���껕���o�GQ�D
�T�*�K}��ЕD$�w��/�w:�*,���7�J�/�F�B\�wPJ�F�j���ר2��u򆙟-�O�{m�)U�8QL�~�?sD|^]�Q�z��T�#�ƂL8� c�D�Q�K��;����?�����g����M*�H�kŐ��6�*]�TƱB�	���#Re��+�����S
�~ϟSΐB(�p�pږ�ފ�F�h@�i�E}��������9B��ԹR ��H��&�8�[	q���r��㚤��t~�S���q7^�L���@�̄��*\�:�ul�=ꖶ�6��b3��zŰ9���hT��7��K�矾+������]����6��
��Vv�{!�'��D�#�&�]��5����T"���w����g#�PJG��
�O��L�r"�)W�:�JO��L������[^\6b�hL�ճZ�~��~��۟�����}�CV�Ԭ�w�E�Vn6��P��w��P$�,�9�	ӻ�ᰛ])~p�0A�-r�w�ɟst ��~����� E�ݫ�7�܌$�s��5�H�H��y�;��N������"w��N�:��ݯ�o�n�������UǺ�b*1��訌��\ܠ���x���6���n[Cq�&-.���J|��*��Fd��Z��f5қ�q�g��@����#}=�1
-�K+�YꢂG����Ukz�pD�(v�k�8� �`�a�J��kw���s��3���q�|���}�h����]�תղ���%�,�	���e2)��G?j��~�>��`��G�P�X,�t�KyG��B���)��>��K���\)X�P�y���"'�E�����q�gY��3��UF���O��o��s�m��"��_]G��H��"X�V ;�q�8~��b�u��\�j7��V���h��U�E]�(�F8j�������՟�Ǉ��|�9�n�PX:�J~<
_�غU`z|պdZ�\����/��NǷ�:iե#�^���~vj���)����	�|��� .�L��į�n��l*m����m���?g)�������[]q#.쐄��;����������X���p6r���J�t8�E{�gϕ���{�sL�������$����zf�"���,!��(W�N�E��k���Zxg�\����?v��G:g�}{l������K�j)�O��޵�M�� I��,�Gm�./r�����bb�ө�H!Ij��m�j	L��x>x�� �EucH�i_�gC��W1)!����~����1')ɘ��E�]���������������w��&��Y�vy�*M�$��y-�4�K��N�{��,��0��w�I��w�8r�%/���Iu�L( /��C�n�2�)1ڈ�	��=�ܘgPγ����iՉ+��Ⱦ3��{}��ʁ_����Ƣ�]E�cA9�E���iX���	k6�b�DD��e�6���F�+�r�S��3�+�{r��`���B�:�r���?�Ϥ�IK�`��G����ԋ{-��XU�.��֬\2��9�+  �z��<�ɸ��40Cw����8���1,3���7�b.R�T�;D#��s)LE��V�:ߠ.s7��[*��}�>����a��_���&�.B�%�^n��< L=�p2I��|��!���z�t�I�5�S���3�0������y�n�J���t=?D:����:�����v��=��'8]�|�J�x�| �*-U�\��?��������h3*�[A�yV�����ˉ�,m���jV�[�d?r߻ݖoye5n�I
���<�����&J�����O��#��Zڦ�u���?��G��_���96���r٤�ҚUKe	��4�J/T�5w�IZ��m<���'�Tu8�A%C��ql�RM<`<w�g���V-�.
%�q���Ժ�0��˜U+����$!��2/s�f�I��#��g�l�_4ϔ��0�L�SV-H:��H�&D�#}�S�NY�¯͒�O�����I<�@��������SP_�+y��\J�Ft:%7��z����^J�!w[T���^�)1����ڿ������Ὲ�zR1���\OJ��k��Ty����6<1��4mr䄍9`|�[����{�RlXYi�2���|�_��f?�2=OtN�)�Ƣ��4��W�h����O��g��ǟ�k��O��>[0�#��[,q�',f�7�'���V����M��W4��E��tr%�x���zU�C��W�i�,�ՔV]�$�K$��1*�8";y�M�kV�R}���'pT*2;k�h�Պy�gR�V��ʉJ�$!%�S612��p2b���IJ�ftS/���q�T�JC%�)æE�`�d�|C%D'5�za��ݹ�F� ��3���DN͉��9��6�΅���Djg%�/���x�ѩ��'sm�ݐ�@Y�,K�Yh�t��Y��:��C9��╈�'�a��j',�#�N:@`55�$	w�@D�S��5��3�Ϗ��K�X�T� �����/S{��4e�F,k���G���?хI{��o����[���8�
���x��K�dS<}~��m�To4c�f8EE�x�����i*Mv(�Ҋ2�*��K�kR��IKj��OZJ!*-c7������D�h������P�S��qI�D�˦J�ty�(���@wz�J�_S�4)�*��S�U�)kN[���TH��1�P�¸śzZ���\���t/�r7�N[�L��Ҫ�G��KJ�8� S�8b剓�;5�V�\���V�O��&$�,Z��X-�r(_���7�7
ċ�&] �X=o���@Y�\��Dx�o����ޭ=D��B�4na�C�lA���-����@Y��L8����\q�EcJu(�g�*OIp$�K1	߈j!>�,sQm�-�O
�l�&�ԦD�&��������� )��U��GY�&]#�a�ͨ�q�b%�*R�K"��@~�챂��w'�΁�	t2�"�HX�?*(�I*aD~S�n�-�뭒���#5��>JF�2爧gd���R�/%�%mV�����PR�J����S�,��wj|lؒ�ȖTGRzP%EI�).,-���J+ŔC��)�5�e����Qzԙ#싎�����Li���3)+݆%MK%I&,�J:?0����ʩdL!ji�i&d����lF�ҵ��S}��oگ�- �W���B2&_�U!��S=�^Hȼ�+���גQ����I�&$��Rzaz�_+�TI:|d�U?�j�H<.�Ht*#�h���)bG��Z�r��':l2�2>d3�)	QAT�]��V�H���K�4���L�P���τ�z���P%�Ÿ����F��Wď�c�5��@��J��y�sy{"(�ԓ�I���\+�����z��$I�0iEi�* ���$}\"�� �0���k��{�Ӯڰ��r�5v�%�l��yv�u[lە���s�]u��qy����hl�Gh�IW �i�I�0���tJ�DBLDH�q�: (e�&�?�OS&lH�"ڔ���1�W�YY)(Oi�J^ޝ<��a�s�(M)@�%��5eǄ%���&;����:��x��׿�H\�N?��i���%T� ��W)��y�pSR^�R���BX�����Ǧ���e���<DWm�w��^D�1!�I�	d��l���4:A���i��+eWn\c~����ۯ�ڶ�����d�����7�{�u�]�n�g^i�,��%��%�#��B�����d2�d��z�[���;����8�؝���n�珂\ހT'8$΋N[�����צ��|S��Ę��V�4j`Z�bH$"I�K�ljR*_�����v��6#.- �^�q�sjW/�e[7���ׯ�4��]m���Q�bNi��L���C˨e�H0UJJ_���N��\�J��k�v\����E$/�M/������eB6�?n3���X�$gX�G*���4+ͽ�ޥA�L%BX�`�LR�Gz"E����Q�\�� x�c���$W{8uϟ�qL��I����[�:ƣ��Q	��3�
�<8�5�~���H�5enG�`(6ޭV�Y��h�V��Ρ����W8��ύ�����\�՘�?bw�t�}��{�ի�Λo�����f��m�l�֮v�|���Y:�C@��עL���M����&��,~���\�����]D���p~��@�"��La)J�	#�O�J����x�Mi"�QI��� @Òx��B~���z\w��+������mݒy6vx���޺�e-N���I���FX���E�(�ƌ��*�R�8���S�;�F�����j��xCLs��YP6������~��~���~�_صWo�	xkVG*+my.ݔ8�'��9�IJ/[S-�l4����1�&^���+�tZ����XS]T��hՊ�xM>'�9�s]w���qD�7��uLw�U�Y���K/�]W����GO����g
�����UQ�mI��{��I�sL�@�ƒ�vS�U��k��.Y4�^������%�ڑ�{�!�eɼyV�����7){ܖ.Y� UR9≄�ȋ��d�*_x��*Ւ���}]��s3S02E!��A�?'�|7tN��G�'VWr��
�e�t]�nW�����O��G��kV��~�[>�Ǭ8�*p�ȸ�T}���>��Z%���x���������,����Q�����ewӱq��l���646n��x��?2dC�����h�J{�'�_r/t�`��I��}�-��J�ē�T�'�|�5�v�ʕ�l�*+�����/�@ �֗�Ə+L��w��v�r�;n��>{��s_x�2�5��i������l��۷�v��c˖�$^�ֺ��;iz���f���N���UG��D����$^�Tz-�������KKq�ĕ��=�I������$��#b�3��Yh����J����]v��a1�D���tkV��|����u��Pi,�u��694i�#���ރ'lRu�c�>��`�=�̷푧�����he�~�g~�.[<`�8(���	WF�1OXNm�HtY=�k���n��?���w��o�_���A�*ߩX"?2U��5���<OtΠ+gs�����UU	�ݓ�y�Qۼv�݊�N�_���-�ɴk��x�-�LY!�Ћ��_~�A���}���ׁ2������[�W&��{�|�;js,���%�$���:q¾����P�[Q� �DjՆ3)������c��/�^��$�J2U��O?j�O�6(�W\a�.��}Rf����H��T�hHZ��?��z�&9l3�ۗ�����_~F�y��kb*�S�E	i�b�hW_}�۔���|�����x��� A;�YϞQ_���<s�1�W�'A�l}B�d�;�!��V�'*Y!����I�#���A�:c������я��Ƞ�#a�]u�����TIN���H)d<���<t�2]3�v1����3*R���~�&���C����/�b�n�IWBO�|w�L{q�>{��mJ<�U1#\�����._*�ы*7����.[�RQYS]�ͨՒ}��w:������M��âJ�x�����T�߯ɥ߽�y��/��/�N_�����x���Ph�L~7�8!���c���Çm��L�j�:���-�R��	�����G����%=X�����l��c�q�I��yv��c���c����_�e#�E�u��=��Nۮ{Ͽ��ܵ[�_u�*�Y\���ߢ'2%	�)�70+�r,J2s��yi����n.�ԛ�'eF�*ʹ��tY�p��Z����u�,��Y�	�I�*�B]L������e˝O�b�J�1�Ͼ���şe�lŖ,Yl��]��������>ui>~sN�<\{� aU�(�G�Jj3�����J���:G�OťK��"��|ȿ*_����ϛnPP	4��=x�=nM�M^���>m��g
�k����2%�fϞo���I�ڱ��m?|����"V��I��]:�訪LM�޽�Wv��CGmϞ�&�c���n���]{�۷_~YǃVR]7�t����-�^a�sI��E1kՙ���'�v�*SE�PՁ�C��3���ɝY`7\�ڢ2�QT��*�j������A����F�q�Fp.�H�� ��xJ����WTa�֠'J���܈��NwY4����+I;M	h8��D�j��ቼ��۔�8Z	�|�n�z(_��43�Y�� �ʘMY�vbt�^޵��9�LO;?%�K������������i��_�����K���W���?ٯ���m�nu�Zw&ee�,ۮ��~�~���o�g��������C�{�n��g~�.\��ܵw�Ť�)ݼ�x�Tp>�=r��Ю%�#���*�oAG��ڈ�d�����[��:r϶���IH����*�L �K|���9��:���C{:.-iޤ�B%mia��:�؋;w�˻w�Z���L������Ҕ-�X�4m�ذ�|�F�U�AS���Q�(7*6:�W*��C����&[m(O����	�B)���j����z�(�R���9��%z���o��C�;&:�t�	2Y&���|3�enU��Ì�HkE3V��X1�����J��
�n�h$mR^�d=._OO���@��e�*J�-�+�^S%V܊*��1wҽ(�, �3�1���Nq��M�J��~`�gT�jt|�A��GOwLcL.RS�K��ފU�-?0,�O�<���e�0t�Έ�E����V��*�S��9<2�~;���*`q��![��~�@}�����9�S�~sd�)��-W�Yh������ރ��L �ڬajU$ԊS��������,�Q���8�m¢X.�f��5�N�����c�C��T�*Z�Xpu�@�y�E�8!�* �e
V��D�'P	����3�bɬL��ԍ�����!���+�+ź-�3[V��Q<�t[8�tJ@
��i���nD��9�t����T��GV�$q�jĝy�_�ÿ���|�f��^3o�e�51}�RUq\~OS&��LJ)���K�t��81ne�8��H�A4��O�t�u�+=z��5�#,$��ňL�t�hi��s�l��EV�����_؉����|�$S�Jv��ٟ|�lfo�T�69r�FO�jq�r��L����SS
ќ-X���ݳ����{^���>�;t��"b2��ۮ��~�}�ZY@��Ƥ�~Bw �����u������59�c���N�i'TR�T  �#>]�R�i [(�.������CG����`9W��D�h.�gP��\��)�B��	�����66%��Jؖ˯�o}�M6����w���	+�e��ϯK{�Ծ����5�*-�=�0�����2���]V��|A�)j��`�U�mZ��r)�kA���,ALz�h/5I-��#e�-{܀�}w\k����X&T�UU�B<[<1U�O�s��p�':7��Th&��v��GUغ^����=��)Wn����a���=v��L؋���#��Q�udX�ö�А����҈9S��	UA5�/�|��� fP<����R�)��q_Gf�D�E�;3g[֮��{l@���'�z���F��0s�V�O��E�얛�Y�b����iSLߪ���j���_ҫ�-�X�,g<�L&'�G>���S��O:!à���sl���b:�i�V#�s�@K������G�y;F����H���ǂ[�SZ_o�͞5�B��j|Ѻ���1�x4!�&��XW.�x]�'�X@���u�c�w5�V>Wٴ�i�s�ʥ�=���! ��}�
�Ӻ�p�B[�|��Qںfαf"#@��u�\��*��Am�Ŋ@+2P*Vy t�A�:a\�I�n差��g+S�684b;���ö���96j����7Gm��۫p`p¶�_��<B��o���l��J+"�OW�Wj�J�q/}���b�5�U0���2��1p6*�����[33������֔
��W�k�=�,�o�PJ�hN�
���LF:]��V%6eJ6d�0+ Ǘ�^�D�:A5��S��O����Ii՞l�f�g-��;�S�rK�h�t:����1jON�g��Ǝ���ÁY)���F��|��ik�9����s�S���qiHf��Z�Y��C꣹Un]�^XA\赎:���L�&	:5x~���`�[�h����:k���ö}�K��s��K/����/�d����u��A;v������L��TJ���T̊��:uBu�CPn`�����$P��&�C*`fә�����ݗ���E��ņ4�_�H���e��I����@�A`F�\���<?([�W�#Ċ��%d^Fs=��[(7�"ݳ]uϕI9Ǣ�s-*^�v͔궺LV&�d3�".D����en�G:'�AQ$�$���!�kY@I ��˟���Y���m\�ք*$/疀3[X*�K�Ukug��%�0qp���I�9ۚ�]�:5�`ƹ�\���a緱,�̀liҎ�i|����/|�>�g_���mhh�u�d����`2Me^���69dC�XMK'�&I-���?c�� �q9���b~����������r�i4GZ҈����g/w�{��	9��w)}|�jW.#�6�rٴ�q1x�9|Іeu�.x�$sD[�Y���	<91f�#C�g�N��f�KͳY3\\&赂>���m!(���������"y*b��=�W��%���>k���?�_��?!��N�?��{jy���L��S�7兯^�p�U侦$�	s�����:%�>V�e"~�,ʜ-��s�s=�%�VQi0��C "�خ[�)�F����7��@��&:�
R����TDU�*�*�\(�YR6��b�����"р�D���l�H���j~]�w+�_	�t��������'�t��T���?j�~�~{���3O?a�}����l�k4�~@FLb�2�#��D�5� �_���qS���)�a�XGS#��RA��@��'�Nk%�2{���0C5��+?�����:�
;~��'�_�n�gPw��ȟ��������c�\~h<�NHsCߙFP���p�w�W��TY��N��{؞x�{���m��OK�M8�Z(y?����߽?�J~��u�0����X:`7�j�]Y5����;pUX���:0q�E�n���A��U�s�C�5��i>q&��t���-�D�tj��������(z����-���۷^b��]��O���/��6{�[m��ٖ�2�=*I�������e����w'-U�a:^*̳L����q1ƫ` :_0Y�bz&1�%��UaY�m�����܊v������dF	m+Q�e�IM��E�&s�Bj\y�҂1gV3-��I��cJ[��NJD�;C��&�����\��_/��e%[�(�32�s2�zz�e���K�1./�%�i�% .�chK�w&��aY�����Jz���2�K2�zgX�L/��z uD�p�3�H��%�`p�A��DC�%,˥^V�T�ݹ��.��Y�g �Ӛ��SU�ū=ɒJ�j�ť͑�RCUH␏4\I��͢ c\��bͲL�H��n�����G޼�~�޷�Ͻ��޷�dkV�S�I��>Ȓ4��ΐ�����T�r^��?'r��p��_�D�C�V�5���ݷ]o?r�����W�[�^go�~�}��[�G��n�z��#,,d����`q
����Ǩ«�Rd�o����1��[��S�P4ϡi��,ʦ%��!H�d
�1�@�5@T�_I� �,��i+AGCBf{^�N�ƀ4��I�0�gZ ����9�zx�^�oH��@4�����1c�Ӫ�d�ˮ�W�g��5B��F�X<s��5�cV�9�8s�̙�4e ��N��-R��H�Y�pAL� �|>�s�]q����}�F\�}SA�j��&�$��nIQ��ͪL���]&�x��mó�����R홬�ۮ��z���]m�n���ڵ��k7�O}����`�Y�	�@)�y=�V�(�3\���ΉKȴ)1�`I�~�k�g\�7)-�����>{�;�[��dss1��Q��Yhr�z#y�b�L���l�ҹV;)����G(��G�J�buU4���L���V�#L�X%?nS��:N"����A^&`B&{WZi2_�Fl�ɡ�*d~4�1�@�vL0 Q"1�1��c��+�z��$���ԙ�8O��=������^b���K0$i{f���q���Ԕ�����\΁�ŝ~� T �|�����L9�&�� ��W05�A珯GN5(��σ��%i�0�O�e���<i�LΥ����,�ٟ��
h��Q��'�Q���ذ�gXVU�J���Bd'*a^�_�˪��1�����[W�%����[�0d�f��"U[ї����a�j뉳~��ڟzq�ɐ����eu"F��w���ݍ۸$�Y9_�V�[�̿KW.��XL��K���>5(�3e����g�����ތL��e�H�����]�V����Ǯ��R۸|��]>���貫6����|��y�Ͷn�
�J�*CRғ����UL��̜g�3f����m�ܹp�|Nz�-��pL��=%�-	s�lܸ��*�w^K`���	Kf�T�N�ə]���6�AQ���n����q�2�͛7�i&�����@H�GZ �w M��>X�FzÅ��=��v&и�F��T3�� ���fϱLW�%�z->c�	*��.�r�(OC�n���%6�+c��Y-�]s�����gK�ϲ93��[n����6��2_ezv��61>h�֭���~��O�x�Q��@S�?�5���Y��m����g�=V���@gQ|%�E�	#��S��R�$�dd�R;I��wR�e���.�o=f�2!�"gUR�81f͒�v�(&m51i+ϱ�3{��F�)Mr��u҂7Z]0Y����&��m������m[���6��s�Mۮ��3��$d�0 =NT���k�z����w�{��~���-۝Q�A4�3̈́�d"��]U�
S��a��;!�a�:uRɌa\G`oIC��Yj��'~�co��O�t��\���ɥ��r�v}��8�l=��t  s 9�#��\�䜜�t�q������n�<d�^���~��v�{�g��'����wXO�)<���#֚FG[��,����6�r�%�e�*7!���x��8��⡪�v�6[�j�����n�I�\>�fkV,�.Y1��Q�W�Vӗ�5GF�įUK�\����^��x�Y�2�]����7IR���;��.�':��tBW ި�����k2Rb�Esf	|!��eYF/���a�&�+s�{%��{�ݯ�gC_�r��x�y;�o�-�v?��f�w��K��W�؄*닟�G��0g��$������R9��T�,Yfk7^f+W]��`ry��6K
!?����؜͘9�Ғ��i+�VCa��1��X���X^�ͺ�fY�Y��$��\��k�	M��B&Ǆ0��Ô���	G\���#, ��1G�1=4?�МԋkK>@B�Z�4��������1�ee�ۂE�m�����֧z���4=�>e��w$�CwMW*a�7�w���\"j�/��5i��͛3Ӻ��v��aw?؆"b3�;)e�:G|�IYS�g�S>I��%.�;G>]0S�N7�W�pi�yh�WSP��B*Rۜ
�LAWkغ�9�����w��e6��&��P� 2�W�3�Z3�b �"��W]~�4h�v����X�TdZ3A2�������c�0/���<`�|�[���=�hkl���qi��S�	�w��YK,�=�j��17�S�
���GFӖ�p�,�헖U�����DM}Dy�2 ��`M�7��D��#�xME�~��?��x�bw���8���i�� �/t�����4�pb���2Am Ht�}}�	7g�.�b)�pi��;^~ɍ����|��'��~�Wm�\����-�����}�S��[n��.߼�22��E7/�b/��x�ty���|:���0�+�:��rG���_[^��	����@�=�Yprh�>d��^��R~Rw���4@7wKZb&E%��&��'���G�|�6l��-R����+���*M�8������*�lǮ�*B�
j�	E�O)s��F%=f'�#�����5� UW�\$%ƪY��d�l���2���	]�(��z����x�͜��©.iְUF�vjQ^�ˋ�
D��O0~��'�	`qɍ�;|���߿�����|1LG�8p��Fٱc��޽����c�rϡ���� �{ b�:�r�Ŕ���PB�L:�yЉB�쮝{lT����`ZV�2��<�ˮ}�՞Gt�5�ۛ��v+�����v��^��N�XY�����$��Z���=)6Z���j%��D6�T6)�'�G�;zR��.Q�03�Ԋs^#�{^���~���V1 FH�2s�����}vT��XA�����f��ۜ�9���0���������L�J(n5��/�;b���?m_z�)��}�3��K��c��������ů|����g���g�m�m�G?jQ�'�H� K�+�`���$�%�Rb$f=���v��X<c�X֢�R}}��]`��o��W�h���6�x�e�ڲK���E�,�5�"�M��Y8�Ъ�T2!�" R��;yM�Z�s� x��9��&�����F���
��a2����>i����nE{L�r��gb����K�s=����'��9JΧ�7�&O��~=}ꐿ�s����$�(]�-���s��)��/�`Oo�n_��C�~��m�᣶c���?}�>�O_���m�����O���Ӗ�@8lR��'��=lW.i�fչ<g����v2�H�|e�AYGG�\c<T�[|U����3&b�dM����s��<Z(�%Swe��>� ��OJ�~����������r~�|9��LVŕ�M�x�h!1h�{�=����?�U�}|�*�4��QiƊ���62&I���.��'�̐��1+�J��"2�����⡊|�~[0[&�>�t�y�Y��/��2MVX_����/��8j��ja�>i��v`�Qۻ�[�����ؾ����[�a��C�����Wv�|P�>��̚)�ݖ-]b�_�A��J�'�v��N�b���a&�)`L�؀������0!	���` ��t��9�'�D�a���>o&�{��3��#�L���O���Z�Y�1���Ȩ=���7h�`�[.K�\Y-���2B�@��Y7�G��s�������xRmw��I�s`��!ök�i�Qe����v�M�f]�7{��ky��z�$�N�!���r}6.k��Д�ͧ�l/�=��U-NM������+WʄCۆ��6'��o�Jľ�:9o��
{�;4re���o���BV���~�>a�?��͜�g�����u[��U�6ڬޙ֛��u�_�s���������VK�Z1�6�}�Z%%hٕ��"�{$ƅ��;&�L�F�
j����L�떨L��)�~�2�WmV2f����箛=/��t�Mn�ࡇ����G:��C;P�q��b
�����B̣�s�N�v�5���e���?�[�|���޻���+Z#��@t���A�̜�@۵k��C4@�~���7!<x\����&!��������y)=�|�Ew�w�𮘴�4����>5�||��V��1��_e2߰믻�n{�;,�P�D�m�x�ya��������t�Β��'�q�P(C�J��m���i�yu��2-�\�FѬp��qӕv���l�7g7d�Դ=���kO�`_�֋�����*������~�V�).��
������+�˲��<�9�.��#ЅЩb^7����c��s;�L��mc���KVڂ9��X��Ͽ�ӭ��e�$�T���&�1�8����OI�9 ]�2 ��L/c2��V�)�[�Y�e3�v��9�,�[TfQ~dȾ�8-J��UW]e��-us݌��1%� �6�����C ��Z
���3���!�y��1���_���t���=��A��z���kջ��O�FJ�sᓑ���Y��I�l:� \0���,������G�>_���n ��t��1�oH,"�q_tǤ� �T��|bv�eWؖ��q�uX�;8)_��v|� +'��E��@3�+�W�T�5�u�(��7jM��
���ss(i��H�ٙ�$��$���������,��wb�^�v;1��b]f
AE���#w�l��7Z."�Jm<J�OkC.yA@�U��_���Cb��n��?���˞x�%��V�z�M%�>��&3�Q��ujLR�l(�6�J�(=cL��i���k<�6�.Vcz�
�_4�SFҌ�<T1���B�Ue����1�4�&S��b���A7�f`��̙�NK�7��y����Ϫ��'O�Ƈ�Sy7F� ���9rȶm��>��(/1Zг��3�?B�U�>�[�j��
��ɻR^@�;��(3�
�f~F�7��3�_��9D|�����:t7 |:t��>^tlL�{��G2�K���[M�����ƛ�w/0�-'�[Tu-�B/�tj2����GWV�:`�c p��-
nV��������������Dʀ��u�+B���ѻ4�nk}��}���?��[�΄�>�-����]P��HT�[S'~�?�Iw2/f�˲��x�&u�e�h��W��g��DΚ�>�l���I)H:E����&n(A�Ѓ�H��P��b&e�I�:vDŻm	ؽYL�*Y� 6c�5���갤��CG��N�/&�$#�nҎ�8l�#����#��v`�^�v{t�o�ԵCv���(��ǎTz�g��<���0ß�3�� ���S�Й@���f  �t8R����y�'N�pG|4�2���>?����<���5�#u�8�~�s�G0��w ��A��2�U�#�[sU�� �8�� ��Ä�r5"*�e)���+��
�&6.��Y�P�{��uJϖQYe+K��������0ď��$��:N��1I��
�
���H���H�%��=3Y��]���l���a��9뚵�"Ո'�R逇�M�4��&��RY��*����vݹa�EO���D:X���(�I��L���A�P�l���j�rѺeJ�������}�BM��T��,�co~�֝��=:;`�}`�	��?л8����&��� .���Ԥ�X�d��$�$�]۝+�Ԭ�lɒ%�ɦm�����`�(�z�G]Ru�2I�{'=w&pO������j�˘Z�n� ���@ӝ�_��߲�� .��	�I�����r�q��}K�}�-�m�Y�Q���0��,|~���j����k��@�8��Ji&��=텥� �*�t*cY*iYc!�ר0h��&������)��T��~}}.��/��;EzqT�T�hٮ]��+���t*斿T�,��5*�8���`FEL�4�2abU�cl�/��CN
�*C�unꙊ�\�ȼL��t�je�2�v :Cd��> �5k�]q�[�j�]�a�mڸ�6o
�u�R��x�u����v�uv�lӥ�lӦ�v٥�2��6��K���͛o��[�֮�b��X��&&ƝY��L��z�,	=�LNs]i�,�YqLv�r��vaV!x���J�I�� �_&�����f��e8Qf��v����"�rts[�T��:�y��|HF�,Q|�b�[b-�1멡��,���g��~ P��I��f��&��S��79:T-X����S�ͤ���:��J�}KA�3�m���8OtΠc�5�vL�!T��|94��L�
cG��m�@�nݺ�n��R�����h��XA~J�����:\c:�Y�biHL"M��㒒HX@��V�QT)������3Ў�+�wRM]��}% tV���1�.��K�)5V�J�)�O�[A�P*KX�B���}&�m�8���6%���Z�rAڴh�¸c(�r\L��OO�q=�33�J"���vu�����b�����e;�� ꘉ�u5�US=�q=�J���`bV�#�\����{�.M�g���̀6���]��=0��:�h/��X����W9��KpF���	Y�8�|���bEY#h�dW��Q�������yS�!Z������-K'ҨC�u HWo�J��S�^����h����mW�ۯ�ܶ�_h�Ɇ@��x
W&�r�du�u����]��It���"��]7N�쏈�a�/=�:1b3�gZ�0a�H���F��-o�۶m������kV8�2o�,;~���8n�tJ�H� �BR���@��w��z�b�����I�r�ߢFpc:b������f�����N9M@wz>?��a��sl�e�O�V���{����}�R v_n�����_�
�G����w���[D�����r:�uL��{���b�ab�HiWf�c#�֓��r\&�j���qγI�i�V:��g*��Gڔ�_:Q�G��6������\zb{ڵ a��o=)�׍J�ӝ��˗Y�w�%�,�;�j�w��c2�F�F,'����l�KO.#5���bɸ�iKf���/WV����1�7��U	�X�h�n^o?����;n�Ү\�ʮ�|���d����6&�w��Ch��s=ok�϶m[V�d�+�ES��7��Ì)�':'Ѝ	t�6�a��~�E;|l���	�z�v���잌�e�'-ڬYO:n�̰�ء��$��:�?���Z2�SC20���`�%0��x~lLڎ���'�IH4-#)�z�t��Pٖ/�k���6����-�m����P�+n�f�ۖ�/�yI���8E0�LE���oU����\g`��o!�kK�;��FMڈ�k�8���� 1�9��@o#�f��mf�p�q$>����������%��^D ���OՉSzo����!{���T2su�����![��r���m���m�(ޚ/H��&���sg�n\�%�Ҫ��(�NX8��$���Lհ,���dݨYUAJ�jv��k��w�nKft[JB)��Ed������.\`���6>:�|�ƄmX���ۼZ��%&���+�������t����\f�A��dҊEs얫�XV/�N��LYO�`�°edO_�a�ݰ�J��>��HO�(��Mv��u��t"�̊F�b}ٜ�m�#���t��5>b��x�̔�4!��Y�t1�I0o;c8�9�|�7
���7Q�:�������s�䩽,\�y������4��4 #�	�$>����M럁��=Qi�uU�^Yh�p���X�(��}�������F�B�1�)&b������t����Vʏ�v�;��>X�G#�2IOV���21>�ɘ�@O�����m��^�U���23�Rڍq�I[=���e�e���cr���#��n��oX�9�����t5��=��9v�f����K�6z�}��l�����[��Zº�����l��a2d5����mW�u�\�c�JV�A�^I���ڮں��RئxH��˖٥�n�g���L)���#�v	�i�ؕ.���zR�2�|``�m�l��wQK괪Ur���ngnr�s�����S���Q�9u�i<wvv:���3ɧ��`(���4@0�|T@�p��JL���Aw�>C
@	� �*Y� ����-G�����o�t\Cc���#�<fe�����[�ؖ�\c㥆����=���4���DR�l�/���-�؊��lÚ�6cf��d�[o�Esg���c����uk���ظ�v���|�mذ��F����p�4��m�o�;��d��'ܜXVLJ���5�8��Ƚ�9g����N?�:\6�^a�]�J|$^�;�B�f˼|�|�����9���Y��>	��\o���&�ֺr�e�Yܞ���	�q듩���џ�Z_w�M��|����౽6�7)����%K��2���{vXNy�Rq�ͤl�҅v���j���.�$f�U i�C�v��I<,�D0-����L�N���$��1R��S���^/�F�
� x�E ���o��
ӛs�H�!�">檟SI}`�R'<q�[	�����'�A���!,K\:%<�!�R�i���W[1��Zd�(_vX(���w����t�V[:�=��6oF����
��^|���m�Υ�q;v���eMYNlV��Y�}�AX� �o�",Jc�Ѧ���zT)�o�ҥ2�뀒K��t#g=;c|�tΠs��!x^a�I����@1y���؝+�ƭɹeC���dF ����c����MY�]��M�sSv��I�3#%GxTi��Rc�������ӽ�w�F>�+����u3�iP:T*�^�穢eʈ�ĩ��`.v�bG1�!�1<g��)0H�s�q�ϕ��M������:=[`��BQ^0>�q ��
�)�ZF^h$��-ӓktJ���>h#��$���k�s+�ݸ%���J�
��с (�!x-�FDPV!���d`��M���*��ҤC��I	�����G����^xѾ��Oٶ�W	�����;p���;�&�ܧ�Y���M:�6������Y>ZL��QflF�UB���JL��
+�:��M{���U?���p�]���� 1�ҍ�U�$�F�bC"�"�t ɻ���y�%[8���YV�,-s�'�ew����붌̈d2�L%zw�خ��=�Fr�,W�1�G��	L���7- ȼ�����Y�=O�����������٘��Ü�� �8�I�Rϔ�g��;�����o�<�ѧ�
����H���T�}��q|g#���\��5T���֬Z���z��Go0�y��=3���?`�vﳉ����y�}���3��$i|�߭Z��V�ZeK/s�S�b��{�cc��zA�1�θ�t�u��%_C� s3����+������Q=������
������A'��ʬ+{>Ԁ��bPaUbUP���m<2&�AfE*k]rx����r��JH�I������q�|���޼0�}���/~����~���ɼˏ1���g��=�����~�x���!�GeRH���Μe[/���Ϛ�6Lu@�gB,C�0a
���U� ي��0+����O�1�Hӧ����>__�qq�u�K@�ی�e��z�%�`2�'�/�zb,�4)��{��=��#���pqζhR�N����a�H"_~���ig�A9'>����|j�m;0����+�[m<�طl��Q{A>�W��M��W�w+I>�����ڪ��l�޽��/|�u�Q9<b�tN<u�S�KM�>��������ؠ5+๽P%�ѣ��к�������AYL�(9?�b�f����z��
�s�H)4��wf¡>)���ן���I����-^0��/�+&)ۤ4X�l��TmZߜ�vl�d�~�{��W,.�ʠ(��d����:fS%Ij��~�%��YQ*L��}{m���np��������hK&N'd�VFm��a:.�{�v��)�*������vŖ-b
����H�a$U�x작 �0+cs\g/L~{&���1������@<����O:\#�35�!R�.}4��P 8N�Y�wߗ� ɗ@y0���6ħ���>OO>�O���z�� H>SJ���?.W�Z��VXgwB��c����I;&����>)��e&����j�CCj�}��.���w䨽�[���~rr�^ޱ�^ٳ�F�&�BY$N�ǎZ�@�z�2K�2n~p6+V��=�`��O}�a{��;uM�C��q�R�v�ji�^'��*��fţ�ӝ���'�3�T�R]XY�{��z�����cÖ�v����<�RKV��tW��(-�l�D�^�w��ꓟ��z����W�2��/���*31��)�~�<��-���T9�|�@^o��ʷ�6+v��n���ö�g���t���%�P�!��4\G��E�0	���xG �y��B|� �q��| LO�xHP���rHѭV��uN�;O=���P��`�v���i=S��\ �G��q�'��P���"�<fq� ��/JhP ��}u�����r�cq����T�a��'�ԓ�4z��ٳ۞�o���/�ޣ�VS['s=�m�X�8Yך�t�K�cvV�WXn�w�N�W�x+/-����V�nt�ibL�۷g�%3Y�̶��q�h�q�P̎O��3>m_z�Y.��şly��v��1Sf�]��pkp����Jޕ�"���*�ܓ/�{[8�t�C����ni��C�vD��w���ȷ�_���t��Ub�m�Z���2W�:�YGكR ���ي:�e�Ё�fO�:S�B1�*Z@eڑ��7T��İՆ�����<?O���$��!�+��¥h %�b*@#y�s�<�Z��̋V$@�:gH��U���u�?A;9fmi���z�?���k�S,�*i�B:Z(�(#q}�����{9�XE�I	!��-�p&���H׃����nL>��zRmP7>b����g+>��(m4㖜9GV��V���RmH˙��\b��Ln���{��,���t�y���	S�t�@�Vq�����m�^صώ�N��c'�����������=���v2/��P�NKSv��Uv��%�`���{�|���V�\�V��3��e11_��3�G!��}��g��o����%�b���#'m�$����!U| �(����:RK�#g�l$��a�� ƻGՈ�g�����ۭ`W@�K�^���HyD�᠕�b�Ҙ���e1 �5x�.�t�}�#Q�`��̐�b�&Ī�vfb�+�`?��5�F��- ���0=@sz&�@<_(��t�����ÁT�q@���ۆx�ۙ���d�ӁD����y+M�	�Ӓg��QV���29�v"�'�J,��"���S9���/���66<f��^�A���m���rn�喬�F�W�I��A�M�����ZAi˂��ɑ4���[��8+��pM\c[�D&!R�@z(+�	�}%Tel��^)�&Pn�xY�x�5�9�O���d��Ȼ�����-�Z0�j�&
��.����*�<���,��{�Ǣ�5n����6^Q�l�u�Yj����֓6f��䬘�j�E�q��*1��	���0�0E�ޮ`M���=��๊l̆�X3�1��>f6��DӖ�ܘ�:`� zN����!ۙ��!��
��a��pj(B̂�a��X�IX�b��G����0	�O�+���`d�v����isDC1ݍݾ����F�H���$0ٺ�����y;r�+�������Q{9^�������I����ɺ�����)��'����|>��Py!I\75�#�B7c*&|�}���b�(a%a$�Ԣb�T֭T/7Sn�g�r6V�[3;�j2)�������Q��T�S�|��K�:4����ܧk,vv*�+q�i��U�CLڏ���^|��I*�M`e'��*�Y�v���*2���l�BQ��Y��T�!WE�eʒ]?ƁP�%۟��:;7�T��z��B`а0L}&Ӹ{���3�g �fe���\�Q���'���}��� �ᙎg�G �9�p�	��k�3ɗ�����Plt� &������Ð/�����6}�2��.>�����'�I>�s%7A]ϐ�0`f����O 0��e_
��ᯤLz�A,.��k4��E���ʣ�		lw]`L��eu噜! �2�҂i���"O�"B����A����H8-�ʭ����[f����PX��^T�������&���	t#��Z���jw�����q�X����h"?)�_qˊӔ6k(K@�j�?��:�k�X*� L'��N�U$��f_B~c�x�]��,p�����Ys��57�`[�m�7�r�mڴ��Ȍ�����$�i�X.`,�y3�w, ��+�3%�
���}�s�k<K^���e<�2���	t�x킁<��o��s�C�I�D��`!�Q&���ƻ�V{��k�ӓ��FD52�άڋN�E���֫��k��Ѷ]�m�9��Rt����rT��Ħ���Bb�~��y��[Hq?X�	�Qw�F`r�TZm&�����傴��k�fd)T\*��ސL�pC�@L��s�]A��ߤs��7�+:��zݮ��@?��%5��	i)�Q�q�a���{\��ebz��$�0C��&��uI�&��j�O�֚z^\㪱��luiGէJ�
���9�/������*�|ޒUv���k���{�=�;�x���~I�J�'�4�����k �ip��"6L]�i(4@	L!ʁ��F��J��T&mݽ=N�3��7��ҳ`z zc�^�up��c+9f�SB�Hp�Z`���H���R�,��x�(�瞸�4�B�u��@��k'?�r|�:H~�ӂ�	Gi�&���xK�������v�]w���~�� �����veOaE�BT�sc���|ڸZ��9��*U���ã��ri�X9�
ME߀��eT7iH�jՂ��p]�{����ټ�9˦��`M�P����g�J��NI�ё#Np�!r��:?/tn��j�;`	׀�W�H�倆lݲ��c��~������Ƚ�s?�^����n�j�-�W�N�9�"�Y�_�yt�ĭP�:�CZ3]��`S!V�5�h|M����
_z�=aϽ��F&K69�v8���$=϶�r������	��+��Ʊ�g�g\�Tv�:0�F� ��`Bb6A>/������5�e39@����v@pε3�ךg�������<G��_�� �ǖ��\�5���:t��ڽ_�5k��!V��-���+-'K�&��I��b�r��ښ�$���b2����)'x�#��0��L���^8��|�V��{�f?���ؿ���ٿ��{��H�̙eSr�-M	��/�JbN�9��<�9��Ό"S
ף�VHSQ��^Z������o�ۯ�`[�ۖ��m���._h������l�̬���dj���L���҅�،���Dq��<�ä�h:��(L��`����h��C.Fd�OL��؞��e��]x�a�p��<^�����y�iX0++���	�(=�0-�>�#e%�r���|!}|?Ҧ\��f陠���$�u��)3���������=�,��ξ4!YA􅨡�,$��|y�n۹w�� .�X����s]b���I�1��LB���/g"K-�fZ�a.%w��:�T��?�HW6#�U�y=i��-7����&�鲕�e�L[=#a[Vβ���
�M�h�l�6�s�����@��SX��ԏ�E���Y�r�s�Xu|�[פ�Λi��z�f�B��)M�-����Q˕�lYwܮݰ®�b���dvH����bɄH٬�����؄eU����;�_��4��$3`�v�B�y�b)V2�@������D� Acr#Ҡ��:���A�o���ɫ��Is����H)/�r����8� ���<�ځ���??�����!5�k_����o�o|��
j��C���n��{_�eJ{%�����N�I��(���;k�c��g1's�(M[T���s6�e��'�����q�R�	K����\�l}ºk���5����7ns{��F�1id)V%�����:7�5��HC�� ��RQ�{>˴,�U�^b��YT/��NY�V���[dj�ҕ���$�K7؀��ެH��v�%K�_����7o���2	��}w�Ůٲ�֬\do��F��?���+�P������ۇ�͚,�}�̀�afO0��ىz�	K��������Ѐ�y���A�Ą�K���3h@�{�@#@���k��4ȏ{>����H��9xޛb�|�������#n�lF�_K��۳��w���S�P����n��kl�%��֫/���,�{�q�}���ڼ�>�b�z��m��{�|�-��g�o��~�#���t���Q����m��_%���RrK��q�T�4x��ǭ/�k�Q���ٰ�V.Y�x���J����<]���]���(@��}�Y[�`�[��J4e���6gمL�¸%e�g���9�6#����[q��6�������W�K�5K�:Uh.�#�ڡ}��f@������X �N\/��Ǒ������.�իV:3&r�9hIu4L ���:�3*��0�]��5gh&��BڤA�0l �<��x�	�'ڐt��yI7?�#,��K���y�8<�ɗ"�/�&.む�@�0&��_#�n>����~���b��Q	M��_s�%A{`��}���t�V{����MR<���lV_�F��7�`�W/���ߺM�v�F>��V/[l�Xqr�܇z�y[�p@�R��Q+���l	Ͳ,$i���������.��K繥d�F����(���q�';C�����^'�e/S ���,�sD=,b�V+I�W����W��
EK��9��֟�Y�Tt��ȏ�uWl���q{���G�ޮ�]&�Ȳ���Ygu��o�1ε���nȤ�c��۝Q̲�LZ�l'
J����ȧ�k�u�� . �<�W�I	0'�"=�����z�s� ���ci��@��z���
��4#�� | ˽�����f���g��1`?߅ŋ��h���8�<��嫭��{=K�܈�{ޕ�p���8���,͚O^9	7�Zsk����/_��9z��y�9ۿ�e:z�>��O8��~�f�|�
�Δ}�o���ؾl�\���C�	��])KK��7OL�����ߢ�g-�*�eţ=QY)g2$����@>�"�<�|_tN�k�:��F���c�ˈ� �����f��@�9�H_f�'�K>Y~��^�,�*�ܹ���t�����#��3���k�v�`F�s����hH��ah>>���i|�K�w�7�������o|�{��9�0�?�䙛����0�ͻ��Hg� h��D �x= �h9�������kM_._~�,���ҥK��`���k�G^S��/�&�^�����G>���&��9cV)V��m_�̧������'>�W���l'��L�;d]��2�?��ϸ��sl��e6C��o�����q�Z�3{@nF���V	�>g���L%�66:h���y�s�K{�e!d��n-]S|@��1�V�����6r�Z���M�)W��8UI"xB~0n�$k��<���;e�h�\Jx�[W6i�]�,LYUwb��)`l$Tj����a���3;���ҕ���mӕW�C�|Ԏ�T��}��������Ba�b��IB�w)�9|�=�����x��Q{�'Ni8���q�����C����73���5��$�@��`T� ip�3��L�9�c�Af��s��mJz�|�\���v�E萁  D@�2r�EK��ɬ?��L�:�y�v"�s	��o4K���%�%�8x�=��#�췾i�<��~�	�?i�Rp�'�>�s���k���{�u�����w�,[�r���t��y��m����/}�v��o[���v�?�zBٮ�=Yῗv춊�d~oU�V<�c�xF���lO����e�ltl�:�\�Q ��Ўg�:�U�&'W�3�{s�@Q�u,��⃏�����!�����Y3m���nJ����D�LɬLf{l�qK{��7�y�T�K6�aH��ʮ���c��]�̳O�����И����а�� ���]LBh�%�6V/��&d*4�\�1����"���\��-��'1`�@E��0��=�8�E�L01�5�����F�y�]Ϲ[A�ʄ<�516��
���L��V�\�ܗ�]W�� <�l���"\�z`RV@X
\��#����9���<C<���ܧl��j�S�=��G{ʭa�9.���M}�u�o[�z�,�b���|���q;)�O*�o�~{���o?o/��c{��G}ܾ�kãc��+;��^���	�(�x����Ɔl��[�p�%d�N�r�.7��R����5�u���}]�Xb������D�W����-�"͉R��x�HX�<ѹk:12��J�x�M�ʫ��V{�����{a�1�fB�NVrL���|��}��G�K�<,[3m5i�Xw�5��a�p<�gbV��a"��Ĕ��+���8M�P f�$���������;s����Ǉ)y�A`^���YZ㨉�LBo��� ��ܧǑ@0���J�8�7C9��|��0j� b�3��w.�����g�fȼ�W|��8,`��ƺ�LM��6��y��Q�ԗ��nNՑ�����~�{6Z�iW�nn2��k	i���dv�č��>^��f؈�1Q���BC&�4�T=lE6|LvY�k�%��o����@T'-ߐU!>�l���j���'�.�Q;
|��7�Ż_y�E������	���.+ԙ�U9P�-�b*�1���s��Fe8]�����99��$a�H�z�e��O~ξ���vx�l��vF+�����>�O����n�$]+Ҙ���|��[��g�(�G1m�&�]2'e~2)Zf
ӥ�N�`�� &(L��0��&|G�8�����B�9"�!��<� �O�{��7����	X�����ǃ�=0}>�O\甇t��bb��a>���Cc�����ג�y�D9��o�g ����}y��I����i��O�I�HV����_��W0��� &�a	id�fjWT!��\�K3�
p�dN���P����8/�����Zn�7����?&ki�d�e�}��oڟ⋶�ؘ��<���-�9;�eJ����_�{�sZO���oOϘ��\^�i�����a_�e��%	6�kC���d�6�;SNmR.3fdȆ��U0+��JȺhʩt|�j���$�*&`F:����L/�Y��.���}�O���y��-4q�ҡ���N��޽�U�������؏��Gd��NhI��i��c|���q�9��| �Ã���4za���g����}�/�F$�z��9B���r*7ѵ�@! DwOZ��s�s�S� �r�K
`!�N�9�Hޑ���mDuV���N����U�������M�Θ+�ד�^�S�f�&Ci��t��H�e<񥧒��+�t~���W*E'�Gc�K�ܖ���qUY}�OJ���Z��ŞY��w�Fw"j�g��Q�bц�5�fm�rV5�	�銣���b?��[,*W�:����Gǧ~}C.���H$����ɧ;>>�*�IߗU�Gh`1�I����xҎ	l��*B�^��$��^n���+d"ԥދb��*+�!��Y�ߧ&t� �xT��ŧ�(���<H<>LO�%��a���c��27�Ya����|��d�*�=0�cɟc|V�o�|�����ivo�)�7�`Z4�q�p��Ayp�����	
3PҨ�@h=��4���|�AE뢵�(���"�%.qо��+���9�`t��N@>^@�R8]c.���j�o�톥����N�����M��n�����l����d�	���G�!C��}�G)��:=�~:z"��[ڨP���3����z����{`A��
�jJ��Ф��)Ygl��YR��.��,�ʔm\6Ƕm^m��W#�F�,�.�O��tN���诤sB��
|�d�z�ш��6U�z����e�\��3-,�V��]���У��8�)IƜL
���u��a�8EzG廸��b�L���Hu�
��D*��k!7�G!&�t�D��G"�<�I��ژ����
�(Z�����e�>�J����,z��ϛ{>�����)�|zޔ�7����u~sD�2懩Iy�=�&M�I����g�K?A�@9�;�������ٮ��$ ٢����+�C���w�۪�);D�T(��ym�]`�
G�bqj���(�v�@|��Ϭ�U�S���f㖌�,�PZ�h�`��A�.�t �X)=`������붢��/%�)��;�̠jV�nj�[7*N׻���~�tN�k)�6уG2૗t��E��P���X!���um�KN���䬆<�����6푤g�OY�sS�H�*�a�ߠ+�df�^S���E��ʪ$����G�����y�9���T`�p��P�9�Y��7L聅V���JZ���_��	�w ˃�32���. ��U>�x���i j��"��}$ t�����M <`��t$.��(+�I��>�ף�՝'V}����Eqk�$d�����m߽�|�q���L��p�|�!�a;�d"�V��z��d6���W�$`���+�J4Yo'W�%_J�]�c�\�%���rI�{LZ�8& ������\'!Ew��it��@��W�Q)B={ N����t��Q-Z\�+KRHb��y�OH
�#��Ś��l��#� Ve�`|O��(�>]Ur��t�/��A�E��8>�*+�E`5>�ES�+��n�6C�>2h����cL.4"�#�(ظ�l�.�=a^�c�A�9�����S��0����dmΜ��*��.sl��9���V�`��Y΄Fh$@F��+�&��VA��i�q�ԙ[=�Q�@�B�)�H��XE���?qԎ;l�cç ���L�����:ϭ�k��"�yA��s'(T�X�5Uf�-�h�C���'F�njjq�7��;,���2��䥵�o�sN+҂��C ~:�q�OS���l�X����|?�l=iř�X�l�i=��}6�eI����2�yR�.����]�[�=���j�+�{�s��XQ8$ ����O����f��fq�r��[6�O��^��x���wٻn���/]`U5*����Uբ����3�0�`���#��(�iL��mq�(I�p��l��&8�މbJI£�OZ���`
�@nB���G����9� `@�A�PN�$A�UbL<�c�1�&�7q}���>��<��" ��_V���g���ƻq��s�r�6�9���,�C�4(��'��s�&׈ �4� �g&l�aX��?Ơ5z�o"��\I����)�;��O:�U�������=��,�DXn��e_�ڕ]q�25K�'l˚���w�a~�[���C��w�bVε�Ԩ��u�Q�JGW2��C�`���y�s��G��E5U&k�p\�zɉ�c�|�l����f?��w��Wo���X��2}�m7�w��[�X2�g$��ٌ^TI���D�������J3>�w�I��A��3]YN��?+3&j�cEI%��)�ʦl��%6o�l�0��iH�K�y�jP�� �jR=ó��	C����g<��`��s�C���s>Ήϳ�M�L��iS&�� ��Ep�U6�&`b�סQI��0)ɛx�����!ι����/�.+�/+�n�2����>e�����6F:�<5��;%��`	����!\ �����7��؎�q8�gK'R�% }��wؿ�~���Z�~�r�v�"{��[��}����[n�\&my�Ied�pWTv���A�^�5�9�i�Os{J�l�$N6i�����5���09h���K��(�ڲ��}�]w���K��[�K��q����`Q��c�l��Q���2Odf��N������u����+J/��z]9�4��7޴������gJ��07yyF�q߈<�?���8�L0�7�(?��k~%�an��x��M$�M����Ngr*䙘g|y�P�0/��?C�<�4!_���σ{��.��Jx:P "e"m��	8o��c{p�D��S�������x��z٥6o�ť�%�$$�e�%s1����ЈM��-�=a���Ĥk{&@(�s�L����܌t�뮶�o�������e��(Yw�`{����n�+6�qf�sSd�5����S�a���#�#�(
� �ax,X%ͥk�]��6�Xh���6#-Q���EO��%�rv���� ��|��|i���g��K�ۚ���'�eK�j������L��E�����=+N�؆�+m�UJBP��x�!`V��g�?��������o}��E��g�����3x" `�yp�����}��
`E���0I131Cy���{r��ty�k$��u4�x�r�A��C��q�g)7qHa ����O��wz�@�g�.??��T�NѸ��I۵c��������;����I��z�u�	��C?"Ss��Ev�6of��&�l�o��zsi�U�U{�Z�̙�h�L"�:V�,_b��F�2��'�Z�:n�F���)K�Ƭ>|�z��۶ڲ��ܷ��Ŭ�<�`����m����p2q_
Nҫ!'��T���sr҇�e�^�Ŗ��Py�z!;y�F��1�q����)�7`;�C'�\�'�����[�+.�-�mp�4��E�C�u�1�M۶	d���9�l�@��_�ʮ��*7>��g�����%e;�{�=���g��W������Yɀc��7]z)m눺�|�ZR\��9	�`h��{4��B�
��`qߛ�4�
�s�̉�s��K�����o@��de�a:���{%phD�M6=✹���/#y�S3@���/�;���u&�F��<����3n߱ݞ|�){Z�w�>hE����e�����X5&+�+.�w��-ⷚ�8rخ��
���w��ҡ�횫m��Ŋ�~UU�����7�t�m^6�j�Ǭ/'��<ac�G�^����,æFY]���Q;r䀅+[�|�]{�Z�K�|*QE�M�\}pV2���y41�IӉ�#ҳ�)d����&;�J�$�r2����M�u	c� �Fej�zIvtR~ ]����v_r�%���O~�����7�s�|�l�aO<�u�D%u%���cb���t�F�:`#�wە������Gf,+��2}��0��f���0x�6���)`��D> ��I�8@��ɂg}|�@���=4����Y�I��ϛ���<D|��׶�� `�d;���rȼs0�fۛ� �w���/��{��z��C�oL4zO٫�<�	+.JŢ��_�t��ˣ�L�t�3�(ȵb�f���M���|�����/����w�׮Xb��1?q���V���}�_Sa˄�����jy�����2�,̘a�h�q�L�i3�ˆXq^�u����UzgY:�w��@�&	��{<0]Ԗ��0!��GI������4�78�����;G��^��� �4<7�@����|�/�%�M�8t��c��T���A�͊�X2צ�OZEדQ���$��<�Ѻ$�z��O1"LJ�S&Q���{��&.G@�r��!��0�O�"o��N�H��\�� 5��3y{Y����I���, �ݜw���~�%�a\�'�#?� B��'_7>���|Y^+��p�u>�L�@2�U;��ۡ<�U@���0t�k������d�/�w�����xh֌Y@d��5��˶��J���u��agf�Y,\�baB�����_��	�~�rcAkU �s��Ô�A�]z#ؿy^�wN���Pf и���Ą���L`6	_��u�IO�]�>��'s 6��40�_q��q���W�j��^�_�n�3S��w�y�=~ܞ�yB8́��5�Q.7�.&��8��ܧ�ܧ��n'�s�@y8�gyO���I��"�`�'mޏsW��~p����0�DZ�����gx�|:�e&�|H� a>s�@>�)����,�צ��9߸��?ȗ�gϬ��"��G���20	�4����tBT�sB��('q�� ϱ>M�u��s�=g�7o����-6o�<7��駟��.�̙۔��8$���R�|���z@Z�M|��~�>�/w��R��+�s��&VG�{��K��	�F�k?a'��%���V���ٌ����h�=N7w���#���O�O�d��+�]�wȾS��c��_zy�=6�v�ݽg��K{n߱����o���#��˯X�X�C����/Y�T��JJ:6lbd��q�հHQa�U ���rI��L۬F��3���sG����	���Ѹ��Z�Fp��t�`)���|�L����)'�8w���`L�r����ע0 L�E   �8r��!<a��� �C�S�D�LM����~��qxΝw�3�3>>!��3Ք��(pR�j�Pܪ��E��~����[YP�I�ґFC!�cq�\�'�������Ĥ�O���cv����q�w��i��*�M����}�9*>��>=}u�=&,��o��˾��S62�7�e�]�Ԯ�l��&i�,������J��ӽ[�'���	ב�X�j��@�/=����������a1@�z�p�%y�c�&�	&Ҷ��	�������ֈ�r�cpx|�`GOY^<�>�,fܹ�5�1��#�g�!�[<�e���ѩ���L�א̗����ꕋ��)�-]�&<��A��|�g��>�}:�c���U�HO@�o<04�������G�`@�D0�P�kć�y>*��׈��$�3u8��*G����к����MY���|� <K����E�����'����N�����{ �.1�[��O[����s�ںl���6w�*럿������j��`|��"���Ę9qR�:f�L��s+ď���)�����r��x�hB ��R��La;���ʕ���Ն���h��I�v=3l��)��7��g���OyJi,_hWnXi��2X�K4��óS����XeI$��(_V4����{ڎ�T�Ꞛwdg�d*gY�T���o>��>�ůً�OX3��c+&��N��j1b2c5&���*���J7�I*�u��t`ש��Y��D���2_ �q����+mْvɲe������YD�?
��Gÿ����Ń	�gЃ�<��@ �g�Bh9����&��+����7�<�'K[ �֨�'=�����]��= �Aa~�s�}����l��״�K|�=|_��M�<��H�՟4U(�cO<%�9��֬]m7�t�-^���Xc��vR @�b�a��\��T6��"[+�$�'��U���h:�WX@a�ʘx�R��E�,�A�F�;q��;�V����\�0��=����W�G_�i��Ҫ�mê�vͥ+,�VT��F�\}xv2���\epΠ���u�V.��bþ�싶���R�q)&�˒L'd
��_�m�w���z�%�}l�"�>YbJ����V�yӅ$!+�奛��zq
���^s�'���;�Jݙ��DT:c�z����Qv?�c`��=t^�8]�\���p��f��w���:S;x��|��gj�\P����V">��*F�y ��Z{9Iۃ5��K��"Ҡ��A9�G>�sp�����/�A�G��z#�e&]���?&!��S��0�}�%k��ڨ��]�G��Є�L�����a��׻OH��/OH�a�PY7��R �5�ߡ"Y������	`���?�����/mw�;<��v����W���HY~��ۈ~�4n[�.���9W��K֢� t���?��=�[
�q�SI�+b�z\v�@Q�fl��o�=n�|{�^�Q���W쩽'�d1f���L�?�,����eI)*��#o&VPe��o$�������.f>,1U�R����L|,_�'���{�}�a8�3����k�R��A�W�9�h���f5�6��o�$��$���B�� �O��4y�#���`J�]��˗��oZx�8�����U�	��q߿��/e�u�z�ә�ܹ�Pca+ʗ��B<�������
��qU��iM�˺�F�l��J� �'����ʹ�L+�c"^������0��qln��|dؾ��K��o>o�?��}��6R��궔ܠ0S�$����5I��ćB��=��+�?�VC��쩫*0��<U>e�s.M�m��L+�{-�3ߚ��l"�m#%�ԥ�l����!���Cg�SH|�13���l3�;.�2��W�Kl�RY�j-I�5,���/���,�!��V�|4�g$�3F;y��4 ��0"�P08��{�m�ɇDw>��~��c�V9H�<Hۃ���9'.y�<��,f. �F�L�Fˑq9R�E�Rv:����=�D��.� ��6�qm�w����&e.J�Fc�\Ԧ�)�qt~QNʞ/Hk���]7$�����&Sa��&=m/%P�sX�	���f͊��	�Y��3��T��ʙYf��lL�I��<_�w2o2�,��-����QJe�N��>�k��6lq�4.f��A���Q��b�<*K�v���^����HV�S��ǔ�rZ�4\>�0��5���@:�>��s����"F�DE#J�	��%-���a:_ �1a6�-���y`ޏ�u �B���Q7̌OG� ���CY`h�130N\?A����Eh[����26�������sy_���4I"nP'�A�9��=�`Z���Lӭ��UʖU]�dSjs�/*���.�N9��+�k8�e�O���nY��&]*�i>f�:`����4��:�`ߜd�&krOL�g,��{�17	ۭ.S���)i��
8�\k�u��e�5T�zU��&�n@:�
az�vT�,����n,��g(Hcxe�K��)=��V�Br��
��r�<�׈A�t[���iTV: .�ؑn�.۴��Β��� �j-׸G�f��-��ѹ��H¤��,*��}�/��k�Ɠ����,�'���������G��.� ����M��aJ��֝�����"L����R����?Z�~����%k�ْ�˭�o�͘9�z���T�������E�4�1�0�+������A��	���;��*�}��w
����l�c|�c
���Ղm��z�y)�����lJPG�	狕Tgpߌs���4A��N�b0	�:6�l����f'9�o�zO�Ҕ޷ac��T�	5Q�.��ׅ����H_��8Ƚ�{��H����\yU$E��H5����N%?&��l��n�f�z���+l�+���-�[uj��&`�gf��:@��9�`c�"�1�Ό@#&cB��2���.�arQ�i��=�ӛ��
Y�g# ��g���i���{�;G��eHX4
�h���h3�m�}:�m|�7e ]�C9H�߾N�Š8,�嚿N\G���^Y��q�9��I�.��Y��7��=�^�׍�/f�!m[R~W_�֝MXo&a�/]+^� �s7����`�$��xt�P>>�fDi,�6�f�\�!<���&��4T��ZT��-*٥���M[��-[7��V�����R�sS� ������6k�P7"�x^�w���B�ةq:��NLU푧���GN�ɺ,R��/�l��2�y���m�ۖ�+l݊���6��j��1�=�֗4boD&��!��b?Ƅ[J��Vޗ�|$�X��dLH:��!����	<���8�a�_U%;����~��}��^��뽼l�&:`l���g ��$���L<3|�`n���@��o�� ��Ѩ�I��R)���1!4N0�|����g��-I0�6e P �.zWF1��r�����Wi�׽+���]|��G$K>}N`F��T�Mnf�0�Ԩ�mxh��8d��?h/�;b�UՇ�h�I	۴4�<��v,*J�6)R�ʪ�[?�]X���abz��r+�"��b�	�q�Z��-���n�Ҷ]��6_���.gw��jC�e ȺP��q����U��
��k,Q+�kߘ�N2���+� ��	S�J�~�T,��$��5P\�ܕ�W�[��kZ6<i�ʰ�I�ly�n�r���M��1LB&D:��������儳�1�BJ�(�-;�2���c�ގFA"�����{`�=v�����|0.�4�!�o��3�3�?G{*���v��1�}'�a�@7�%>q ꊴ��;c��Y��ک=�����y��?�t����'>��!�� �H/&�%�B\ʀ&�t�rμ��"��cT D6��~�a�}���>��ƃ�w�� �M����
zi\\�ai`B��|'�e��C��+/����zYZm��}�q��jLX�:n]�	[&��Vۻn��6�^�/$����)`�Ƀw9՛r~��@'�4���x����0�̄5K��M֢^�G,gK7��1���F�6�Xl[7�S��a4%;��
;n}�[�j�-�;�����볅�l�$R���2?�\-�������@L��%љmB�vgs�&�f��1aR�wo{��F��i�V�K�eeR*(��L^i��	���' ]��9�=�7:��#=@��qe4�E�\��!@��Ǒ�<�;A0m�>����]�#���C�\#ݾ�3l��Y6{�\�9���������^7LB�f�t�>�Bg��~?aC�U%7�Y����˷٣�T�����s�"����Nۊs݊�t"bsf��/�,�3`�P���1۲~��W��ۢ��mْ�֥vo��Y_W��P�[o�b+�v��P��)K5��&�:x���l��v��M�S�x��΀
��cS@I�)�
d����kl���-�ZFrid��ǭ8t\/,G�0f)��U�o�Y��K/�d(�����m���yۛ�k��Y����mW^fKf��[�t��{�[�:���z�����]!�d��e��s���|�᥾��T&]؀�<3�������I ���9��0:D�h8�c���8�Y����T����χ �t��� &������1�dg� N�,> ��~��2�ڎ@���� �����x����z~�w����Xc"�/�ʗ��T�n��M��7�nw��F	�^���+���-�(#_l��u�Ͷm˥΅Y�t���w�<	g>�澼S)X\��e�J[<�Ǣ�)7a"$`�ɊB�w�#��U�̏�ƕ�lŢ�r���.Ca�8�p��n�NZ�iW�2�`:��K�)0��V�<�z��Œ�
e֓XR���JV�ٹt�z��J�n��|��-��o/?���=`7l�܎��c�A>�O�L�z�����m��9�X =~���fq�I�$_�d�P�[%/�@�����B��!��>x�_�!`j�㜊���:r���4�Q<L�`洧M�O@ F_4�B ����L|&�}&>�!.�L͐L߄�)_g|l�Ș��"��� BLJ�E�`���/����Q�B½�x��W�L��*&�! �tU~�!]y��g���m�>۷�e�̠M�8h�\��*�G���n��2����2IYV��PE�C|��A�`�W��V~�27�7&���K�d�L�R�v*gI㊇�G"��U�4��)���=�9�N�v���F#��|��J����25T�>��<�ԧd����7�,�T5�X.MZ�\�C��ZJ�352*�t҆������?~䠽�ⷭ05�C4�[�!U׌���b�
[�b��]��1�7� �� ��C����j���&-��#�Hσ�s�g<�N<�A�p��Y05}وC|���{<�=�$ a@�Wb��!.�A\����<@I�9�=��sZG�yG�-��3��k��Fy��3�6+m��նx�*�9`��ī*�f��}��\��M����	;|h�u��6t�?�߭طk�}�s����.�����$�%�C��"VLX���v
�ƭ��g�)�,+�k⹌����m���yW������|�9���Bô3�F�7;sqƤ���C���0K�(�t'����[n�'�|�.�|��۰���w�_Wv�y~9wD$ F�a83r�&��0IS.��.������r�*�j��u�T�l˶d[�gF�&p��Ð"� 	�A���~9�~?��^w�����vU��������sO����4�>���_qLH���}���cT���뒒Mg� �i�6��_��}��_��w=���M �r��l|�/J5	�s=��@�l��}�M�`��/@�0 !�x�`�>��>����k:L.H����ob�)i	��G�x5x�Gg'�x���$S�B�k�������0HC HG���ϙ�́��o۱�>��/���e��GI�W�_�W�JPwu��s�n>�z��;{��"�����|L��{���vn��/��˄L��O������L�����9�v�7�$-f�Sޣ�a݈;u��ե�G�E1��<���P��$"���q?��V�	��#_��KZ�l�UƉ(�z�ҙ�]��)��L˴���po8�<&�?m��߯�̞y�E;���vql�^}�M;�Fx���lR&�[�cO��y�)��9s��E�)��0Q��L_�'H f� CB�Z =1��\��&���a6*���M�Y�g��NXV~��L:�@�-	��d7nt��w��7�C =�SW����H�a�f�{�@;���4�dX� bL:�"<v�b��-����|e5
���6iD&/�n�����O?gG����}������{��!+�Z���~ �&f��^{�ɧ읣�[���̓��nj�+�vF�g�+ǚ�.�r>LP��3����Q�׺�o!|I �+Y�'�İ�q����A�j_7\iً��s��[�U,��VPc�y��d�w���3��
;=R�o��9{����f�66Y�\:��:���<n�\���=#D�#�6U�ۻ�S���&G��ԅ!;��I��5��J�ݐ�Jъx���S���o�w,ˬm��V�;<���	U�%Ƨ�/�H�� � �D����y��⃁ ~��ȓ �y�A)�qho���1AI�:?�ߔ�����FT��@>[��x�Ҡ�� s���P����ĘpV���*���j�Wf!��Cy�Ku{���x�z�t�u�.+J�9}���}��R�u1�
�ݑ�޳���JxNYIm{����M�d+��S�쵷[Yy���>rⴝ9?�R`���/+ϟ�U]Y۽s���'Fm���}�b�l�B���~��?x�w���>�����o�j�J�Xb��l?�:��0N'�~K��w�F�@�H�t��.�N�w�z���-1K�a㵆%{����Y-��#g��ۏ��:j�4{�$��o�줤��!�'���s���ή>k�2,���U�-�0߻�>#�%rҤα�{�U�
r�9�spd��^ ('�΂R��R���a��E��&X�~�o L�Ϲ�c�a�SF�5?ߚ�l�hN�Cs�s	��ӅL�;0$Z�y����F�7[�A�@@W-�� �� XN'
�o�7��8OX&_�١;�ve�$��3j��57�xYZ(�m�_�����z]���H���11�8�d��O��=��glx�b9��tE�lS�0S��ɲ�Տ~b/���n��[K'�LaYk3��yuq	a�+�w�bqi:�PQ�"�=��KvQ�sd�ONۉ�j��I�4�4�11�GN�������5b9k�9�bi�`YOZ��Uz�X���K�2'YK����䔈�����*k��x�&�!M˄��b�ĕ]�]�w�l����[��PhIa	��8D��.v����V�F+�,H��݉%���\�w���0q�Oa&b:S���$Dӱ���bUt��2����0�.3ļ�G ��HOO-Ke����3"J@c��j���1�����~��U �FP^�kz�l�����EgF�֭^c[�n������b�ܲ�ڮ*|zgG�&|t��2�e��2CU���"[�0.��T41��'.�"��x=�F��hJ陫�3��nz�]iB�=����	��ç��O<��a�*��L���O�k�VkU�R(��b�v�9�ܚ\fI�kX����a���i��~�H�ץ��O�S/�m������?�7����m���z�^:tܪ�$VZ��2	Z���ɪL�Z��cr���L5��od���#ӡ�4���� I�T7��+�!�R�6o��}��Z	bD �0\C�!��B�~hs�������\���g���k��o Ԁa��^�0[xp?ia:xh��OZ��f���#O��f���7����zŕ�J���n۵s��*N���|�vf���\�d:8���4QM���Zh3�q���Ov�����A�h���5V�v�o���߷������������_�O�h]����hH��P	k6I�錷���G�Ea�/;��  �@�F������D֒�6m+G{���`��z�5���)�r
�#��NE�V��a ?iEH���������Ji�X������(�����|�v�ΈH�ukȗÏ��.؍;�ۖ��a��oBB �0̿+�϶a���{��������U�"*�Y�<C�ѓ��������A(�l�%Pz)����}X�{�`!o�w0_éb�WY���������S+ze��H��b ��� P�@X�/ho�}aìf����:>I�0e�}�?'W�b�_yj�c��$cU?S�b��)aL?�LN��N��j�$w�ۦ�T2rG�7Z1��[]6�\e3+�Zt�&k���0n�ﲕ�q����yk�uYjX�A��zNZ
��2&���s3n&�8eL� 0]�fd$cS�j��(�RY�2Lj�w:�7 ���Y�(�º���
���d+���Ό��f՚b⣇؋��w|�;}�d�ê��N ��W
�`�J����X��51�||�+��߉�O~���=�!vޡ\�	M���ތ�c	��zC�N�y�wa
p������z�"!	��*�څ�L�zz}/P��E���֭�I+�ͫՕx>��Ĕ5���&�����7�}��A{��A}��l� ?Q��,��P*W�<�$I�c*�"
��B�ԋ�o�z��0^mT}ZۦZ��FJS<oK�D�i�e}
#�_�]�K���ǅ�r�	~IaQL�5ַ�,�`��T}F�L�!W�|�a�&d4���$y���L���
��ef�[b��)�x���"`!�Y.iK��C�01c"Ρk�)E��YX�3)�Ӗl��c����~Ӟ}�q{��'�'��I	�F����,c)�D���~$��|�5~3���!M�5u\�1�=m'&`Rs���W��%_��[|�P��uMo_�u:�1�w�"�����luH ��X���ŭ����6����=,�)�!C!0	ڑqC�����%(7i���F/��G%��5�;v���_�3O?i���o�K�>���.���n¥�谋d���i��j6)�@��_��jONs���Cl
�p,�zs��x&&�n��Ye���&h*!Z��*2)�o)-�RK�ba����d�K�v�Q��i&"�� S�����lVK�6Ӗ��l�@�﮴qU�ugT�ڴE��.i&*�FC��bs"$W(�����`���U%�
�ni���%fVk����`��%k��m�/<A8�Jr����)$>�8��B(����q����]�t�!�@c%4s)�3�xNg es�*�������"=�K�P;���i�v܈U2�KNl����H �hÐ9W�X,���qt5�an�F�O`���
~�n�(a��P([8pM]+U��ȓ�o�O'�k#�C���A�l�xQ1�Lj��)1+�����i�l�mMO�nٱ�nں��v�,Z�����20�k���ڭ!��b�M�D!hϥ�E1����#�	�fgdKg�L�V9i�}��ؗ>u�}�K������?��W�o�����;n��9I�1I7	�Z��Y�kU?���=3蝒�Q����帕�5'��|FNj��"1�Bc�xԶ:�J��!�֙��p�Rߡ!!R��s� ����J䀊T<? 0X����D<i�\�R����K�;ދ�4�
�o��M�/O���&�^]B�4�kH��zQ���z�w8Lqb�h�Jǜ���~����^B�q�Rї�y���y���ĳQU��@�,��k�XMr�VO�ؒoޖ�����R�&sR�G�0�8=�Uo�#���-:��z!V��-�i�����o�����q��_}�����E����}k'�.�c���A0*>�����E1�>	��0�,���n^�t�,�v��i�=��O��?~��۱�6���M�������~�!{����$���tF��_�a$ͦ��t�(ҍ��,�,0�!.����j��
��b�)��Қ�U��7(R��ĥ���p�K`�ف@�- '��ǳ[t��ء�x�w��脰��H:H\�	BmE��\��)̃��>�2�S )��t��7�7����Ĝ�t�����W;|��1{iك���ޗ��ȅ�څ��t��▅��3�0i�8�K��d�wIX�=�J��1�	��c~oW>�6�{�e�V�u]r�/���ڢ�Vt�o~�a1�}�wC��Z���ɚ�H�/=r���g?i;6���S����2B#�3u��.1����K�&��� ��d���W����m7oZc���YuĪ�g�9z���Q��[�O�y�=p�^_nі���fV����/�Ic�Y*N�/�^��	��zY���Pm*X��r{:Y�2��,�i�!��d�� �wF�εt�H�P���8#),"vT:!vbx@�B3�1�G�L޶ܰ�V�����>�¢Lҵ"-�.&`��B��z{�m���q��w�ɱʞ20A�̀�!*L���������,k�l�Z�e�Ĥ�v	8�[P��L�&���=�!����J�:0�1)��U�]M���Y/��3��C�E�?c�gN�*[R~��Ƞ�"�jIڿh��xV�15h%�z���I���U����o}���s������E˷��/V����dm��u�}��o�����_�HXX�І�����Wh	a������׳�+&��,�Z�^z��]Ve#��=���}7���Vu\H�]-�6!�w�wa�OK���]i�uY���Ysݳo�}�c�����ٓ�햛w�ß��ݰq�]<o{o��>��0��bU{��Oچ�l|b�J��
Y�����Y�m���j�V��m[lݚ�6!��'���+W��7�A��q:�A�0`�����R��\^�y�4��������<�/Q�� DO����7��hAb�l"��m�l��. uD{�!Ԕ�&�|�|x�<ю^7�KX���4W� �3u��Sj�o���p����릛��;l��]ֽig�W��ں����^{�_�]�w�W��>_��#�o�ͮ����/U�i��^���>��'m��;w�L1)�aS�pמ����7[srȧa�Q��gY߹[�\���[aG�?f��bnk���7�-;�YF���fkQ�	�yzM>�bt	��tH�� �
�!���WZ�e<���m߸�f��u˨���1UfrD����$H\�c5���~�%G]u�ļ{�	���g����~�����A��l�6�����f��[�l�]�7ڙ�G�cҪ7޸E�ZE&�\9X����s�}��|���+�/
]�D��f���z��i�=\��|F� p�Y��0:�.)i�Gzʭ�����I	"��L��ob֣�|b� 1'.��3gNK�1���?L^�Ѳ�1���K����rL�,��2/�����u'��ҳ��q1�f����O�����=b�rTm��0Y'b{���y[�Oz'�΍��(k����� ܺn��Sm]��O�ݷg��-	#�4��Ϊv�έ6���_sN��ؤ�;����L�P�&]�W����-��;Ⱥ�c� D�?m����E1]H���M�΄TzZ�ę`�TL���2n���t*aIє')G�*	��e�pN��)(S��Ǐ�kO��q[��W�:h��|�ΞzOZtF�����@&X�.^<mo��ߎ�wX�T�z��IF�1��Sv��Ii@�I2; �&��!d~C�U�����k��IK9�f��H�_�.z�N��ߤ% \��1y7�fe���\�~��̬����#@Z4-���འ^pM5�\Z~E�u|n���g!`����v��Y{�7}��}�����ݿ~Lnäo�p��{������i[��Ϟx���ǿc���aw�v�]�9:t�̈��5џ8���/��/�｛�?���`W�����~­���J�̰�3h1�(}�Y�C0�	����@!A�hEf�obF ��3�t�����[�2.�M����;}JS6���ҜH���j�g�Ng���o|�^�o�m=�}*���Zӆ�'��v��1t&0����~QF�M��z �����8�?C`�On��I.��=|��|Y�<b�6E,\����ChP��{av.z�;AF����+o�N=T��;�Gj�y���I���6�<CX^�?��ⷧQ>l}����!6�.}��|��#v��9+1CEߢ�3���`���ҝ�̤�����d)�9]�t�޹��~����^C፭�=s�J��Gb�Ù?\C'~^:ڎꃣ%�E3]!�zϢ�npp����R�.� ۡQ�`][Uҕ+��+lLf��Ș��,\��N�='�p�EY_3�m�n}(j[�l�J�"�6l���1{��w|haͺ"Ԍ�e��6&"nZ2��uu3���ʜ��Y�&� u�pt2�_�{�MxvdSb��Y��S��%�5�l��/������	ǊCM3?=�B��ZA):�����1��ς� ��ͥE��ć�tN h[ӷ\-9��lh@,fm�a��U>�v_�a������k�۳?y���q�mؼ;��������=�����;GlZL6]�Z��%혬��#t��Y��ˤ���D�-	z�y�:?�3�ʕ���4Wf� �D�����Ho�>��E�XWA0��Y;SI�������?p����l�@������m�e2ʩG�7c�\�/n�͸}��w��o�ޕnj0�ң�b��)K"�|.k� ̀�t���9�:)7Ǆ0��T����0��-���-�*پ-k���lzt������&����n�i���o��$3h�����ge -���wU`ro��д���}�{�j���ĝ�B�}��[X���^N���#���3顄�=��i�x��6Zl�G��{#5k�
ކ�ڏjT;3Wd�!�����,N��V/�E3Q_�̒-���$M�%ga���T��~�A�K>�2-�F�����nĬ�[i���}��g}��Ly�~�����/ZD�#Ѷ�3�r������:���K!�} �(@�w:��,���0aʎ��`?����?8jEi�t�ߗM��9k&�vn�hϾ���Ŕ~j�l�l�@��*-���I�����3�'�X$���rÎ?#{�GfdۦJ��!�:Y�u��$ە�]�w������rlH��C�Ks��: $� �qb�����G�=q-]��MŮI�d=cH �F�נ�>�Z�]-0��05`�����7dD<;̡k&'0q3��,�ڨW%�fl�lӦ�����$H'�e�8����5;]��I	�V,X+W��7��m��dQ���E(�;AM�����^�����=���3[�h,�n��_V��/�.Z���V���2��=�5�)d�?U- �%�E1��nRAB��n���b�T�^>��=&���OߴC'.�Pi�NMT��7�w_������vN��L,-D%%E�m�eI*5`"��YؒI���k��&%�L���Ya�Se���Y�����g�[�aB�ٹ]Z_#"�U�"�-��%ܧ��~Ǘ`�Qb	���C��3�G�g�K�6_��\;#��R��>#}{^���c6]z}�4�G�y������e����B���P�2O��,)�z��t�:	D�*��"�=����]�V�<U��9��B�hDB��b���dE�Y\���`o�a&M�:��9o��Gn��߷׏���e;3Y��?��S������0j�L��ʗ5.L�/�9�D��l�%e8`���ه����L !��;UJؿ�wj/<��wY6ڲ�Đug㖑Y�A��p�Y�##V��D�%r2�Ү!�z;+��c���^iv�] &��h5��%�stb܉3!�ӳ]+�i-��ʸ�4�{�3�~��IISf�4���`۶lvS���pR��?��ó%��n�� Ӓ��A��9Ӭqi�\=�^��c�����~ ��w\#�`�#G��zL�=ݶv��G�VN�m*�gr7�3	��Ba��I&�Z �]��x8��M��1������:�b�Q��E����D�82h+��ϱ];�	ќ�%�p���YbU�/GG��9�����ޣ���L�W�d'�3��o���F�p�b��Sb�'W�[%�m
i��i�'��?���s-��%�&��ʴl�(�(c�VU1\ݏ�m2������2wl骭��~�� ��!=��;�f��Ф�F�@�-=P�z��m����ïX!����R���.A����'m�p L6�11�y�>
0^�G+�mLV����J2�ܣ}/��Q�����%����`�Y��aB����a]��E���0��>&S�,<�Ħﱁ�����oN�΍F�sP��xGm.넉�t����x�89*-�l�y���n�3V+4�ҹ�/p������|?zɋ��w���>nGgV^�:u�����~�s��*�:�lf�63�;{W��=��3�"!h�aw1�8�����=U$�0Fdc�$���hu�߬��YE���LX�JWz��+K�1��Se}��B`ƶ�	S�L��1���R�Z����Y����ɤZAt4���ů��Y3���vf	RЇ�rΙ(����x�Z�vNf�{��G׿o�R9��Y�Ib7EU.�&�7���A`s^Bn���)A�Kc��G�A�^1������}����c2�o��3�]'��>1�pa{x)�ejr\�$�}�����s�Ɉ�w�]0&Y,�����JE'U�v�E$MǪ0�V.�尔��)�n�F�_,˝IuY3�e�b�i���o��vnӧ���;��[�˵ZB��t��-
1ߤ�� �xo���l�l�*��J�����d��$"��4]�U�z_�l0�i5���4�н���,.�KQ�F%���*���,�*��L���4>�qSN�şSѼ�������ѽ� ���ix$!C�o��7�	��>_�Ο1�Hͥj:P��E����D�ܷ�Z���4E���P�ؚ�N?���wm����'�ڬ����R=��>����>2i$�<����]��}}��o��� Bf�����S�h'��&_��x����U�^-	g���J��K�,K��5�1� g� �M����L�=Zպ�LF�lR������3�vi#}�C0� ������6��p��Z�_��˴�=��З[���i��Q�,L�(o�A�_�Z��Ǩ���gs��6����D��ƬqC�:i�cC2IՌ�YU���r��h7���h	I>6��]�|Ii-�)af9�k�c]��߻��tJ��ly0`E�`%_��r���*3f�5Q�a#|{p�s^`5{w��up��w;��3+v�U��d1��T�s	P%�)̇�H�>���!��-�
�/;��{l	���ZT�Y`+t��A������c�k���a���6j@т���,���N��g3-��`�4-�)%���ԅ���C�Ppfn
�<g�8Z0�$z�쌬"	�vq�b��hQ�U���+0L*����}�G�,9�-j������Zs�׳l5%�f���Z�~��;y~��L�UF�[Q���{v�����k�����-��I+M�Ik�Ʉ5_�#�F$���eM	� 5VC��i��BNĩI�F�;�s1,c2L��*�ct�Ȭ(�O��p0f�
��~1R��k�[qT�!�6iɿ�|6�}��<Z�-��rv��N��NX�s������Il�g���z�w6�S�
�_g{'�@H@��]�O��~|���Ӹ�cQ�����q
���'�M<?0����W��@:�f��`nVL��|��d�y����Đ�鵈La)J�$��#)���mdP�9�=�cU�Y���@(�$�J���������V��V؃�v��ݲ��y�m�a�h���U�)��񒖒صi��y�_z��L$K��3�s�W�����:R�=���J��	a�����6��;����ֱ���o��1۹y��+f۳{�w�sȟ�:J��8;hϼ�����a�,rE�,����{5_�Ȱb3Yf�W|����Ϭ,�*�� aV�˄⭒�T�`c�N
iUG"D�u�8��P���ɼ8$G q�{�a_��|<b�ҽ�%�&As;��% �8��H�&:vİ"�/�!��F<
��oqcr�D�.�;�ɔ/f�_��'`��u���T�HA���T�הG�P�N�ಡ6�{H����a�%��ݬF�`~����q�[0�-���5$:a+Vny��� ȱ���Ț}�;�[n����;�B��)5���_�K��2�!����k�˟�x[ZQ����Gc�|�����J,,��F��ģ�(L����j�����{��y���-�������u�nIm��9�Q��lrw�僝������k��#]p۟}/07��lL�dw�k�,Hy�>�`V���c�,Hg�s2��fG�h�h��A+�]�.cV?�4�|�ڵ� m 6s��v)�Aȁ�D�-����R:�_��;!S��4+4W�|`$H S)s����;�ahF�VB��0��! r�_��=>��}JW��S��{3��K���a
jt�ا�ׂ��^51B�-��g���]VX��"��j�Q�%f�m,��*������ǅ�d�TJ��~3k:m�A����Nد<t�=r�>��fy�V��%3�"ٽچ�)�֓�۳���?=b_����[�􈬶)��a�X<�޼��?Q���E1��3��5~�2�EU����dq��տ�c{��{�#t�ޛ��O�z�Q+N��:/z�2j{TyeF��o�=�3�xUv�>�O�$�z� H̉��W٪�+%զ�����v�6l�#G��s����Z˯��a�1>��"�KJZ��yxpy�dF*"�¿�2'�����LxZ�K�߂�|��f�c)�j��^)�60Y��=�K�ғ�_���>�r�q��ls~�O��.���/r7Ԥ8�t=?B��_{ FsSW�e"+�0�ƫ���.�\�k��Q�T:!:�J1۶e��[��Ξ<ii������
�c؀����	��u|��f��o]�c��k������E�	�5uYN���+��c�E��?�3�1f	�z_��]�~�6Sg�1]�P<��?����àVK����ӕ����J�F�a�*3	��W^���[%��؝7۶u�6S��i�ҏsߴ��ec���+�J���ਝ�8,�&�\��C��c�֯��[7YD�a�Z�/}�S��̤�~��}���`�l��бr�؅�Aw�GOTD�Ì�j3�v��J(�n%�.�ۉ�~g}̑!�f<'ӃXRS��]!�{a>J�׌���TFi	y�\�=kz�u\���[�+f��j���U������z���q�Lȩ��ʗg�C��S��ޣ��{~�kb�WS\S:�L�)�����=3�7um��$�v�c�/���PO�KL�M�A~�y'�oΨ���l��4�̌����j�;nޥv�������){�s�}l�u�{n�i�7�`+Ew�֮���!?�+�4,��o�c�ˏ�M��v鎈N857����tޙ庺�Թ�64x^>o�nܺ����%�e@"�x���4���@(��	�f�<$U$S�i=Hj���͉TXN�lK�T��֝��K#�_�ԫYO>���|@�W��P K�_}�y{��g��f��}��?j�O�/�L:CL��c�
�ŔS�#�ݼO�;d��IZN�,��?��1+ь�Z,uY\S\W����.�B�<�:���U�XIR�2���|��B�~U��W�&������4�%߄1˺��a ��1#�B�j�`P��QQ�j;i��6�P���;k%�S��<��wN>�|�V��R��	m�8X���2�	�jͦku+J��Jʻb	�O�RV�(/I�g��*ktO��<�ң���@�<Hs]�r�mJ���p9��!_�����!�Ї�GD��D�[��F��EMFm��땟�i�J��$lr��=�����m�:��S��x�6�[����l&�vb�m 1�c��<[��H�oZ���I����3��^���aQL��W����4�E��Ӿ���+�:!do3���ZU�(&a�]��%/��%�a`;�J�~��VXY����t�$��~��xL#JI��8����S�u�f?��df[��)x�%@`�ja<?ЯrIE���1�>iU���T��=z�B���bҵ�^��O��0B�ӕK�={wڮM2���uU�6�Glǚ�mY��M��m��s���x'�%��Bz�VfTD��^�ߣt��歫m�@¶�m���m_��]Y۵���i�ݶ{�� �vq�-�!`�� ��\I��\�й�i煠�s�9S���b�����	L�`H$	i��LJ��R�����ׇ��}���	l�N���.�e$\K%��E���[��[Äxv����w hl�,za�����'�w��E�N����E��'�6�Z�_ω��E���e{�#6<6a�l�6I�o\�¢b���<mqj\�&f��)K��醽���6V*[&�s6l�޽���,)Dx󐯱{���������Q_c�k�;~����ݢɌ�;w����T�� &i
�Mgx��B��\{�N䄢��N,b��q2���;h�:��OV����+B�Ͳ̥����<l[2�k���)۲*o�{s���`7n�j�ɼM��	�0c�)�e�g�(3F�t�������~�6�L[o�*�M���=ʯG��m�@����(!��Ο=+b*I�!��	�FQ9�P�'<�^Qƾ����T1�=��s�\�ͅ8���@
z<�߈eRq�	@���M�Y�}ᚎ��;���-��ןr�|���';D��7m���{��]�;�4��r���m����d�_��<`f@e��6Qm�v~�̓v��iw�{��U�/*SS��)�,�wyfu>��v�`q>�����	h1���7�����V��fM�l�]y���e������L�x����u�^y��̩`��Uϟ���Q{�����[�X��c�x��'S�:w���{���MeI�c�Oر�'�!d�=���*Ӂج5��Zt.��M�7.��]_-̥��dt��T�i���xC�=|�NK��X��a�i�X_�dٶ��V��"��k|g����S���'Ǔ �T�l�a�ƴݶu��޽��c'�|�u�'-��|k�2z�Oq*�N�ʬ|�ͷlB�LLma�^�*����:���1]{�;�˙��0�3��܄��!�G�-�F��� -�d""奲���q��G�6x�^&�6::n.��م�/���3��h���S���vah��s��'�b$��rq��uYV�6����]"	�g�~�8-"7(�u����ځc��'��m㥊oF�g�b�j����d��ğӽ�.�f �|!����}K�a�&�U��Wߴ�rݺV��iI:5�;���xa����{慗}�;c*1�pJ>ȁw�ڙ�I����b�B�����v�C#������d��<q�L�<��;�=���W{�;�Ü���o��悮тj8��y��(�C(sXL�i�[��b�DC�F]��<?v�bpB��0�1X�����,������-DET3e��3#�-�4bZ	��rZ3&�ƶ�l�Yl
ޮ�w���X�ʁI��8�K�~X�ފ� ��%$=��h2uU?I�� h9!�)Hځ�G�(}jh�;�FE_�F&�,���g%�g,߽ҪM��u� ���8f�~�)YuK�e��,�풖��Z�%$�<*A������شE�}�U/�dPQ�Ѭ�C*��¢��r�� �)����Dtb0$���/�cO>o'.N�L��ڙ>��5vN�����/�����0bMe�:z�*̥�&s]��L�����%{Ĩ]�6,3�ްt�
}#�	�蝴�[�U��|rf��z�'a��'�}�u����g���i�{�gkf#��it����<��j<VK�DD��V�b\�e=���C	��n�u�	�["%&���o��"��|u��S��Ku�h,-���EP)	��e����i�?�9��܌:qfr����v?VL�%ù����q���A�&*�_迹&�hKך�Ø>~4�N2�>��Vl�橌/jm�q"�J<%Ry�6��9mf�(��Y{��s��������c��6&7��,X#�k��ٟ���v��	����cJ���L	g���%Xr��?���3.W�XM��$/���������wO��db-�=��%m����2�XNQ���̅1;74ic�e����8/��?��Ü7��=b��|>+DN��48��Ä��!&cz�"��u���ˀ:Ӆ�&�2f 1b>p-�꾊�>��~_m慃�DB���@c���(o�-��R��]W�'��c���6y��������[n�-�������3/�풝Ż�<R��ʛ��x�h�l]kwʯ�M2縥E�lxDU��t���v������lH��I��h}�'i�M3c$P#��Y���|0�b����Iq�� ��&�t5e���At	(m@{|C1v'�Q$6��u��@발���dA�W�,������N������(�Ȣڰ�ߧ"2���3���X���~J槄OL������о�eA��j���h<������3R�>u�c��~�*&�j7�t9;U�ٿ��������@U4-KK�U��}[>Y���j�DNRk��#��F���P��_�`�jZHdژ�e��uΦ�y*s��`Z� %Ee>F�}i[�Y%B���t���OA�C$L�Iʡs>�'�������}ރ��k�U��ZIμn�&��"�FI�Z.Y�h"�᥶p&B��H[(4����P��Bf�iF�XLffN~��	�
32@ab}_�@�,F�$ӌqB���nVbr*	y(?X-�OPf���w����0|�J���M�<W��M��\��`�,��@%l���+��ZQ4�*��葖�#&d&=��T�B��s��X�*�+�I�u��"X	��Dsz�������Q)3�	��C?g_�҃��TT>Yo���D2�O��Y}�g�9��3��?X��3���?S�ؿ��o�O�x�Ry�K2}'���7���F׷L�������fAw�4����r��1����+|쉕��4S��9|���`:7��dH>��`J&�r�Q��u#����'����� ��Xi<���T��a3��	I�2LhfL�-.�4+Np̢G맺z�����B���`z��������IY�Z2v�N	͜��j��.�8�iGڴ��e�aBM��`��ލ���Ƞԍ�q�NO�o��]	:��,\���Z��?�R��\�X'Ѓ_�*+�4�ͱ
pkG��9nѸ��i�)�`�BNע����h��<`�h���&�'��$ ��E��?��{���W�:=�hh���s��?�e����Ǘ�t����O���S�V쉲W�ZlZ���;��{�.H�,��W��D"6��<7��
��baC�f�eX����pY�d�g�������0B��2ۂ"��������q"���9��5�) �@���U�G�� �|�N>F���|���:~��~��������q�FE��b�R<��2��B���� ���^�b���
��}?N�]Kw�1u��f��5�vˎ��g�6�nJd�D�������+�&xci`QL|��7�p�w��F͘�ڒ��s�BK�L �0��Ml�$(��u�\��o�sf���?(��w�b�5;-�1�4�Ůp��5��]�}�������k=�\��׎���P�,�Iz����q�cY>#DD�Ֆ�*<��jJŢ�-D2�eQ�^����L�ب�p��U�{>w��������sn���?]�׳+À�*CoZC��O�e�w�{�0��ha^L1s�ݤ����}�xa�c6ɽ���ﻦ���x!�^�#��Z�Zp�հ �|	�t������ʁ�v��&
�������4��fa��:�����Y8G�-͇�ѐPJ�t�f��m6<扖�t�kG�=zar�wV���gP�V���[R��$�v���F$W�������C<�L�рs���%1LM|%3���Y�/� ��6�FK\>�|�y�?�`��5�_��-򵛢Yi��c2`��Z<r��n�����D,F���b:୓�>q��������N&Vf�I�銟��J&'#��L¢�hC�h1���SA����]�wј��ye�v�%�y�{0!Y^����\r�/��K��P����N�f�F�C��S�/d*b��|��~�x 
]����/Gj)��@�f�������a1�R�f"������0(I�c&���3��ݰN���`���g�ee��{����<��WJ�!�2 !Q�h"i)f�����j��n6��˝���u6����K��z��>uqh����J���@Ή��!�X��l�S�6�xG�jK�A^Po��Ɍ�4(�/�:��
� f����z9�/Ѓίk�ӱr�"z>A+��,�:*R��;�C�τ)bk.f^�����Y�b'ߠ�07��>��x�}��3�X����#P���ς��'r���_�%��]��c�B�N�������D���L.�����a��CPN�^�w��}�<�t~�����z��t ���yٳ+B�����s˧�y�uOaۏZCz-�Kb6���`_>�ֆ��W{����O@�u~�� fL�6n�堒��! �pv���R0���e��e�/�J{\	���s���J�0͵���	���a���`�a�#,3�2,�u�e�[�e�ΰ�t˰���n��:�2�-�2\gXf�eX���L��p�a��a�3,3�2,�u�e�[�e�ΰ�t˰���n��:�2�-�2\gXf�eX���L��p�a��a�3,3�2,�u�e�[�e�ΰ�t˰���?^��(�    IEND�B`�PK
     ��ZJ��F�  �  /   images/1348d1eb-e6ae-43d4-937f-d455f2ad4bcd.png�PNG

   IHDR   �  ,   G}�   gAMA  ���a   	pHYs  �  ��o�d  �IDATx��y�\�u'v�~{}�@�$@��Nq�(Q2EQeɒ��Lkl�cg<I�)g��#���JR�+qR��8�*UM<��Y�dm)��HQ��W������������~�a�~�{�f��}�.��;��~�R�
)�����TH!��L� ]!���� ]!���� ]!���� ]!���� ]!���� ]!���� �I�$~�T)I����M��SE�a���_Ķa��aD�i�eu��M'�@��p���|�i�w�D[<��	�˯-�X�i�%�F��]Fᒣ���$��i��f@�l
)@��ҍ���^��i��߸JMՉ&L2*��a�lc���y�4��VJ�%�Z�f˲>�&��t��^�B�^
�m�DI��t����n�hk2�\6+�C"��٩Mf�)2�3<���n}z�Vo(��1��i��v����G���� ��t�Y���*ن���	k��\������t�	����Q�"o����N8a��[���a��	*d�� �X�2�g:�k´-7I�ec-f�r�%:97� 3d&[q�����K��3��w��K��_�Ӷ�W}�����6���Vh��t a���U��7���G��*=����_��:��:��PI31Ń�X�1Ӥԁ;S��>q����m��C;&��f��45L�Z��t I���coe�Hq'�r�J�s�����3ϒW�)�d����ㄭ;��mRb�������t��+��%�!ˎ9�Hk��>2�R�n�Ag�.��-���<�R�f�e��v�S�1݌�-��M�m3�d ���┵o]��k�Mǉ��P!C-�6@Xw��57�<fʚ,�r�B��̧��|���&�%�~,�c�J��&��B��㟤w�|%L5}&�A�~�
�ͥB�Z
�m�0[4��$���f��>�~������$I��5M ��A ]�tإ�A #a<9�Ci	
��&}��_���9*�<Fe7Ň)(�������{>D���N�#�N89S�L*d�� �FH��K�a����\�����`8�̴��[컁m54e�2�R�n��bh�IL���J���:}�������1�Z�>�P�rP���G覛n���>�Q��B��6��� Q��z�.Z��r��Z-��Nn��To�6)@��
̶lJ�8��V����/����t�uVF��o~����E���K�	:BQ�]A/�\
�m�0�0�-�y`YL9m˥0�(R1k���5��eZ��&U**���lQ�;T��
�n� ��c��M'i`l�m߾���>z�G?���%��4��?x2S��<�������z���,l���A7g!C)�6Ft}��2,�PH���@d��~j���K<///S�ە�A3Ơ��^�r� �H�a�l����.��.��633C�jY������2�рS�{��}쾏��}�Q;h��ҢM��K��6��Ei2մ%�v�%����eFIB�kd��I����-[�Uy�����f��z)@�1�\�P���R��]$��t~�������aG`���A�����t�u�I�@Ebt������ 1$�l1i�'��`�As9���mHk��4eLBqH2�A�v)@�A�c�4Π�V+�%�,�$�Δz�J�@@X!�r/�3A�s���~�>��_���]J�^�,֌(/���a�t$LS)ڱ�>eܹs'9�#��Sr/ek��Bh�ЮO��JU�O�<��l)@�bJj{Ҙ��(
izz�~�3���{��{�|ۗf��H��v���r��ҍ7�(�Mo'67�}C.�6Nx&*IR
��^{�5ZYY�N����_]����9����T�f�t$�V�iQ��s\:y|���H�n˖)����X{�L1d2�z%��~��������
�D:H^��6���Q�����b�Z����z�{�V��~����:���C��rH���4�y����~���ͯ}U��� vC*�j�%@���[�]�z��J$>�J�
n)@�A2��V�E���q,��u>9r�������8َM��Zn�H�dQ"ɹ�x��5ɵ�t:��o[�+��h���t�?�8���t��WQ����*v��� �	���m�a�!��R���������M�{�P���w�^ڱcG�#���Q�+d�� �*Ǳ0����z�.MLL�m��'O�c����o�p�=����H]�#�P!C-�6P �0�_*��J�x�:~�8��K�+�Z�3�<C�o���$塞yP�&z)@�A'�aۖx-���f��{�,äDi�fU�k[��j쩧���G��mw�JA/��1֍�I�E����a�]C�D4R�H70��\z�� �0��ҝ��.߷O�/�-�*�?�mP����� �h��P�B�v:4::J�����G���>$���Z\o����w�I7�|��_�֥�s�?+@7�R�n�D��$�j�Vz衇$Tse��i��Xl�W^y�.�b9e�fH*U�E��a�t$�i���b=�0�������M��e��~e���^x�^~�eq�,��%+��6TZ�nȥ �I�0�����,r���}�t��?�4��>)1k/�ﰞ+��@��ޞ={ĞC�L	��֨�B�R
�m�T,S!��dP%QH##5z�i_���?�?s�l��-�g�4��d�RK��K��"4��<�Pt�.�6H:����KV�e����"6z��K%ꅱ��ÿ~��l�h5���}��������/$YӮ�tC.�6HlK��S�ףJ�"�:�iH|v���U{�R+0Si;�9}��<�:88hP[�^��� ��3�
�c
��*z���G�~�b�0�	X��V[�.����ڵK ����-{F�6�R�n��l3H�"�t��1�\����irz�N�<�h���3������=R\���v���+�2�R�n���h���Ģ�����o|Cr/%�2_{\j��.�J�{�<M�t�^�NIb{�[Z����� )c:�G�+�_������z�G�ԁ��9�hb��{V:	1�����a�t$a��u�<���^"��'l�u�m�;��k�̥+4�[�#m�R����, 7�R�n�]S�X�T�K��� *W+��u֦�7�5�L�K�NNN��N��2����K�a�Y=���b������z�rI��n�{����c�=&C^�c�hK�+���^���QҷY�L���#2J�{�y��z��x�f�,]G�_��t�Y,	�m�e��,�� �6H�2�J�R�$�=h��O}�zE��<�?��r ����$!�HE�E~������K���1�+&�����yl��D�_׭y0l۶mTib���=����W�nȥ ��J���ZY*�ii~I�)O�:E�j������y�i�~�������S��+d�� ���^�^�ش-�� �B��5�)���/��SeKcYt��IY@)`q�E�cKp�4�b�!�t%� ��8��-Wl�g�z�bw�����>h:��;�H}�{�뮥�ףVs��X��rȥ �F	�ǳYKE������5�Ϝ���Zә�&���eHe<����Z}�ϖNb&9.�Q��5�R�nD�0����N�<�VV����]�'���2}��Vy�@�\�җ�$	ϟ�Ľ�tA:YW� ݐK��%�q�PE�A�xݱcǨ�h���i�{��(&bvif��)�n�&.�aL]�4���� �vJ�V�iaDT������g %��<B�֨��Dϲ�Ę���t$�aw�2OТ�Ȓ_��{�����Q=c���[�l!�u)�B�~�%��(bz)@��t�$�����G���t��: ��_�g��)Q��|�Y۽�����d�Vɒ`;LE*d�� �	�d坻E+lˡ?J��$wtTW��Iκ�l?�Ph�v�M���SqQ�3�R�nDnD��t;戩�֭[鳟�,=�ԓ���Ȉ�����8"��Ib�,x/�G�� U���E��!�t ��6$NL�d����ڦ�Ozl�%�^���\KY���י����� j{/ҩ���r)@�1��(U�ً���xl�-з��-��*�*�ǔ�^(`�LE�v@k;,:U�裏J=ݮ��}V\�\�o�X@d� ���F�q$>�~
��抰��8�r>I�iD���q�z���U��8�����^��� �M3h$�3��T���������������铤A]�\�����@��ߤ��aBb+LAZ�q��2�R�n��:�+�C[&F��YÅ�.�~E�#�vl�vs�������E��b�X�uzm��w��|����i�]4=="`z	�%�|�+M����t ��Y�j�G�4��j5��ے?���k�����џ�ٟI��R�DK�Җ�F�'�rbm;�T��hg��}~�c��B�Z
�m�L�k�qf��Wl���Ҽn7$�6��nR�V�Nr.ٞC&3�w�d�Jk��r�?q�-����Ŵ��ӥ���k��%*d�� ���ё�+Q���]0/���ó�IK����m���ΠI�_��=g 2Πs�9�A*L(�l�l���4ۙ[�7WM�<C����@�bj�WN�҉��|�%�Vj�d�x�����T��L����Ex�fJo�O����ɱ/��آB�^
�m��UJ��[<��6�5vX�!�C�;U�:�~��<0�N��~g��
��&�t,#��\B�� Iz�A'0�ة��ydy���	W��I�v��5�+<��H
�m�������������6��怆�H�B���0&��%pbZ�Q!�F
�m�0�L�hRT��I,E:9�4֦�?^0�Y-J����Z|I��0�$M�N���4���Pr��_mNSN%)a=��A�m�6���`��9�N,����H/��p��R��l���#YA>)�n")@7� JP9��1y��︀�@9�4ͦ�ߪG�5���*��6��A�!M��B(b]i6i�V��3�NK�8��-Y�A��,�REg��$�A�O�U� r2A1QL<��}2��j�B�m:)@7�����u��3ga}ˍl�c��c-�1�^�ۉ}.7���]�:@}M��I�6�vh͇m~�0���a���$�@��/��o�NW^y%���}�{ߥ^|�~��_��~�z�U�$�H�_���^n*)@7´�'����۳k7��?�Cz���������t�]wR�mɂ"��2�4l�B�_
��$�,���9h�nR�R"3apEL7�@Z�ix�����XI�h�W o�H�!��(M��2����%-9�p���dG	9�0Ƕ(	���t��,Qh&�5�p�I
����`�c�z�������$+��֞pP��2sJ9�e�)�K
���)m�ԙKL�c��u�<�;U�w�d/�W%B����r����ǪNv��LR�ndK��E��t���_+��K�6�y�PB<A��&&�zay�������b[���M%�D������i?c8�B/�9�I^��T�V��5�R-����JE�M(�Hʾ*1���:d�P��
�̫RY�y�8��T��lN)@7D����ԨUQ�*�=��:uYG0,ԓ��J!�R
���61U�x+u[u�bb�,%9_	�=�k����&�H�O	3N�1���A�sD���lL�P) �9� ݐ�JÔLL�￯3-u�ΔKbmR)@7L�t��V}1׽��	� ���2tx@k���	�*���Vnn)@7D"�OLi�AǏ�j&f�cuF�#�Pv�T
��(��9w4t�3iՖ0�"K�s�J�!�H���HW�Yb�4#�Y��T�h��R�n�Q��԰2�Xo�)醳�lN)@7L�Ȱ�aZ�j�0��F�k8:@Ο�Tt�Y
��HY��D�wP�+�X��|Ud�lN)@7$��*�,#�O�t�:3t�A���@��tC$��`i�H�%ԛ���%��I� �	3L3A#>ǥ$�|�lC�;E!�M+�I�T�AY%�_] ����*4ݦ�t(�V�V�%�_����%Uޜ9_��Ț�S�33���zQrń�<��7M����N�M+��!a���Q<��{�{Ub�h�R�Y��&Biʰ�����q��h���hS�����;:�[MTB�ԬZ�����I�ޞ�"~#�I�y�K�9DE۽�*��I'�B^�b:��z�-ʣQ�X�<�m�G[@ed%�Y��t�2���{���S�xK�e��;�J];JL�L)1�QL͕U\�J���+�#J<��꼉� ݀�è~(�~ׯ�~�F������61 +1�̯� $�fE�H���;�vB�$*�;Vb-e��jMX��N��:�B �?#�=rJ��=�=9C���4Z�}:d��"��U�2�)� ]&A�v{��׫�����i��N���:������-���ZHCj}$�F�iJy-�h�ٺsǔ�^Od��6���^-�b֕Aџ�ɟЏ�x�~���1m�~	�{���i�z�
ٔR�.��v�z�^���a\Q��b�3U�W�B���
���P��m��j��zqke��/M��5�S�\��f]O�nŐ��o�٠��%��o'�f���ң?x���v���T��P������ha�4g��M)�XA0����W&�l��6���(�/������O��^~�%E3�d��ئ,E|6ɣgh�=+f��(��$K0(MJĲc�F�p�:Ӓ��[���������]ӻ��X�ƊIc��Je�
ٔR���h�y����{K��&���Q����?��?���)����}�t�N�h�ҫ����/�ʉg�������$N#J+��͠�z�U{�+�Ee�N1���[�����,�/ˎӢB6��܃.�?H�.
��g�&Ky�w����B5�����?�}��ǚ/f0�YJ��C��M���n;[��xU���yn�`"�ޒ]�L1ۡ�P���Js��t�rlz��i��t�0�mo��oWU;$��ӗ��5z�����M���BKYu���;-h�Z�{,s��(����Y� �A-�$�0a�ɚ���Q�R��ՙ���[�+~���_��}vn[Ȧ��{�EqR�l��Z�����9>7ۉ���K^�LQ�K��r)�+2f�E��5��tꖙ�Рܒú�vF-��%-ҳ�͆��é"'J�8柣�nt����,���vɣe�-h�&��{�%i��q,�p@�X��e2����k@X|�|��':rz�DH�Ur�X)�L�L\�`��&��
F��w��
������)����HQa�&�B��jw��v��Ɩz�+WLO�`�V;N��g!?����-��Cs)d���؆#�٦
�V�(\(��/,=��8�﷎�>��B���6#�LSe�*__G���V�y�>�4��1k�7C�+���c���#aəll��a�fB��g#?��c�b�f�pA	��F�� 2-�"�hĶ=w���x�
)䧔�{СEBB���~w���m�?�l��|�
be*۶,��TH!�@~�A��-F��7��z.��
9Ķ�VRK���F�����Bށ�3��VF n�!ŀKRKR��c�b��6E�*C/�-Ӊ��Bށ�܃.[�M�"�	�Pk���"**��i�Q���Q!����S�.IS;H�r���K4Y����O�=y"ڣ�V�;�J�Ymd�l��F���w����W|�1&?�4u�����c�mo)6��t�J$Ԇ�����X�an;�m�eZ֣l݅��e�/�v�uT��4��)v�X%/���[�ݼˬ��2�'�TO��_3V����[�����k�����?~i�/���~Og���D*W�8�lG!��yUo�[d��&.���� ��T΁:�,�M?y۠���u{�f��W��{�m��<>]�ۣ�4J"E��K6p�/���ٶ�Wcg�8{-�T��m�\e�����U�7߲Uy||gɤ���_b{�LٖK$���X��6�VT�,y��<�_�4͹T��][[�}� �9!)�{ӱ$s�g��;�`|f*�`�����a��X"|�C�,���\���/�]]��*	ϟ�k���տ#kY�f k+�պ}��*:��h�)�9����B7p­�4����Vʔ�چ\c�YV�M��W�\��k�=����nU_m�?����*�ֺa԰.���-0��ý?;��R��C_ɔt��TNټ7��q>I��H�Կ�?y�PY+ִ����߈V�	�]��q��F�BDN�I{��T�J�G<<e 2���?�$�]۝����mM���T����Q���]�C���a}'ˁg��Z�n�4���Y�����D��V�cR)J�@r�5�#Zz�V�u�5'�t���y(��[Y����s�1|�����w*�73՟#�%b��.�]6�7S)�7dw�.D�y*�T��[i�����k��&E]�b�ۖ���R�|gK��1ϝ� y[�{����5>�/Gc����F!Y<Gؒ��1��i�Hteh�5�0��\C�9�Q���݋l�7��^$�`��{�X���Ղ��������F�MOl�zU*%�<�������Ð:AH���(�8-��N����@��,Mb�Q.�\�b��k���V��^� ��ղ!,��k�����h�yA���N���?�|B^������!<��F����q�15_���Xi��jG9�^xLS\�2�nJ^h�Jj�;���8Y;�0�ú���E��|�s�3>�;<���j|�.�����r��^ޥ��w]t|v-q�����k�`��[O>���Skp���ȇ�%��n)�	��Y�%N�R�L͞ZrkuJ�2��x X�M䯯_8�uz�M�^�64Ӂ�ٶT]k-������Ȋޡ\��y�l�g�.�<?����[��r��O�TO`��+J�� .И��^"��S��\��O�"��n&�~a�Tz�����:xd�Z���;��T�yTc&2�^!���Ĕ�S��,K_�Vz��/}�e�� Fŵ%ϒ�/����fN}�\f=���H'GfJ�w(�d�M��+43��mJtxf��>�:5�,)�o���_����!��&����V���A���g�btZY�k�6��)���
����vO�o�S*:�3�OG�O�L�ҥs3��L���(;l�쿯��K��`��T[�6�F��G6kE'�Q�����$;4���t�4a����;^-Ӗ�qRݶ�j�[���f�U�u/j����m��r��S��]=��������S/��ʹBt��&u4h����ۿ� @�$Jx�R�@�7�Զ�a��Qg���i�����/(k�����.�
�М����"�jLM�y+���R�t������k<IO��Ls�&%<���y|^(�Q����&�T~���|�؜��i"h�}Ǆ*�C@G�_BKæ}-N�گ�;�u�G��A��X�<�T��|�>d��*6p��T�ȹD�I�d�e�K�T��U��Wu�D�l,���B9���sوK:�؊�J*�O�s7����Ju��Z�Ԏ�(�|C@%��:�6��B���dv�t�GG�i|�DSc�4���aL�F�rY���)�$��&S�n��J�M���g.n@6+����&����fp�oL�*�fK=����p��Г"qBd4w��/S�Gao�ۗ������,XnR��Z̫���'�À�J�����E����Ϙ�f� ����2����y%���6���}�qՅ�4�Ȁ�<�b�#~�[���{�8���ɔ�0>xr��Aq�R0�lx�-e���l��*3�A��h��	�N���"�m��(��@�)a Z�I�E	�4giv�Zd��T!?+�Պ3���~��Gt�@�0�g�L�O,���>�ρ��LhۖQ�'��vN��K�q,�<�,�ko�El�L���W��y���Þ��%E��;(�<I�J,���n�F����+a{���|j�zrmrD��2�N�F��L)��1PIv�Lq�Mn���F�����r6�,QcqQ�̍33�{���Dk�B���=�	�A�"ހ�NQj'u"2���8;�\/: ��3�>]7���Wk<����<���F鹌�\��)�]�]pt\���s���h������-Tڶ��2�*�S̆�œn,c�b���0$����`|8e�/`Mi�	���b���}Oy������.����Dj�gү/v�~|k>�J���3��������5	˨�#����'ðFY.tI�K�%�I "�|�B/$�O���d3��� th�c��إH�E�Ϻ����G��-�Us�#�~.d��$�~l�l�U�l;�h�Rf
�,�����<SƬ�<�9
�4����aV���.k3��a��ͣ��cM��P|�ha�i��c��H�u�t)��Em�e��9����&�]��	��0�Ģ� 0�Z0�I�[ya�%��^ˬs��|���^�m��t뽽k����u��!��SV�5�Ɍ'��-�n� ��@O;0,8�X�ҏ0�@�v�7��`��X�&����7�x1�l6jyLqE)�3v��X����	2�|�o����w�d���@��92�ϑ��;C��7{]�\�R�,�2m�ٔ�i���d�5�W�-�.\�v"����1*�-�|��hi�I[ʖ��q���-e3b�d�]�Y����^�]5yP��9�!�f���Z�qxv5l̖�˩�{��$�X)e�0u��h�c�T�g�kx�����5'B�ut�ل�Bi.�f��3�0�x�~�L��Bg����3����N��ؽP�5�`�=.T��[�����V�1�}Ɉ�x�xH�.3�X'����� ���3qܥ�g���Q��3�pe��j5��a�n��Q��l0b��c<�hJ�����P119�0-�Њ1�@�)E�<�^�n�� �BHK�@��^�Z��^�
��U��`�� J��dY��I(T��m6P]�Ȇ[�����D����{�{o�)���x�5��
�앥e�y�^q�LLm���8F�<�Trc6�y��|�R�`�%�&m,U��+1��ulh�O&8MC4j�����-*.|j����1�T	h$��\�C^Y�|�n�@5�%_�3,b��%yn`
ne6ؠ5�]�#⬃zu�$J������w�Y��D�y�z��َ3��7Z�[��,QhL�6��'4�)8~�Af1�D�'�b�0%L��Z٢��G;vL�©ST6\Z�_b;l�F'�P�M�������/��`+�<�omB��o�^�)�SGԷhh.kה��mf�w�d���&��E��rA��ܹ���l�t�6��<b̠YXSuT_��f�V�Q�Lc��l��|��D�_�[o��n��Jj,�ҩ�����h|�z�ߥk���B�`������C������Yr�G�s���^�5KhH�7S����6_����-lAT�1e�45�v{b{���}f�7�5_ͥfץj����<�t��sH�Zp2��Λl��?����`�P� ��`��<���Q�����{�6�ϒ�|����7��T�QI�F����(Ww��g�q̵�@G3҇؁�l[29�9a��}1�2��<!��������cM)qݰE�_-}�Λ�������������C�����y�)��_����$N��zQ�phk���!���]��i��OX�Uhzګ��C�m�↤�Z͚{�!��ra�[7���o�J	�e�@3d��?`ש�� �����kČ�i7ٖ�A�f�\~9;�
_�tͥ�i��Q�>r]�o��5X�|�[��~�ў�;�գ�������D����������ƅWY&@��.h��žx���{��c��J�=��>��^ܢ[�?�����&�n�sH���U�����*�z�l�(�ńv���ۼw}�.�PL���Y� U���:G��=�}�t�.Ϙ�n�6�����)z�\�h��"��a`�L�}f;	Ov)��]�	}>0�X{��^��إ�w�K?9��iХ;/���^��;�Х۷S�٠�F���B����t٥;�O>FnݣQ��p�Y���+ �[ ��	�OtB�N2U�G��f�Һ���,�B���E��t����ee�G�}�Nqi�K|�p�X�� 6��Y!��4�9�h�[h��$^����*Yt����GѳН� �>3Of�I��v��N�Ex��H�V�}6�ȣm۳�v]}9���<��z��'<�ڿ?��
�0�GF&���	���\�Ŏ�4��５�}���|�j�q��6-/u�R�����χ h�'�j�NG��Ç�О����k��z�*��9��<������׃i�Yc�a�������V�:y� �1�6פk���1��d9.�,ӣ��P��M�=�vѻ���'3��N3�I�M�a�%�*Y�6���:����Z��ڷ���Mz���t�n�׎͊V����})�������l�o�.�oJ��uh]���Ȳ�,���he�n��@�uG��r�)J�u���02z�)�!��GJ>�<���b{�\؈O�.|�hsW�������|����x�ң�N�r���֝�dM�k�n:v��z�Mm�	�g�T\�����v��ڽ4�PԣS՗^z��<���1R��_r����01XKU�5l��W���
5ﺑ�7O��Ӓ��X���b�x-���<6��.��=w���4=����<I�������sҿs���l��,�軙��V�Kʳ���@e��n5��;��_X:��d��NӁ���������Iw�����(��LϠ��H����J�rN�N[�z�<����]��H�S�tใ���^z� �^�x�8���ᕣt��b�%̪P�e�W�Ь�5i�M�Fڶ���~�H�O�Vd$���`l�5����y/X�J�58΢���V)�$�OQ��d��e���p�G8C�]IRt .�t��r���ߢ�g�k?�i�O^;��}JlA� �(dޝ�Ă0��e����饣'i�x�����ۧr6�e|A-ǖ�@��|�?&���_���1E��і�:ӡ��?�xH۷M�/|�=&>�|��v��>u:�Ʒ�E��v�v^��?��;₩�;or��\�rc�	E�X:�jʣ�1�i9�g9[R���f�H���0��i@g�dgO�ʏ	�|�}ˣ�J��{I<����nH�ئ�3stp�Is+<��%�Dbt��I�4{z���C�f�ߨ�����*�GSB4��[�xJ�?&���;X&YPK8�*%/��Y���������ki'��G��b	e!�S�|�wo/tCE��6�u�4(��tK�K,y����3S��G�� �+���"�Iy�c��b�M����F�V���7\�D���:�a�ƹ��E:��:���Y5n,R�c��O�]�Ց@=��c'$M����K�c|.�N� K��|�m�E:u�ua;im�ϭ��O�ϿQ�9��rE��G��F?y�y�g�����;���;���Y��X� ߷�5��R�갇^E��S<�\}ݏ�I*��AE��'�}�^_O3̵ [=s����9�H�BBy;�eN��<��/:H�ZԵyL�e�����b��RI��K)a'�'�k�X�>V��m�_6�A��!����v�V��C�*Ip�a(�@ ^2�ro��*m����c����~W�D%�+��6�nV�._�;������~���#���IS�� O����Y��2W�y����Q����|>�%���|��@���~"=U: 4��$���+� �T+[�T��e�8�+gt��Elk&a��g��J�:�.5x�F��Jĳi�)��Ⲯ.ς�r��|��)�����7��竮�j�a��J;"t�i�k(_���ILK�c1�Aa"����i�Ӊ6��aI�Sv�k'{�
������L��"F��u�N���N�ͳf*K9�w:�Ul�<���K���aZ@�!q6�pm9[���(;y�p�8~�m<x�y��l$^u=I��_R=Ycl�0�+#2v�S L��`c���Eoir�;�P�T>Xt��Ń'���,�ǯ~�*p��G���e�G�fԁ5M���ҋo����Y$B+��Y�*+ߌʘY	#(��y�R)���x,m�M�k����� ��?4�c!��GJX����d�:\�a4��8CKg�Q�]��=��#l'4�g�e֖;w_I�-�?���(k�3����1h0A���������<���!������Ck���T��d�!�}�[���k��YUG��Ck ����d��Z�%�T;��"~��Rf����ۚ�e<�`�B�g�lK��Ħ-[���|CkÓm�@�	���C$RYv�v���dehw0�8��1x?�[��i88_������Ζ�"#����ͩ���G�B3�@̒2�[��-2�p-6�{Iڷ�E���%�YH�:��Q��#d��H��KA(��Tv�W$��TǨ�.�d�$h��*���ͳ^Nqr��0-3$��Z+*5��ߙ���/�I[��G��^9#v l�
Sy��;2Pz�Y�>�K�g����'O�)�A&�?V]	1�a�N�|���8G&v�~ڒʊ�㖵g�А�۱�<�{u�fUpr!��p˹:��)5Hur7�B^h���եj�*ǂ*7 zL88g�x*\K��/����A�L�WV�#���6�i�k�]�Ax#��Q��Deny�]�m�n4�djR�'.���8x9'��~��7�=3O/����\��H�@r*aMF����g��a {%�2�qںY��x��0�'_:�S�T�x�0����M�A�4�Z�)��$��ۋm���=��I�Me�E.t��P�KHz9_���8Cp�"h6�ʚ-�6b3�[� VْP<�<��%�[)���*�ng@b��İt���|��^�K�,�j#���*�E�Y��V}�2Q�*o�ZzD��XT`�\�j�g{��3�A�O�a����K=K'X�|�G���M~m�
���q�㬏�b���ۅr\�2A�AY�@V��ס�@� R}�v�g���5�$��fjjRr6�M�+O�<A�VK4/4�����Єx�u�Vm-�j�hyyY��m��Y\�4X�6\Ncs���*#/�A��Ĕ[oe�4wƫ�t��2�`�nnq�Ǒ-Y*By��� �	-��B�h��B֊ru���k���G%�/N���Y�>V	p�b7�A�;j����	HG��"i��	�cg��N�"��K[��!�jP�IH�Y����ƚ���f۵$߆��Đ,:��ơ�d��5=Q�ڕ"ɕmÔ�)վF$�RR�Az����T(���t�J�4��zx�y��ϊR���e���֋�5f��������i��z"A}؉�T �1�c�tg ����p�&�졒�i�4���bib��<�x��y��$�֜%�.���x��Zy����Д��r��̏��F0[躽Α��qve{lsf�������$MOMP�V���%�n[ )�8蹤5A�uM�"m��^'�&/�i\(�G�J��\�L]w���8U�Ð�3ߋ�v��[�n���R���I����<I�L_;H[ln�̤��U�b�d�m�Ц8�R���y:����Б������@'QqK�[gu[�]��EhX��񀏙r�˾�Õ��1�W�ݎ�n�}:�@������!�4s�Dߚ�6��$�Ւ����ҩ�������� ��Hm�m��\PXh`�AhڐRr-q�`6���<A�"`-`�͍�w\�H|���[����A'���^�ˇe=K���5U��$�T����ѯ!8~��G����"k��|�'�vr�s�Z����`�fS�c�Y|?�W�}�1�����k{��n�� �z����i:����<xF�Q��2Q��v��Y#��Ĺ��9t�W��-L�Jg��_�A9f��W���X�r���Z��	;�|0_xr`GJ���\�r�D� 5���r��R;5b�THt+�M��� � <��<�۳�.ݵ���|�d"`��~�$�|�9q�5@E��Zh��f�ZRu.K���L��-M����KU�S9��K"�l�(��ulU�m����_0�?�2�`[����z��;;�Mӑ����2�J4�u!�>��1��Þm7���⁤�A�zJf ���K��gUK�W���>y�D�LA1�Q&��3g0+����|G���1P$p�tʹ�$���e$��jm۶���&��,�,�d���@%�Y��:��r����S����da�FK�옷��<jF�<`:�j L)X����.^Muá
�o�I0">�Hi3���K���sar��b�nE<�%7l���.��&�U�:����+���c'��zT�P���BP��0���7�^&�E�u��d�J�]�j�=�j�v���E7^}9��)����5t���=�4���I�,�aP$�GYf��x�M�&l+[2�;�&՘��ր�=R�B��NL_%o���@�ϼ�Z.SZ��~Ig���)5���h/���E�1SA޷����`E�L,�� R&CR�Rє�2:�D��%����u�� l/PA�?77�%��g�zO��ceZM�a���O{�u��A����|�o���s�@[�Y5۠�U��0L�
�2�H�Ce�S�Sl�So��M��,L%	nǝ�hA�κv���?(<�!��-�q}O��+MtyJgۗ��_�ؽt�5��2[%�;��+��=7҃����qj��xr_a`iV%����$v�2��ź���l!R��N����1u�ɇ�Y^����_��zݥl<��ى/X�U��S�[���z�}��vÏ_8��tE�(|�_���O�^75�ǐ3���n#�:E\,s��*5IG����昞� �ޚ����V��2K{�/�0M=[#��C,ې� E���8�)>�|��D�t�I &?�qz�<C �_�;_s�3���P˅�+WV����ct:S���ҒN�q|������A���&� >8e0�u�D]Xs�|�w���*��>\N�mFB��A�{�D	9F0��2,}����	֜w�=W����� e�Mi��OD���Y��/�E���J���vx��S�ƭ��GGh��R��D���|�=�����w���>�N4�6~֠S�tPe����w�g%�5�D7��K���I�Hv�t�O$�A�[��B	���G>�::3C��*��^�)�-��v���k�ŗQ7%鰽2O�w�r��U:r�5:~��ؕ|�Q��k3+ٱK4=��y|[|Y$��2C:�V�{y��S34xBI�k߹�h]�,��+h\�w�H��#�K���?�`�BCa"��v�3L+! >l0�$1�! �<��i9ޗ�Y�NL�~�)�gK�Q��<y�v��)���Ϟ��,�M��qԪu��1�<A�"�H��2Q�`
�E�Ӏ��S�8�n�J��
��=I��.�#G�е7_G�/��{�G2�_w���z���+�\j,�������i�a��Rc�e20}4�j�Ю��������׎�J���D+a����q��B+�#4#,2�d���Ve�v5�r����ao�����d3_�ƩD����F�L����Qry�SL�n������/�H~o�>���oF����{��P[�{v^B�y�A:y�C ve�;K�����7�E6�M�����_��,6��:�B��,��fgY<gW7ʃ�.���8ՓM�g�k�<�[��V����A��@��yn��xU�Y��+|�30��zM��@E��� ����	�0�/%^�Y5�hWx4��R�o�������D�kUd�_y�Utݍ7�iQ��2EǺ=��	�k�����ۮ�s���q���>L�>�Mn�����n��z��K��]�pM0~���4k��gf,����/�:����*1��O�%�N>�{�GW};�ґ���]���`D��J���oא�]g�c�_�n/�F���ma�����/Jf
�m1��*է.�_�1ߥ�ъ�v@
�ݻ�_F���Ͳ&�39N+'_�˯��n���C4Mz�;ү����mj��86��)IR���n!+��?T���{xBX��
UZMFV✁?[(�_�ɩm��m�-�I��P�u	�n/�V�Gn�N#�[hdr�8M�;qM�i��|z����Z�Dmh���r;L�rp����X;K�` �bl�S�^v���t�7�aAas�f��5��6M�g����s�
��PJ�*���Sb��J��U�$d��uf7]���<�D5Ϧ�{vҫ��DA�I۷]G#�*=��R?Y��������L[l���&�{��3$[9T�u�N�g�]�l��3��\gMZ�8G
Yɇdh��.Z�+c���+L�V�6�6�0� F+&�T`��j�z��Qk0�
A�^���]���}Օt�g�W^|�.��J:yzN�%�&��8Z\iH�� H�ȱ7�'i�%�t�tEe3.�]���혈�����)F��'b��D=	�#I�$�Lձ-46�Ե:!���Gh����&�r����-9����y@[�tP�S����J�:�S\_�۰=��"���  ��k@Y����b�.lG�>�ڹZޣ�u���xⰑR���'Lv���h�B�S�������ULg|�^y�E*1�.߻���7C�?�(����t��q����43{�>|�}ҥ��g���؂�鄤+��	K[�+%	��̮ʕ��$:E��!�Az�k�L7פ�%�H1W��LILFk$#���؉�t�U�R�Z�g �TM�Ypx���H�x/�yM]��*vُ�|�>ǔ2i7��@�8?���Z�62��t�~�W~�N�/�+��Z��|q��'��L]�p��)���F2{/Ϛ�d��Z=}�����E��V��}-/������Cg0��_��	�pl��Uf�j
�$���:�t5�}��uoK0X0�1ـ���b�|x@�S���`B^#@@�6˿�s�)"br۷o�����2X��� <���F%Y��Ύ���������}mz��Z
�ʗƵ�FF�����
Ę��z�ueSd׾K�뮥K�n�N�M�N���ôm�n:����1���Bq�؎(*v：#��Q#UO���nCrZ)6;L�+.�<����z�8gā��?��o`Ȁ���]�q4 ��f�j���׎��h�S��9�A����J�n��B �d08O���O�Q7��5腣3����hz�N�:� ��y��1������nݦ���U�ѩ��I嗅t)�z�e
�����uIZ2���,�|e�-L��J�;�CK���2�#�i1.�����=��hGe�^E��K���e�p%���Ά�
��DI΀�{"]�ď�}<��� x��P�ZEc� ��a��3�j����屦��Nm�Ӹ�ؔ `����66�~����y�V`g�&AI�˄�>���n�����|����bz��Gi���{������c�kϥ�̃��t�͒�2�����O>MG��^#3i�����Q���w�y�G'�W�1;:��:���[��d��?@%���%X?�\`F��Rtɍv��]�!�e�����K��Gj��J�	��Lx0,6��cU^���~����ߣ3�M��<���x{A�;A�!���Vap�Ȋ_lJ�\J����6/�gT�)f�$��}�N6�G4�B�5V���Mztݵ7�V5M�f���'���p�J�i���!P.-�L�~�v�ɗ�K�GF���|C���}�I��7� b�0\[�3(o�&2wt�Y0zЦ����'t(T3��0P��D0`����h%�/0 ���~���jw��,R}+���I ��q��ţ�l�t�nZ:�L�N�BέT�z�@M�b������Q�ɹE��ˬ]i���S�PutLF#=�mlhR$`�/�����>���F�wL�b�u��dט�w�a����!�*��%9_/UL�=��{/iC)����۲�,�3f�%i[g�}jD-z��?a�DtǍ�Ӗ�)���E��S���o=�|��p�R��:��Mi�f����C����-u�&%�[/�FD����:]{�^3���O
�n���n3��8�#�<B��_��y��I���@j�L�����|K��$���������;�Kc�u)�A+��)_����t��.�Y�xl3���s-�;TtH$/tM��K|�)�.Q߻�v���U��w��]���h���)o�?��uP=�\Zda.O��/�K���>�*u z�DJ{UQ�Ó���@Nm�$��k[�ȹ�hM8�v9�]h��XC
�% ���?��[���;&���C��4���ez���ӓ/f�ƶ.��V'\ct[����k�\.tF�Pl{�t����o#Y�Gd��"�����C�i��2��<�ใ�h�g6��H2�"��E������8wD(c��m*nb��/Wuv���K�i���#�73ף��|?�޲z�ڳ�2ih#)u�^Y��T�![f��A�8�3�'������Ę�ĵ� ��~�g���	�\��.�<�?����(�\x:�hb@�W�{��`��>���<�y!Z.��CF�|�>���f(qkl����L�W��,���/&����B`9�R��~w�fz�v��GV�1t�	�ْ?ɓ�?A_����3/���vҮ[)`0�]�^���OdN]��a�������t4}ߤ�`�R]�-0��ӳF!x[=�NI#����g__�72ѝ�R�DN�N��IA"��ԥ=(�ɼLR��}6d!����@��ЬP�C)����z�⳯��~�**�*fYhs:��/�s��S��e����|�����N�C$�k߲*�|M�n�-1���lj5W4}C����.½�e�I�|Nq﷧�����&0 8�K�IG�΁�g����fݺ����jۅOe~M������?vT�ˢ1f,c����o�`��D+�B��N�ѭ��F$nx�����I��QV�Hb�%ݱ:H�gJE�<�ʺ(V%��3�s(�$�~¿{��L�	߳kK�!�d���,5��T���!N;4POw�2Qry[��𔭓��N��v�g�*��G+��.��r�4�P�f#��B	.K�g����]�A�+ P�SW:�������.6E��A��!���b�Hĝc��cd6 t�G�F(��`���lWl����V�U�݂8H��P�z�&	}��������c��0�-M��r��8��$�HeM�6�R��i�<Ԑk��;���{�~�1� u�g��ΊY���8��9v�8��,�����hB#�1r�'}j�!��`[?�X�Q���!C�Ʉ�;�I�i*Xۨ��=֔6���B�5ͪ������0�q*��f�AH<7[���(Љr XF�7��(z��%�N�V��"���������wm?�?����B���#8D�mt���{�?!.@*��z�$�ڰ� ��vV%mD��9|re��d�LM]���uE�ܵ�>���J+�(ʝٌ��m7��0��L۩�ŝ4�����k|"+��$
H�r}q�XD�f^�����x��\w a��Yr2p&q������yh`���N��Jv�]��.�@ɓ�򁲙��\�4`8<�T*�!/ʦ�&�BS]	�_B�9���b�e����ŵG6��V'�����E���2�I��y��+�|�0S)Ñ�]ԑ�i�Gh���}�ƴU�Hi�A�v���QQf2=:I�g��(3�Vi�D�[�I!a7�#Za�3u���e���2�ݿ�j 8��&�\�*���b�y[�̪�#��hK�֛o���d^�o��$Q}M��Wco�t��$��du�����_\��Q�ё.�yӥ��z:��e���j����ox.�-Җ ��hWIDϊ/��K?u+��r ��` �$߯"gׁV���o+�<��/8BXV8��R��l)4e��v�!6v�ԎI�v<��o���]e�����I�i�����p��8����C��Q��$x��(�����Pe�#���5�!�#�t`F���K���{q���._�S:&i-O~y���yVD�
_�哄�Z{�G��}W�.PL}�N�-Q�S}|�V���!�l��9��?�٬�"�� U�X�ڞ-}V^�����.�.Ӌ2.<���=�����1u��c��yJL5���Ƒҵ��~��5W��}i%��ϒ�mp�6�m�V%�6փm}�z�)~�m�I{�'���I���t�n ��tƅ��kS(�^TE����$ؓy8�,! ���Ӛ��e���kf�Ia�k�(M�$xSj����2�Մ�Em�+ѥ9�I�72EK�%���T�w�PV�.��O&��"8Kk)F��L=��%�$�gH�H�Y z�$�-�XK�Dln�a�M�l�]w镴u˄8��ϝ����M.ۓ*q�@�7���}��n��k�V��2P-���Nr�^�`�SB�O~��t�uW�����1�G���ˇ����q��+uI@��=�R#sq�<{g�ϲ��h�*+I�L�謒Rv�P������ݤCS[���������:u���^L}ʚ��Fy�hO��j�<�:?H��g���-@k�u�{[�x H�8 &��4�-����3ŅZfݸ�$[f6���ry�_�-��|���4?'I
���kh�\����lf���5{|���6M�ԅ~G�O�ȥo
K�	���-�����85����֪�Z\����2�ZG�>����p{������뼮��/���9$� �(��$J�e�R+̸��^3�C��G�?�Z��=�m�$�DKI�b� AD"犨�r~w�>�=��*�dQ�.WU/�����}�	Hh��EQ�]|����?�sl�PT�Q�n.Vqiv�|����'�g'$c:�p^�*o����֣k�����7OC�M3���M������7�B���^����1�}0��^������9WQ.f��պR�kS��c�Q@K�Ly�!(�����B�+�q0gH�;��e#����{�|��� �*���0;=�_����g�igs�b�A,�`�uF��Cl�k�2������k�d	�4��D�aI�3[o�AWA4��̴�8T�B^O(?�B833��v�d}Va��������=������r�� �
_Cb\�G���ڰ����}[i��q\k���G�p}v		�!��NE���Vk�n�qE���H�eS4��k�dI粨�]���kj��s��o��X?,��.�j�_#{Q��HqD'<�9{��x�!�SO��no�eA��=s/Wh����s���{�#(��>r�[�$7�m&�-~��F\��8���{A��6Z�eD���"(ʥ��[rټx��V�X���ou��<V��Sz���1ij~6;�lѣ��,�7/��K������mf����˒#����m뼜d������2 <���q�F]���i��T�=���Z�c#�����DC�����7��J���;V
�ʃg��h�h,�Q!���E�3�w=,V�"@mp�QV����b�ϩ"��תb8�G/����X��kG�rv��"���V:h4C,o����E|��O���Q,ެ)���,`��D�:�j�ߴ�{�+�~�'X�_�Ǧ�[C�Q�\�]?V��|�#J(�0}�!q��|�~l�:?��h����z��b��!�8J����}x'�th 9�wmߊGy#������8��#/lTާ;�5�p��)lھo��6���c���G�d�d^�3*=����x��.3�0K���P������k�r��U�h��i�X��j(��\��A���p��5�U����3��.Z,kb5+�Y�^',j[�<J\�p��Z��:Ǚ��APu4�k�����u�|7��������o~\�'o\�GW��v�"Og
����<'��)1lQ��EU�����$~�ʿ���"�q�����:����J�������5���z�ѧ�w�LߜB&��:��������˪T�8�o�۳GKK:K��+�?�2p�:�IxR����G�ĨIĶ��X��woW��L���8|���$��:>�&�P��1.�И������X�fc��|�M�b�T�#m��(j��h_�x;w>�b6%B�Ş�[�v�VT����d�;������Y��0""�AMύG�֋�%���`���9�.{�L�Y����76ܔ�v��t �ՙ�QP�uŰ�v�=�C�Һ�m�73-���2
&(�|��a�G���;���v�Qm�%%½Ck'��)�?�
���(��2M�Q�l���~	fE���{vno��2�~�i��/�[�lƿ��ݸtA,S�����p��yǰMܫX�u�c���+!p�Y[�f\�Yzں5"�H~ֽ;w�ر�|�l)G������Z��FUOa������y�r���甗��7>_!�d�T]q#(�l�eb�Y"NZ�"$Q^��8p���l����9��Ŝ�M�J2Yrb\�p���,f���_+�_]'� ����$ω+â. �I�T�Q.0��v�{,��¤	������aT��t_D}�VL�ǂ��6>�Q����1p�,	:�}Az_�T]W`�ׄ�^"]z���H��a�n�ɚ�C��JKjm?<�w�
�t�4�rs����l�+�K)��1�xlE��IB�5�7�+���o���3�q����ʳ��=����SW��T��Y�"+�2�'1$.)�Fő!,�����

^.�B��9��zG�i�ZS'L���@Ga���Ǧ�������$(U�ܰ��iٷ�JCi��Ar_v���&�]�i^�Ù�ɏ��\������ �3��h���/��"�u2�T�߰o�����oazfIݎ�n��r��26��hL5��U���!4CC��`��,�f�[��Sy���N�&�_���f�n�&t��u{!��Gc�B���R�]֑��S���(���Ԕ�CDJpz�Z�y�Ifus��6�kذo�v��Z�8��F��I;����~���(�H�ؼy3������L��%��I���۽G���ܾ5��]��?�c
/\�/�(�%�6���2�<�T໲=μ�=;:��L�Ǒn^�ё(�>�h����g�����czC;��+�,7����]؋;�������7���U�z��;q��o�i�\��g�冱m���7/��'W���*5�>f�֬_��"`��NU�կ�����ܕ�t�6e�6�Y�'܇a���'�h~��Z�8i���ԗ��Q4������'+@�����e+QDS��
��n�0+��\E�]@����؛���޶�۷k�KEԠ �.$O�����˗��%b���.,��[����%q��E�_����Zr�d���k1��?��q�1T����}�0�%��7�ǭrCk��l�����%�l�*U��q����/`~����ỄS��h�覜gI�0�+�U�h7����c���0!��Ѫ� ֭�7іk���y"����9��pE�J�+!H��=$��[nޏ�����}!�R>�t��V[�8q�q=q��Ñ��D;/ꠎ5�D��#s�؆�87]���>�՛�H��kV��g�]��+��X�M��P�/~�k-���]����Dp€ʯ��Rɼc��oI ��'+b��!FbM�]���!�A*u�me7@<�;�\]�7�}�=gBg�X�a�Lʄ��k�֨�Z��1]M�MW�3��JZAg�z�b0�E��.>��(�z�vL���ҍ�BV��F�+s-�M���c��}�zC�le4fOJ(Бj�Tb�l[[���.�Ө���h���a��(kb-I���rsJ��
v���g��������� [Ƞ�4��*�"[>^|�\�rS�(N�[�WG����$Rb˘?������G���5Y����w�pO�/�n]�~ŴJ�sW�ߟ	�~t#��X"g<7
�Ң�K͎�U��m4��.1s=Nt���788����o<Ȗ]<{g'�K�P���q`�V���Q+���~l9gvt���
/^�ս�2��: r���!C�H�VpEl����X5�~����13Gύ�Y�N�7&�Q������D��v^&p6�'"ʄ	���q
�gT)�����&V]I�����	\�rE�"���Cwd2wch�V=t�$��F'���ÖD��3G����ISb�k�}Oa�L�qY8�&ϖ�^?���Hrx��G�n�xI_��x^�*��ko���>�J+�u�VgIc\�G2��ϲ�����|:��h��;�����i,��oq��Y�ٱM�K^C/^����?���:�te�������J$�E��WR!$�k�np�=��Q����^q���9�J]�H�%D���tV6�hz�p�EQ������Y�A����V�p=o�$�{�H�4n>sUy%� uo�tW�^^���,!�(-���xS��`��]Br"{���̐�\C��)�jk'V#x �k�{ʶ/�
�C��XL׿Wzt�`# ���x��ڂNW�U��^�<�/����&xJ����\O6)*��_��7x�����Ѽ��_ZĻGO��d�������BF /�R���{��)n��O�yD3E���Xi�Xq�2C�Qi��ob�ڋ���6�dA>Qܲp���~ �u \�A���ӎ�Oa}O��xG�-�%��<�$�[r9�'��7���<O-�B�d��SD�x��T_D%��!��Y�e�e<�V�x��g�� ���9��E[u���ԤNw9��,�	�<h�(,ti���(+'�lW�wQ��ҁ�%���U�a<��CM��}g�,�Jj/?�����&���}�P"�Z�:j�4��N�y�[�Aa�Ʉ�z��5#�kROg�{���.�[��q��<R>ף��Sjɿ�q�3E��)Rr��f���s�?��J�X�����}�1"	�^r��G\���bCL�Ccm6Wq�3M���ZGPD#��'�Hr�'5he,���m�Lߊ�Ӎ�G`Q�@xnE��h�B�u6�=.�ѭ%P�ˋ#�����	��l#2��������a����G���=���)'�(���>������� �"g]�j�z&������f�e2+�����	,>t%/lP�����;(|��(����^���}�j�:�H���㶵��Y��Q�+��Ik���ֺ}GR���A�]Rε���ĸj��n|�u�Ow\�o3���dFY�	�Φ���:1���t3��IZuc:C��ktmO�la�XN'�қ�3��sͶi�YhSY�\�駣��}���M�� M@`k���`4�c���nxl�h��21��s��:n�!�wF�9S�.C".��A2����Hw��ٱ��Bw���T��\#���۽����*w�s�<���y�ڂ�Ʌ��mĕ��AI$��m��a7)c&���2��I�"��q������N����c��nrl5Í�X��L�j��3�D�|1ה�j�]�R��xfUym</����0ƽ;~�j6��{87���]׷)����,�˷$ncg a}���P�Si�ؽ@�N��'��x>���]��n�LRyv�M��mB�R����g'-��}�v.nך��a�e6F�$^�u��2�cUB�Pkl�r;u`� ��3ͨ [N�ds�$�-�*:W��2;�{�(L�s!R�F��x*h�����]~\�ݔ�n�=���r0\�IM��ulٸ	���#'N���-�q��iW+�ݸ�X�kh]���5��4d �y)��ϥ���8�I>n�@��zŝ��x�j`&�]�Z>�4*|�L�K��-ڜ�c@4��c.�@GF�w��j�8
���T�rRj:�¶͛�a��cY4�CXJ��L��Fh�]"��r�S6Wp�7�=wN�d\C�L'>�(�S�H^��`��괈	�"˒F�����heSrOޓ�$4���T��N�:�?]P��D
��ym8n���h,Z�biZ�*RI�L�׊���#�Әi�5`�+nY��\4g��`>�N���x��u�0wj$ܴ�:N�%����O��cӎx���H��9"7}v�&��f0==��B�\���9�H1G��HL�qW4&TL���L
�+�׃�'����e�9�b���1�hʊ̱[��r��Mߡ��-ߛ/�&,W�w�s	�eVv���p3��1ϔB�u4)��c�RG��ou�e[ 
p���q�Ωy*l���ǚ�V�ܵ_��7E�������>^x�j5��!!PW�y*�X��D��;���J:>�od�b�����Ѫk���t�~���}b	�U/�X ���a?�l���(���GFQ���L�ͫ�>g��ө�~��g]~`t�"��s��D�gd!<����{vm�S�?���6ia�/Bsuj�9�c'>���l�!�j_5W[�MbDY$�
8�J51S��7�-�Y����#G�=#BE�H�P17������سnL��tJ��h5+.����mdI� �D���gf�h�_����;c� -���,
D���%ea�,�	��ǝ��
�ghG�˺,u���e�hQ����b��q�E�P�FV��O-L��dS�����*��r��B������e��(w�J��N)�q_�	1d7BmQ?'�iM�ID���Ǝ����;�o��IlN:���:�\��7����Ye��D��դ�Nf�xﰗ�E�WPJ ��&*�2
Ve,��C��S����[1�p]]�X�6m��mؿq~�o/kU*?*7��4:��@������#J�1$9Od�u��h�<�u���\$�����J���8u�x���l�<J��A3g4&���Gc�ґ[��n�X*KFpcr���L �):xC,:c����0~����ڎh����ve�
C�غ"�^4�2�������+b%��fJ�N`�/|(����tٔ��YiQ�%qO���ss�ʵH��B>C᪡ߨbH6W�4���YbHg<�e}��Z�c'��ܖ1Q��Z3+�t�$�f!�ElZ;��������(�$�'ҷ����"܄u������
&g�4;�p�t��=�^~
2��;V�{�/�ibC�]di9��,��Mk�����c`/Ӯ��P-e�b�� uhn-,��W�A�$�	6vl��Ky�,E�&����)������o���E⡖g�q?행,P#H�#�z������~�mD�"Z�7��Z�\欧�xlߵ2]o����k��4Ƅ�qñeV��NE���Ν�A�V"b��n��+���h,�oky�n�ϸ�s����o-��ʋ�!V���=Y�I\� 3��FE��\/���EyqJT:W��ɖd�^�ס�=u��H0���o�m|��mH�-��f��(�x�+K|�zj�(��ߟ=�{��C��#�ְw�H��c���~,���d��3wt�ɤT��cT6Γ�;���d�6���>)� �JP+n�zqӞ~��;z�5�њ(�;x��N<��Ӹv�*�y��ٻ{wm�嫗pczx�lř����[o9�N�i�0��W�%�M��s'bѢ4rF�s�c���Q
��࿖�0A�m���,'�m���aF�Đ Q�W4��{��_	��1�Y=�h�3��R�<���,_T��ߐ�(��?�N�&�0��RyP8;\�%)�۸�7�{6E
�
�l�"v�����1u�<���^x�wؿkؿ�$x��W�^��Ï?��/��7ߒXXV~�"tO<� ��݂�����;h�B?`ld�X[qI�cx��n���\w��p%�&��k���/��< ���y��,[c��ܲyN�iV�����[5xD��%�ө��7�cB,��P�ōK ��G��OD �k���~H�n^���7g�s�n�i\�vEyOH��دb&���x:���#عfH�]�ͪ�5a����r���?�on��L7��j#�lJ����,?��fD��a��������~�s�c(���)S��wBԨ���83J�g��f*�3�8n1��}vw���LZ� �a߭��T۶mC��É��h��Ts���׾��:�d=�&���b�Xs������"�~���!��_y�A\�yE�q;.]��d�yq����޺㜊%�^�]�M�B�U�$Z����"�m��;7���J�a�6ɠ*��f�{�^� �E�)�gb�9�An�X�������&gxsri�Y;��Hn��5(b��8�s3�6��ѯ-�ˏ���4N|�Z�%|�/�X���W��dhtT;���JyZNP~Ɏ�y�A΋�\��R��Ejn}��WpG6p߭�esܸ	I�㦘�����Fd�q,���Z0��g�>�3�)|��5E�ŀv�!�_^��%~8�8�[ìdp���B�aV3Z��X�,���<��Z�?.���<�6���<@!��Ȏ����hl?=wK�y�IܞϥuF���5\��T%~k�~���������g�xD���(ԟ��������g�ں�/�C*&��w�v(��-�����Vb��SZ�^���z�>F��̐4�Ў�ÿW1]T�u��S3z��R�����Lj�䚆��>�p,̜3��l����C�S���LJ3���}"��q6���>�����p��Y-��s���,�{A�C�D��[w�t��WO��. K��VS7��¸��=���Bi4u�n^�!P�0/se-˩��K�y� �l?@��񋷼���*E[���=D��l`#���-�.�c��-k7�a�o�
7E�?ʳ�t,�q&Fm�:�1ʕ:�#��!�cXlŐ�ǐ�Ɍ��;�C�Fnڼ�%�H�)(����������QÐ�(�o뛘�ÉO�:H�\^>���✬�Y��N��ҕX�\!�	A���]D\�U[/�l�=G�4&Gd��W�ū����{��'9��qX�3���Y��A��bV�~O�R�"���.jF�K9"�X?�k��8w�:�(��܋��!�۽���>9;��;��щ�J@�؀L�q���Ď�n]���ɛ8w�d=q9��tD��4Eo�jI&p*��lޝP�M$(ع��p�07���2,k��F���@��-���f��g��<~��-Ȃ�桃 o����de+��3yڟ75ƭ<7Z�;�1ݶ"υ��1��<f����$�'g�I��要�-����úv���;���/kFz���#Y��Y�{�b��-�_��ܥ�x�w/����/}o�<+�]�nR���w����{R�٭�ʏ�կ)��%��Ra����7ú��κ����'��Y���Z�~�Hiqñ�(B�ya��l�#",�ʂ.�����:V�X�X��K���g��7]a�FK�Ҙ6/�'��o^T�0�����%�V���(�꼫�4"[H6�Ү��"�r#S�e�1�u�!&<�F$�0�Z������8�Od?7��yD�Q��.�	I%��Xi�E,�Y�o�;MpC��~?�]tPdt�͆c��>Ǯ�@�|�nn���	�0����.*����v��2,�q�C��=�����ݠ"D._���v�W��ˈ5k���{�%��[\��~��ofz�ꝺt�W�F�S��J7�S"����ǧ��C�d��u_���XL�i4%$*����{���q�������y=:R�s��G,�S�ʱzK��V0�U��B�ku7����Y<��o �*vo��W��1ͭG�������o�8*�f]"ϵ�ƒQ>UԹ�,E�.����6抜���R ]�x����؝L���k�C&b/�b,�
V�ɾ��`$��M��MR0@���V�8�utmA�s�x(��s��(�s�@x������)�l||L_��qM��&����\H��[Ik�½�w�hBe���w��WZ:;Xlfm��G;FD���ry�4�{�P���\z<�=���B[�m��^#�s����"�i�����z�t�9Z4�(��V}?���HgSؿg��3S��-�����}��I����F�4��J\�#k�N�
P6��1��t��8���2P�m����ډ�z��X��+O<��;v"��kAojNb���������|��u�2͞�q�i���wV5$�XB��*�I�xn�ڏ�T4�Tڡb�#��}smMUS�g%^d�5��,��w�n6&�����W*˭P���znh�,W:�β�jxΰXȨ�s@�݂YH]���VƪV�l�9�U��v���_�i�L�-��)+��6����e���$~:�pXK�(䄦��͞f�[}7"�3��q*;v��� �-[A[O-��e��Q�L�.��gp��4��O����<x�^	u��Jl7W����Ŀ���*觇P�I����j�΁��6���^��`��FW,[ ����r]�乷�\��k�X;�Fܽ��j��~K⾶�����\{_CRY�"��ML������G�J��ϙ��Jh���t۶�B.�A.�Ҭ����+N���n𼵻���q�޵Rx�J�=����9jp�L�1�BbTy��r�	��H�ظ�I��5�⺩��abǒ3</��X��~�30�eZ"�N�i�:F�NTHJ?��n�Q~��ёq4�*�J�5*\�.���8[_Z9�ֵ=�9��3'8�@xqI˒�����
0	¹�}�Ɉ��˙*������g�c8��扵 3��B�Z],��,[$�]삸�:���S~�s`x���_��8V�^����nv�۶�'�G�|f�Ь�E�n�9ilR%�9?���	�
xa��,�q�0!�4�@؞#ޡ[�u�1��L�D�� DD&$���?��w��� �b�������Y�Z\�s���j���,�`1YԽ�a�dI�N�n{��u��kx�%��nB��F��j����~F�b���=tGGj�1�>���>���zD7C��W
�&�Ҍ!q��h�w�KH�ҭŇ0�����P��5�uk+���&!|�L浜@��R+�4}MJ�28[9.[FC���R����Sʌ�,��ĵy9�4<�le1�|F9z����h��8I�������^Y����R/-�1��%�M��~R�/~�X���a���sI�X�'��ν��阪~\�AJ���%nDZ��|�2qWWQ6)dy��ҕ���43��/X*�Q�Ɇ��5�빸%�et5v���i��o+��������Jf��00���u$1��Ab$�=�؊�l4o��l��q��;�dh�L�X�ZgW�w�,w���0&O��d�"@���y��õZq�+��3�{d/d�I.T�=E���ql�Z���+��:|��un�5�ﻹs�hu�5qB:�+m	I�:���9��)K�4��u���6�:jKq��*$!��EQ��{��o�֦چ�6�m���x�!ʚ�m\�������U���a��rYt4��Y`:R.���u��(�	v�%�*꿧�~��F]�����:~W�\:q��+3_��R��2i��.t
M]��M���|�����@u	�܀|�Ca_w�.Q�ܸMs�o�{��9�l��ʁ�e��N�Ng��h��@��*H�d%���i�`R��o�i�T��g�M���{����/&d�t�Z1���"���J,�\�MQ�s�X���)$���_�e�������/�K�WC60��T���U+��6z5�nn�aG��M�N���
c6Ӌ��)�Zl%�Ǭ��r�K�������a�������&�ܱ{1�G3)=���=�Z��,z^[�.~��c�,<_����9rR�&o�wY;Μ�{.� Su���kc�Y��\P�L������.*�	�%~L�.B�'b���8�	��7n�a����5�Q�@���N;������C���V0憦;�^O�"��0�ZNN���;�
�Үn�hO���\0��|78_gc^�����	�Sk����\Z�UQ�BS\6k��Vgb[�����XCT�v�oF�&�'ݰ�Ė�^������+K���~q�7�+s5C��O8^�f��}˺��vԝ���w�ɫ��F�-VETE!0Jg�kK������+_��r�H��h"�)Iqyf^����JՒ��,(J��E��Q�!Vm�V���C$�A�&R|W5te
���9���Oc�&#���#��{eA<�/ߜ��sWq��emB�X�,��%�4�R|'9*�F�,7}|ֻ�r�:GG�݃ے��[m��c�tr������,��W��,�s�g�H+F������T*�g	,������(/K��A������t~<\�c�Y��v��;�>f2Z7,�	���\?ş�[a�id��O��[�Q�X�~����%�	a{mq������_N䥐J��ih�V��6��QHڝNx�(�4�fL���6��Mz����i�/��}��ȡ���k3�x��)�8wM�gQ'@uu�A\�+��T�7��ޣ&�XYłL��Ǵ��UsSسe3����������t�)�:���\�����S�$�fP���9���`G�&�R[*(ZS�F�I6�����؀I�ʒ�/��
_V>b��lں>t��܃�X8�FA>p-�����gR���X*ګf�~��M��:�^�M�0�ΐ-<Vn�h�2���6p��-�u�i�d���"�͆�eV�t��-�̟uD=j�"�37<���Vp��jؿǯ,��bC��(���k��ڎp(���8CJ��X�a��IAa��X��snzC�����ɵI��K��������_�pN@��8QP���KG�/�������REλ��+�>:��覘�;�$��ҥ}�P�^0���l1�L!���s��c�ѭ�6��4N��uOe��a���-�OGO_�
X��.��x�tl��!�N]#� ��L��3�5R֩.,t&8�`dT|�2겑w�[�g?�l��1qoo5+�b#��wꪾ�#���L��=u�bJ�?����f#l!�p����V�21���J۲�_̷N��f։2���`�q�eW4Z>-a9=5��' �"����Eq��wD�&Q��:�@'Xwm��od{a���x��y\��s�=�+��3�TaI̵tkA��Ƨ���>��sc�*�Z�^1��9.���|���7�Ÿ�����і�������0��?<���«�j���Z<?�.p��=CJ��c��� {�hԘ�Ȓ�L�qF����=[��}(Oc�HQi�c�[�TmbǺx�у8~���S����7gw��1���t��ځ�QGNs��y�ڶ	��>�˗.ai~��߫٩Sg��<�T\6'�i��3�?D���4+�!�1�����2Kg�{l�԰��O�w+�P�@X�+Z���o�$bg���F
ktxэ���}v�y�"8�9�����&�𳢊�Z}o2��"��|��nM��?e+�5��0�%�b=vi׵����Q�{{��94�o��b�������j�S�,1ޮ��D��ڵk�����a׬߀�7n(����[�ar�&����E0ؽ��Ƴ��W�����B>�BN�j�z��m·��.^��+�.��rM�\���J�Ǫ,�=V��Ը�� 0������6P���رYf��K�]☾vQ��s�
b���Ø_����۱s�f|p�#�]�u����oS��_��J���k�8qZ��|�i��3vcj�&�o܄-;v㵷�����/0�~�����1�{��}���b�gǘ&/V�_����hv.:�����QBY�5e�s�SЩ�m�.t |�B>������/�(	����n�	�%_�s��F	�T�M�-���D�k'�Audk�A��,U��1B���M�w��yTZr��<�߄ܦ�ȮقY�<a"��+�����7����'X���ǿ�u<��38�F�ݳo�fH��|����XEN��#��!���8���2�ߚ�Q�X,����z,��o�(�oY��k�%j+~�K��U;�'��ʩ=�Uzn>1�Y�RD��9oLn�X1+��h9�t��[j��Ž��Q]��0�$r��qeM&Relb*s�:5�7?��X�1|��'�������a����E{������_�[��:��ԃx烣X��?��{^nRcIrg���Vkh���u��l�0�"Z��J릿��MТ��Y1
U������1s%s�Ϡ�Gd��
�z
��Ӆ�]�
�5k���GPQ)_L ��`���ϧ�)L�b�]S��VRA��~^�`eTt����=�T�Z��<BR�SIk	E\f�9u��t�R���d�S]S��]Q7/���%��e�����܇/?~�������'(���}حְ~������'.vJּ[C�2��o�lN�'4�s k2qbŋ��eL��x�܌{ILdx���j�a��D��L�B`rc�H@���<��FG�������A6�,��!2˅�9�P�����Iɭ�c�h����ƞ1=?�d��H>%.fC���C�w(����v�v[�f�.� ���oO\$B�+�,�A΍n�q�u-�$u�S�X��<(���&|l�'�E(@Ƙ+gd1 ך��̈́��ۊ���"ݹ�~9L|��劖(��}eM��	��wSK��0��NB��Y]�u��ΤեfS2nr�+^�>�~�W��ē=�nbD�����ћ���ؖ�hV\�|�s0�J٨7�ͥ�L���œ�(�E�M<+�fJ֣��!��k� ΋�w����d��e�x�©��NP�	�;+����iM��@�0��R5,�j��w���t�/����ǖ-[����Ӛ@�����ɩ�������nB�j���9+h=��:�[��v�¶m�5�Z^_�¹8J��	���=�ʁ?�ٖ��hH~cl�q{?�<�7ج��nnf㬧ι��0��ϡ`Ń�� f��	_˄
_cTZ���a}���&hF�|Ye�Q�fS��t���D �)�t��0]�=$���kٹg���|�%�cǎ�ȑ#�힞���˗u���Ç�L��i�^��իׁ�;�EӞ��(�X1�c��P_�87�s�U�9�jZ�{��~��U�t1?�%x�Bō���nN���'އ�k�P�wr|�R��94�5��=n�8yBgI�X������{G1���о�Ŋ�F��?�	��<�^����l�"�m�:J�ؾs�"� Ap[\�&���JO�Y����ĵ�~[�-z}�����`�GyC�	�	5��3ĈYC�xfm�i�6�[X]��uZ	��{i]�|7��)Z:siM�L@������(�:g�r�œ�nd��Έ?�p瞐0�\yWr"2)�JXZJ(���/�vk��h��_{Ǐ��OK�ƹ�7&�pmjε�g-�[�d���;�7ݏ]��C���ŭ_��J:qc�E||�N_���2ɴ�mT�w�!��wO:ǣ�A�9L�)&�.]W,۩�W��w?��� ֏��޸6�ф����w]�2�w�~�J�	?]ԛBA<E\
�i�K+a�\AM�5�)�2_�����#x��s��1�X���Z��_�u�܈��w�c���ĉr�]�̒���G,+�[�Md��@�a���ϱ,#ZX�Ӵ#l�I$C��eZ60���A
��)�}T!�M�nnCF���8��,/�#���wxMZJ��Q���Þ[	*������y}���i�Flٹ])�xeq��D�0-^����]΃��<5�kӳ
���Z�)���񜲌�,2��c�TF)���L�F09��_��6���������1����a^(�ޘǅ�^��<./T�e��ҕ��=�a���ah������ҽ$4���j�����(]���^|�(�*e|�ч�s��֡Ԩ�pTp������p��h�̈j\"�9-%�ʁ���и\<��L(4�w��HO^���zy��%����:q��6q���$E�o،gڃ��Cr�d�����X�����|�7�6��)h�Ԗ��a��	|��F�.Z�#Z��R��F�6�u)�4�,��9��`�`x���X0w�(���ː+����:�e�e���Yǝp���PBGX���0��g�h$
�����ӗP�p�C-d�>�^_�8tʮ����>+����)2E�V��jQ>��ζ`����T&��?:�D�_{��ٱA��nm�b���_�q�}rU��Dʴ�t����a(����t�����,S�)(�`d9���
}�k�5̿�1>�pF�0!?���U�.�gjI�5�6���8^<�K��)�
�NY!d}��;z,^��yv�Vf?!c��
f[�R��Mb�hC�t8�ެ�J��;����u���-�[ˎ�ܑ^����;5�������A6��b?ÄZ��v����ٌK,�@�^�G�Z�2��]y~��A�̱fGI�$
+��z[��ʵ�"O���u����y���YYy^,��U�P$�b|F�l��a��g�T�Պ�>�V:!��n�,`��	Ӿ�q��G�b��������h|w8Q�e��qwq(�c��qϝY���k��M�~�f��8Cw�ߏ/M�bbJ3VJR��Ě��&�h��Pi~���Z<�W��_��!�
SF)���6��C���>���e���5��5:�����ݵ�ŭ���D:�9(�i�O���q#�0Y��ì�k���h�h��fAV�:��(�2�D�C�0�~����%�rqk4ƌ&]���X�f���h�;P X������:s�øL������gq'��8~�.Ί ĳ
r��UE�$�e��,#b��`��k����J#�{�ΕQ`@;���lt�'p��<.M� ��
$��9�;��+̬'�l��<��uB�M�����j�. �{a���֞\���;�������գ���o�t��*my���V�5EuU�CW�Tj*���0��E�$Z]$�ӯ����5J���Tɔ,RS�jW1a��4�*�� �Q����ǂ���ܰܬ��i�@��3��DG��8K��b�����Fٗl�+���j�w3��h�ȱ���G&4Q��	�^Բժ˄.����. ����{��wF�7�*M�7q�6gr���4���ƍ��u$���fҫ;���7d3���1[.�1���3�)ػ�L%QO�¨��4��%���	��igK_�0'V6)��#8�����S ��Mk����ez!������� � �>3���%�u���9�]��8��7�4~��R���yts�}���m�5u����g�#_� �H~b�e-B�D��b���
m��`n��`���-�N� ������b��l�mnhKr�p��΄�h�(č`�$?��+If2��)B�5�/Jo��h�1J4��2
[0F�bNsy�w��Vs|��|?R^�/���<������츁������-^E���V�v��8�ƈ��]�}0:�V�rD�����)�]U$I�{���|nBb�J��?�Ԧg�2,0O�ݤ*�X�ۺ�)n[�c�����۬�,ǔ�\]"NR'f������'2z����1�r�y��A�Hߵ8�Vߥ�e����2�R�u6�g�q�iH��qv��x
��mA�5c�$v�8`/ս�,��`��\[��p��	�x�����dS�N�97f7I,�ZP��Y�M�K*p56�&��l(�޹���T�M��=�z�[���~����^�zv8w��q��]�^R�����T�h�O�é�ɴ��h�y���r�nGx�B�V�
��`RA��Ҳ�9KRqE)<r�n$�-ᓩ9�G~V�5s�p�L�W1��:�S�/)J\���R6���z�SZ�㜵���)����)�U7����2���%I�nU�n�Q��Rh4�:ƭ��+Ҳw�X%���\�A���`m1լ�SXڵ%��01��[ί*ϳ�����H �'U+(�݆��H��h����o^g�qXt�:� H��3{�_eCw/-n�ډ5�w��P�Q"�Z�q+
���K]-H�S�
�Dt
-M��Ŭ�u�|���2��D�m�!3�oC������t�J�0��}�YR�=���Y2C��9�S�T�r�e3�"�}��m�<�j��*k���a��<t?�O���ݜ��o�T^	��W�\A[�������U�U�k�d�5�ڲ��Fy�D�P0۵
�	�|tL��Ʌ
�NN�"
�^YRF�XW�uݍCv�òP����|�Z��A.:�-E�!n܆��x����.ܿk��╚�N�>:q�;���g$���T�L.8.�Z�j�ʢ�p{,�t�mM�M>���k���M��J���Fl|�tk�z�&J7�!ݭ#O��XC�Tݵ���?����h�L��e���iH�(/K��f�=�p"Lz�wF�a%=��O�N�1~�N�L�<�u��(���>5;�\� ��� �V	���3wħd�u(l���A.T�����ne�W�Y�c�Eʤ3(���(jX��Z��P�rTq\-����R6�\�:�H�rM%-��(��c��[����3OĮm���y泥�ݜ��N���O��<�MЗ�x/��8	7ft��ղ��l|Y�`���G!֎c�?����cX?���)!&���M)���ㇰ~|��_^��y�8e5�6::�ri^~��|��rURt
��眼�!�W��Z;v$�Ŀ�t�
Z�N�9�F����8�=	o�f7G tњ�
2��m׹��5�Ld�*X\gβ���K���i�͵G�a���W$#UfQY��8�,j�-bBc�����6 +X��Fb
�� �w>��˻���skw�s��u\o�'��0Y�q�?�b٤�"�v}�fJ�E��캱�L�s>�I�q�hV��/�u�N�VK�vpr^�sO<����l\+��)#�I�G�8^��u��n���1��c���8�@w����]<bJ�lN���hu��&�pߎ���ֶQ��7Q�2&��D���Cxd�v\~����o�Ԭ����i����MZ�r�֯�!�bB�� MR��kW�74��&����;)7w�P���d��Զ7��l���[�gҦQo��ot{�!���h�:�\LN����l�BK��a���<�H.�ZsYo��9$\�����p΍H���(���aw'N���cE�&zOc"$%/"������P�;�s���L���'����n��x,���Ȩ�_Ogc�S�S-뵬�q��6�J���,��ĵ��1�Kb��]���q��14<����^�Mk��ܱnDn/i�e�FFV\�ZY\����(޽��xW�;�T��\�6ޢ�����������n|BM �G��Ō�2�D���BC���n����%v+f�䣇�މS(Oψ��Q�e<u�ˢ�ֈ/��яO)(��?�Ν;�c�>��G�� ���p��Q����oLkccW�O�ժu��%9�s�(�\5���
�U#]NnF��1������u�X�`Sv��hnd2>�I��6������E�h&Q�v�E�5H�B��-Ǿ��6ZD~�a+Y��j��~�2�q�sg��;����oY`/���ZPm�|��˵�60�l�Z���.簸T�~ ��!<t����_������#-B[H%$���K_��}��I)�
|ΰ��p��^l�Kt*��axI�	�C�IP۬-���۰g�f?uF�_:5V��`+�Op�J�xZ��T�������l�5#��K*ti���h|2Kĵ������Qj�Q��12�Eb^.�1�|�����8��[رm7��ȣ���?�Z����������ޫ/��'����q,N_�����7ʈ���H����r~��g���2�&�YQW�3��lEp�31�T������}����抄�m@'0�Ii)6A��Fb�h��	��E�؏m	���/��)�T�� f7y �bO������)�� ��yV�NGL� �4�X����� g\V��H%�KSq���غu;6��峧q`�Z�g��Ͼ��&���g����>N����\Z����}a*��e�쇶ι닥(5ɽ�%O��e%�ـ��Fq�D[�|���1R{~8���p�{��tj �&���Ԯߖ�21kĴ--WBܮ��Y�o܎lZ\�{���h��~�&.��L�:�_��};�GuaK�fqk�:r�am����q<~�0�o^C�QÃ�fu�dA6[�ٰ8�F����z�6ғ|��5�^�?@]4sT[�%3f��Ec��f�n�h�,���q�]�.p������
佀Nb��t։VҮ��h�@�f�����ie* Z���������Oy����g7���Z�LL���2,/�Y�kif5�r��1�4fn^��������N�p���o\Q����gqsr�{\�ʅs�E��ѩ7Tu޽f���)L�P�XZ	����`Te��q��Q���*��n_{��=<,�e�lR$��C��h����[�.�ia�F��d�Z&H��n��&����x��x��A�N�8��l���O#gI��(�Kظm:�����Y���}�n<��Y�8���Iޟ��?)�zt�Yg��@�b\�`�������T0<o�(g���a��i�c�GK�X����{���Y��<}��3
cCZ(K�0�g4{�yXЧed�Œ/��9���XT��)e��Z��#��0e����/���{��}��sh$�"ty�~��o-"?4��q��0����kM�������Çq��qQ�cO<�M;v����r_�ߦ�eI��Y^ʥBP8�'�rI�\�ņyb�A�1��|97�ܔ��2��Hb��4��"���S��l���E
�z��Wb��8\T��f�:��V�+`F��$m2�Q����$>�ſo�N|��Y�<y	{����[������%|��ǲI�8yR�?s�\��`[b(q�R�7� qX�q��3�Z���^�P.�V�tz�L�B-B�@�L����o��N�;���DE,�����2��[�p�;���v��4���:��z˂ZK�N
�Ϟl�j�m�;Z?���YQ��h|�$�� ����?�ʫ;$�=�'DPB�v,�r���x8�7�H��Ǯ�w��� #.1�oɚg�����~Ͽ�
�*�;?4�^�-��7(��o^x7�ߐ���s늝<y�������l�K%4������4�-�(���_����y4��p#��E0�o9��|��8��XhBx�u�󦝽to=�g@aMN7N��6`ʩgs�<W�+�����*��Z�+`$7��E�.(�2#�O�3��m��)��rSmׯ�����S�E�D�=}���*����sطq�6mp������N
&�H1�ɒ,^����,�	�J�~BlyC�D�<f�9nnD��������b�R��|h)i�L)X���5/�]�B�/��[�h�P��Ւ~6�2�e��=Q0+�N����J
�	��Z�|m\�Eݗ0��������Ԓ��Ή2fO�_�O�7���F����ז����-\��o�eK���C%_{�#����8����֏�ѹ�rɡq̈�C���3
�'pP=&u8`�m?��M�<��z����ʱ��R��!L�/��/��7�о-HŻGW��s�.ޘů_y�N�G"?*~�/~�ڍ��HC��#c�=.����V)d�9/nȈ��ǒH粨��_��\�p*��ׇ��]���P�9��v���b.]��b��E�����yD�x��悚�5fWpGX W��}���k"�1&ׇ�ǃ}�|�P����~Q�IL!�>@;�h6U_�	����"۸>�J�ir�@,�j��5�����J��BI�NV�c򟒡��Ι�L-{d�n��b�8���u	�|��.h�E�XQ��.�y�<��C��/�U��<}c�+��R��c|�T��o�����|>G�l[��1��-S$���R��Y\.%B��!
��pnr�Ͽ��C����*��us5|p�<N]��~�J�[b�Z-_.:�^���k���;����>���γ�[,I��C��@\��Ęn$GlJ�$;4�l&��K�b49aqV���َ����`�C71��BŚ���+��c4��G<Uu�ĭfY,ia��,��>��P
����4�od+vӺ1����
?Ǭ�#4rJ�*B��L裟I���� b6����������NW[��79m��:zIW�Z��¨Xd&=�C
��\�8L�\*�(v1UD��E:�(�cHK��
��I5����/Ib�C�O��X�㵣'p����&D9�>!B��ۈ+�&�&��"�3��}fs �9����m��q���['��;GŜ��Ũ�9�]6Xq�m�����xFۢf#	�;�/�f�(���!	�7j:/Z[SX�m6B�E �5N����=�˹֗Jl0R�;��6��Tw
a,I�2�2yr�#�ZgUT~�����,B�*I	�Z�uZC.]@���A7�:�լ]PſJlW��0L�)�BK��`*����`M��ZV����0��ۃ��y�w<���z�Q��r�0d;nQ��T~=Z)����B���&[\./��5�;μ(�x7)oo���\BQb��S�퉵L�@H�����*�����r��2���U�t��)ee��U�
����grÊ��{y�
)m�g�>�Hi��L����W���5�к�32qǓ��K����iml���-�L(7D�%�}$p�5��c|������ڜX��b��E�gYǁ{y[lX(8�.	Jf"R�[)x~�_�����6;�C7����PZTg��/�z��2�X��%3�F��L%��<��i��@�x.�F%���
�D�L�����s�M���/"q���#�X�6,O�;���m�osI�\�VC���z�!M��G%P��Ck�����62����!.%A�I�p�)N��E.�F�ի�?j��D@c�C��1%d�ؕT����g�/� k�vw�u���9 c-�\ ��h_g��u2KI[.���A���@2�p��و(gPm�����^N�u���ß���5��BR
n:�D�K H��G�<�������p���<���h���Z��^�P.�c�W������)��u�c��_�(���3	���A:#nL��
D��B},g3���5�#����͘��|�q-M�K	�N�f`W����b���(�(yn\�vEa�\pD���Q��Ӿ��[�8}���"4�1Lu��M��1����v ��IX����R��N<3��:�yw]����)p��u��4��x�q���l��{��QZv]�7i2���� �m�(���ڼ|�@�:��.�ު'�B����h��b��N�c��v��C.rL�$7�'(��*-�Ih�8!��쭌u�)t�Tq�h�ɫ��S@*�<�5�U�9j�D\,]�V�Y웺v�,N��i���]�5�P`7�j� }A���m����D4�v�w5Y� G9)7��trJ/�s�U\���S�����:��W..��͎�q��~��LFҸ,6psb�^
7eyq�ѹ�ehU+���h�G�_r��D��+�+̌��4D
�ͪ���Xsk��c��6!2
�5s/kJ��:�/^<���/��H<ڕ!�����ψ���%���~L�$��Ύٻ3�ңzI\E��#�>�J���u�~/%���{�G%f&K�)�v����v୵e����
��a��t�_�y�����`�q`� ��Q���v�vE�b����4�xb���:�]*�iC�#_���i�p:��1��`�P�I���Z��L]r�k�2���
�1�_ΦF�z� OnJ��n��Z��h��9�j%� ;����՞�׻�u�F�9�ĉҞ�c#��i
�
Z9�����hlh�zF^kނ��%n�86��hTk�yN&qh��`��l&��U����C�jV���2���S��{JR���(�R$Di���;Lȉ�H�Y�F�����_���Q�=�1�뜡]�f�	�f�I��!MoC�gl�����\Ӗj�$%n���ת���5^$^83��Kw�X�{��Ǟ����(x�<٤\�����w�����uVA�K�%�I���ǧ�љXZ�%����k��pt�X�q�n�{L9��h2��ZՁ��\�~[]:�Ht\��7����)����e�)��
�QݴJ�_^�YH+�V_�tv��K�ԷvNm`mqԓh��Z���W���(ߊb��R��1��D����Ni�c�FK���u�p�9�Uז-CdV׌lYZؗ����u��� �C�y�^bPg�W�/�[�X0(4��mV��r��z���b����SB�]��&�j��f��SɄ�O�ڰ���rJd�y�f�>�SnG�o�����q���f;S:��r��^ě�K7f�K@&M��񠻙��Ě���$�`�M��|��b�/ϔ.������o����s�>�� '�'�!�I���	�ݲ��n��x��:�#��#F~�Z+�1�
V���$u6c�O�A�\Gw��D��v�����HP�����ltu�xC�0E�y�K���e���e�Zy����_-)D���<�;��kt�(tx�ˈ��A����,�Y5nFB�X>`|-�s�9��h������ �y��Fi�+9�rI�a-$x,��;�渞*/Gg�������{>�f���Z!A�X�%��.iE�+����J�W�r����7+Ðʏ�=k˾�61����7q��]:�)�y��׮Mc����i�&��Wq�ڴ6Ew"��v����Eߛ:]Rk�2 �u���'qՎ�����<���o@�J\�����z�T�]��#��F)�wo~ �h���\V�]iA�*A3*IU���W�Ep�ݹ�i
T���z������� w$N��.6�q��֊�sckv��Q��E�`�ޱU�kZ߂8�i��=�c�ˀ��-���ޔHk֐xOm��8Jr%����݀�baXDi*��f��
�X�^� x�w;��<	"�W�tx̜�6̥��9�Z\�G&x�יּ��F�V؆�Ѿo�fS9�#1{W�-U�
`)C����uU�Y9'򛔖naH�%����%�F*�v�;
��qz���$/����pd�v�[U�/�r���3�{�n����P�0��z�c�t$��Ȑ�sf;v/�t�K8G����b�Ţ�y��~���W���iWO�i\���:^Z��*��=�O��L��L�%<q�0�ۻK7�+���<��<�������g�v�={�7���)nio��JK(�2�KܲM^���V���n���*���JE�<��o��l�E}��������6݈G�nH�:��7�TQ����@���ڏ��se��{�"�΁�Z��Q�く��l���b�1p�W�V��x��31-�C˲q+i�e/��(yC�o�T�2�^7>�o}��n\�pKs���w��L1��}�i����V���7ޖ�+��x%��y�=q�}�i�by���عa�:(rX{�֌&��t���%J��v�����`�Tܩ�V�GQ,p�6��q/Z{\���ZW���v�cE�ٺQזX�2�%�Y�U_;%��"{nj	��������J�=�M�������x��>lY�]���o�˚丮�Nf�^����4b#A �M���YK#ylO8�Eo~�_p����Oh"�p������,98Z(��� ���F���]{Uf�|�ܛ�U����Q7DU�*++��=�l������������`��E���4Mߘ���� [���/�?���������Iݳ���Qʰ����
��W�\��z��Ҧ��X�ֹs���hݚY1c=�4���>s��^�ftpN���Yw ����,�Y��,iQ���A�`ZKcF��5� A���|,�t�B3�""�����+��,�#zt�9��dk������_�c��A��Rm����3*D��~�5��;�P*�Б}�w������9yhl�ǎ�իפ��4����>����#�_��G��@�Z%t�e���~`�о��e��Y4hlhP
�o^�H	��@�4�B�ꊶ��4�	��d�ʼ�Ng�U:�^Iqej�K�5Ԣ$���檼���S��_���B>K�\F�-Mޙ�,��/���U���w���̧ts�08ߜ�B���W����t���p�2}�$�AJfS�/�_^��ׯ��l���vk,���=�a���ҡ��<�p�v�3�?D%<�&]�<)�4w��6ri��Zf�p.��T�:峹�8�1^�n��V��s�U*[!�5-�c�
67�(6Qh����Y�KK�4SY�Kw�
�2�-5?{�~�ӟҟ����u4q�"?���ܠ�#C�?�1����L�}�������%��A�.��5���θ�PP 8#�7h��׷�Q���6�P�FI�U�,#r*6�C���������� � �I!�� j4_e�:�� I�V��I��Yx>H}���+r�`�9�B�<&��G�K�`?�я���gg�����LK�w3���9֮z��Z������qe������h8ǆ�m�cK�n�a/2w��Q��w��f-Zp���HЪy��Z[�G��
�6�;wf����MR�g�1����;
;F�	}9�|����Ʋ�<8��zdl���I���!�YC�sjsl@�_�t��+�k��/ ����>:�����i+�={v	ǧTM:r����������Q:s�,�_U۷�K�FQS\�$��E����B�%�`Y�-g�] 
�)�؆���@�=i:� $�����Kȣ����ybKҊ6�;9��;��"��I��4;� �<
��t���{Ḋ߲�~��'�A<x�N�<��m��|�m���d����ZX�c�<G�Μ���\���&�<.U*�@\�&�/Ipe��y3�9[c��Ռ��2N��,�yd�q�"D�F�L�v����|uk(�?�v~n��k@���D��A�"V*@��?�³C��k 	��{t?�:�9-����#�i`x�Fv����Cz��W��Z����/���:��Q*��U2�_�
�Y����Co=i�"3���� ����6\\.�� �JYK�
��(/J���>�R�X��&t���@Fk����d{��鳴o�:~x�t@-� �����+���%h����'?e�x�Y ��Ԩ��~r�>���A����_���*	��r�nN��8O3�7�$�����6�P��#�Ë�TO�Z]dD0��d��3�WIB�#j���u���'�*=8�^'�RNk�9Ko����\í$��������:>m��m��ޛ��"t 3��H&x���]�Fhe�NMO�
�ᅾ��J?���!��*P�y��o~NM�$YC"��ť�Gr�Rk��gg�����(D�b����/�'N�KON�V�|Fs}���,遗�gOх��p�z�Q�_����=�Ɩ�f�AKC�M�7 ]v��Neh|����S�/di�����A� ��J�hjf�N��J����vF:�����	��j�!��X���U�W���<^�t��%�Uص���la@������tht��v��(�Lx%ݤr�;f�ߔ�ڨ��w���P���kh�s�w���z~�}mm�)*Bg��[�v��� 4�j�s�L���h�}�k��t۔�NAnR�pd�a�ǁ��R�P�s7n�4���2��X���tg�&fw����.j9]�ͱ ��yI���0�f�$�t�*�z�2t��~J�:��
�)�,��>��<��ST���p�0l���<7����xR�$;��-D8��^B�2����
�X�|d���� #�qӗ&���	:}a������!No�F�\Q sh��&�.�ܚ�l6t�w�\�*��I�`z�l��Bfs��c�\�'^���e�.l!"�ޒ�
��3R,�k��D�l=9�&Y�s �fC�X�(@"t��7X�E(�X9�&��F`7_u�D2���|�����\�D�m_L����]uW�xH~��Z*�G#l�Գ	�23G�@{S�9����Rl�(�	@'�vg j�r�cK�O"�&eڴ#Ĵ�-�x)�rr�n���N�<�4���Q������M:wm�>:�&f˔eA+�S��/y�V��~8��H�	�F�EP@Z�jW�� �s�w�e�]:�:��w'�<�ڪЭ�9�����E��(�SI���ˁz�w*)�@�>0���S^⦳B�P?$2�[ZM�̲��/�WD�&�]��O~Iay�2^(�v�ς�	�;Ｃuk	�l.ŊVeؾ�ӊ�m��P�I��$u��L4������:v�
�J�Һ���t+�*�e�X?%"��ĸ�� '���� ;\�x�J�
5�U�ZIQ��&�I�#�ʗ��Rf���ͼ���#u����T��!����vS�[ +��@���zl:��)	>�d�(��z��8��<����%K�-Q���>%e
�;��v�W
?�(Wq�/9��sڧ_Xk�{j ��3�7/��!9��n貺0��Yc��sjs7�m6�uX�(ؙ���4��{I�;�hF��M_�ìEM��*�(��"�Yn3��,�g�>��vX_��AK{���_\���+�}��g�O2��D��ܽ�D$JkP,4�����2��B�m�RG����D�D/��Y��Ē
d:��Y��c�b�*<�h$h����k�=@�p�ͦ+�e�������x�BP� $Gɔ���D!�a�B��*w���;,��K֖J�K5l
i�%�[��R�-)�5�^}��Б�ߡ���i�h.0��[��l�UJUApׂ�8ӄI�I����8��1�H�Y�c�~���{����wQ��n6-�V �=v�\^��������uR��VY���%�Ӓ�
��g���� �9��*�֨�%�ms��@�ט'=�
�E'�/`q���P�mԮ���7:7�F�U'�6�<~���l%%��g��J��K7\�k���X�
�����9a�eey�r�$���-�j����s���-]�*e�G&�T؈S��+�ݨ�&A��_�F=HS�G�-O���[�d��4���x`hk�%�l&)�0���ܬ�pJ{x���B��H�w�	��`���_E�Yl�{)���Dր�d�'o����=����ƌ�ҡ%d3uq 2�<�@M4��)YX���������C��R�#�F-H�-M�NRn�5�}�.��$�����$���u8
ǻRk��19&=�4�S_�O�`%x���z>���&��̧�\�-�i���ܶ8V���DG�+>���j�s5����ԗ:C�r"�R$�1�I������S�h��Z��R��E_:�`�P�-G��W�y�H��Y��Ңr��F�ϕD0E��I�L\��[-v?X��R6�|q�*ͪ4���
���5�c٨\3on�A��2�l^�����g!ee�啝�n�4؎�7L��8H�\�Md�	���b�e1Č�����C�N�;vѝ�ɹ�C�|��ؼ�5�|�IN��-ixؒ3h
=Bݝ�x�Rk��JN<�����u}�y(kJ!kG`ړ%���{6bD�]mC[�cܱ���lԺ��H8\��I��&"���&��{�gj����Uд��w�����[F8���i�����\�.��	�h�շ���ҩWA�Hd�����ʫ���~�H@�4������L�~ �_87��	t������L�lphU����ڄќ�vpŒ��xl{ɻ(։��8�5�hUa�
فM���g�@O<����b?��5��o/��.��,�7Rbn�lU�D%u(�r��& O|=Lb�V]\Z�5"�E��,�0e���J)��-\��d��nDy��VQ5��(�8���Z����6�yc�	��|�5aEn���ȋBJ�lj�DcY����/��H�̞�u����7[?�j�z�]yۍ�(!�X�B/UG�Q�����f-���v�N�l�"6,҄�RZ4H���b�PJt��p\!*���S9a�J����YP�2����ך�)�fjX[�~�������H0|ͳ����q�2� �%�\�����$��2�kZ��l�(�	m�O�"ЂP�2�wA���:r`/���q:��a	�#�+� A/}�������9���lk�Ќ���l^i�bB�ာ��sPW��KA0x�Xq�e�����$燝�vR:z�+��6�I�:b>_|�k�6Λ����U)I�ϱ���m3����}�Ւ�캢Q ��T�Q���E��_��c��T~_��D�f�g��k��Bsr	]�5scy;�o� ځ�R�dLN>�!�堓��[��8��@h�Ō�yf�dB`�+#@�V(��V
W�}�@
6!w��o�J/=���#/h��l�����c���_�/?<%�fɶX9H@ρ���cyh�Ɛ:�rA�},n�W��=����"�t�I� Pޕ�)�R�Q�\*C����ܛTf������ħ��F]*���̤��W+-���V�Z�%���Ε$jY%	�> �};��DW%k$u'�m����Ys�*����T�l�q�n�$� ��K��>i�c�������:�(B��*�@Ϧ�E��`L@�{]?�(f�Z��\���[��ۍ|>��5��E�1=n��l����i�z*,�������W�o|f<��8��S#��,L����K���ו��x�$��锫���ty���/��r�Rl�4n�Ρ"U�*�����}�W�^i�o?9#���H�nl���#t����$/&��@������G����(V��2��|~���7��"��W����ܡŚ�^��K��=J���$z��u�1��v��ˉ��422L��G/^�����˿WX�	EdwR�Mݔgso���i���A&z��֩h������SHɱa;�n�R��B���oP0�1���g�^�,i���ф��|���0^H���� &pF[SP�Mt(��R��s�ũH+)S�����u��y��W�W�{W����kt�4�s'ݼ~]Z�-�/P3����iv3�4tbbB
�lY��
�3J�=���uieyC.�P�-��ÖSؠ�l�����|���]U�Q=4�!�ү� �v�c�'�؁}	uH��,=yp/�_���DH%���y*�����Eu'I��a{������6��d���WiLŅ>`�5��H��+t��Oȫ�/<+q�`�Ξ���C����7y�Z����i�A�!0�qN�#N���h'���Mb���]����i5����s-�|1��2����[e+���<��4��v�
�	�X�1Ў���K5[<�ѕ�f����F�P�:T{E�!P&�z.t���}��3��	0�l1=�f���ղ.}��ߡ��2��������6`P��U��9E�dZ�D�?@{wSm�A3 �~gi�����V���*�����Յ[�f�6�lf��Y��1��鰨�E�0�J�K����a��ǧ*�X?���%*/͑�/��5���Ɗ����f��ɏޣ�L��x��o������i����y���_�����? �ՠ��9���h��Np]Z��;:�Df��5^����K!R?H4�ێ�!�:���٨�(q�8��JZX��0!�����<i.-t�	��"�V!b�{;"�h���A����/�rh�U��=	h�C�D�FõE��k����ʀ:�x�8B��� �g,R�U]!�	�����ݰ�y#�5B�3�t�� F�&i׮]��d�45{��?�	���[t��ݼt^�ae��d��7�\6-�aK++��`e���s(�.�GK��߽�N��S�d�ɂZ���5R^�?���4�(�>�-z: ^�ة�B�o):/]����٦��t�\���f�9i�����Ta�U�0]��R�!�c�_XxQ���Aiu�>@�Ϝ�\_Ձ���z��b�=4���c`1�W5�D����h2�}?T�0�����=�y�tnR|#M�4��9z�w���;�.���4���R���aJ����/Α�BR9�����gT�����9H{wR��H��9ٕ��%�y��D�
l���B.^��ڠ)WH��i�l����3��V��k]73֘�]��Յ}�D��m����{������L��XK��e6���"�8r��g�f���K��7^���7$H74P�|6+��lb�����p �2)�[�Hs��C����D��Y���4�\YEI]&wI��ت�3U��p��%��Z曒2w~� �vA�>˚-+�ͳ�ej�,V�Y#�D@IZX^�7�z[��>=s�?�b��N��}ҷ��te��k�<���RP8 4�&p��	G�U���]8�j�	��}:��"�_ޏ��������2�7؇hұ����~�-���B��8I؎��!P�aax�=�<oL)����+wn#��"_�@U��衽�����N^�k�?'jԄ�(߈������t���J%�>u[���	���P}�̅�f�ܮܡ��n�N�a�#��@r��t��
�k���֬pa�~�%���1�90LWǯ���K�`�c�D����x�nݾ;�%I; ��d��qs��姴K^����tB��m;6[�R�����
��k�$ S����G������f���v��?
X��{�}�g�8H�Y���N�fJy;�Z���]'��la���~I���0+�����}�c�ru��Xǯݤ'?B��"qaa�����˄���	�����ifnN����d{���].��T�{�l��]�l�޿��v�eJ���ZU*zUz�Pa�De�%��X6'�~�R�oT+�L)�\�ϵ�م��k$�Y�E�z�v���3��c��B��6q��a3�0BC�-gxSĮ�B餑ViJ�G�\�1-/%EP(��t�wO�w���1뱴PI�����H�{�/�Ke���A�u��\ `���2�I�Ы5�;s�Į#"�`��4q�&o���{��Va[���L´�N����c}pn�Ƨf�,MIu��x���aѷW�0�.pŁ�N�4x/<0�I:���}���hx�^Z]^�����~�Y�����I�lB8"�@���|�M��X����k3�B���`� -�nT��M��,�1g�W�d��\N|91Od�$DҊC-dlu��c����5��Zv���iVX#�ȩ-S��DY�.kRϕ&��~G��+���[B!��俇HK,�����)�:5�M��B�F9Js�$�ا)��iаŞa������#�"O��+Jښ����zkv��-0�f����0����kAĝF�}�l]�1C7��$E4wg����W��S!��g�7h4)�H
�������_�����������R�.���t}z���oꂘr��]�H�r��n��=�{ <������j9���ES �y�-����׿A��(@�1��J��\�����3�~�}�� O��{���1����z�J���4�fk6��(/>a�?G3-�H�O|����B���E$�#��%L�gf��Z<m�y�X�q,O��5j*hW�[����EM���A�� ?�U!˕����/�|��G+Z�<�J ��~9��<)�{��Z ���MR��j����k����U�z!o�n'Kzi�,��*i9Js����J	~嘜��1U�&����7���jQ�2&ۧT�%����¦й�ĩh-�3�1�УΗ{���W���?�+���/ӓ����R���x����OЙ�"�o�5�az��psŦv��alM�4B�qH�!�{�.�=����%�=Z�ޘ��G���Jo��[4ug�*l7�a3��z6tA�;�p:k�I
�-������e����h��s"aZf���l��]��&$���;jS�wY��|��e���p�Ji�jR�3�4�)g%Д��>�^����T��N�Ӭ���r�"�q���x�ս-7XS��G`J�C���	�8��K�w�g����˷haj�7�������?�{Z�'i��$����G�Ǒ�$ $�p�4Ռ�)�5�G?�פ3�ճ�;2���Xsյ�>nYӡ��:�B�����^`��jBƄ�pa.�O�s�w޴S�X_`�9��3�gX��K���G^�ter���4S��g�Ӱs ���.E���Z�n\nYӱq�d��)��F��D&ǻm�w�eV�Eɗ]��a�}V6�*v�$�s��7�(�pa��  >{�#�sW٤�	�W���MNh�F --��E��WrNM�M���:���\�ɋyf���"f^-g���ȼD����4e������y}���6i�#�ͤ/�x�KvVv;�L* �BK����� jȢrst����4Ay�S�Y�dBM!�Q ��&�N�k�~*����ͱ%�6��`sճ��f:&�oZ�4KsVN�U˰b`����%�ՍA��·��Q4_*�6¬�/k��`�RU���L
�o����Ʉ���A��(!�o���Se�hr�6?�i����h"r�&&��F�F9
�\h'���JH�7h�ރ_nI�RI��sP�7���b	��b���� ]T�s#=��$�EYP(�I{9~�$�h�CO2�.�����_f��QlEuq�����旚Td�+�d�[��(����Eyp-C~��ozf;djDCn܌�4;3y<�;�g�&a���.�;�
jd��gG(?��b��7YUx�����Xe� %��Ҿ�\���q"�Ϧ��=�2p��� � k1_2�[(����i�`w�Α�ִ�i)��:%��vq�6��o�؞�x�G�<��j;�~��?R	� Z)�V��v5��t�4/|�M�b�cM�SD9NX��g. [HIm񌚱t*M��'t�T�����D}��ȳ��0w|L>�G����,�V�qK�ǖ�nG_����S��GF�ѶS	��?|�i:���>���n�w&^4 �EIH�$��y��l�8���M���Jb�>X��9�~�!sq����F�6O��~[�B�3!�^���P5�a� ,b�I�7� �6��܉ �A�<v�����o��#�9jGn-ȹ�m+��5?r�ȊXk�����~���Uk�w��z���#��}�E��� CIj�����вՕ,8�l��u�Iz�cKB7�W�ɤ�'n�X*Hb�_}�qz��	��k��	-�e:�JE��Ά�`3��z������Q�n���p}��`��e�C���׍u��p�nW �k�~�D����?�.v�~Ks���p����W2����`�X�B��쪤Q:6�&k;WS�et�)d�˫+���y���r��ɱ��pf|�����' ��`� ـz7ٰ�ӡ3��6�߈X�9�����U/��N�Ɵ�p����ھ�V���5Ts�tm����!m62w�p�b]��xa|�u^8���_�f��W�pp�h϶е�U��,\���S"��r�_I'�r����<�,t��v�\���[�+�f����zEkQ�PR�j��R
����LG��h �K`t����6�6;��b�M�Ưoz~���l_��f�V��n�������6�Z�e�{�X�����*?� �;:��]j�������Y<�Z��!z#��z���?�:�히�^x����������3���W|�?WɁb�^�J�t6��%�!*����|d�m�ω�q8
���+u�jq��e�G���q�5�����aA���jq[����u�붗���b�[r�Z���R&�FOʢ����MU����v$�s���n�1o��&f��㬹��1�-�
��{�U�9kwg���^'٘Ut�[e�1@��z�ox�!�0(p4>)iM�Rk��fj��\:��/?��I�k��0�����扽cNܾs����K�˫��	�HVM��~���_�S��O���I���Č-���F��F����2Q����Z�0W�	ǉΣO�かE��j�j\��k^�]w`|V�b��O�)���3�(W�����[p"G��������Q�
6T/��t��ʫ":"c��o�L�����b��Ub-F�9��4���f��T�,cǷ�넴��덮�B-�>��r��'���e�e�C 1�M?pU4	l��33T�~p����}�[�5�{:�T"Q{ll�I���j��6n�_C��v��>�?�n �]#~��	E���M�������|��{�{��l�����}	�F���N����Q���l���9��xX��5�*t���q�����m=���������m=���������m=���������m=���������m=���������m=���������m=���������m=���������m=���������m��$�Ժ�r�    IEND�B`�PK
     ��Z���S� � /   images/0795b188-35ce-4b4d-8dd5-08667f88bf32.png�PNG

   IHDR  �  k   Wԕ^  iiCCPICC Profile  x�}��Ka��ʆ����h�J� �5�"谂��<O�����-ZC�?Ƞ9hH"Z��!��&�������3��ޏ����󾼼�?�1V�P2+��K+�U)�
=�4�f1U������/{7&f5����^�tz������՛5l��/RXg��dbu�a�w��,Z��"8�����gnf)� �!��%n˙?������Al4��E1�4���Cʐ�"�G~��'�A�2,�ˣ �zb�	�,L��L� LRĝ[��o�On{�/�t�s~����������F��@p]c���Vɟ�o�@���5;Q��q���� p 4+�rެR�pi~)j�^� �   	pHYs     ��  eXIfII*            (                  �    
   �       �       �   1    �   2    �   < 
   �       �         i�      %�    
      Apple iPhone XR H      H      18.3.1 2025:03:10 13:59:46 iPhone XR H      H      # "�       '�    }    �    0232�     �       	�       ��    359 ��    359  �    0100�    ��  �    �  �    k  �       �       �        �        �       �        ��    �  ��    �  �    �  �    �  �    �  �    �  �    �  �
      �    
  �
      �
      
�    "  �    *  |� �  2  2�    �	  3�    �	  4� #   �	         1   	      2025:03:10 13:59:46 2025:03:10 13:59:46 +01:00 +01:00 +01:00 "�  3  '�  E~  �  %O               ���2Apple iOS  MM )  	                   h     	        	      �  	      �  	        
     h  
     �  	        	         	        	      
     H  �       �  	             �  	             %  � ! 
      # 	      %       & 	       ' 
     # ( 	       +    %  + - 	     a . 	       / 	      � 6 	     e 7 	       ; 	        < 	       A 	        J 	       M    .  P N    y  ~ O    +  � S    +  " U    +  M X    ,  x    " # # " #           �  "   " # # !         � ! " ! # # !          � �! # ! " ! %�*"�"� � �" ! ! " " Z�|� � � ��� � �" # ! !  � -� Y h � U%� � �" ! ! !  � �C� � � 9� | �! # !   �� � i � IG� � �  ! ! !   � 	� w _ g 8� � �" ! !    � � � � Q Q � � �" " "    � � | i _ E.� q �$ " !  ! � � x 3 ` (	� i �$ # "   " � =� I ) : ?� c �# # $ " # � ByA8�!� W �# % $ $ % � >��/��o : /% % & $ & � '��2 ��;J  | bplist00�UflagsUvalueYtimescaleUepoch  �e<���;��  '-/8=             	               ?  � �e���G )E���=  n`  �        bplist00_Ab0ADS86MCAjpKaa8LFhJJlP1mqK                            '     �  q900n C4B2F7DA-8462-48A4-BA2A-55C71892FB82             6    @� +E  �CB48AC14-E04A-4371-B2C5-73D7213C0CAE bplist00"A�                              bplist00�Q1Q2 �
�	S2.1S2.2#        #@=      �S2.1S2.2#@3      #,5:>B                            Kbplist00                             
bplist00                            
bplist00                             
bplist00                                        	      	      Apple iPhone XR back camera 4.25mm f/1.8       N        E                 K        T        T        �
       �
       �
       �
       �
       �
      /      +        d               i  d   � �         OO H  OO H  zQ��  ��IDATx���Y�$�y%v}�-#�ʥ��^�D� �� %�̓l�>��$����?Pf�IF��J3C9�F@@4��}���r���w�wι~3��AQ�1�����|�������W}�;��(қ�Oz����\�}������>ܾ��y���jo�8�?�M�u����z��+���/�_<z��ɓ'�y]��Ţi{o����i+{�$�y��I��M�;�'v{S��h4������,��ri�۶�<�~�{�������4��,��֞b�������(�� �,�_e�OĐ��ǐ�(�l6�>���O�s��.N����/g�TEݶ����>o��?�Lhy�v�}nC���c�[ق������7v�}���c���؝�b��]9��{�e���y�W��~n��f�Qf7�O�&v��0���Ӊ=]Kd�̝����]�ߺ�K;�a�F��ԆiW�E�}Ĩ��y���)֧�1���m����)��b�|�7ê���j]�����dd�5eo�d��n��¨Kz[��#|��t�(+cö;�Ol�Zm��ę]`���޵�Ʀ�S��F���A-]�a���g݁����nqO�����͍��n}k]�;D�"�C�7�p���4G���pM�o{Wbl��٥1��V�����]-�9w�h�6�(��Ӎ#�V��8ύ��,�G'in����;��Q�OFi&���4U�kț)(��%����{<�۴��ܷ��4m�x��O������,Y���nQljϲii�>Z���5� �>iqO#L�A8�^܍Flb��YIf�_Gs]�G��D���v
�m���A<h��}��䷈k�������w��
�h�{�b�'����'"{�-��qF�;z��Ư D��k��K��K�IW��y�o��>Y:�:��2$j7�j<5�h�q�.���$�N/^�0akolvvO�\쉍k�Q��;LbL�]�oew��D�<�U������dH�2��oˮ�3�*��=����y�jeF���I`e�M��D;��AQ6F�f������$$�7��;�*�G.3=b�^�Ϳ^������F�۞�^�L�F��O�`��H�M���*�� �'��	��bk�,B��;|k�G2�$����6�҈��h<Ч6)�M�A{�rH�,���NQ2�n�R8�Bc�n;E��w=����m�8�
<h�L��89g*.T��l�2A`Oi�UKU�+S�NB��a�}]��M�py��L�p�H]�*i�Ob�a��zm���7&
��M*���9W�1{ �ʘ�H�"�7v7�W��Lp�3�ڀP�{#�������l���v�*y��7���Ķ�ل3�#'�HP�2�Ed����}b�*	d�d�\�G��͸�E�M��)2�l��VX���%�7�}����h#U[O�a�Sh\���,�+Z)%5D�x�c�5�UX|�l�M���1��+���j�D�j��ʚ�ޏ[�X2�����M��8k*���t����͆�(�,jn��r.=�_Z0h�^<3��{]�`3�8F�l+׫�>��N1���8��K]nn4��8��v�f'9�/yP^~��ڈʆd#��<�m$�%����2ʷ[�����T��{*�MJ��Ʒ4��aMUڷUk����ڨ��+�����v������S��7Ҁ��}k',���V>����l�e{�4m��&�������a�օ��\kh��m%�ȧ0\��2K՞s�6���"�ݜK'z��F�����6��v�=N*�6#����(����2�����/ �f��ld��nq��t4���[�Y��¦0���tA�!42�lF� �q �nt1��(*N�������H%�i�:���N�:��3��<�_#`���KZ�Mϵ�L;8���KrO�|��g�M�D����uލ�kf2-���E��8[-�I�6Q�}3��S��c���]\\���0mk���0O�5���|:��R�6�^�ET+}���,�ζ��VJ����Ǵ��+6��|�#�WҪǘMk�
�1����W'''���1eB�G�1	��re�4�`]۲���lv;�qA��4�"����\QIE��f��k�|�称!G���~jK�Ory�6����h��C/.���D���.�g�]�PlT��l) T�fgo"�AN�4��\,D�� ��=&u�n��ʓ�(��[G���1a�P���IZ�g���&k��م-�h��е��.æ��bÁ�]�6�WZ�ղ�on#�}��fwv���Ç< ���5gW��l�N�.^�y/�RB,��uS�*�@cQ,�k��v�(�f?�%�N���Ft�)�ᕣ�L<�d/齞�@P�^���<��&o%[� 50|E�#m�&cj���X�����[�>��� b�a�o!B����]��*A�rN��l���l���1'�A������{;ʞ^l���zy��)��H�k0�A�%,JS��.��(���ƫ���io��M"�T�* 1�P.���m�G��L;��ˮw_������cy7��zZ�����*\�v3ob~����u(�{��5۷����z}��D�����?��O��_�{��a�Ƹ޳�ѱ�:�&X�<�N��8l
��
�&I�R��M%a�?�x/���9Iy^Z������Z'����+Y��$���L��3���#�/�i��SE4ݖ7��]�(R3fd � ���7竅&�n�*6�4�d{�HS�o�+O�9�u�	;���ı����®��Z�M��������}�'B�ecJ�sg<^o.�z���=tg::<�7��{�9�"rw�XN%W�w�/a-�����f��� ������c��)�$�k3���e�;�R���x�E���Wu��v6�%a���6�	���l�Uo��ų$O��BDf1p�i6�M_�ڦ��Zp4ɵwj��5�];��VA@Ogc�I+�W��P]G{�V&����aJ�����t�v0I�B�;����p2�	�5��`j��mM�-����I�/�z����	V>�
c��!���+G�X�`6�[r���<s��I +e��O���O��#h�Z�	A�AԸ159˅�pm9٫�kLJ8`�a�m�0��=����(.0����V"�2�1Yl�d��?����fVŹ��w�Y���:���0�t)
7�o��z|'����S��e!��xp;���@�j��8G��C�hQ�;��_2Bm�ʆj��M֨ˮ�Od��{���1����H��i_I$�Ӕ�`��LR�F�
FL��_�*�	m)�R�z����� -�&=w��7���$�ˢ�O	Kn ,���Z�<�oӵ���IѰ�����I�~�0*8?i{}�X�]q��^kH�ϴ�S;��D�,OE�m넰(��+��D��D��F��/�"H-��`:�o�7�y����b��qDn����EES4�C3�w�j/hj�ɦ�xODA ���)�XF�4!����+��z(�zv����R�$��c��l�ɧޯV�M�lV�'(er�IíD��O[mt���GcLp�M���ij����}�i`�3JW�
zD��eR�J�5�� �%h:�8n���;/(0�UL�^8��޺a,-q��c��m�9����*�I��&D#�+����.����D�~%���p]���m�x�H��n���~���;H�n�X/�ō!E@!��tY>�RN��ǟ�h%B]10�MS����L�`���R&i�,ȱ�զ��ґC���G�6	�F�	9�e4(��aC�7�
:BD��f40������r�9`Li�0V��� ]���2m���� g�m	)��ם݃���M#\�;c�O�m5"��w�ѯ�z�&h�5;@"�H��߂�8T 1���`�b�J�{-ȏ7����T�"�p�mcO���Gay��{�9�`�~�=����[�;ߧ..;�����������U�1't	lv6)E˼U�H�p�>�*����K��pt��@p�YQ��ީ'���V��V���aK��{�O@F�=��H9�h�j�����޾�N�� �Z4��q������.�{�G��~{xtvr�I����]�����?Ob�E벒���6{8�
�����uU2���}Բ��-ղse�s�"�n�� 
2�<^��<����5]oR�F�q89�n�Ĝ�'�2��@�FK��D�f���Ƹ��߇h�jy��gS|Ri�@({���-J	:�.��
B�/�����a�/�;FqR���-E�	%m��...z�xNh�;#ʷ���v�`0��4�'�lL���J.�2B�e�$]�k�l
�p�Y>y����b�g�߽{���"ާM��yjZjK�o�!U��a ��՗Б�2Nv���wO�\0����p
�����b��y�2<��.���/�Bt��{��(�ԍ@�p���#�y7�����v@"�@}���$��/�St����.������I0���Fig=:� UWS��W�tw#9ä�ӷe�)H�k�̛�3��*i�[c��|���g������ a�J��|�^��NhX�$ ���W��$;�� ���?��}>��}����Ǳ�0�MxK4�LF���?���������F`�G�e2_�l�����㯁�A�Ů(M1K�
&�HW�[�	Rzkʔ���O7���p�\# >6�7S|���T��Wg�^8P�TFIƁ���ވ��~#q�"_��6�Kא LL&�]�y$Of*�و2����1�G�D�A��ֳ���*�b�@��	��P���?���^^�k �j�zة6�،Zxg)fmK�6 �<���`�.��bn� Ц��1�gyGؼ�ߟ�����"c���è�����K&��Hf�)k�ؿ !O�m3�a>d*�aȅ �7Ƀ3,��ŋv��ϟ/��_��]�8�v��>���ӆ�/�xd�~���S�5��&.1�]�p�F������zk?)���'Mb{�D�8���8�������������n Z�6>x^TF��4�l�{��tv��]�X,#�M#�n>��eE	���5�Yo�����_]\.o�1��c�c2��JF�r���2���8$!q8R�
)J�,��	�i(q�h
$4�i)2�k������V�&h���	�(+P�Υ�r�V] R7&TW��MB�P˨��}�p���Eh�s�bќhBJuv7�8i�4B��ݰ3˺Y^o �	���_-���9��+�m䡴2U>f��Nb�8ݖ�I��o��4�"�=���f�ew�*��$�Aԕ9Dr��`����
�h��5�2|M^��ֺ�ɡH��73�f��0��^_���W����/������|f��4��)Q^$[�eSWzt|�RP�	'n=�aVq����h�Ј�ht��ue�P�	����K!\�U��*;#N!�H۩,+�2�fG_�
x7r��j�f�B>�z�^����j�qU(�o0��D�d�*(�JE�u͢���ԝ���l�b ��^��%[� 7�1j�ˤ����������B� ��gP�
T��m�dgAi�5mM�D|D�)%�%!�㋫�$oV���Df5����f2����7x�N<\ �,�M�f�g*as���1�o&D!O���$�u>���)>Bӱ�c)D9TR��g�Z�;Sܢf�y��,W@Q�����C��s��Iƫ��#O�g��R���u�t�ً}Jf'��k:�����73� j��Ք5��saU���H��r��$�%h����\<{?ʠ+��*?��c��":�S���iT$��ϓ��F�ڔZ�29������`�_+φ�����3W��	�>񓂹u���-WD���K� ��t̢WB�LC�j�������$@�O�6U��L�h#���)@M�d�1�hS������2�#�GEԀ�ֆFZ�'PQ4�ed
ʍ\ DHz���}ʲ�e�9wX����l�a����4�l�G��pU�₏gs��HJA��{(>��lC�/E��ײ-;�k#3-�
dS[�2�2��Iof�g�$8KрGC�{L��JW��!��x�(AT�4���{�ŬŔh4���md���I�8e)�#s[�&����?A���0*U�t�i��^�8��Xh�8���Mƶ_�9X�uU�v�V��b����PgLnW��D��*����#7DG4A#v��K��I�%i4 �P3�`7��$���<b2�rR���5w���ø�����߁�HuB�d�D4Iۆ�VivÉ�7���h+�������: �{{s��*�C�/_��ϟ&��K7���_��̻VڟBI�7�!�OЍc�I�L=Xo�[�C��k;)�9&Q'�D���0�EAB&O��ͪ_3jxS��1Vm�ג	�a�xP���-h;D��Ӗ��7bP$MgԤ���q����&,DL��(��<o#�<e�M��rm�R�[3 ؅�Xw0�R�JHo���M]�4��!cz<'�1s#�+1S��'�A�f�uCM��Ǟ�g���$���l��(gӘ3��M�>�[�P�����؇�kyv�+�A���%K��a���TUE�h)eA�w��19��3��e�h�S���y�q��,� �V�rx��O?� ��;T[��tkI�V�e<�����E�ݐv� �d0�8�&�-w���� �Ce����>�E:�=6��H�(��@����m�HR��Z��&$Z�MpF�����H�%���݀���;	M��S�Ƴ��ײ)E�HvP����%�?8<b:�H(�2��F��x���
n��)���5�7�^0ݿ�J��u_	�}�+��ko��o�_a���۠ �F���>|�w~��>~|��f��/���z��CVD�y�����q���IF��^�gjZ�gg�Z����\�h`Gs�k n� 
TCFLقi�hB�D5��q.Ж��MA֋^�P�]Ȁ��P�nt�k�lȽ�$���萣բ8<+D֬k�%x�T�M�jY��ő�]B:���J��F��- �V��ݹ���ٙ��>�81���X\�s��g΀��ٹ��4n�XV�W7f��;e`ٰ���L�,��J�-Ūa���R��8�q�a��T��o̠L��%����Z�jIT�e�ۨ�����<xP3���줋�|.C���H
��,v�t�y	"�#����pfy���ƹ�:/
���Wr���7ٙ�W_��[���=}��xh����RT2�� ��D@Zj����gϞ	#H|�4AlhzȦ��6e��c��z�����)v���'O�>5^��R�V̢r ��{����渾x�����,
[�����۳����e.�ƺ^��A�W��E�ꘅ7�sdQԦ\���������|n�L�2���Ye��2�|��B���MF�s.$�*/i��$�i��{خ +#��ri�� ?�i���#�S�D�OɃ0=��K#�[c2�ɧ>�3�#�sCnB߹��a7��b=Y�l��S�@"-cg3�:�s	�+i��&����������ق�"�
K��$b]#����ؗ��.��S��x+�'�!�l�:fV�O�Ҿ�(���|p�Ν7�|S�a���mZ���=�,R�:@�!�B�w��8Θw,=O��eͩ����0�U�ʇ��N��Z!�t2^��z�B��|�-�T	M:l�:',�k�7��2P{�uL�״SF�xz�]��eTV`��9�!aR���D�[�<�7�$�O����{ +�+�-1&�q�d�F7u7�o�<`F"�c�P1�z���8�X����ֿ�?D��TA:mo$�ug��4��	zD�F����Y����Ll�Y�k���5�t`�ei�pG�պ}9�L:}6���\�\ޣ��`o(����xȲ�)�ʪ �vco��q���Oi�^4z���%3^K���f�m�40�\��(�#n5 �ԖP�hHM�e�3���&�Y���$U)�M�j[&�����<D5�h�-�ھ�}rU�۾�f�S-�T�rQ}� QW�R^_���)�Lլ]�A��+"Ij���}��X�O���dl�Ć|�tNIv�@�`�q^�~DN����⇭�KL�@��ŀ=r��#���KbG$怀�^Y����ym	�X�U� 2f�zǒUޑ� ��|I�81F�����B��ܰ�낫VU�F�]�4�PBe7�n���tػ�	��;�z	혜Ѷ7I%�P����ge:�܅|[�G���	�\֬4T5hʶ6��:�����J�d򅜚`�݆�u�ii{�В?�	���*H��8V��}�33Xq�Z"�o����u��Ib�l\$e���'w�p�	+�|�sn�� �zQ��	�h�Ȑ�qڮ�D�`�J7����l-z��y�3�AΈm��$�){}Iv����B�w�EDIh�Kħޭ��	{	�uQ�w����Ь�$�� �-j��'`�ݵ��h�$U�*�a0� %PiP|6>͕�ô&�����P�7D�c?�]�J��=�F;^r/�:�Y�:x[��z��o��HH沢���H�)O_�Q��;M�K�E�f�y�&�?u�:��%�R;n0^8�h���w�CID<d����.e`9�CZ�6��!�?a������7W�n($�L�PX@VwL�BQ�N���� +/v�R��/�����:Ix��ǀ�� ���n����H0��`��\�|�K'(��"02��҅��#qCEj7���#�f7���C��7�A2�H�ޔx?��l�g>�%�Bl�vHnz�Hn���x�;o�uCm��=�@>�>A>l��2�D��P^�Ś������{4�(J�n{�	�1�-I5|uSgqX�"��JIg53W���q<h:�b��ݶy�����Amѯ���%��W�y�s9��!�=��~�K��=)�����/�~xm�=~����n)�4�?~�����?��?|��Y��,BL,���%K$v�ݝl:��X��7����w�������j77_]M�$M�[d�*��z��],������}�hP������.�1�˨A�H��TR �Ft�M�5p�PB�)l^���xHC��|5Ah��$�(���D��ns��	�a��l�tl��*���ɵa]F�J!d���aN�i���	�!�6�G����DÇ	|`mP�Rya����!!�vo������/`�ui���[֕=5I�k��i(@���u��s��R��]\��t6Ÿj��1[Al��xW�~2��䲩�5�*[*��K�(o]���Efʩ��h��0��:��gO�϶~��7��Y���^�_��7��H�kG���O>�a�Ε�����欚G�*_�AUl�^QW���g�3V�L ��&�'yV5�E����zy}}�X\�6�jfT�l�����ãc{8����z��R���J�\D%6��P�GF�e�T-�������3�y a�l�y�h����fhg�]]/�
��zZv�^�����G���;w�.��_}���Y�L6����%�B�擹�p�5(���� ���3�u3%����F��P�˖<��z����Y��U��-VoB�f���K�>��b�ZA��� J5���а�&1�V�b�>t�BÜ�>��/�X���h������u!4���k��n�����O-W�ϋWo���I����Ǐ��z~�|뭷����ذ�ڻ�����o�����A�B��}`��|�����g��ݳˀ��񚖙��^��;#��:��`�۳���G�l��b_�M̌!�W(	T.L������Jګe�
���8��=;��?~��n��o~���R�X��?��Î�:;;���M�==���|������G}���9FNO���S$Wv����_	��`�|jT����߼ͩ^(��x�\��O'p���&n�F.I�L�}v}�T]��,�U\{߉�V	k�c���9XVQQn�͆�Cg�i+c�]����3˯�=y:ʧT+�Y�(�k�B�M&>�o�`^+p���cq})w��h`�*I�U!��)|�J��I={v�9_���L�`/�e�}����r�2���!���b)�uq���ٞ��d<GV �@VW@(�<�٩��*��eC9�{n��9��)1�k��r�L�_+q.�ؽ��b��f܈��jYɒ!�Ϧ
�6�eD�����*�e4�w`��h��_[Y���`�H��PkG��^�
��j��U�7�MG� ZW*x�r��}D��4��`�dܤ����T�B,��^?����aj��eb�����$HNZ�Nj�Ŷ�m��]��
�Η��k�Q�#K�9���P�T��F����b�1n�J"�Rh��H �c}��R�i�O֥hF�y�0��l�����ԭ/.�.Y���5��V��n����'M⻦MS~1�v�1����в��L$^]_֥����7���k!q��,�񺹶%�k���+�v/�sZm�[�:�1A��WyT�2�:�{�!9e�Ɗ�;�J���,E�j�M@�#��=����	;b�"��v��`d��I�+ֲ,V+f���@@!��i,S��)���F�b�7�0F��b�H�n{���k:b˶��bߥ�'��^�#��v�B�W�~���th��o9�mc;�XW�&�|8!ez?���v]$�-�<��7%�f1�' L�2�4R5��K�)n.Ԁ��!m��4\��b��	`Y�0�*ul%Io�Z	Pl���<"L��ocE[���Ģ�g�>>��Wz.1DG "�	��;�3u�z�K�XY�94�~+7�3�Q�wM�bS�w�*��Fk�CN�t�%_'T�H��%i��s�?��H6����6�f��=�i3�Sd�����;߽�QNFqԴ>��+��,��o.pu���	5Q��l	=�f��픕ҊkR8]�����)A���fBa\H?ڐ�>H�Ģ�A�Q�6dx傷e峰S�PA8Ž�t�Ca��^�7�ވ����~�I@���+Bc4\�Qg#����Y���Y���Ⱥ����x��5�3�	y�	��V��ݨi��t�R<��"u�K��c%*c(���m��<�Ea<SX#�U��n�(�Q<ߨ1�۸�~�Sr�;�W�O8��`�ǲ��j
}�*cT��c�l���y&�����Wq��ֈ6N�I0���%N��Q����Eޭ�sMੑ�#Z�=��GYO�:a5���$� ��R=����������ת'XO<zŎ�yZ�!�V�E$/���d�)�8H�@{}{��/R�@��'��!۩�q��\��8O�������V�w�2�Ŕi�S��
� [�� ѯ��%/��o�݀o�6��A�2��o��Wz�����m�a?�ͣ!�`����w�}����>���d~��*��|oo������~ס���򝝝�X�������䦁��d��m�0K�2�^������g�`��p�./v��Պ��T���*�����2�S��Ag6v�A�G���c�>qTQR~���Jtc��M�Q��j�Կs7�����!G�P��,b�[�5h�"WB����p�@�� �)�������:��"!�
�S:�/��[�������{��Ν���)��H��(kXGVu-�Wlۯ��>^����t`�&�E���vՆM�v������ɣ�<����~;����p���_]�=zdC��G�"LP*�im#�C����f��,Zȴ�fl�2L%���1TT���/.Vf#�x�>}j�<�2Mv���4VTj��s	@-�Ś&5���b��:���->��x�/UOj�(G �		iZ&�p����Sߍu�g��,�;�c�_|��k��2޻w�\�IYN�VF?����հ����'��Ǩ�&,�H2��QE��$F/�5��4Hjq%x���6%h��� �VJ�})G:�(� q�x�KFc[�I���9PBm�E�}����/����9�����S���N*4PϹw��[���痗�FH�?�M� �G������={�.9�ay���{�G� +��?���b@iv���u��ꪚ�"����˹B�,����MF������o�%��`�]]]���cɕ�K��nW�-��J=ȓ�7�C7tRNDz���~�Ń�?���5���6zN>��3[�������m���?l�!�.�`�Q�nho��O������c���w� �fM�S(!߰�4G^����ַ~k2G�������d<o2�n�?^)��Ue��A�@�T@i#�D��A��x�Iݔ�ɔ�gc�G߹s�l����D.������ѣ'(��(�`�fo����M[�@Yu�ٟ�6��,�s�K���X�D����th07�f�4B;L���*�F�^%]%ֻ�PsOP1ͅ���<�~�����|86'��{���(��������}!%�~y��'�������]�ك=��w��'�~d�����s<n�ƫ�|*1w1&��P0F8>�W�Q:t%3j��TI�a�Q�:PU���T�w�P���t'�b��߇F����j�t�	Ҝy�� ڡ�E~�Q)2mY�)gL��H��k32Y}qq!���!47/��n�#P�x��C/v�ro�<b���g�QK����)w�y;�E����Y�A�;�xE��4�\h�P��$m'W��MI�:��	��v�MsC��^�$4��s� �|�o3����,�~��+-��)�S_��Ok6���x�"9�'U蜥�x�5Y-J\6c.^�EFd%QΣP��w_����Tц^Q���hGB���UYPAn�C1�7j��b�����@N9����Ϗ�o1��QG�1u1U��rW�5Aqۇ�)�7����&)S5�޴�S��UM:�)jJ�NL'��OS�$ _�#Y��XeS6��ǲ�B[�	Ál Q���S1�z��������ʧ����J�
n��u-�8��F��8c4�s��~�uw.X˚i4T.�������~8�~��|���ۑ�=��d?�nȺ�����M����KV4�FJ�6 L7�"EN�ܷ6����|�Ce�.%�f��[i|�%�����^�l�n��X��r8}�m��'R��xP�@9�A��/�v�ӷjr{����v�l8�a�\�wa�>��5NX��E5i)8B��]��?j�&��ZЪ�fT0������E�����x���ۜ�8�=@��DS�KF9�o��!���Ε݌P1���	�yvG��K��@�x(� �� ���U�Sb�]xV4�ݓ�x[�xuC�Z?�7�9��0��~ �K�9e��G�]�b��s�^�:zsT^��n6���U˟x�J�����q��![9Z�5٦�.�(&74���(��E��x#%
�
i�T�0��p��g=u[�y� �`T�?�e����!a0z�	���ehn@����X���{��b���M>���&>H��}*`�S¡���>��َ�*C0�6 &՚�g��m^�_�3�6�n�&-2�.�q�<܂U�.�Yu�P{���~K����Կ�[��wU�_�J��h��>�j�U;\6!�y�&�[=��ڭ�L/`�>W�� ��!�"�������(sf�O�y�pDZ�6�z���o��o�G@ں
q��R�w(�ϳTA�����d9C�"���|M�''�:�����2S��rI�ޘ����//W�D��54)�����g���㑲�6�g�<�
�k��A���Z��,��+����
�1��a�8���*d㌧[��n]��r�r�A�JD�V:����)G�t<�)m	`��(PL���0�K�(z�*�DGm�+@Y^.���Cơ;;3c�����lFK�<d4�G�E ��{{��������qZ��&�a��s��M��*��ޣ�]��8I�c�$��s�=2�WG�����R�+�[�m����ܨ;��ϳ������yۮx}c.�-�m�tǶ����9��d�"ɴNL%s�		XR�c�PkIpY��b�p /���'�]j;8��3�˒,M̡Ǯ-����M&MQ�M9�C�^��bQ.ˢj�]�NfԔ��Mq�)j�8�N��&��|kdTC��0ϒl�6j��
1dr:��蠜t1�׌&uIg�����U}]<yn����V����d����g��,��?�������eQuF�e�{q�kR���.�}R^�O�9k;a���.���LfƘ��ͯ���E�7�����_�uo2�f�Q�1A�瑦�69����4���5�'S�ԛu��u��1E�'"^�q�ij����a���+��,�q��������rf�4����9Z�X��ڱ�q�}������ۯ����ɭ��i��<�������{��;����e�Y�����g��Żr�?Z�~ɲ�?��w���M�
W��ė��=�ܨ�9>9�Gن>p�7]���%���':��P	��8ۮ���^.i�uh��~8���H��յ�q<ɐ��w��آ�pFA�\5���{��l��ƣtw�7� �2���f�x�=[.��P*�vr����B��~Qv�?v�ǧ'�~��w<<��'�ѷn3Ѿ8�}�����}g�&���S7Gif}s~�<�y��j�m���F�8a�EU��P�h�vYYEEa,�c�l#�u<�2(�g>-\��)6�lX)L��EN����u���ʪ����w߳�lf�ptr�e��m�{�t�4��Vpm�v�s��gO�/JX�����L��kؕ]�p<�����?����''ǯ�9B����G�b:xԳ�-6b�p�h��;�ST���2�!���ڨ2�o��T%�(��A��Z0�fi���HL2��@���ӏ>=;��D���������o���#tYH?���?���} [�ׯ�rj���j�`�p�[{���j�����mY���{:�O�9�/vv��lww���f����Ç�<摲(���;.K}�\&�w��8K{����;�>�������x�.j[�U�j�[���5�N'��4�f�{{b������Wl�VK4`��{�w�����-{ e[�4�(e5�v*�My���72�$$�ƩƵ���ڜP����gH,��bM&����B;���1�d�͆������*"�ӫ�d��:������RS#O|2�y�c�3a��д$���3ƙr�p�􋳧v7�pq���=��2�F+�)ۡ��|i�ƄMQt�j�XdI��f�����OǪ��<�ڞ�F3�����g�p��$�q-� �m�Y��%�kVr�<D���B9�@m �5�O�V���I.�	�����C�~�Б#ik�5ڷ�W��,��WV�� N4R&���C�wzn%���h���2`��t�R!v����R�`ob�1�1���I��f���eq��N�ݳjw8�C�b$H��cU��ڣ�̆+ؾR�0�����+�|�����?Fp���W�w����(FĖ�1c�
��,�vh��\�zp�P#�q(Ǎ�&�FeF6%^ϰ4�U���O�Y�f��`LST�$[4���^��_ƿn�HV��C:�ub� �=:��"��u/��|L���]�������2Y��l�6iB�ݶ�1B/4RRV'���"������8�{��[ߛ[ZꮫH���+=��(����!F�\l�%R��Ta�U�gv:�t#���f�y��RԹ�Iq4}�-���u[�$)��
>��)��6Ń�ӝ�.��
���h(�ƀAt[��1��g�5mG�#}6�����y�#��������d���6L��r���6j��^Y�h�{�%.JjxE亻I8��q�ǃ8��u3"Y5�1���a�ѫA$�Z����@t�g:m$q�du����Ng0"�WY��aw��~)�@�Ȉ�2��L�#h�ح�2l��2��E�1��t� YF�R�Đ����Q\SU�Z��]����'z���.���X�T2�p�n�S^�U���tC*��|ͣc�p,/CӂV�ѵ_L�혌�0⏍��-i����p�P���3ھLܿ��-40��[���K0� �Q9���͹�PY�=�h8�i�M�C�@;$�E��[`^��f���w��9��p,�H�G5ny@,XN��zr7�c I�A�������p��\Y��
����������E�QǇ+��!AD���I����y_�m�і>�� �s_��zw,��2��5�|]u��#"沙�����}�� "+�Ld3m���޽{f���o��ʰ83���a0*���"���
������o7�"A۱s�Wo���0��������dw~h?�6ˇ�.5�nȤKR���L����Y[�۬UDq(�H�0Z���������Q5ñ}*�I��RA�~����h͓�����yŖ�p��>�p
�|Z{sqq�<�c%t�J�LF�|"���o4�uh{������_�Ν����C;���\�0��hWi���َ��C���ή&k���gF	����+�9nVct<��i���ꫫ��<���>3SՈJ�5RW��_|aV��VqK���P���$�?W�aoH��'�EkX3�c2����v״�.//�jl�l�9	F����w��1Fi&(���a)�P��ٕ���0E�¼SOn����������I��IV�t��0�n3��q}��e�{���%�v?��󇫕yD>J����l:��d���X����$CQ��i�f&C$��d�	;j��!ob:�
4^�ݝ��o��2��M����cE� 4k�n�F$��3y6h�mE��1��n��2�-Vw<޸�����͈ ��zv`1��I�_��%}?m�|<�-�s���ɓ��G�=2��a�k����ᘳm���_��w��|x�}�;�1'_��@o>k�f�j77{z���ɥ���U����ՕT�Q���̃u��aG��Ұ��S�6������POOO����x���x\�Oe�z�������HF����mm��nb^`�,�������ݞ��>R�n߾��[�"��q�e�+��L����7��0�o+V�5.a�M���p���Ch�D>ц-!M	J���k�P �?��=z`�u�a~h�,��H���F9O�������Y�Js6�����b��5'��[�ٌ>������)؂����_%�������<�<�}V��S�Fl���|�8H�N��rQ��gp��=�;u��t8�/qU#Q��
�d�[H��H/Ә4�"�B�@�Lw�>F�F]	�P���6E�[#����ߨ��p���<��я��G�}���󍷌�l���-b�4H3���a�S�9r����V�Q�ϣ�x�����ψ!&�1/n8/{�XJ*�t[|h�v��Ν;�;�y#�	Y��5�.�$ț�}r|��ѷ���Zg�������i�/��l�W�g/Ό��������h�����DVl4$�&1ٿ����@�Ɓ�UQ�V���|h��6v��Y�߇��=�Z��/����Ւ��/c�����g;��(�1(��:����M��ޟQ&^��OEr)�d�K0>���7��ɷ�]�?kh+`����MПt��O4�訁Y���@)E�t뵊�O��:vK��?{f;�`�� �߿k�`O�R�=d����+؄�$3Ri�y�|h�)������u���(/d��^�6Х��R���(W���i�����Q-���x�s�l�v�>�����<�<W�5@U�;<������Ʉ�V�z�^"I�Xn�6j|���R�X����%���,<����1�llr���x�Hf���^=�F��.�#��`]4���8��߶_}�駶e?��υR�� "Mgr̦̊��J�m6 ���/#���8le��p�eK-�ʌ�5^K��[s�[�N��{L�'CkB���G�G33Y��C�e��2������_�O�,�L�>�E�dqm˲fu�I#��CkU�
�l��o��^\���\�xH�	�P�u�.�+y�Fl�`�LWKP��d��ڐ9+���$���@�����Y��.
Tm���EU��.t�N��u@�G�5����
=��)��=�$9N��j��N;�.�챥�P��.�	'u���|�p�(OOTT9xaf��et��ox�;CT�]b:����r��y�l�����Nè���w����N��֡m�����>�ٔ¿�2��3�q��ľ�����i6���&��ё|�.X}q
�>��oJ2h�e���);�7�?�U�ː=���G{�T�3e�WUʖ�oG<�^ܫ�a�A�� �s�lA!#�w�e�ϘŬ���I�8`�AԐiX���M?6<-@�[���I���<P7�|羫�ñ�fv���t`�eQ�`t��πU�ZR"8ѢL)PqA���xV��Ĺx���Hi��H��'I$�������߾�L�m� ��&[�ʹ����|D�
̴Cw� ����79��97������dH�n��+^�0��{	�+�m�u�&,�!S�1��[����z7K�tC��o���Mz,	F���9��
��p	P��ьA����Ͱa)fj�p<����*c.�r8HZ�K[��� 9���K�L�?��0���h+���}u�~���|�𔇹K���L�C^-�>z����d���ę!�Y/L��̎����m����������D��Z�b��m�Yg��B�^�PX*��Rc�MS� �L7���Y��hShR{�L��qU�����9?O��1����@�,���2]z���l��rf�#I	Jh���v@?T.��Cۘ���Ό���r	��4&�v��D���~+ե"�9a�aQC���E3����L�F�p�6J����l��N�"������6H`9���S���_ޑ�ѠRk���OQ�^]\���4�dU����@�<����ML9������i�6��K��_�Y��צ?"�7�'q4*6m>vY>a(���\]],W�B���Kʑh9�۵��_��6�g���s�W��ج�ttp0�u�Ԧ���&ɂ�G�l��Ū����q�ҿ�������q{x���/��&��k�v4���T���)��PPMeq���/������68p pv������-&�<�ai>U��7..��D3W_TE)�q���Ng��ۦ�Wk�iU��F� �ZU!Ys]F-r�f�<Ϣl\��Mݚ<����ޔ����t�gq;�w禁���//.��.���z�F����ژ��;7u�b��12VU��+38���!�u���?	�Q����>��7���o�Ñ;p�l-F�����0�ǟ��Ḥ-��w��q�N$�Y�QF�d,�9N��̷/ʅpҝ��Fup�4͞<}�V�t�ɽ}��q����k�O����,c�{U3����lgb�g���������}���������^,.�����/~�K)c�v쎳YB���͠��<��U��ڍ��� ������u��*�*�{֭����=�Z��F��V�c4?�i�'��)���y�>� �̾l����m0�
g'�)��zy��E�y��z3��G����������k����W^�^^\њ�s���O>���ۄ��Qq0���+�}������S�}0��%�SM��m&��rq}��G3'����,�[w�t�{��{@�	��$%�Vn��.��8Z0���n����+��G.e-A��IL���_����ڠ�2e_��0�1Qu�$��Sg��=9:���{��9Zf8OyC7�˔OY�H�E��$��hy�\�_�����n������Wc�<�Ƽ�5;<���gfΙ������ࠌ��y>�Ǚ�@�{����1@=S(w���T�<\�.L��C��	4W�εE�ئt����:��hze�yxN�ov���œ/�뚄=+w�s�8M�7��o��En��{�-.��_��?�O���ac]�v���
�$���sD�fӽ����}��|���ӧOM���.���c��S��&�Kl�k���:MW{G��]�f�OC�����e�V�bŴn3jܝ��޹{φ��^0���)A&}�#kiWxSj��]��S��*R�L��>?<0�;V���B4=��T&���h>6 B۩�_�4sd)�F{l;����^�S`8�(Z+d��6z*mv�����$��p}�6����̤��Wv����"I����q}����O�3�tP2����wfȫ�{����Qt��7�ه��(X#㻯�vl���qjb�'i�u�F����I>>���_}��ϟ]�"7��}�w�U���|�b1l�Ln�>9>��Gn=��W�08?)0*���ʌD{&��=�;?���fe�(a�ٺ6޿�\S��{���]sE�/���^A��WD۶�^��n��!��՘��EA5 ��}7�$����Q�\ףQ�j�ǋ��X���܌�E�V��8N�q�PP#WuS�s�7����l0�z�$��`��ӪBoH�+p�zmc�1s�7~����_�(�8�b��1{m��l >��H���<(��wv֫v@� ':�@�����f��}?�m&�NT/髣��r��M'������䉍�4����ųV�,�O2&���?����N>y��j�]�/�rqU�XGb֦}��B���j�&�|b���)ح�׵�x|6�^�y�� ��888X\,pRSSW���^o���*3Ѷt�.��e2��b�c�`� y�?	!���\0 3��A�m�ceh�� �7v�2��S�tA�0�\l6������탇Oa�Ѹ�c:��'�f�f������ݽ{W�B~M�uV�+$YG��
��'��0xo(X���x2�Y�#���Og��`����l�pII���K�e��4�V.s�8u�h�Ry�7�4܊F�HB=�X����g��v�����x����'��z뭝�]��D��}���ԱQ�N�P��0��uQE�F�=ł=U9�;�iQf��k�&� ڝW��8<<��Cq��*��
�g�d$�(�LǛ4�mX-低�رG4@��l�w+ƮLm�]^^�.!1&3�W�1<��L;�EU�}���?c�~2��o�-�b�3U˼���?�� �����vtt�yf���
�V����<��OiP�n���ٽ��L�v�����'&�̒3�u}uŮ�<��c+>m�56�.M=���8��p���*��G_<���ZF�/��.��f��م��qӉ]ٰ���z�˱�^�M9w��e㷽�:��<y���U	�Ao����Q��b��T9#А�UY�Q���ۆD��,BW��*��Ñ�f��X���p���\qVLgw�T=[X ��8�j���*;�y.�mٌ%�k��!��#5z,I?�1���ڙ�+�\��B������ۈ���d8H�j���<���[E�=l_NKt�m����}�Z�^��G���7���xرz���Fs���I����p���gt�j�����t���[����˙\�V��F��l6�!�8����.%�MF��+c�!�S�;��OK�ߙ��� $�f��황6Ķ;8i�Vz"�:-ș P�,�?{<�����/�����m����}� ��WpC��_�����_�'� �j����؈���� �G��E�tϷ��	�����(�SӎdvC{s2c$i�:�T��)��M��4څG����p�@|Oe���k��$�o���/��v��5N���y|q�E��RM�k��f8^�Nވ�wF�d�*��F��x�C�J�-jV'����1� ɇ�Ƴ*���놴��Ce9�zK���[.WfRP����%Q2�|�u�DEl�+��\�~�Le��f*��O��v�ݓ�&�gJ�饘UYAF��@(眲�L��+�BH�J�
���9S����7�{��]��*C�(��/����[��ɶ�k�k_�u��=�[�(J��bY�.V�Q�_��L��n�ܵ�?��#G�^��o}�[�)b�>R�&J�6��?]�,�nEZm������^���p
)BVQ̈�V�Q���j�H�?��Cm�Q���|X)3u�0���yy���s��p�PL�ݻ�Y;;�1�Z%�C��n�C��Htذ�f5�־5���w��ӓ�Ք����$C�f���|�4�0��^c�/�F!p��c���A3�[G�I
�h�X��^\�Խ�C���net�܄��ӧ/&s�vy�J�gƏ����l����v�f�����̈AjOW?|���&a��Ñ�AE��F����wvܝ;���w��=���x�Q�z"^����xcd�koڍI��&�V6�}Sưą�n#<�ΖB�
��Fg(["���?��?����gLɱk�?{a�x�7�2��,�ꫯ�d�2��W�͆m���XBbD���w6}�ΐ���;��n�j�Z����;f�9�k	fw10�['w�~�F�༂_��FTF�'���I�+�p��:����c�;�N����r͙z�i�DXA�G��q���g�?�˿��G��?u�����f+���9ң>�����o��?��:<����gO�BG����~��:8��<��\Z�[���#n�NJm]�5(F-��f�RO3���)̑�!O���M��6�&t�u>,�q���)�)^�xnW�����W_92;���߳��y:��~I�9��?�#���1��� �����Ҟ&jD�{Y_]-���h�{n
p�Yy�o�bv�O�:á�Y���HA?��֜h�$�jL9C�RS���`N���曯���%q�'O�����uF��w@�]��v�'W���T���D��������������I��c��u��6 ��}�7�t�^��ƹ�;cDK��r�Ŷ��XL�GKs��Ϟ=-K'���C�5���W>�u�X2��i�2l��gm!B���t����4-	���k��7�Il�T��wh}&^b4� �˄�����p[ԃ߾����i66��� &W���{��W??W���=#q�Ԧ���l��+h���iح��K�}��*;:pF?�t��/�I�� ��O����w�`����r�Y���	5�K����1�*>��[��k�TL;�G[޽{n�6�������r2�{ڒJq�W����=O/i���|��.6���"F�Zv�Q�8��1}]~�a?��6>���:i2]�P+���c�sp8��_�u�>��W��U64X�������o߻�������5��я����x�?z�h:��\��2M]�����B]�ӳ�Z��HU������7�ꍩ�%W�׈���޽�2�I�vg3T���}X����jr|�W��Éd����Fi6���LnV<ۡ��0G&>G霯�W����#n�ޒX-#m�e�(F�\�w��q��ɇ~�R�x(��=fW�\b+<��MV/h�{��y_I�+�L��!j�E�b�e]�K���󬌆�w-��<�lF����L`>%V��i��տ���Ƅ�f]Ҵ�~���W姟~���|��~�X�������PD��uv��vk�(���֖�#��lm�ggv��9��Ϧ����^����XQW��uL_yF�
�^7�\/5Ds[}�{�82+��Vf��T�b�kN"��&tJ���1[�j���>:c�j�V,Gxe*����͆Uǉ�[5���	���
g4iN�`]4�����i����\���\�k����A��OY�$s:��r�L�0��o�+�<��Ҝ�O>��)˛��K�97m�1r4B�����pWbGSb0�Bg��v3�����d�|�gV�m�-����.�7*_��
g�������Vx�� ��7������L�\�7=�77��JH�k����m��LEl�B�c^jH�Ї���P��d7�U��1s���GOM!���d��C/�Ԉ4`�����'��Ip@�Q�'4[�
DCޱ��9˞��^�<��'�J��%��Л<�Z��Ý�ut�{��.�8�� ��Z�;��Z"�k�)`	\^��d�R'�E\j�jwqC�G3�2_G�݉Yz�[9/+���Re<��9��eu�<O�k�T�c&3NQ²�jێãcӼ���eUQȘ���4u�H��P��G%C�� <�
�E��������ޞ��W1�]L�5����}u���� 2�MP���L���vS������������k�Og��y��3gwUt@.q��K����!Y�j�4Y3?�tzoTeJ%�9n�]TM3��Zo,9�Rr��#Iփzr4N��6" u�|�g�u���������?��g��o�p�u�������
�W;��L]mp9X�6c�,�Ю�ʵ�ͿDϗQ�!�,�%�SU�nQ�C����k�m2FJ�'*Պ,:Gg"d���F�]ҷ������c�N�8?7cG��zw�l�Z��:�2S�����ǯ����7^g6��g3��A;��I7�n���|��Ƽ)�-�3y����e_1�'�o횾�u{qqe�B��mq~����$�������
������QQ��lb�nE�����ν7�K򓟜�=b�������p�<�#�/f�EG��Q��-��]��պX\]0��M}��IКe���f�-7��x��+����~��\�Vˋ��oNw�|��DH�w�s p�%#��sf8�&`�Ml��TŃL�\��N�cˢ0�R�Hӏq�)�Y;iG�^�:�d�٬����W�n��:�۽{��Vl�,�1K���t>G����E�V,����
�)��8ί}����`s��K�ۛ�d���$�ٳv���#<�㓣o}��;w��jDP��2K�l�,��$7�K�q<�����Gv���q�RY�.���jg���uQ�u�|���gw�V����&F��d4������������
�a��b=i�.�q���U�(��|��K�$�>��Ib&�r2�n�}g:���&BG��u4��߅}l�\���D3��L����m���mSN�� ��8�����l��<��%! 42Y���O���9t>O���X�������Q6�����3����0���w����}��y5:�a���ې�jOV�����t6��4���){�&M��J,���k����F����� ��(���DP�dk��7�p̕n�tii"�px�]Pc�T�
�,jH�C��@�� �M��v7z��Z�5�L��<�Y���
U����7��Y�s�"z�i�l	,��d2���IC	g�L��%a��-�N�QA�uZ����p��
#�ą�~���1�����z��2�,/UYj��N'��աsq�9)�6��̬֬��^[
o���,�pr��"5K�B�x�2��3e��(1��|��k>qi�#�W_���ጕ/ס��!�>eβ}iؓY���w-{y}eww��r8�L^�a|�Mxk�J��ZC��܌Q���x���%�x��ڒ�@49ͣ9�aX<�5N<B4�n�2iQ�KcL�$���W��)Ɠ����'�i���?����S��-��oL�p���.K�<��`�|h<!����;K�q�e�l�"(�-b?��@�pF]�aت��}�u��Ã�������𨬩�-A��/ٷ�ܛ��Z���IZ#����x�Q�r��O<�����߿Y�V</+�w=��^V
Z��C�|N���+��KΈ��������*�Z�l��� ���p��+�����if!�	?�m{Y��'M��w󬊣'N�Ap��O���D�l<��ʀ�]�}�"2� [v��hz��6��0�#p�|�$p�}�̐<_U�Y��Aط��R�y[��p�$��\���$���X�Z^�EU$�����V?��?�䇱�������ܼ~����t���O�I��B��;G7}�Y���9-nE��q��p�2=8:Z�xdI�9Q�	n1��<1N�����"��vo\5tɥ!�ӹh�e
v��o�x�4�d�I:�\��pKj�� ���ʹ"V��U�Y�'z�a�)����.�^c0�	�2�/D�k��<����w8_$�� �Ƕ��d����^[0�5ii1��?wwwarŏ��N�Od WWx���ׁi���d�n��N�<þ��E�&�b|����#��~�
B�MJ�!��)�9R���Is�Dq��3��F+��&l/����=A������=��ܿ����g�w��޼��'ׯ�GD���擊���>��tO�@洁��G����Σ� 	km��boa7K�xNf���5����{�kSn1#DzJ�����0"�'`M3ϐT���P��6��Epp`am�,c�!"������S}�*�˳��t�*6&��L.�ȩM��	�0��Ν;�f0\��)iM�t�sB�Fv�4�y2+���B��5y)��e�C�l�<�̭M�Ra�5�tuy0��i?��Ct��h0�i����R�Go��]4����AUJ�֓�h�AE��kJ�dJx��Vhw��wU\�H�خ�y䑧�~���T/y k|wg�V��_��t�����r>���ȨH�R��0Y��t�ngw��;�\�ؖ���y�{�^��å_&�1Y�f���Kir����q��A������QO�
�O�<�2��O�:gMSل�zUۛG���o-ا�^��M)*�G3���po�0�(�y@��ՒJ�UK($��U��8��DꃳR�.W�TP�E4��A,1�R���Y��	)#ymW�)�JO�S��B���� �duy����~�̙3��J��ݡ�X�G����Y��J<S���
��Y1�~��_��*�t�ݠ3���9�̰~
��:E�`�ED�Ad�[���j�7XF�|�<p�H�xj��:��������GW;X�y�H�!�e���E�֌�a1O�.!��8Y����_��ٮB��� �2����uSq,@jmi}ҳqk���Ȥ���YI�'�.�Ft�����<� ��lJs�-��1�nb0锣>'�p_��%���RF˽f,���!��]���B眠3N���>쿢��B�^b1ו�C(�!t��8�
/�g�LԖ�q��E���8͏%*��(�Ʒ����+׆����{��Q���Z�ɋP���A�j9�����a�dQ�\pS�0���-R�[]�hP_f��\�V����?Y.�)4)�`�-I�n��2`�ǖ��Q����\ر�8�5�wv�[,��z��&���;և���Ȗ-�-
u�nU'kt���ϯ�U��� S� �j��s?Tw�ɿ�s�������d��㪘6~_~��;w�G�SO=uv{��FmQ3}�]�w�Y��i���{��L�0�i�Q��V�
:[R§��8=޺Y�䡥|�"�����d�������M�q����<զS7���X�E"�-�*�S�Y�p�ͪ���֮~���<��v��
�	u�詑�=��Z)/Dv֥p��ԕj�)�H%P�S�6���z[8����{'�hl o�`�����N/����Ga�����2�F�kd?�BXE
Y�#��>�0N�,�TL�0��"�L��zr$�2U(3>�`��Ct�D<�P6!����O����.6��g�y/N3�F�]C+&Oz�q>o"ը(�gR�R�	���������l�.[��Ar]Uz)�V�%�3œ���J�î#qy��K{v�h�;�Y	Wv�j#������ i�q�gN��^��4�U���nd�Pft��;�!��b^��4��u:]=h�;e�R�2/����oZ��l�d����s<^}���LLoH$]���PH��re�J9��b�-"r�,f__T,��~������B���Ϧ�����("���M\�b�bW0���(&����|o��ft0�n0_ Ϊ<=,fM ������XV�5[�9�T�*�/^^�Ai��-VWz�?���S�r�ukQ"���2��,��g���`B}�~��*��6��d���րT(\.�ŉ11�.�.�	�CrW����	 ������ߟ��G�~lss��k�qp�(p�P�.]B��ԫ���r7�]~�L�E��i���}����� �e8��Y�i`�.._a�� ǹf���A�6��t6gTa��Ov����
��$CpmphNOP���Kw�SIC|$���A�������|�El<|��J��P�YA��a�ʄ�JJ��(�A�9�C�g�)uz=�g*M+ǣ!���Ga��q�W�$4�Qa��U[���q~�����5�S��6�X~x��.-//��q�8����}��_]Y�����o���S��x:�v������?~�.��ٳk�j�,=�
S�ƄP����/N�_�r^���]G0�")��V����
2`��7n�I)Fv��Z(2W�?���?�$�VT���ͮI�t�G�9"�cT`��uEKX����,ս!�孷�BZ��I�'ث�0r�\g�߇qV��Jc�q�HQ��)u�1r5�ˏ���ż�G+G���p�P�
4���X	��9�c��k�hVE�T��%Ŕ��,(0z��T<�Q��ʮ�,W�B#I�F��T���]0g��o��o>��O���_��_�J��~���H��K��h(�5b�}։1�QG!��V@*C�vY�.}|����_x��08�-�,�K�ʪ{����bѦL����`f{1m8n4 m+�W���/~M4��Z�^+��

��ZrLlaJ�9�[�0�*�G��v�]^�rN����!�իW�mnݺ�s����C��8\d����3�8oo�9w�?Rf��,��r@�ڄ�Ԏ]�0�gԈ�
��m�DB)�!]��f��.�S���/��/cg��p�rj�����_���`�Φ1^s��}�p�\�Y��3���Q M��:����cJ�4u�&Oe�̪P�F\ۙ�=�}�aĸ�dmr��t�N�5���n�5�����Mq�j��m.���j��X
�l �/��(UO����<�[�����K/�t����!k[K�jy���t���/�͆
!>҃�H�V�F�a�4��G��-�O�����A��B�IY-/��2��'�E Q�.�ӌ��N�z.�#ꝭ���X���5��~��_ENw�&�����6�����\Π�����
yyt�M��� XY�"ڿv�]ܬΒ�	��x1C���(�0�h����iʿ���ac��7\����Tfql�7�Y{�m)P���T�@����a�Z����u5#ӕ�o,[D�`:M�J�P�9�|��JIe�G�UԶ��|�����i�NC�!��GQ�'R����1�Y[5j�%�KU����h��(ш�u,�����ӧH�g��ǂJܒ�q�Y��+R!#@�G�-���J ��U#r�'V'���f�03�锱�Nl��w�V�5CQ�3\��7�_�q<9�EdS��g�}vu�Vt:�����4f�N����R�L�8��:1s*<���|�u7�[D�Ѹ�-p����hM��xī��QG�mE��`wVq�H���b�o�	u����CQ��VںAGT�ٟ�G��	<�Ԭ��C��sKi�j�~5�SǨ�T��섢Hy�U�8�.}����6
�v�9�/�Ғ\�(�����\�"��V~@_��p�ܮ�^�㬦OU���A�N�k!o ۺh�pPh�g]�[$�d8u�f+�l1�)�@�u8��A��F���l��ʕ��u1�����Y�Pa4�r���B�>��|?H��FW�?^�s�
n��JM8(�A;J̞��۟\G����������Q�J�w�Իo���o}k6=<wvt���.<\�%)�Fe��w���0v!#շiQ%�tH~?���Yi�t]O�-��d�bS�Q�J(�[w��
-2ay����.�a�I�W����e�bN�������� N{��^���e ɶ�$Z$��-T��j(��X#ѥ�yO�%I�Z2�b;�vE=����u`7C�����e�vSc�h�`C��L����d3k�l?V���8uG��������k- �;�������{;EV�����q��L���m[��l//�y>O��FU\Ӏ_!��� ���YD<G�İ�'ĿO�aU�Z/6h]���΅W�1�O���&2��Aw(uDϰ���>��+WѴ?�/����&�}��o���Sv;�!VoyyY�sYۏ�f����°١�X
����>�1<]�u�f�/?���<+㻁T����3	�ȋ�B0���ܦz�"+���Wj=�6
��!#Wi�ؘ�☹-�
D&>��. i�.F&Rپ�� d����Ss���!��HQ��atg�hz4ꅞMv3/��í��7o���;D�� ws�����F`�ZP�읻��Q�����b�zeŜ
bum�}f�?���M(���0N�(��Q;�x:��Ƴ���Y4�;LnaZ�F�k����V� �@�'B�N{d枰&�Oc����Z���t��ՍNw0>��D^�m�m�w���O_����^�/��s�A�����h�K6XHF��?Z��u�;�ju���[�&��g,�6O���0�/kep\��*UP��M(��õ8���3]���T�=I`
���;�Z!��B�X�ആ�l�ʂ=dC�����I������(�7n"�����|���w��/|�_"��ҿ�ۿ��׾&A��k׮��'?q���D�����w��e������F�s]��X�+�O~�#�k�g$ZU&]�E�2�d��]7�O���M�M*�
<_�TY>�tE�O<YMZ��3�}X��Q�ήI�i�=��S	S;{�o���O<���O^�1�1#�V��v��JGMP2Y,vWVoF�Wv0�.//#��D�sl���x�ã$�]gѨ=~z퓟��g�t0N+St�E���r�1�}��)��/1-~��;�Q��tk��b�LВ�� Zǽ9����kK���WR�Y���$q�����/�3gΜ��������ڵ����w�g��h���휟@9?v�9��M5S2��YJD�����^�	�
���e8S���S��T�S���x�
��y���|ޱ]a�L���3��'=[Ǧ��#��ރ�Z�&��UG�pq�� ��d�5��Idw����!�2l>1��OD���L���|�x��[���{Pa�v9���Ϊ���r*V��������斃�ɰY���T��ND��J�V�������>=�O.r8� x���ٳg]ah5+ �	τ+Ky/mg/����'Ri�o�ˑ��R4[�"�h0��4�J)�
�xNy�4�k�p�c� ��D��yTN3�(�O�����o�?���_����W��g++�ء:�7
�c�'�2k�aG��+��0�	��Q�YN�%���o�"u�Ps6NT$(����*30R�:R�GE��Ҷ*e8@�9  'J�iF5���ݳ;��!%`:�^|�Qb�&?�����GZ��v=v'�.Lߵw�#�8qZ�I���>ϦTI���%�x�p���N��$���͍3�L��<"�|vHq�����><w��c�>�� )r��5^=I-��E�i���#o�*/PG����W%��)�l�R�W\�c���
� ��A������ۿ��^x�r�!!&b�۷o�O�|���'�xbyu�c���{����tp�PAF���0�ApY8���I�z�� '��4�e��FFs��f�c��!��[�W�������� 4��)���"�p�`lS3OmR{X��F"4i�묵D���PK�aQ��l��,r4�b�Ι~�.�mŜ�P*��cm���ˣ���/\����'>�`��h~x��� \���t��9��-�����cᾐ���g[h527�M��K���\:�q:�\���k���?��2�D��}'����#�������!ȡ�hD��m���YjC2��g��B��۪We��2G��l"�xR���lF�`��o~�/����v�/>��S�k�p�����!-�&�Y/�7��bA\|�h�����jq��%���S\���zV��
�G&c�	���rG`���pDv�F]���䑾{��A�s�RO���Q����J�`�8�d7�h��Z�%�I�d���1����x&9%�Xh�ZK��9,O�Yǻ�p.l?�1]�*5y'T�`�a:�\����jd.��I@[�`�RR�O��s�ݥ���-"��d��9-�����	7-c%M�ᨿ�����ÿ a#D�x���l6��ٕ��o��f➸�`H�܌��������i�?�+�'�\��HK�Y.��é�y��()���qL�n��9�����1lfĬf963��͛�����b����p���D^��NPn��,�B	�F��<��q:+MgX��C`��!o$
sF'������*��++�.r������A�_�>�D7��"��r(�!�lo��X�b��@�</�s2���A�4��>��d �#gsƗړ^��<��`�5kn6�]��佔�C ���!����#OM���B���ybX�H���g�% [�He�) ��L7�&5�H�4\wM�Ȼ�`��?͒�l_�-%(����i'��N��\5����V?�N��9�35�!)�RIӨ�&<���'�2K����FG�_?<c��%�,�����p�eG��iz���Ν{�sm{{��\�`��b:֢��ޚV_s1N���E����DY�lt;���6d�V����@��:�*x��?����}�?V�<yqfC '�ݏ��{��i���G���N>�y�𲚑X��|Ƃ�2b<Q<��^z	>�vwwW����Z�Ëaz���EZ_��Y?�C�ٻ����m��	׍U�ˈB�.u�Lr=x���~zc�<6���DE��x�_�m�82C�5R���݆9RSS�A/mtg�h�?���-+����+4dE��o6fo��bw�zM[�w�X�W����9���?+#*�[��ۣѐ8�9u�}��x�g�����ͫה��[t��#�H�	�X__�I�γ��M!Je�2	�kMM��q��b{�^��/�/�ʴ+���� O5�:�(�ցL6CX�v��EeRG���~�?���G̈́x�����;;s�ARJ���`0�Z5J��[�\�^©�R�Kac MnZ����qO[�}|#>���	�j%쿎t���Z�ڼ`W�0}i�Ħ���aV(����:�v�l����E�� C7�vQm'�ݔ�Pd�а��Kb�?�J�Ta}�N�0����lnR+s6U$��;����%m��U���:�i�`��;�\��(�1˴�#�Xj>d�Eֶ��T�xf�[aJ�����Qk`i��8��j�B5����ew	ǖW���Ci��������k�����
��ã�
�;�X6�l
�gZR��<M��U8_&[��G�hcc	>�lt�3�y���!�Ʊ������De��b����Q-��C��(4���0X�E���"o�[[+��YӒ�Qvɫ�I���³�R����s�=w��Y���|뭷�F���_�S���om��t5v�8l#�i7" DG���%�X'`ܶ��$y mN�O�V��zk�B_���-8�S+d�����V���HE-�b���W(]}S	�mܦ�Oe-�&�[�y��r���;j!�7���/�=J5?h���<5,���p�R?��E���Wd,��!�a��ʡ���\cW�z�D��R^�|`:Yhm�>4��_�M��eJ��5�l�Q�u�E�4��m+W�햩�Po�Uԯ}�k���g?�������ο�w��o��Y��~�H���m��.`���lU��D�hDK���^<n�w;���ב/��35㌡R9*�؎��-���[9C
�����>�<�U�Y+��=\�tE�y�1��:J=�8?ς�kC8*T��^lڛ7oN��x@x�����94��pJ�i��J�s5�.%yn�p{|5�pPzJK;�Oi�L���ז�5��q���Fr�S]�XfB�Z�E�5�W�c��=KlB��t��O��/� �葺X�꯹u�6�@����J�W�C ��o}�ӟ�4��g��ɏ
ˀ��:u
K���)S��/�mM�u7"A`Ra+��hٯtz7c��u�.<r�1F"Q�b�\iCi|,(�zv3m��45��m_wD��Nl�Y��j�-�j�<W%�+�L/U^v+��A�`p���Ν�I�,6L_o@Z+e�*rj��E-	���o��+p!�vFO7�#A{Ue"���._:����{[,-.�sǖ'�L��S�X�RJᐱ�ٹ8�L�����Zµ�5h��2�S�n�/!M��ٟa'<��/��/~;��o~��޻u�����˸��|�#�����I�YM�U#�,��Vb���T������0�W�Xu�����mm-+�Lw2)d�(�3�c�kk~��mJbY?���He�ZC��Nm�B`�A<EඛJ�O�=�0JD�"�ˢ�ƨV3dW4��:�V6�&->Z��D�a�V��\�a��f��z�O�.cB_���=�"6î�9�}��	5�m�T�*��,��Z���Eآ�aDS	�̨��T�3�v�\���~Z�w����|�z���ס�w�Z�q��%1���c/�	�ل��Sv)�E�=�'��ݮ)�gA��Y5��F����೶k�c��)d�ĵ��ͲQ-ХsU��~��)�Hq�p��)8���"1�>��c���fW�Y��4�-�+!�2A��WU7�h�Oz%���G�r!��|�#s6\gEҩ�7Zq���C��N�|�(�����9�&rQS'K�?�`�#<���%��R4���.����s�Y@��Y���Â���U�#K��d����1��S��������ߦO�� �]Y�H�d)�_�9��2�+�a�v��4bѹ7��<��gԐ�lf��ij�ނ��\Wv�|T�V6JZv�z&�����J�ݻ{ʡ��
�9X�K�?��0�:!��7��j�5z��53�ޅ&��Hbb��Z�����55)j��6��-��:1q�+�����D�h�B�� ��\&'�GQ�ɞ�t�j
=��3���Q����+�i�� �-���{V3�W�|жs,_ՔU=S��[�)�{{DzNav�D�eH<�#i�H*dWr���":*��+'ۄ[|YL�.�$]�E��7�|��ٳ�}h�F}j���z��K���9غ�ꤊ��ˈ'���(���B��ߛ�<���ʠ�|�?�#�������3ے\�v.��+�W^y���?�P��k+�T���F��)��fbI4�֜�:k�H5�O`�����!\�x����K�~!�j/��$��%6�i�^�=;-�S�����HH�Fo�Ɂ4H#�ǘ�x��uN98�r�h����Ø�E�R�1\�BXk
��NSVgJYFJ쥄h�(e�9^V�9>��L�q��T��^�I���v�8�ztk�|5|t%Z��Qzh��'pA�Ma6I}����{)WD��;7o_���˗�y/<���k�$4������ah>�ԓ[�f����[��N4O�G�t�E�\4���'���<�i<aX��f����p�v��đ�d�
K��~%�.3�l[�A�b�)�fw:�t��9H#�y�C�gΌ��/��"(�\�h-�C������P�3bD&�N���b�L't
��:����.���b^Vʘ�����<������㮮|�ee�鼞Nj��9�W{1�-��ȧܒ���JZ����BH]�I�*��ښ��0:ґ�ʚmP"~�#����N�b��\1�og^'D$��Ed�q��2G�1������t<��N2�:�2ܤi�F����Z^�Č�I��G")�d
��W ��H$`�[��]+��ӏ��TA��1@�D�1���k��D ��/�!s�2�5�E�="����Q���8&nǭ4\Q�����a.G2+��.��i�-8�\x-<��Q��9������&�����j!�'�yi����ͥ�\"����*%� ��M�"�7Ϝ9����m9��#�W�7��T������>�F{"���𛶡�}��U�{�v�j5F4��Bj_"�8���VK)����Q���4���Z͵>������Z�z�#/�>}Z����ƍ��U*��ljh��zd �?����F�EE�ܾw;K���l������F���b�'X�d9R��RjCO��"bs[S��	a"!lݱ/�\�)H�J�v#�q�z2�N�`�RlZ�%`d6���ͦ�P!�ʑy��A&�qQR�����wo=�Х�:��H�p ˬt����B,`��V������第)wh�-���ѴP���I��uΜ����z�F2�<#%����D��4�������D5�I� ZBik3;�?���3zkeR�aXHMĪT�=�UHCs�_|Ѳ�_��_����o~��_�%J�A6Z�XZY�-��fp�2$e��jI����8/��(}'��l��������&Q���/��ej�ʒ��`O8zK#+�����L�gv�?�޼y����t�1�hb�
K)'���芶`8�DK�����*A�RnH��}����Ia��?��^~��K�h>�`�m��@�d#z�Љf��7���E��aJ F0���.e>�%��9j���y+#��g����t�a8���iXfX䖤���.Eêb��+c�f.oe7"Nuk�2K� 
�4�ܶ�
LR`��ف�٢8�>���ĸ8��������?�������^Ն�V+��h��y��{OG�َԘV���h�`�2(��x���g�yf4𱐮�\1;��f�o��������3$���ҁ�zz���\ɬ	=��@� �Bs�� ����tr_z���#�ĭi"i����#sȫ��Ʃ�$������iF�����"YH��93�vE�l�h_���C�8�!�b�!j�Y��}sk���ʒ��м�>.(7T	m1�$��aH���a��6�G�a53���Gt3��QU`*�d��t�Zf����&GQ��f�w���g-����W��yp0y衇SI��عw� �D���R���4���UK�`y@<K�T*Rla%���4w[[[0�"� 8�H���J���넶�k@�R4MP;i踠�S5ٮ�P�Q��j
y��6K�e�ӵyYX슱����{U����bF˧��777�Σ<−��^����~)�9>�	�<B�;�uWXV-ʔ� ͹s��v���?²,-�g�lG� 9��Z����>�|s��wn��e��|ZŦ	�$�5t1*e��������*��JY�Y$]I\���5c(��V�9<+6�f�	;d!<�W^�r����~'<���t'كbVT����`y��WQ�H�1s'���W��3\Z^Zބ�G����[�]QT8���Щ[�+�ΰ�~j���Vw �K�v<CR��\H΀߲9���3X���2j�e���O�s�j	�(��QzY��_�������0Ґ�bS
�ɈZ��.��=e�5�Q���ɳ�������Z�BRX�:��]��a�3D�H躧�<��d���9��,��N��W3��|q4^�()��Ϫ�������B�I��j�*t�����ے��BY����i��t°�]UF�a�c3f������H �6yQ!v�� ST� �ue^����T��d��s�"�H~#�uu������2d�Rʒ	r\�"*XZy��(�BL�b���T2V��ω>�P~�<�R����ּC���<�u6��ԗҕ/O΋Z�H���8����<!y���)Dԇf��1 �t�(���	�ق�B6���֕e+"�BVP"�V߄;+��'���@�(C�����WZZU���ݻw�WiK�<���J:Q�M3�8Y����*2�|����l:���=x����=��.�צ����%�}����
��%d)q��6����D&�n�H��3�v�Q�+�����f�ͣ�t\�e�J��~��G���A�!~Gz��A�Y���Ww��s<���C ��t��k����͛�x�N9� KţN��X�Aֽ
�ь6j��	ҿ�/�>G�B��1m�:�������_��DO��<Q��@�R;E��_}�շ�~{uuU���_����_w�G#HN��E�����7�PP6+���
��-�T�Ot����{��Y��!z7x6u,Ҁ�ڶ�䖹ۨ�h]_��R�2q�Y2����?P�p�/�GC3$~7����l��i��U�d�Љ{ԩ#c�����m�|�V�:��}����=ٛR��ަ��(-�*�5v�P�;�
o�h�d��`�����?��?`�ҋK3���}��� @�6�5����>6��l.�/�۩q%z#��`�Y��l����r��M[�G�Ũ(VC��zB0����8wW��	��Yd�rz)�X8M|�O}��xR_����!PÇ<��c�/_z啫q�s#h(�K�w�d~�/�푢̬��ȑaV�Ɣ1�c8~�a��/��֍Q��D�xa
��Zߔ�b�G"'K �H�.���K2+Z����s��4C�}ri^�D�Ԭ���p!yM�ưOyj����t;���ˆ���j�P��X4�Ӫ�V1��ID7,�d��da&��]� �����EFH�/#�A^`5��m�Z�Qy�-��?-����z�gGsNE ��+ǁ+��-0�(,E2�h���˳�/�p�����;�Sr��G�Q�ծʐo^{�Ep�Pm��y��5�4ݐ�a���	���EDu.��Q&̌�ƿ�)�4��Ȥ��q"��曂M*�y������-`�l:��*�ɅI�%�9[��p�ʂ��'>��|���S�G�q���ݪ~og��Z����L��� �1����G#^��:j��Y��ų6<&[Ŝ㎣x�w��	�~�&9�����+m��M�c���� ���I�Ƈb��,�����0�#X�sY�zSx/N�d��͍0�Є^Oyn�k�Lժ���j�-��nf��ĥK��+�	�Bάjsg�Lg��&�z���E�.C����f3�v���4�i4�E��n�%Z��=V1�m4�����?�����?����������y��L���ן}���ׯg	u���F�.s����V�
.0��E�D�7�3MG5qO�Z�PP�m���Q�yr�#[��C��B$��U���H�&i�
�#�-j[�*d5��U���"�j�u��QU���6joܺI��%���C�D
�Q�kXy��2�U7�Wg�m�ů$�Z,�#�ɪܗ���'�"�YZ�KԚ��Z�"��$UN1��b�����-jU�U�����.E)LlD�(G�Yxܟ7<>\ɅU��Q�<�XHدHe���~��_��G^x�s;�?��+W��Tp��丢W�V��Q��'5����B�*v���,�	L训���^ow�+6gA+�!ܥ���zV��bǴܺJZ����N��Յ!S�X���^�����E��KѮ��+G&���	���R��y<ǡ0�ZK�ͺ[�����~Sg��.#j�"�C!�֠-��jkNƬ6M�/���e�RE�$hsa�MAK���NI�x��#�k"
3X��}�d����/�N_��'�V>��!Tn/č���+W^C`|0MA�Qk�H�輘�?u�(�	��ȼ+�!6����`c����ƩS����r�����橜,.i��2���RC���o*��IY̲u�f+Q�n4���=��Ã��!t���}`��K���T��N��&Tk�r5�ж�x"c�u���lQ�.��/x@� 7l���V/jw�G����p�tL�Ku�-�c2�O&<��X?˖�\V�7:�C<Ѩ�j`e��B/T0��9y�Lآ��l$��%�Д$�q2㼂�f�j76�������.�:��y��;�w���ݿ����
,��q J���=o���O3�U�F�L��JV@��3��S�U60ع�W�g��H�I��K���;�L�M�l���������И.�� ��v�Qka�W��bM�ɽn�sa5D�w9��������N�)�3F3���백�N�+��T��0�8he9,��OMXJ�@�h���Zc[���s��շ*���h]z��k]���nЄv#�\F4��uڊ86�%�\^�B�'�L���K0c&�<��L�&�'�b��!�ڬ����p�,���z:�7?��[�JÔ��:��s�;�9V��]D�2o����P*��&q�Z�D��/��l��R�e6�
��:��Rx+ ����RPh���Q��v�E'X˅DԷw؀�����ձ��"ܻw���s���ȭ)$E�:��ZY�\`;��$�OJh��(NP�^����*A��s��J}���v�"��L��c���ŋD�,�e��!���#��3?�>�ܩ�Gͬ=��<�ҹ�`W�o^5�9mɾ�ȓ�}�e�T�������A|��w����p<Q��`-�]h.iK]������������ar�_06�h�tDj-G��FD��J]4�Q��3E�IC&������#�m�����S���X���g��!��^�����e�����V�<�� 7�^��x�^���;7��~�c�X5A(�g���+����0?,(,������w���?��9�����e/V��1	���ŋ�|8-
MoɕI�`8Ȇ��l���ѺR8�$342�DBD��T�r0,Ew��΅�C�_y�2#�8����'�o�u�~��{{��,�"�u*�*��b��D�\l��E�G�g9�M3)te��D;�6s:�_|�3�0��k0���k�2)����J���v3�å#Q�����Y+�3��r�3�II���"�Ì��
�+�� |��w�~�r�X�����d������I7|���<s1�ۤ� +��=XK���ޡT���D�@��cCtz��2D���Pɐrdr��pc���e�P�?l [ҽ��\�s��AӠ�̢E.����ާiv�x<��.��G�4���;��1��b��w�mĲ�����9����S;�"�C�ā��i)hx�Q�h`y�������X_�a�We2ǔ�Bd����I���(����sR5�|�J�m����A��L����Ȳ�QWj
s����I��b�����":b;\S�Ȱp-Uf��d٠�S���R�E"�������iao�gS���:TOgbI~\�ٔit^����q�ގ�f�!+���������������M�f��!c��Hkeʩ$u��̺>�[D���o��1v)4��MۊD�
�]�(=�2���dՎ[8vY�mp�Ic� �� ���<��w��k���L�"����?���}<�7�����Ye]���|�(;���sǡ�eb�)����N�d23MlX�����S���q���|�8��Q�.����{@��A� ���?PP�v�Na[�����!�$sY]*E���yAB��[��2V��iHaYJr��$?��pJx�2t�q�8::����|yUr7�k���"d����(XK�`�DkR�>{�_���{�<�����y�Α/�2������Q�|qZ�JCN"f��-n�;8��Y�K���d׮,l�L#~)�u�����(�0���t�V��@� �*�ȿ&��5wa��39e8���Xj�xc��b����Gy��]d���k����|%���g�Gi�V�]�$��PO&�jW+e&�1�+a� #��&�;�{1��H�Cy��p
aay��,t��;{�"�p��q �r*��QYg�ss��D�\2�R�M�^�a�ˢ����,2u~�(l�b"
QH=��wy�l9���	2��/�������CO�O����?����Շ�����e$O]~�����_����qJ����66�	R�b0썖V(�k.��{����eI�����H�WI�}��Y0LX�(Na{a�E�	��W	��i��K�7O���oܺ!�cxo����%
x��g� LB��(��?�4G/��
�1�TxW՗8����.V��a%���=��t2ẎܥeOS��3�H�˴���|2�`��f� ��kDď�MaϙN,ۇG��.6��OoM����6K��I��"�2� Ŭ�Lg�x<��'\�q}�<�P�S��J�"�b�E1��vK�ɍ�l� �x�h�ǭYӛ.{3I��+��v�㏲؜L�,f����3[��z�"�n��֏𽧞z�0�Yt���u�t|��P��p�� WǱ}f�{ ?��S��g1;-�t�2�*I&�C>�q?��Z<��t��liK�k��#��l��"����������hd��]��b�/iS����I�`��%ʖ��Ǫ��L��f�DK�p�� o�L����,<yË��t�"AFj�����sg�ڵk�^{OJ%Βk�ݥ��b�,j�6Myl4�D���E
��p4��:����0�����M�����L�at���t;��7lf2�t������M��/�nUdU��a�:��	lYgZ-f����RB�(
�������җ�Dḧ����a�K�ϯ^����z4;�^�s�F!.�u��bÉ�lB��J<��4m*Ϊ0��hii}�@��diy�ĥǶ�����V���9��he�R_�*?`�d�'�d�Ęwq ���N$MR�P �ٖxt�D�d-�f�p���Kh���иL�Xų��D���� 4�$�Ƌh-�o�G���D� ZP��4��l�z�$:�C����eDȐ��Y�l()Yb���"�� ? &ƚ#=��*�&�4RǮ����F0�H_g��{��^���WI���(k%�u�8��q�SIYY�*�N;0��]�*���-E��>W����9k��ɷ=��}ͪXA
�(�wv�\�	G�+�X�7���y'f˃=��Dws��OV+�/=�����LA�e,����>�G�t��[�哑�b9<׌0sA����<���k_��b���-�܂���ab8���@�Q�2�k3�:ߥ2;�$�X����U
'����J]ۃ�A�����_�ŅJ��6X'�J�JJLFy��?�pS8;1�̡udZ<��0A�Ʌg#��z%;��cޢ,PH��%yfe��a��X��3-��x-֚ӏ��K��)�tefpāµP/[)>d�������JM�B��{w��X�	EE1���ٚ��;�d|8>����Ly�~w���"�<+`����H�X��V��|y��p�������w��ӛK�~�7ay�0����{�o�	:dQ�� �4G���k[
�l9�GX�b�K�I��G�Z��U6���
^F�<�X� �s��?+RvL�%��6�#�"����u���1����)��WrGhQB�Jc�o�Έ��\�Hw�����]t#�OJ�9�NE�0���Dq��Fލh�U�����-����k�Z��P9|NĒ1B	]W�%�'���<ޒ��$��ǀL����ܗ��Y=� �2~'t�}�+�al���/y�"��u]ڙN����3X!����M:`͌��p徖�ԟ*|J����ZmȂ�� ��������G�\��:c�n�ź�Q<����E�>::��f�����{��������;������8��C<��
�%����c������_n4�M|�JLboIj�!�q�L�ld'�%�J���VE�#qEe�d���J��:kɯ.(�u@��Q0ޏ�����е�a��&��ח5�Πi�`��r�YVJ%�Rh_1�+�Z�ǲ���f�~�r'&oĺ⏍.1���g��i�Q©S�����'��}�0�K�ǐ��������Uҟܨu�c�If�po�5����N���OM�+W���M:�zTUb8���Xٖ�����pı�]�=�tfjT�~��k�������Ik�dW{#�	�(�QoI[ک�,�v����{��OO�V��}�{�{�ɋ��Upl�@�Ai�1�u6՗`ѐ%��
o��^y��(֏Fx��;w�O���fB�\���y 3�Z��%���@�6�2���!�ɔ/r<�٫���z衭'�{�ﾉ�w��u\�������'�R�K�Y@����Ą��q�S.�����iQ�{>7|���'�i��K����)q��6p�e�-(��5G����E��:?�����MA.�zBمp*�$��-�	F�� E�U�Y��L����L '�1n��t4�̀��HZ����׍ꉊ�vmy�Aξ��gc�����)�ʮΝ�>�ݫ��b%�*�=�0\��QB
�8�.�i)GU�l���>�*TW��1)���E$0X�i4�j3���'��f�k�
q���ŋ�������H��x��H��Ic���H��Q�!�0{=�,p(OG�RAf�yd�?1����t1�*T*;��|ge�}Y�ML�W���D��݅G����!l_�u�D1Y	t=���)��J��ڍ7��Jq��W+|˰�w�<�knݺ���@WR!IeS�l��v��姞zwt��O�y�e>x��äZYw����T��V�5���J��.�6\����y�`�n�m����k(���E9�#�j�-ʉ�v4�҉Ϊ֨m�
��1�������$��/���W_���{^vMi��@�ݢQ��$�{{�4��a���1���>�q/���+û����wI$7�z�:+<�1w�=֌6K�q�5�5��p0��]-���u}������Y��w�ת`��l�C�������'�}����1��^xᅫW��R���ʧ>)qX��ˌ��,��e��d7�7�(�<�Q��_�z|ϤF�����z�5��=N�ه�O�eDܖ	�.��*%�l��h�ֹ+"�C�S��Ԓ�2�h{VK"��NY�k�����P�yqI��a�$.�����b�jX�1�Q�\/�����zT,qD�N���xr�%��bwN�/�tR��ݽ#��C�c�a������KMAan
"�W	)�Ǵ��&�+o�h%�2o���|0&����}x�S�V �o�5����g?�Y�Ep�x�:���~{w���L�XYKa��ꨓU4���*��w3N ��me���Y㋔�A<nn��ݛ�gc׹+���{(�{�q�u����4U~�J���@=k�H:�6�����AC2b���8����P%�)Ʋ������	e#j�?�_��%��ID�pd�}<_�*�QU)��2��"	Zg0"?�#{lި���ʨ�H�<8iԏ��dj�O�'
�Q��������O#�>u
A8��M"ѣ�~���<�[�J<�Nا�AJɈ[7�謺�"����퀳�Lq��9�.;a�t����%�1�_�HO�X��dJ��\'BV��8'4���	V��cнQce���m'���E���d�vy�:�+��~�D��?���k;8G���*^���@8C��m�C����LHV������F�YO���Vu:ˈ��ꊧԬ-�.c�gQ��l
D������I�`��d4mMӷ�Yx[yJJHY*�Xҍ�M��8ʼd���~�G�/�Y����)Bዌ�S�X�(Y���zzF�ۍ7�\Y������N�WVV4��c�4r2v�!w���$�873�R#�d�F�z���?��tOw�"��$n��X�:h�M�[$}�#� ��B�áo�J�	�TK-��;,��Ta\��M�<�g�QfKiǳ�����NM�#�N<5HH?P��yeͅ'^�~�nB�7�o�9�1[)�H*J��Z�]�d��^
��!��5Ǯ|���Y���(Z6�e��F���8%������N��Ҋ�����"w񰖵)?�?݀�Vwf��r�j�nYd}��y�òa�~^��5���VJ�J�tA�4��������� �`�d�O�?�����wv�ڼ��M:��P��5�^�b��Z]%�u���w=�����x&�+ѭ"�V�|�kX� 7��Í�*K�4?jʆ�T��$��3���L6kd�-ˡ��lv��m|���Uʮ��__]�E�\+�4t���+P��h�Ż2t�J��R��;�����nІjZU��T�Wl�� _�� �CV*�ÑƱ�4�p���q�X��$9[��gG�ӂ����CЎ߻v�N���>dwwW�:N��BmhB���55�&����Hq+l�x�P��,��� ����ZK�:�Q6�_�#���`��������F��h��A��[��p��?���;��엖G<t(F���6J��'!���8ʐ{����w��!���!����3ń��;8�X����Ξ�:s�a���|�&B���:�Rk��!ͭj��c|��~C�ǿ[�h��p�k:��T����p�3�:����< 9cVE����-~H�i��)��N�|�ZE��h)��	M-�Wʂ!?m�OM��*c9�f�X�H�cF3��ޚ�X0Cb���5��XO������922��=�dl�޾}��K���	��=x�759XC�<�#����buy�̙��Sk[�7.]��~�#��}����.��,��gz��J֚6B"dz�l--�kW��HFj%N���Ї����߻;nnmn8y���|�ꃝ]D�ao���'�����׵�n�֛��� �T}o�4��.<��
:��d��r8�<7�N�g
Y�f�*C�G�6�f��fn�tM�,ZkP+�����rxH��4a��l�7 ����ɜٔtZ�[�@)��$��J�_����V�.������q�MV�/����<���E����'Re���駞z
���W^9�<�MY��۰�F�k�j;A(��H�z*!ڲ*�޽�r�^�#�@�C�N��G���ʣ�(,5kg�xq��O+�n�ƑCzAk+�� pB�q*͆0c�	'�P/$jq�ҳ�E��"�%#�c¤ln=�:�k�n޼cϩ���)3���)�{���7)RT���e�5�"=����t�7FK,RkEC��2�D�cjڢ�|�2	{��0�="׸�v���{k)rDzI*_
�ӱ�8�:A�d��h��V�^tZα윊dr�ͮy_:z`ɬ�����Ba#z��Vu7�a7���Ԍk		�����?�������ރ?�яv �IJ؝��׺�/�_YYrm�H�����OӣY$�<#E5��Cb��Ҿ���^Ydt�9�8H��"�K�v��W)ѿ�<�D/h_9R[D��d^"L�ʧ��u�hG+-o6�|:�.���k_�җ�r��=�l�X����V�{ꚣ: � ��d {�Pq��E�|mu�%����O�����">؟�����9������Zc�ԛ�L����S9L�,�qa�p󫊮 ajb��a`�=I�S|�:�4�_���o�{���������s�c�i���5k�y�S��|�F;�{K]9˜F)fD��`���O�nj ���BTJvi����0�Z�Z�u0~�Η�H�7�]�ҹ��z���]̣0��q�a�.h$m4��H)\��)a:R/6k^���Kʉ�1]N/�E��-;�����R�n���~���{���߻wsmezp@+���gUq>��X�@4.�R�r���rA|l��U&ʛŨ��\���y�$��kT���a�P��G�QA��Q3^��|2s,���I^#�!_Vn��f����)��`�J�<)TJ�-g0\��h6[����[�a�|��{v���o}�?��O\���k�ݘ_�1��+XE������k%��42>�꼤�� �2Sij�_/�j�f���pm}�)�u�3%�{���?�R:�X�P�h�+5�'���ɃF����j�PF��=9���Mc��I(j-�^fu��88"Ff\�t!�B��>�O�Z%0�,��{�J��7Մ
�G�k(�"1�Y�w��B��O?9�3-셖0XyV�	|�yez^�c5���Ne�ّ`I�]�ó,��i'�׀�Ԧڈ�/���[
��券�ӂxG!�O~���_��3�<�C�x+ϸm���]]]={v���[��O����'D�F9`g�F:�V.��+% S����wX�2��|�*�F�ip�xQ���(8qB3�ң#N�����)<��P��<�e�;�6t�W���U���ce�T�ZzQ�����if��m���i���[XK�l�l�	Rw��'��'�}2M�~�Q��v�啑��Ei2�Mg㉖M5��N���f�u_{�]��f{��\�t���V/�CS��%��X�?�b7� ������~�e�|�����3�E���琱���}+	��!Y���]�0��z�`��:9�tkq�B�2��
�A�ŋ���{�1Ċ�˥��ٳg%#��,Ȯ0f�7%�۽u�b�A����	bi�Tx�`6��6a�N�Ĝm���(��~o�T�ôL�r!�(5=E��z�$�J�z������T�ɟ��eʯj ��hy[G��wE�)�b[�%%�����AR�/<q�:�öBZ��-=DK��s��1�o?��F_Q�A����mK�j�w�w��qE�"��L!v�W>�����Y��oM?������n1�F.O&Vrl˶7n(U(�D���9bC��D�7��7��Muq
LW�~��%e���E=�F�3^*�/~I`�)3�Yqm/]<���Օ�u�ct
�m���v\ߕ|<��P.r=���H�� �P�t����s0���aMcZ��q�r}d
RQI�T�+�GPJ��A.��c-c���>k�E�(���J���i�4"|~>'��c�l�0Qp�YՁ5�o� ����h�9{Z+�M!ڔߴX_�T�-��2�|�2���HK�H��kӾ� ��6�4�yS�=Y�+��tCm��kŎ`!�v8(�nb��E4�����lx�3�ڬ`vB�P�Y Ae�6��;���8����[l�ԎN!�����Mh6�e~j�^%����|%�̬F�ն�f��nllln��VGc��W���B�Y�0t�E����,^`=�����ra���Rv>,!�&��Y(V�4��X�Eݚ�}<�� $�c���=˟��M���k�zua�g^�������ɿ�]�O��$�����_}�'������V�l�(95�R�����b���/���u8�����+ĺ�~AF)�6xZ���g�N�Um|�6��Fe�����\pk=�����.��8Ab�$#���#���u���t=�����?���5<8��b�*�_�0av73�����-�ַ%Kr�FTq(U�&��
��Y���P{�E��I�m��茶��_����J�.E'�Po����ˏ*�"oK��%01�5|��X��x��"�����[o��I�S�W~D$�6�U	��J!�,)�ƣ��w{����2.�*��ؾ�
~L�!YpE�wqU����Z�i�~}�����1�lM��*�0I�2�,O���ǉ�zå�
���'��G�=W��F�Ϫj�<�Ǎcq^E~�'��x����e��]�؝0�ܸqc*r�!�y�[Iqŀ�<��TM��y:5�qL!L�{�陼�)��=�\i�g��>\�Ѓ�=7�2�*�nT�L[/�<�裸}�w�	/���������`�=}RHz� ]�����������,ͮ�N����*���Μf�3�4�,�-,�-�� �7�U�MR�(�"�!G=��ΡbW|9�|�=�k�uΩ�t��p��������Q��*���]]V~��iŵ���@�0ǖ�%��'��i]���	��CCX%|6ױ��	���������Ŝ��;�+��?�'�������8lz�Jq-+ZVr�
�!�#!�^f��)B�	ŕ2�4��m���n��*фG�*�q֦�6�We�c=�K�X��$���(j�;� Ds��Y5NT����
z���:�&��0 �����k׮e�����tBbs���&�5���������ʫo��B������O	F(�P�(�a�y:U��Z:u0|zzf1�q�eF����6�W��*|{������D3^����*�'�;6�Y�X�,��Ј�	��2

���5Z���g6��ܹsx���`
��r�8w�"�E�[Q��8�5<��q��&0X�^�L�����l�xh�ѡ2zXfcG��H�d�e/G�zE"�aoL*Q�W#�4j-���	�2o%Z�s|���!�୷����w>�����3|&� 46��wgˬG����Om�L������6�m2e�����y`1OPb����*t%�Zf��� 44A&��!V�[�]t0k�{֪җ�$�J��L���ٳ��O��X����vu�X��_4Kh�9m��p���Ԭ�{��c���j7=z����c�6w�e{���O����)f��B�-�gd.R�:&Zv�5��ƉLV��y����.M�Xg����6�vr��l�F��u���+�n+S��0IZ���K�=������?o�z�#t������I���?�z��=ł5LV���E�('��2�"��vvv�D$���:�H��ͦ �;K2�)~Z��Jx�\�H(��(5��A�ÜC����3.�^x����'�!;���.��O���cLa�^ܞ{��9Z>�?�G�U�j�ڀ87!0S���M���@8#p@|�f�rc��ȑ9��D��:{M|�W]�X�������z:I��ߣ�mL���{��
�~)�x�U�q�������7n�l#��{μ\Z[Rp�?a��XXo��"V��њq
�H	���<ePZ����nߛ>y�����:��N����I+*+������o�2�[/�]+W������r�T��V4Qy!�Nxm7��2b��&��S6�2�鴗�g�\�X�!�2O�)�X��f.�^Y��������x�U==9&������鴞W"����p�E��@h�i��2�޼�F����uv|���/��+;�i5s�֟��*^f_��/8�`�J�d���������dpZ^��ܼy3+�H0X��^�#vz:�DT��4�����Г�N0�\�"tց��5��Y���x�CH���R5Fi�\Rbf7��Ղԡ���]��Q����b}9���G�V��jt$�O��Oy��mfdp��!G�3��±	0+x�݃r:AB���S�N�
%SX��-f^����I<����XvĭJy5�t�S���y�6Z�V��J�6ժL�W�Xf����2/7���L��黚�k�cX�,ɍ���Ȯ�ݟ�i5T7��;�9�$
�������� � �T�Նa4�'b�I�	d�p�C7m�:l�1N�E�k�9#�W�"����$��J %�ϡ����g�h�,��_��kzOiD,?��IAub�,�����Z�d��G�i
�sx�N�N�jA��S����G�⸗�,+Q�� �k3%shN��Y�;��,��\yC���&oJ�PgE*�V��r��--���b���[m�
u�H�kc�M���p�I �5��i�d�W3�K��$�귕����W��,m��W���<��W�ryU����R7Y��OI.ދ�vu�];�����s�,Ϙ?�nw�[D�;�St :K܅�I��ml��O
���k�t�Sa�jCV������N�
��_�^6o��v+�H�w����󃼊j0�QT��_z� k�Y�J�~1�st��ɓ�>��������xd��D6���z.=�Ã��4�{��tJD�x�,!SoIV�:��Մ�Î���{��+�B�ꀹ��Z�UE��GΒ�y�\����̈�/wU�Oi^�йf����5���luR?�jupa���ؙ��t�V�W��|��_|���h��������q�U/��uwO^1}��W
��!��_�o�=7,����"ɱ�D7�
�EEn���mei0R�G�����rN�;0Y$�naeu�k���N�W׀2M3w6Ǯ�|�(h�`x;���,��K�a�_�/�_����S��T�K˫P[���ˁ1�?z�n�t��0��ޤt�[�*����戱E�
�&���q���J�)�Đ�J���)������������v:���l�s��)4kk�0f�$�؛�|�;�M7���Jѿ����;�l��P0�lD����t�'_�$rR��p�N��XZZY�/�j���8lll���������>۷��xF_��:����)Vײx�����B���F�&i�V��N9��c��ֽ��h���G���dDؚ�d}��w��ß�ӄo����?8<��#E�7���l�ӧ�������c�[�޻���ɓ'�����2����]$�6������0	ϕ� ���$�0��+�4c_�!th��]/��f���dN�D�,ۂ�N��l���
7��CY�̄�1�k�.syP`~^8�^w�h~1�#��%�u�pYf���r�)Ĝr8�s"�-ҥy�[~׉��ɎN������o���a�~����H�T�D;�̨&6wH���<}��Y2����u�snb��_�v�-ZyƾH�o�9��Z�[�+�5���`��p�f�Ԩ�!�hȐ j�<脰ՀC���q���l��a�+VMm6#�t<g}c�N����$h��j����c��awVW�ᔝ�Bf��s�O��O�y��.8L��8��#��\縊���e6�cI���'�03)����6���YQ�Q2}j��J67����������ܹG&��C"���{x��s���U`�R��&��M�oyV�!-R,�#�����P�f�_�+�޾�����u����>��Ν��b�ȹ�~�G�Z!�^�6"�<~��ln.����f#,�NG�8�X}-T�=<�g�4ϖ�W[d�ب�Xr"q �J�J��fs����\���������@�#u���Fa�����Y�G��~�����_}��c��Y�`������"~N��@����~�擏��ɳ�u����j�SI�:'�x��Nj^h�ZY�0"KR@YBA�c���,Ƀ���(���`0<#+%eղ~����L��(4��#���!���� �Y6�a�����՚�H���Uړt�^�co�Va��<��$~��`����������}��\��N��g2��|�����xb�d�����R���k"=@ 0��d� F�on�cc'��)�����Fd}�f��.���b�$�����&6�y�Zb]hv�B9[d�x)���v��1`���,k6�zr�c��?�ɯ�گA ~�����]|�?�p8��X��D߶��cyu�)�fh����H�ي��WڍM�>�A���[�,���4�Љj�E��&4��,�`y`1�=y��2��;F�v�x6�A��b>Đ��k h'+'����z�]�j�<K�DF�ID��]\"hl�L���t��eD+�g����u���̨j��Ym5�
dԑ����֖��j@��i���󈉜Nƾ�d���g��ȒG�1�h�r\�xL����&t/|f]�	�ׅc����)8�A��"���d�/���W�"���Xk!ޗ9�^�j���9�vwo>�u��k�����t�Ɂ�v���m����	�A�Ǝ�7�F���U,�s�'6��c��<x���0@��}��;�($�|���Rə�n�r�!�B�R��X�U�����害����0F"95.�*�b՝D��!X�h9C0�W�C���sr:��5	�	�o�I2����̞��p�Kc����3lLl���ɻoh,���\ؼ�$�=t����!��W���#�b�$-�B�`����b����ʲ����,B4��;��
�҆�>9�:���C��#p�Gc����.�#�}cop�]��@\��Oҵ��PH0�PӪ��U��쓏?���N5˥�n<��т��|��ؠ��_^�A��<y��O�>�E��lnl���k?��_����'����G	����4[���Lg�po��P�3\�h�,����U���'jM+G:��!�zV���kX{w�2]��1�P#6�{��	J�
C��?�6n�;��B���Am��͓,1��Xx�np�R�̧p�P�l�1K��{Մ�,��kF��(,�pD}�=��a��#,]�9��;��^�P�i���y�[�nA�2m��<��J1�$%Gn��ک��e�i�(��> �l0�'�Y��m]pL{F�l6���`�l=�t[˫+�A���d�}	���~wI�0m��[;{� �F���JRm@C��:%>��[�R�K��,TzW+�[Ok��7+�(�/[��[6f3��p�!
�eB�y�4���@7�j�a���,2���2�e�������A��l��;cW[Tc�T��]&	�� �y6�GC� ?�\�x��˗/�C666���7�C�pZ,,J�"Z ��+�����W.��r+���sqz~��7*X⍃�r|�����f�7�	!����+2e�-!bI�r\���3����K�%��l��S�2'�0F^���;�aooo:}V�I��H��ʙ^�z��#ț%�N���O�f԰���>���ՋK+͟}���m�g��ӓCr\�7����C�SUOs�'�h�On�z]Z���考�-Ɉ ��1������Ζ�a=�2�Ps�j ��h���#��ܗ�\n51��a���(���UJ�מ��5Y&TՎ9�O>���ݻ��+W��k/�,�f( �|nSF�_|��waEx9���fp����%��6�g����߂U����<y��ǩg�KL���L����/���-�/�X]ӋU���:<�g{�D�u�{�m^^�۴PE��x��e��e��9�,�*5�U�V��,�/جD�ݑ�U+�Kg9]7eX_�p�&�������R�D��.1�Y=���8[�}:Po�/$D�3�/�]��K��6�!�k�n��:��իW������Jی-�-��y���w�}7�vg����<����|#��K85e�@�����fE�B�\Q��3��Tj�TF���+���������X�r{{׹��e]6���F�~�����NER&�$�5���*MF��._#���Ȟr��R^���dP��������vwu^L΅?r*���b��� ����pVdԍT�EB?s�jg] <G�Bs����ׯ����A�YbB���_ڪ�5�9ƴ��g0���?7�&�i(U�71�S�%Ԃgc�N��&�F�V5`ܾ�帉��.�F}^��e'K��Ç�S��8����i�GH�#�,�$E��˪%���O�K iQ��	� 7�d��G�z�Sf���?k�xJ��+��X����C�lff����� ,�AINⲃ�X�F�7j��&�7�x��ן<��h�,���t���o�qΜ����>}����+���x���XJC7�vFX� �^ɢ]���KZТ��hՆm�s(��{��ƚ��o���|�mcb"�n����4�D��Y��%��&S�Q�,�8�,�X�/��}a��)H�p�+�����������
FG�[�,�eF�A�V�
z4ָj�����H�:a�:bw����1�t=mR��d ����a��@:������xv~3�|�u���l�Δ����"l�r2��OjE�Ttf�IR�z�PA�B�,���'b�YE��J^�K��rFjN0)6Z-���<�����<30=c�`��f�u��%�GH�M��s��={�z����K��/spp��z��p��|�%��ȬYU6e�-RVV4�j��c[�`J��xi��n)RQ����@$ո�~���CT0w����_�,��!�ejxd׭8���E��J�V�G��)2���O��U�/���������	�
�����������h����#�b|�s��*DZ�8��*Q��<��%����j���(�b=W�Lu���T�Ws���T7�K=��v¼�r����:Qg����*�9���Z��ꫯB��l}��=��ız�c��Y|+a�gǜ,����'�}�D����H��TJ���^4N����@�!:�2�uzm;��xK��*C��p�4�M��Q<7.��\cQ��]jfPT��?�HȬIa��"��1�ZZ����0�쐾�˯�����4���UG!nS`m��Db�`=3�N�kK����~/���̒��66��w��Y��RJ
~d���x��	�Ps�կ7����l�������4"�����gϞ�F�fM�U@�z��?�|�@�T�.��b|�NsK��ܦT�עt�����̟�JXƈ�_�F��MB����)�&ZN�w��%4c�5�_ȶ��nV.��l��O5fں�"�_�/���I�����7�����1����g�?N̢�з����ԑn��qJNUZ�9��l���:�Q�(ϊ���}�WA���d�� �p!��"^����4B�+o��k�)�`�P	����E	�8��Tъ1|)ob�N V%�2^yvj���r�"�ᴱ�A�Ճ4A��
���%5=��?
���j��!@@�(L��/�^��W4J�v�f�3^�Am+u��VTK]���:�{9B�_z(�WI.���%�-[+�L擼����W��k���x�S�ENLc��z�7��� �Ў#�;��W3�d�N��+�M]�S����Hvͳ���6�a�BYo)��*��'�ԓ�n1�/��P��ډHm��&�n��mZ����9ICƟ���Q��{��3��{R+�Y�`���h5�BG�C�O���;����A�j���(N_V܇W�"�'d�	hpS�W�t�d�>$N#���p�硕�#���v[��3}���cѫ���%U����K��H&&�S�(37x�wmu�Ш2-�#�[�'+�	�c��7�����ٕ��e��d�~r�޽�����"j݀��_��L�;���_l�}S�{(�#��6��C��nsD���Q�2�x��1$��2�EaK�`fs2G�jw�p��%��¿8��)��-N�Z9<x�¸�G?��F�� :�B\��j�
R�;w�]�Mr�Γ�P{�����waݦ.��o�/�N�����n��)� ��_f3^t�d_B��`uqWH&!�yټv��j �e~�$�ˉ���Cǳ�:������]������6|��2b��6�|�4cR�c�<b}�o>�7��o�zi��F��(zK���N��w�w�<��O>��l��G�+'--D�Ml6}e��1�����>.�q�8ny���Nŋ,EV�(zy�t��̞9%J�[�XQ�W����XT�b�r�(�����zK�V�� I�|k}��˗/>x��οo�@j��:t#���e���2)k��SP5����8z=��Ə+�XI�[���J����a��� 2s�P��̩45�IhC�X�_y�S(n��P��Y�x��(��^������!)~����|�0p������s緸�a���G����_�4��g1<܂[�n�Q�����������1�-�`0��9nI^l�d>��l���ī�-�Ncg{2:���yN�"���N�<;۾��������v�V�X�����=�;��j����:6�	W{|�ސ�`�T˕m��'�z6כ��vy�n�z�f�՜j�E�Bӫ��I�p�"� zWɜ�1=�
'\�"�ú�}���������]��",ijY�}O��zv=��!����	�MB��9>�lf@K����j��������E�o�wZ9	n�aY&#� 'x��������ϟ7���_�E�6NX�
r�F�ks���^h�ˀ�60�w���
��LF\j�?u�^�u��4������׉�n?���/������f������7�����-ìL
�֨j�K;����o���ꜝ�zA?�8�����٬��q `�vp��vCm����}W�_>�5����4)K�_��-[�����}����^)��"�v���4�h8���z���qڶ6ׇ���V��5E�̌�������	�`OR~��&���$s�$U� ���X�^(C��B�e%M�suT����hE+�K~�|�6��:LˎFS���A��8�	�+��!^�lo��`���ŋ�l�s�^�X'U�y.rhƜ�t�{	G�ښ����i>"��ͥ�������[׿����]����[�˫+�#ϟ��)Nc��iD������H3=����iC�g��Pc9aɑ8E�/8o0�tz���s�x1���/]����
Gpows0�;�m�w�u0-g�2���M�zY�y	8Cu�		[0 ����t'=e���2yĚ��`IW#�ޯ�K ؜�g��ZZ�v높t�!�Kr��ژ���.-l����4y#�?�жyE�מM�P8�A��l��1��G��^�|��Wn�y!�Q��p7��`�?y4O(�p�a>y�����88<��ب���"���^�v:z@V�L$�,9'�3i�l�s8��3���g��W	AA�7�������_e�N�^��*i��1��v��Ba�V�
չ��W��S��<'.���2_��4�u�B�B��%|��,i�i�K~��ッq�ִ2�e<w��[o��x���"a���"ĖSrS�6"o}m	�lF�@E�=�ƻ���`��~ee:j8�FdA"����Kc��Sva���,�b`Y ��;O��\,"�Σ���^��c[[��B�O.6w����>,�mKGj<��~�I����_|y���7N�Oq�f�1��l6:V�q���+����J��SQȴM�e�AS��C�����p�8��믾��x!6w�ѓ����t�a���'�QL��X������ƃ8��J�c�=��Y<��]�<���d��a��#�U߈�Z\g�3N����Ӟyki��x17�1y�����:�����r
G9���V�2�H�rì�MuH��AmD#�H�4W�^�u�?͓!��xx��C�q�+��g��i���Sk.aN��������4�[�ȭϙ�j���W9��H��9��b�@���iA�ej�+,�`8L�aA+���lY�#D#Q��nݾy��+�_|�f�F�ji�}���a��,�U���%����a�H<�"�-�ܹ�^���:���d%^���4�.���5����c�遠h~V�_s��M�p7�2��^6�Nl=�Jۍ���-�$��[�蔝\l�T��������x���C�Xۄ�.K�to�jGiB[��d�#t��P0�$t�'�$*9��[#���_mP�lw���6䪂8�D	s�q���#��� r�E ����[��z�7V67�h84�H��,��7L d��;>d,.#�T5�r8�����!�zYH
B��]���4✙A��f�hM>���x����#�ó�c�'���,6�G7_}}ccK��8;gg'�n�\_������� |2���h���&̑-�%���6�Pad愂��T!$^ŹTT��e��,��r���0�p_��^[��/�h"bb�l
K��߰{�t/�Ž��yR�7��|�bȐ�ԃ�C]��1!OӬ�?��c1ᴾr��+W
�yT�O����{C�6����gRcm�Zhb��a~}�vҕ#*��P:y9�"w��,��ha�i�=mSj�v��r��� 
C 8�Q�y������\^'G�{����x��UP�)tUB����р�1���rfkpv�Bo�z���S��i<��O�M�Gt�,���N��_F���:I9��^�d6��Q���Բ^e��*��|>��lZ�A��j��vG��H�0����)#�81�BS�u�s�	v�	�������o5�u�&|�\�$B�lq2�P��<��6��d��������/��rww5��~�駿������Y��n6-����[���) ly�k��iՈ���9<�5���2�jZ�ۅoA�l��=j�y��#��-|��GJf�N�;�Ѥ6X�$aB�&2��I�,�#��NVU"/5,d��ť�i�3�@g3���g����'4��#�������c�VPM��3�
�1�uG뀿NG�Qln��e�����e�|��2`�_���t:�(�x6W���l�-��e���x4 )��k;X<(H9�'��)`/3�Ks��3�r�j��{)XU�~)���?�)��o]�?�o_D�
��z���|�u���U|U���`�8R�y�TH�����������s�(�ȬN�t|���{�ƍ��"�J�F�Ö+��Da�0>�j�Izc�y� z��֝�|�I}<ܒdī��Z^D�k�w���	X���lф9i���$�ha�r�E�ZV��^5RU��]V��r � -n�iT�ڄ_��^ɗ�Hj�Ia�D��Z�RC(d�ƪՊ,qN��l�s��-H*���b�)�1�O����T	{���H�p�ty�����su�ʈ�]�,��;����q�����GGpjIGE��0_ӪIph���r"V�J�+=Cz�V��+nQ�UQ�6!�ҩ��s��/�<�m�"܄P�_?>"����+�~�������ϐx��ѣG�I(��+�5����!L��02n��M6�q����f����%=x�@���m�J,-��ɽ{�zP�"%E���S�\q.�f�zN}��Wfm,{��7�5�ZԔ7xV�0>)�1F�������n�����0����0���M�Ј�i�d�	�N�����)	�f���]�v"ۀw={�u��U���b1 hBM8q�z������!��/��/ON�����h���HCKQW��V��pQ2-�d��g_L��F�}�b́Z[���o~}�1^����YZ�a��
2����ׯ�&������w���O>�'�?a7I�j���UD��#�3k�Af��ܬvʒ&6�&���8k%���q0S/�ol�d�p8�ſ�W�'���y��9��v߲$�]^�Vɝu�ֽ��G� �-�ɤ��?���`��B��\35PK|Bc�-�:�`��C�X�7n]���l\π���ų�LƊH����f�)K;AE��e��M_/�PX�ѐ.���緶�^{�&������g�!!r��b-�	�|D_�9D�N������hF�<r��ܥ6�����_}��g��Ǫ�l˩bo�FS�2����X �q`�',,�|���Q"�5��S���&�R�6��bE\��}����<����@,X�`U�Ν;���'�MA���u����S��}c<QkC���������l�O�m1'&é���'O� �4Wu���LRd�a!?�ݞ�Z�.����Ÿ
&��D��0S��p���=)����8�fd�A�u���������MZ��� '�m	6B�8m�=���ݎE��<�:�ԍ���J��ē�ϦS������.��޽{�=4��k�!��Ѱ��؃��X��[
��J��,+�Z
����.e���i�ۉ�Jc�������L�w�m	�͛7��~oc{�0�;>'��*�SF�)l֣�{��+B�Df�T2�H6�����q.��~��"��\��9H�1��O���BZN��k{�����YE�3�i�M��1�1� ����I!O�&�b���cq�y��K��&��3t�0�L9U�Z��mO�y	a�*H [�{�K~�+OMl�y�$��T8%mK��F!qS�������gX�o��cA��/>?-�$��s;A0d)^�&Jy� etHB�'Tʟe��M�e�Y�I�j��9&cX��[M��\[Y���Z���]��o�߳�2s�m΋�i�&��*�Hh�}@����];��`)��6"f�t��X`w��B!��3���O����8ګ6q�����R=fW �&����f8�te�̻�[��֑
�����?{6���Kj�B�(�Jy�GaHa���a��A���Щ��[��T.��0��x0�n�h��N3�����z��%��0v��h�c�R=���g*ȗ$d>ˌM��73��=`m�!��m��Ji4pJ@��#c��#/���͖�99:1KQ��Tnv�'u�Hv\Z��E�GN�$��;<�0��E���&�EP��)���qz6ßԧ�[b�~ng8 �����͆�>��^���\ I��0�bS����OU[3�͌���j#{�RTO�(X[� ��K��A�$���mI^�Kk��R�c������S�}�s��Ǧ�;=R|���'���9��(�]���s�����Ɋ�
���o�ܕ�c��|]騬�s�維NY�H��VXG�� ���9�>�;ۄ�|Qn�5[xu�A���D���+��4 �#�ь5��Z�T��5�~Φ��feu	V���M��vͳF�-��$�R��U����Z����6��\URسt�SM��ar�u��i��o5"��"������dL�dجو��h8W�M;eشyR�-Wߋ�7�=�?�E��X� �X<���b�������,��h
����[kZ��J��\3�?e�U�NV�#�A�[uJ��3��H�B��`��Er��PA�vsZ�����*uٙ���H�|�@�Gƛ~oݪ���81�:;˚�-%��O^���X�| fE67Ձ�A%�����"�&���=F�(��XÔ�F��M+m�-�+-��W�9�bV�2���K�x��:��K���è6��;�Tb��裏�W��T�����s�\{֧��@�)	Q6��/xP���
")'��`1i�	9qZ������.I��DC���
��T�FԉA8#:b��o���N`�#;]b^l�%]��� �h��w����ׅq��b�x�X�m���#&�76��7����[��F�ts�R����թ	�k"e���TR�ƹ�kj/�o����&���] f�dJΪ린	~���l�._��z����0��wp��{G�w��[i#�7<�9J~a�[M<�^���D�n�D�,,�TC=\<�X�TDU�T r�fC����W�P���9|��&鮲\3Xr�a̓��i{��>_̮\���i�$�+א(@6r�d��<���'g�/fw2�K�>y��dG��h���g�͛��v.����g����w��ĺw�����J*_G ����}u[m���2��a�1�<����s�A�q�[:�W�CY��㎧���g{��>���}�sʕ�|t���/�	�FX���|�b�%�?�>��� �Z^��$?Ɍ~"�B���é�za�V�V��tp�:��n7�#0���1�(�x�4�s�=�a���[A��씽�073�/�FGш����`�t���p��.e���)���^��d؊�XZ7����OÀ}'��ՍU?\K�dns�O�������ɲT�+��9�"�67�ϟ��������k���v��Nw��B�o`O��鐝�%�Wo����؝��S�}�ϗVVieS�߰::Y�)lM1�o�I��V`���g��.��έ6�˺�V��hZ8MS�WG?����M[Ͷ�x"qN�
N1<;�:�%�_yNme�',�pΝ�INFN��8��sZ�p�{�6���p'��؉�&ϳ��ib[�Q?K��_�6�[Xi%�v��������oΆ\I�EH������#;�^]Z��M�f�B�Ϥ�Ec�ۇ��`����얓%�	e����2� �7Mb�9A�9ˤ����&�-&��2����qFc�(��˽�Q�,�C���F�nD���m,��;_,u�}�K��v'h����ذ����	�N�K�.���2'��T��mk����dVZ�\bS�"1��[��=�e�jw&é2���x:����"�P����*�����/b�)��3�v'��W���+�^��1T,y�rg5�����Z2�ワ����)L?cie	��la�șB c�ub;�|:���7^�R�C�w�ƭ�ʊc�9NZ\�x�܅���Cc�R�Ǒ�C&FQ�R{D�Ujs���bBD��]�v�ƍ�k�%=:>D�;����r=z��(79��Z��OΆ��$������{�y�ٱ�~�s"h��(NpaG������"�)Ǭ+d���������3eYk=�
F	4��|�;����ݏ~��<8:��?��Ǐ��ni@�������y>m�Ʃ��2dC4�'��a�k�E� ��g��gSO+����o�0�:���<y�D-�p�ݶ��f���@,ҵ+�{��Sd�37nG��Q��K���ۅO��܉>���M�F-�
�Μ�M�x8䜻$N�6�7��9\�ͦ�����t|�[�����׮]:��@�����ot�(ǡc��Ɋ�$>]XSDB���{���+�ݾ�k򩕸����������Y����rO��<��f�������3���S`�lm��?`�O�m���m��}����RE��'�d��lSZ���믿���ϼ8j�x6����'�⒞=�G���/X4�K�a�'�F%��Fx�X��7�A�����"�79�aD�E����{���o�D��jNx㾂�6�����;)2V+���rڭpO������
e�m�CT:����J=��Y'ZS�PV�v�C�f����Bx9�`ds��]w�n��
�j�78�������ׯ����z0ɁdcEݜl��x6�_ȉ��nN���8�?�䳯n�vcyi�s(��g�}���f�������~�_<{~D�`�u�~�2�]�+Z��;E����X�t�����]''"[K�þ�w2�&qK5C7��Ҏ�d#�(K�#�z�gǩ�қDǏbr���\�����-���w�<~fՔu��,�w��O������hc���'"j;��,X�!c\��g%%�ǌ�[�|, �FW�%�>���h�`�e�l�P��@p���im9������.n����%��kr4��rp�ڊ!o�>����8�)4*�޻w������Ӵ������t��u�b��uw�����_��%��#u�_����9�0��0L�Z��  ��IDATn��k�*
R���e)��>��wacC�����!a��7铏?U�'�[ˎ1'0P���L��glqśaؒr��������ϧ3��0����ee���D�@�u?�0��n�lx]�A�fyFˁb�G����F�%i1sJx��7�����������%gɲYt��O�DHB[\�R]�I��jxe�im���r��:hYZ�Q����yMg�R+��ް��bwW�+T�kջ�����/b0��n����a�/^�p�еLt��qrx����ei��7��-��WV&�����j~�Ѱa�;Og����,ۖ���n��xj��с~�h=�k��X!	��,�+(:vSd�!�7�1$.�̱5�N��DGUL��YD�����_��ٷ�iK�����ރ� �����um����!tF��(��(��CN��S|R#jI/�T�ی��݄Y�I𰿬��pH��p-�/��+Vt[�&����'d����S��#������zM��"�<�%�ʙ3���P�����9/�H�h�c3�8�A�$�ĈN���o�����\_o2'fоQ�5Ч'�8��̺���pFz�����y��Lb�~�c�O�$�+���<K���l�n�K����I��=���o_�rC<`�<x�{ϟ?�޺Pp���l8�/�^/��F�V��>|�λo0�kq١����J���v;�x4p��!K��2G!\����!l��I��S����Bv��C�1�ji~׼��I3#?ȭ���%���YH�L����T�V�'^��60{д� O�$6+�L>4bV��j֫T���ҹs�T�w�G]�s_B�N�p���{?��>}�c�T#��dKu������{��}��}B|�$VV�8�(�*\̕�׈��*�y��^��q���bN.M����ոɷ���!�;y�J(��SIY��&d������#/\����߂
#p��Մ��N����ll��\�"/�%򅃹�{���+PE$���ԩ]o�W�9�j$�}���s��W&.+�ODl��A�������"���G/�R8�f�XH�H*�mHu�P-�uV+p�׻{��q����*��rI�m��cV�r�i޾�YfZ-܏cn;�J���aUkr+:�y�e<�rNPT'�+X�y����C�{����S]�	A��E�8>:�*!�&ɷ�`;N�'Ɋ�/q��է<v���3�:��ؠ��t\�>t#�`Upл`���@Ob�t��E�6��p��`Ȝ;^ƙVf*b�oZvF\G=R/�_ezY�1W�RQ�[���O��=@�6�MNN&#sIi��\s]��km*�s��i��@��-_ޕ�ש��RDIE���y�MӋ���u��r��y�I$�X?��'! �?���v7�W"�Ļ��Q�B�����-�gr�ǵ�+)�pyb��` ���'?`��ۤHG���R�rL�f\l���Y@�]��z�V�S�m\�K�2k�ilB���W�`+<W�_��~�����/_<琰�h�+�f$�U�	���O��o�2��Z����)�Q[ް)�Pb�3�Z2�M-���j@!���{>R��+|!n�$�̂��Q�1{n�E��%�~-�6u� M@����A(N��!���ʛ`a6ᤦK�.]�v��i^3�!�{ǐ��[�.����r3;,����Y�臷_br�	@��& ��Syɜ���iK�z�iSpN���*>�Er{X�:�%��JHEf`����%~�䄤�G'<�i��i9M� �4x��UEwƖد�����w*8D�
�ZK8uVV^{�5��`0�)e%tB#׷|FPЫt�
��d8���]�UPI�l�Sv��L�X��7U��S"YR{��_����I��U�k���Nz*\.���#�Y�+���%|Nʸ�:\d��ggg���s�����2�����������G��2�8�y�&oz��W8A�+,ͩ��2UD���boמ�o,�d����q��>�t6�Am"ԏc< ���`��w�1����G2j�|j��K��j&�1���&�qem.V��<�L�\U�g%�'N�+��WUߝ�Y�C�!��E��h�6������S��4[X��J�⭋�ۋ�;}�Vduְ$ɂz����r)�ܒz�y������ v���BP��:�	��τ㎳,M)g��2���/���+4b�	�
"�������;�� K��ӓc\s�-�Ii�~k�٣�q(����:�(���?-sՌ.�I����zUg�����.�txX;x�J��MI�غ�6p�re�g�qhɣ���-]�S�[�ϣө��F3�/.��k��T^=Qv�{����N�g�0l?��������e�킗��'_�j��k�w�~�w
�~�r�-���s���Օ-���މUF�G���onloo�yyww��O?�o_��8��Ϝq�N�Y�ty�������[U����#L�q���Lg���sq�<��H?`+w��C���bV�e��+Oo޹s�lx�{T���%J����WR�v
J��ؐs	?�j3�����Wɩ���\XR8
<�ote�M�G��c!������7��uL��z�S_�?����m�lɁ\����x����o���`@ڒ���[o���[�ol��Ƈ��Ǌ��jЄU�}�+(%�`%U�x"^3�{�^��9|��0L�ĕ{�#��C#��SƧmm,�[s�#>zG�P��zf ���ֳ�p�����C��Y��&+C��F/� ç��`<�	��(�T�T����jz��O[������M2;���+��T9�i�hR�eT}� h�T�жP���֪�j���i�Bl-�2mc�{�H�oiC�Ij��+jE݅�L�a]G5'��܅�S�q~Gg�ҷ�0��)�-ㅌ��:w:��u�.�u�X�m����)�e�e^k+��v��*9�lޗ�K;��c�J�}��\/9W�C�?T�+�Y;)���L�-��z5$6E�q(�U�[X�w�x���VI�ǆϋG4̓�Sh�yүn�_a��ƓX�u,2$��pF���S��|��?���m(d��v�)~�#���ͷґ[O��j�v���ܛ(���%�S^3�ܫx9�
�9���`��-DUK�y8-�_�җ:�A��s;`�v�F�.:~�9�d/}AwV��j7�}is_E9=O�
#Ȇ����[?:ƙ��i��5ϳ$���q����p`E�Q�$�pj�3�JDТ~	ߊ�Q������)�n��_jA��P�8�x�D]�=�/F\�T�:�����@��T󈝿�E0�N��*�o�*�H���ƺ��>��i\r�K��͆8���M�[q+�z_���Ff��|��'���������6Nt���������9<8�����?��M���� �s�;�������w��ޯ]�~U]�KN	�)l"���憹�N,��htu�ϼy1{�C6�{����ڷm��[,��DU��W�^��-ס�
��6��5�:�������F�N>�u���z�	�X��X�7D��g���V���d*�TC���[eI^�����HI���H����^����ƴs)7��h8{�g\��;�˝ϛV�14H�[�yr����)+*I������6*��$�d2����������v/_��^ɦ���o�����Š��cc���x|��}�w�ӳ��T�NAZu7�u;rb8�e��!Mx��s�3C�T�9�a�{��!�v��..^�����<{��Q�k��'1ƾ�)�����+��;�DQ�9/��t��X�˸1+(�S��T�Z�ڭ�mS�6T�&ؚfSdX.��9sa|�ⓗ�0����*�X6ӹ���/s��j�XQOn)*����a�Y�m%o����?�/H��˘rJ��$��,��Q�T�z2F:��vfT|��&i<G�i�NS�V۲��BH,b��vۭ�C�w�6�$���<��ľ'TxN�?�����O���~�h��l(;B���
!�ܠ�xa�ߵsd��wӪ���r7'B�):�Y�&8E�ܻ��U�9�$|���<�!Ξ��U_h�*�Z�����k�����^5�ޛ�q��V�ݾjxD���O�/,W o���8�Ά�3�ۇ�����u�-|!�l?�!/�)��t2����5�6= .R���։��R��K%N�i`���P��a�hQ���>�{��{�h��%�k�����f�����N׏�T;k�;:�F��*ʸ��i�V�(-�R�TU���ֆ_�}��׃Ql�i��^��+7��l���������>g���xucss��~�����^�qu�8�h����?{�X\�����r>�:n��308;�cA���~�?��E����R�����CU�
5��$�ݴ�Q�I�������b&��F����?b�%���y�4�~����X}n[ޡx ��M��X���h���GPR�Q�H��O?y�w�z��Ғ!�3=4�$4<�]���8x74���9�����8/x'����|ee>44
|����bp|p�	�,rgccey}�u4b�t�(H��¹�( }��0�G�5�]/�L�>'>�d2J1,�2G�op|��j<'�I6�&�$]���\a_Wf+�s�D��~�姧gG�.]�O�ʕ+�^����Uh�V�_�?��pȞ?;�c|A�0�U�޿ar�%�.���z@��AP}+�(ȃ3�I�쳻��1Ӊ]��eI������"�;�h<�@����۲,,�&S���`��pn���_]��t����2?k�qlDe+ql�b��F##�@c h���������M�s�"����ŹH������S��w:�#�<�(�^!\<���P����d��t�½1s@���I&��tn�IFt��j:��ML�1G+:q�qW���}�W�Ddޮ��9����'w6�i���MgSQQ6�r���I�.��1����ssi`۽���^Y^�>}��awwW�Jv@��2کHej��3��5��%���E_�k���"��>��Q8p�ͯ�ez4XRm��Y��T���~����N~@�����:nt+j��]�WxsV�j��,�JI����}��t�h�u�gD�QIwګ+D�E^qv��������\e�7t�xH;p����F�(�f��l�fn�!]D��U��E���yĞ>?XZ���mw��f����8t>�GG�����s:�����Wob�����l�ャ#��Z\P�p�΋����W7��egsjf��g����&ں�Q8ƲM�#�V�`V=�k�V{:�������z_~����P/��謬����'Y���_��ʥ�מ>}�q��]Nx�?���~�T��� Zԅ�p��@�1J�Y���;�6b1]$o
�o�;�1�{7k�V 8;����Ni������s��˟�9��~b�hU3H]�+H8|6{��4wY����� ޾u�������>�럨�z�wO;��T<y띷�7֡����cI��hpzz�ωg��	�Y�ݤ�&�^��ѳ��R
��B�6�W>��K8O�Ԧ3��a@ @�Jb��k2��H7��u�+69g����YI���Oh�l��e�2�d���$��0�3��Ɣ<Xl�T��g�ܠm�/\8w���7�|S���1Mgf�Fp��޽k�dj��A_?lw�)���`OsΖ�$�rY`P%uH^��`�<�����;�0+FP!Vp�yD��Ya�����j����q�қr��˂oJ>w'%8�4�tR����hF@���@��j%*�Xcq[Y]�Ϭ�4��P�%&	\#h�n�p:mL&����������j�S�F%(M^ƕ<�~���^�ą7g8zYn�l�>���d��%������F��Gx�*��v�;5�Ba��<��BG#�)�,]���^�hf9{�"��tqr�{��ScP��*!�2HN�#�z��-�/����2�nT u,��7�6�=��&���v��W��u�����.�x�楇[1Ϗ�%�hVbl��`dTr�&L�wx*��iu�o�z�h�KY�����Xa2Ę���PA�PDJ�
<h���(����T	h���z��mz6[	��֪�c���)W�F�%�=�d�0ӽ�c�l���n��Ր��s�ˌ����1�i��� ^� �E]�r�V�f�������/�x�aI׷��Vל�8�B���]��m��gb~k��R���[Va7� ����f;&i5u�h�k�7޼� e��!pf�aLL7��3Q�%J��B�-���Xv?��������PA'RzCr�*w��f�>�����F��:�)EV�4�Zy��0�Jo��T����y`=Ͳ`�Q��ƂWì�l��RH$v9|����LBSH�ؑ55L4�K����Ν;<6�1A6��f����N��W��ox��w/_�\�|���fi�-o۴d��(�˨��U,H���D	���c��o{)�~	�W�o�>�ٛ��/����
X��t��e���ꫯ�`�Nu����Pp�3ý��wե��"e������DЈ��B��(�T<�vO���HK9f��)�]�e�A������\��YXr�HA��5�Gs��V�����8:�A�Xp�T:n:h�O.��j�-�Da_�p,�!�&�p�8��:�%�ʶ�`�XT�Ģ��
q1+tR^����VC.����J��}�jaItk">0�.��~uބ�g�xQN�6� y	s���q�UK�l�%�����(�f÷D�So:��l<�֘WN>���UCN�:
^�E7�êP��|@&8�FQ��N�ɭV�*9(yk�&��5����\��;M��4�r5Ħ{�e�{�������vt�
�r���ki�7�2�*�.!G��c����� 
���+׮]��?U��I@��ʣh��"ƿ��ǐ9��ݠ�h[;;�2XY�2>��VCŏ�"�-�;8ڗ�� �o��V�<�o��M���3�SU�^��1B%dN���o�����Q5F\e=�?V��_Ϊ�wY�挛�>�����ڂ:Bp�g�g��ʭ����7�6��x.�5,���/��B5	�4�Dر�]^�%N����͈v��xU�Qɺ(�'k�I����tlej��t&
*[F���	��nFh�I2L��[1|�X��dU�%b�x����R����om�3<8�n�z���|��+�(��a��Jw<�k�[��M�7_}y:��D�r[E;�c�x�xj�rd������,�P��ґ��_f��mp���?t�Tl��bO���>~"��)ň
`��APr �F�昆�����c���\��d t35$*�i�+�w����I�q&j��G�7����7�q	�|��0���Tu��hY��j�Tm�40�C	��o��l����t}eW���9�������/!
\C�l2BGO/D0MX��t�8E�B������E4��\���D+PC�U_Y��g�ւ����E����/����!	/^�G9^��������d�WX\{�RT� ;�L/��$��n`k��$~x%]\ң�����5�!2˾�04�#�3�\���o���?�~庥2U�z�pv{�q=�%���n��Qӟ��b�Q�[�Ss�����߫:Mȏ6a�i� K�ǅ8D�?Ƃ����I�I�8��XX���)�u�8�6�O���C}Z��L9�9�)"��.��P/6�B�T��glWlGğ��6j��@!RS�\Ve� �%�Z#�t��8)����'����fp�y�}(��ׯ�Xݾ}�38=�����cz��d�h�Q���j ���QWd�KU�2Y�4#}���7��ӣ��Aԁ'+�+81G?���i`�����`�t�o�7o޼p�BS����z6���4v�nś�Z'�,�<m]�Zyn��ǒ"�;�%޿���Sx����_e\mN�X�a��)g2�Uk���
��
ݩ'�d�9���4�
l>��ý����!�r��|b���k�U�.�Y#	mzu�:�����xt���:�͜����Z���@w'�;�<I�7���%i��B)\[� ����h0���i���c�.ǤzW^y����;�������o�	��8ܠ��5���]YO��F`�(�¢�4�M9���H<��`%�V�5�4d�"�h����r���X��͸2iٲ#	��@��s����?��|�"�/Ue�+�A���/�<�� s�NHI�_}#V�ZO\5BO_��B�39[�6eEo���p���6���G�S8*�I,?�N�g�����MOZ�7d�ʥu����~C�1�c���VIl>���k��o�Z=D�Df�G��y2�H|���������Q��M&��x!�����3qaf2�Ø���f5�F��6�p^�R�F�'�1o����8[�/-u�[�df����o��\��ߏ.��dOu"�
�V��N�n	|�UKfU:�NV�Uۭ��"��Rrt�_����D�D�s�X+�C�3�<���S��lFx��SN	=��w�j�Ȕ��n#Tt����ׯ���T����!�oʭ\��h�Xf�!Ǌ`+�� 7�f��ޛ-M���t�����:ܻN;/�۹��_)Rś�1���P�)���R�u4jm}���Q��nc}N.��Q���[�tϦ�F�����123(����p+�Z�8V�$u1aS�#��WE�(JqiKƼiy�*���˼d^��׽+���uJ�[GЕ�#y%���Y�,�,��Ĕ��Zo+���s��+U�������,��E�=�<���.�2�a�\2���#}�4��*A2<A�馊nOJRګW>�L�(h`e6|��P�����>�ի�o4���vØ=X�x��!�`<R��P�T��%���a<!��W�������|���y��Zg����7M?�mA���F���8g���6�2�/7��_��Ad�r��ˏ|9V�c]5R�0�y���n��l�Y2�'U�&V���/`����<��Y���/���\xQ��{�K���D�tX6�=²r`���[��M�e��j����Xd��x�kS�rh��ٳ݋O��z����~}���W��K�^�ń��(�����@�2�j.S������&d �j7Z�gS�t������%UGP�6�O��f��Q)���3Bt	_^��+ly�u�5co��gϪ�\8�NQ�-,v��eI�`��c$<�?�H������>G?bA��x��Uc#j�O�E��~u������zF���N����{�����=5�4�c����~����F;M�G�C�c�]�����S[ސ�I�y�h�x8�@����㳓�'s·� D��&ǶΞ�&՗�K ?��)�/u;]���0A�y��Uh
�A����	
<\PC�2/[A�����t�O>��"����z�&���J��Ý2��9�
U@���D5[�ڊf(v8�p8�_l�2?��'*�~E�I��(�ŚQ@�r@f��̃�����mgT���g����q�m����>l�V����3��3�B1�e1�a��u�%���`��S��*��9=՞
��]�)V��m����	�M��F>�k����W��d�Y,~��_?;>���,c�Q6 ����n��T�E*o��<�x��d`Ɯ�o�z���������7?���!/��àO�5��=�I��!kG�v˽�.t��� �<�vp��&|�4�JϚ��]�0 �E�L�)�ʚ�J��������9܌�n��i�7��������J�d��O����4p��^{�7�#��*o�u�9������=�¾Np�&@)A��X<���X>����Ǐ��gx���N�#�=d��9���i2��4��-f�i��xњ ����j���/�8�U�0E�t���E��~(<#�f�t���X��w}�7XB��u��7��H��+�\,$��p�ţ�҃�z=�NAf���G/�`�%���vQ�?��{4�D�B���[�|��
'>��D	����]y����lC�^�u<$����,���Z�dcSFlg���k�\���Uʠ�"��V�	��ȭ����ӫ��s�ǂ�� v�@L�	��5���$�5�/���jG��S'sFE�ߛ�۟/ף�p0�Џ���%O�/�J��`�?����?����Q��;_��Z�?�>����������>��O~rz�&6���B5v�0�,W�d:2�����V��������ǫ�c��J^�ܼ	��&� 3�CM_��d�������vY#�{�Q��hs2�!��9���乓>��O+/פ.�nnlCJ�ܔ�-���E�P7Q�Vin��x���י)�"�"g�q�`��7�7Ϟ?����~�)�9��y�P���[�9�pM�F3���I"&���a	��,��q�sD�g�o~NV�r��"��X��G�)@N�̞,���bJ��w0��@X�(��L�xl�&��N�?<8��y�\�
��O�9k� �JnVf�G���|�ܔ�U�W��Mrϱ�.��C{d%ia�b5�-pR�J�0��)q��ՉqjҬ��A�dŧ!uh���,������lx�(i��,�@���ᕦJ�Ra���q���#���12��x�d�)�|�GQ�|�Z|�Iw����#��^�����6[�UYOۓ�^��&��7mn�����ξ��@Z��,��V�
;?c8�K�Y"�Íjx#Q��#"�������m�n�3}͎����	P9��HS��������������	�.;x���P��9�2&�n�S"Q+�i�F�������1}D�b��ټ~/pl3Z.``�W��y���4��4�l��8�v6���яRVb�8ͅ�����	�L�7�f ���^l��bA��#.\��흳��b��^�L�>y~
WH�[bF6�,Y�\/�#��=_L{N�r�6.��F�.�OV�j��BOpX��1�(.���;���p�z��D³Qy�Zfi�O6����{�̏&5�Ъ�uG�{��{�0�����,'�z���,�e�C�0��
FQg2�`��p?+h.W�<��x���Kv��8����	�{2�����m��=7Iv�:�]!'���G��8uMJ�*�\�	#?}��j.]�UYL�a�˅��FC���$�9zMX?�����G}KZ������V�T$h��M湎}�k*��ll�p$E&�,�����n����J����q~~���#ش�l���dW��j0I"����n��J��	�-�u�����8���-�M� �2i8Mx�4B�H�JV&�B.�+���p����kO�\�5fE9鲢�.�~xtt�-w���I^���*�I$�9����m&�������5.�|w6'k�Rc%YoӶ/Ըp��[w�����?��xv���Y��(�5�K"�=�#$ג��AU�k�h[����:x$��Ѯ�`�P k�a ��������_�u�?X(���e��1I{o��_M�>}:��+�Ƴ�dj{}J6���7~qy%�?��`�ƴ�<y�������xGq��B����:N:�B�oxήY5�}�V�������>�qb(�� ���L�U�r�U��T^å�J�q� ��d7cI�Rf�˺���!vO���O�����?�C�q�D;����.J�e�P�F�n{}5�	�_�N�� �\ە��z���I\2qnR&��8��+�w!~K��/�.�_�ڜ�-F��*���5���4�����
+��e��r3�V{{{�k�^�%9�Z���-��(y���6���V<��!
�&h� "�Z��|����Y�n�MY0;�묹&�a4M�vW$֌�����G���h�l��No�4�lCb{f����V�2n���:��{���筷�����D5��ѵ��I��-�h��!�H�
m$i�BK\�
OO:��O��$�[愚��vV�ˡw;ҵ����Ԡ��K���3�5sd��/���j-�|�Z4�ii]�3ʖ�K M�g�l��z���Tk	?>�B�F*d����!"a���_���]�{]ي�'���5�����ֻ�7�����Xe���x;����q��.c�!�v�d������ql�0�XV����!h����/���9���w߮���B
���^�N�r�1s|[r�t��:"�_1G�����/��PH��!W^Kv���õ$��ue(�J_9oY�LN�w;� � ­�P����+W���B�#/Z�.�)t�B�V�ʗ#V�� \���ZR����@���@�&{�縊�q^����	4sxq͋/����ͮ��}����!�����a>�D������U���y��	�Y����p�C>�#*�(Yq���C� �?&#��a����ԜE(�e5N*��]"�$�� ?{��-�lP.&�Z�cUF9Ԓ�b��D�IK�9)\��b��
�q ����d�0�&qy��׍�R�����0���vt]6��k����%����B��"N�~9�-��� #���������I�ӣ	n��U;nғ�o�����	׫IsG�-Z��,h�^��ׯ_D���A�դQ�r��J=y}��]h������v�v:� &Ew��*�J�)s+������-GC!��4>}z�����yˍ��--�=�3[�BU��j��);�olt�a23�G�:�j�Kı��s��.	�����z#A��_��c�^G�%������h8�Ge�d�T^Uxb7�h�b } ��[ic/!o�p������N�������ؤx�%'���������RN�RV�K�6���Ľ�@�`MBY<I���M�Q?moQ4�-8�[����ńl�Ҭ����>��|���w�}���ot��)fA)&wD'-�tz)�����R��
�y-bLv�]O��
x��(2Zϗ>F%=w^;�T��᪂1�n6�b��@�j)���Ǐ�|M�e�Rc��J#B���l:�`i"xO���Z�dc~�ϟୱ84˗� 
x҂���Smѱl�"��7��>�H��/��u�/��V��/��)�T�*=���8�=Ay�k�b�N�vV��w����F�2r���B��^�r�Ng�$�4D\�\�A�?�L5���:��	�#�����>1.��o�V�����	$h�gZ�\����)�E����p*4����?�*^��D@�Z�.j���o�����+HAZ�j�Ք����;��i�����a���1ʘ%t"�䰨�!9}Id������5�8�@T���A]0V�-u,�D��K��2��B��;/E�v �Wx��Y�M�%�[����J=	_0�����@I�͋�DMMr�6���=~;*'��}��]�L���Ta�2V�������X�)�!J�J�"'�����߿���v�y<ݜ�f&��bs֢��8���j:�n���"2|�� �VC��}��g�<J
��y��{��ޭ[��>d�I�m, "���]���Y�xi�^�w]�7������9��{��1����{�T��l��<�������1H���+I����v܎!+,�h�&��]P���U��NO]k\�F��-$��_�"}��R˴�2��8�<!�F��_լ��%�k�s"��a�� IF�o��6r�툘�Yo[w��8��H�Ӹܮ��ka�`*��K�!DF�����S��H���ϼ#�b�uƲMm���#�C72 �	�1ދJ5� O��m9'����=��Ė/
�~�l$!��LD)�ǫ�q��?�h�sQz��ZE���;;Lx��R����u)y�G����[�-���P��Fj6�6)��/�˴�F�qk]2����S64%��Ufե���� �lq��Y��\�/��:���!����A��B*j�5�����G�Ե����a�u�H{e>��38C����gZP��
d���{�Dz��qF0	�Eo�IO����I���q��:ʇC^����k1�]sv�������hw"��#L�ʪ�:�֜r�%�PB\H0�}W� Dl�Ӯd�ux}�(��I�%S�_Q�i��ˋa�9JKj
����\8ز�-�ވ��ɉ�V<ݥʆD�=IKZ��ֽ�1��ܘ���Xi�+�̈��E+�+������8�s�ӋѶsU%OeQ6~+�׈���\AC�#u��j)�	S#��?W��vwZ҂��5ӷo�~뭷��z��r����WbW������kl=<<x��"���A^�~b+�N�8�!�n��%��Fℨ'��5��P=M�68�	����T�������h_�~#�'���}k���o#��qD.���5�3�J�,��mM6��Yi>�&:�l�����\�6+F��I�l-�x.�W��s�v�Sf|5�Z���	����xIMwv��&��f!��r�q�_�l������し�
S4��陜	a;)_�OF-I����7n`#t�� ���'GtB�)�-�~Q�����ڵk�ZL�h@�O��z_��VlX�,�|���laFC+N7KA�:F����Jյ�*���)+��%�\!��
ګ۝��[wM����I/�7o����C�.!cD�gl��������w�Ԉ#c��_����q����o�	�����?<�.��Oh�8(F��٘S5W"`�f�EȐ�a�h�,y�V�8��������B]��+�n�Z�N8W��R��A�]Ú8�AF�83���W���4A&��g�{�̰!�߸q=#�Đ���dg�.��N��OP���]��;;h���]��UK�ɍ�����'����t�
�r���1Day����@�>��On4�r#/��Ng���4��ʌF��ƴ�V��E����\����ԉ2�����/>GD�C���;i^<~z�9�5��ƓM�rdb����k"�Z�fp�:��B=�;�^��2Bx�D�[Kת��5�Vm��q�	qfsօ ��GJ��hJc�->�,$l�|I�G�Z:�_�Y���+|�5����pYC�H�'8j�'Q���V$���~<�4"8kNB��ׯCO��+�b���S����K�u$�bN���#��v����J6W���Y-Y��N�R�8n�r*	I�sW1w�JK�Oc�a�����;%j�^�u�[�dY�!reI�z%.5�'�l��b1�v \���ş�ٟ�Q�LM�u�޵cN����k8�7��O?z�ZF���^K�Cv�U�<~��7�9�LX��j9ȯ��Rz"��T� Օ�g�!��4��u��}d:QG� H�&�%ը�MO�z��l|롼9]� K�^ϳ��+q����`��p�pL�(��>���{{���[��v���C�������7М���9�_�%�޷w���'�z��lS$\oH>������¯�h�\�)�:��V%+��T���\���Ě{a��tvv	�̻��d5y�J����5��°����(<e�1�fK�	�P�-�![�M��,G�]#�W�[f��l��@"�"�;؎�j�N����+X�j���bT���4Y1m^\�b�ЧOv92e��X1s �U�{$�H/�3ܠw��̒�!�E�Lx,��,��MzH�l�����%�O����������8�&�׫��M�q�W�/�z�YHH�$T�k8]JN�	ۑ���{������j����01�;�ׄ�����G�_?>>���o��*��� &�jRW���8�8J8I��&�L~���$���;)$v �J"�>}�ඬNOϽ�`��T�Z;�Yt�p�C��B��x�X�z��Х��`��㱹9���n�����Zj��wS(��4�^����J#�n:��������q�|�����o��&﫯��w��'���ԕ��6m�	AiW�Wg4�$cUf����wY���V�Z挝�Ӹ4�#A[�Ӆ`���3V/n	����/��/$_P�{PI���燚���z1d�� �/5ǖϧJW'0���D9���=����~{�h�xF^Y<[��/�l��%<N�+smVБ�̂�D3�yκ���N;�K2�$���u�>|R)���jR����"$��`8J�$���B/s^Դj�t�b������/����J��$��s{4@8�	E�W�{�d�-+'&o߂b)e0=�#��%m�l���`KO��XB�Q���T��oz��5.���tƢ�SUڎ���Oq�a�7�6��SA���/����g_|�9vR�2i,{��m�ϫ����-�x,��Χ�7l:�����:�����Y� -���!�ۙ��x���vW���nh����f�3S+zR���N�3B��`+ÕZ�;>���=$9d�v>]\]L>8~�����"��f�@���ں����e.���+ݲW7�jԹ&�:DVZ�����8&3L��ɐ���z&����֟UR�,���b_�po{���t�x�0�Ր]1��iz|,�I�@A��A�0������{�ݰ�bʌ2v�ل�x+��:���'?[&Z��i~b[��4�7r����
ޱQ��?)u�:}$��B�̤ڕ�I�gl$J
����b9ݞ�p����ƴ��ŕ&zċ�j���ᔸy�9^HR����b�����VY�P���P����$�MmRޖ�K�Z�Ln��?���ޓK��B2����p��}�-ۖ�J�"ڂ�q��[4��A�-Ke7�1��;.\k��9{,�Zj���3[�R��P5ծA�4�\
����'YL9�T��<G�����p�=�sj�_��TzGM ��g��J�%gy�z�W��⩆��5�2�fQ}x��<՞�3Щ�����+�R}��#�;Ќ�(@��4�Ҽ�F
��K��Y�c�~Q�� �n��u��	<)a{w�"�e�p-M���M�zV�H�5��HR;:=���P��5��vQ���ݯ�Zj��l�x)��P"u�.�)�ak���f����#�^F������X�� /����ݸ�B+p��E'Ж��t��Z���@]�~�d���>z�w� �R�#�q����d� �YAf�ԩe<�Cl��ä�V��S]K�z~0"6�[�����K�#(+��u8!���M�������M5�M�l�po�W����kD*��q}�HP�YN�f�y.�����qqِ�_����4'�����[R�䠞(�A*6<�Ze&DL� &{sk��G�0"0Ӓ |�*-�^����4}~�S��t�N�#��֠�酤T�V�	M���qUZtź�����xH'�骔Cd{��?Tp�â���q
Y�k)-Z��=zb�ϲ����Z��OX�^]2B$��.�z@�[S=jXG��"5e\N=�����_�x&S�Um6y�$�e�9Ӭ�iXMV����(C��h��f��'��'���c����t2�ʮ̈́}RV�+l���u�SSQ:�Y_���
B���ҋ|��W��}�G��c>5Z�8{i��G����PG@BV��ڠ$v���UՊ�fֻ�&���x{��R���RRюnЅ�p1��(�&��iQ��fav����j�h� ���2N���믗�+��K��5�'��%zԭ��6-=�O*�%lYp�ke�꫿^��1��P�S�
�g3vR$H�Q�9�̇�n�썶�n��t)vH����؞@
�|1���uit*�,VA�+�������k�E�jh�Q+�0�ܠ��\�^*�ٗw�U�<==�b�b�(�?���_q��"uY�F���;ۦt�5u<�?����GM���Ń^���<�_~�(Z��G� ��0e
��DC�@�܁x�����BדQpf���De����κ<��8tsG=R]@��;w,�E�I�R��,صkG����w���V:�W	�l���R-J�l�.�>�*gM����e�Ϣf^�/��Q%�ԃ��,k^~�� �@��/t��!�I/��D�,E��l�<b��R3��ذ��
��l��X�q��o�a��j�>X���K��b����������Z1,d�/\JI�V4T��\�$2�[vS<$����)��rٖrP��=)q��~{J�&��h�yu55^�)�Em�2���&�ڣ֤��K"�H=���Π,&A,Ļ����D��aqNN��C�GcW�Uq��/Y���+��#M�Æ�sn� Vi�U6�h�S%A��tJ�^-�!�?	�d5Cc���Б�^��K����ɠ�b�V����
ԕ;2���L��h��7������b:ة�%��R��.B�50Pd�F�>y�������c���5��S���vS.Ȧݯ
?��}�Z����{B��둩�,S}�\�YN�&�FU��ٙ�M�+�K��ц�ł׮�*���]l�`��¶�@�;�ǁM��I$7�^�T�F�r�jG�{�����o���O�x7o��*iF��k�?����p���\h�O����E�i'*�����H�%�'[���c�}�R>����<�/Ma�4(C�ʒݎ�I(���U�(}%��h�B�Ttׯ_ד9��Ν��gD}.e��ZG��.3�ȹ)�6S���5<��dRt$��O��?~�������=i�Jz���J1ʈ��>$�)�L��z$5��^g��X�ED���)X6kF~�+���Q�1���7ߴ���#�Y���j�ԃ��Q\Foh���	 � �ђ�-�>,�k��>�Ov��"M���qp�����8���D
���tkgt��@U�p�D���X ��l�%ǿJ�g-�B��]�P�8ѐ�۷�(��V\� áF�c�������-x�vd={p	t����3�^7���3iO���^��[�%�tؒ,���{8���nƉ��-�on�į���$�n������Rjv�8=��lY3����A5[J���_B�=}JH���3�Z���T=j�@�7D�T�	o:�'���6pipe%�Z�~���Q��ݦ�T� q8���5� e�J!��@���y�P��G-��Ԕ�B�XI�������:Wh<×_���ݾ�Y�q]j�3yXe	Cg��ޱ��T!`�_񦆄�L��F��~@�&�)��9�['e�u�MZ��P��%-h�����{���e]��C�`��$}_�*/�c^g�ϻ���0��U��cW2�5&�����^�!���(Oڜ��ܵig�3)�y�(^n�T�*�Hj���ɜ0w6���/�3��� 4d����̊b�d�@U$������u�)|�KJ�I8�4�T�/[�L�."�5���]Թ��K�'_�.�]N]w|�g�f��<���Y��-U�Oh~X�$�]������T�%vi�R�$b2!�F^AO:���!i�`6]�W��f8nޯ��Q����:��a���<����5帤芙���첝ϩ�kӢ�C�iߡ2����E�G�y��|�?�;�y�ظ�F|�O>A��������/��4H�\�e�a��|	 ��~�o�ls���\>��{��)��ƹ�K<cՒ�Q�&I�J��p&П� ���%NI���?|X]}K��D\-�R�e���7I(�aȄ�\0"��U��G����	��Y	n��*�xG��LB?P!�ޭ%�R���ũvJE�^C���t�쫶D�K)�T�!U �v0��x��ĈbWB6D(P�x�݃	�n��d�Y�@���LUz�
`u>��k�pX�|���~F�x�$#s/,[�Z}Z6I����
,��0�I?y��H�-��VRV'_)}e6����H{E����^V�:x2<X���-{��oC���jck��llc_�C��u���4ݢNۈ�g#pMT��z���jrE�:l�6��<���,�[K���
�
����fk���dg}l��l��pTH�.1�'���r��I{J�y��X*�~G	?k�f���k��2iJ;n��OIS"ڑEG�#<��y��E��Jk�l���J6�@/tmχ�#�&Y�a��h1�2*��tl3�x� �8��8㶈�}��Ы.PԒ��<QN��.������m ��a���Ve�f�Ҙi�k.��j���t>�m��_*]()ד���H����2���n�~�"A%�[V�m�����<�p�I��t׌=�ʫ��|>�3KT��oZi���8dD`,���c�$�S�0�:!&������j�īi��\6\Em��$%�n�_j4Ճ�~�N]�q��u|�����,���[�����l���h�B�/_�G�C]q�"3O��ާԔ���̾H�	Y�p�/������A�%�^�K&U���)��3��vG]#��^��C)^�:��'�V��eIi���NvAp�c1��/�S�*M�7���t�^��؜/V�Ϙݸ�.�j�ng�.N�D�6��a�N���˳sx��� K�خ���������Ӆ�����&��`���4��A9y=��UEz>�
�fI�1x{N%NN�����r͉�&4O�vRJh��p�%)sB7�e5���p�~nZ��.��Uf�dB�B���D����16ne�p�P�&	R��Ƌ���:��.`���`{�@�����o~��Z�ur|������!,�Nko"dS��U�̥�g[e�	�5�1��]*�h>�^E���.��n8�
���ic��3_���D8��	+���UEP5Z@$��g�}+.W�u� �u,��Q��t�n�q>��w�q��熠�\����O4�j#�$)��i��*����[Q��&�8����$�jv�� ��L�2u8"Z"�j'}�,����t�d�#��y�zA�j��J���j��9��%�CL4�m�J�b�x@8��/��S��[')�"��ӓ��w{������x-�g��2����,�b5����X,��0���9}�p5����~�3s��xY�f��LL��\%��������eU� ��c��Bl� �ȳ�s�U�@����-uJ���)�|��z5��T,6b�(bꝷ?�ꫯ�~��#؜�H���7βJ���`hO�[�Cũ�h��i�ZL����#��l�E��f�D�̘ĦV����V� �wu~y��8Z.�����?;y����n6'�C�����~���q;����?�kZl3�ƆV��>�ka�����oL$�#z�7�CӤ'Jz�!2.|�9��1�by�+�u�����3���!\E,W��+��Ԭ��»r��CZ�哳&�4�9�;���j��� -�yKi�b��Y�N,Q����p����H%y���� �c'�����K81l�!�צV�R:R��b5���*�7a�<:�������U�V������J�Q	{��rj�C�]�]���^-����>yv�c�}�pW�,�����lq�A.�84U��dQI?L�a/�s� ���Ž��'��Z�!���xwA��d��a8����tڦg��]Zn�ZB�����t΅��	/F?諃��ן<y�t{��a�jaaZ�^?Z�Զ �x��y�֡���`�P���}�	�}xrr���b��2��M'o���|s�$�LK�VEF��>Q���>1�VuT25`��e��N�z,I:���������A�ص�J��iR,�h�\�En��� ��C���r����rL���{�8w�#��[8�xhlۿ<�x��9�9���G��U�_�OV���i"��p�����{������u�f�'u���Qϟ��8
�H��Mw%!�"v�q�`j�v�J�(�� �3�|?�D(��FE�A��`)�.,��e&�8�K���Ǆ�總 �l�57]f�G����c���놻��`
���_k��^Ç,Śx����0�h��`=��h2��B�=ɋ��ȰT#2O�E��j%�Q�^���1����ɓ�/��r1�Yo��#d��~����M�f}�3�-x(�qQ�~Z2�?��-쫴L��;���S��f���`o�hz%���h���t�Vć�!HHb�GH�)�5쯴��/���h<;9�jZ*��`4�+�Oe��R���醶�:�o�&���l�l{F����f����#�y�Ě�C��BO ��I�X�e���v�ⷊ�g�>td(���k�\�o�7���6�a9_B+����O�-�����oo3b��7w��^/�V��	�)�Ζ���ʦzg܁@Đ�����7�����2�dR��E�pDR8iQ��g:����d�j��X:Yz������$-o٨����:�H9Rp�eY^]%�M���k#�n���p�ۜ o�!�z��S��~l#o8������q��U�Y�d̼<��H|�� ������Z]�W��ϓx�_�k����T�<a���b��r�(��::i�쟫��.�8p��H\2��Y�	�ʧ=���|�t=���}'�e�jSɦd�y�:p�IHY���bQ蜐�v��@$W��Ζ	̟-)������#�D��n�-���<�Y��2�{nxX̪�8���˦荑/��� {������֨�G��_DÃ��*�d(Q.�^8*�)N�|8n�;��$g-�J�<��?�X��;*�W��I��ʔ3>����Gw�hi�Ơ?f�~��t
]g�o���q��pk3�u�wwH ����ƍ��{��b���)-4�����l7#�2f�#��R+-��j!�~�^(���\+�b�]-׋`�7p�9�Wh����IW�<����q]\\!B]F�8���h�ch����?�T������o����ٌX0Ǘ�1�u�J��o��$"�0�&���vd6��Br�]/�cd��yeZ���} �p�9�:�G�-bV*����	"{<�b)G[��0��RIĔ��n�ng�/./N��7��	�NK<x�ftȝ��ˤ��9X�*�|Fq��|y9���5pC�e�YN�����NE�=�B@?0�6^���l�0[ΖV��^����������C�|Ȁ��ikaPeA���lg�h"j^3��ŷ����f���ɟM��LFKq�"Y?��������&��+��L7؂�{p����ۜ8��Z�����_��)ӖL;]C�b���K�ą���4. �e�j�P�b�6����T�ٰ4(wd��ji:N�.���.3��e�fm:.�R!h��;�yW����ݽ{�",���'9k�s��<[�.n޼���.�r�9�[}�7�_^Ɓ��r9��LH�"AM1.��T���P����_��}�٩�B�D�:���^c���a��x%8 ���j���
��Zv���R�\�� ��5��Q�	`��-��u;oH��*bNGQ�&)�%]"�A��3D�gg������V��ee�#� �y�މc����!W�98����G��vWO�^�n�EW��u}Y�3��-�|n�:�j�m����fu||�ѵ��eۣ�L�qy���C�@1�@1�J�U;�V�i���.'��Z�����k����%?����yRKN-�P<�H$�2�J�Ζ�leO���b%��_���i�L��Wfz
�Q��o�Z��2�:�T��A�p�K6���:�0�U�+a�k\�y�Cv��0����H�OjQ!�v��2�IᲴ�#(C;*+S�՘ϖ�w��R��ztuIT��j��i/mYj�Q&=�T�U)��V!���"C�P��2+���+�/V����j�[�VK7Z��fn-�6EQÓ2>q@�6a��k*G�$X�Ms����>�Y��C���Y_S�^�V��vp��cU��~wG���»MZo�f#�x",�"�:��f�}:%-@)�`M^[�.��k�L1��֜:�1�il3��_�o�R���Z(�J��%��s���m��r���^5���wDt�*�Z���$kf�V���}BurB4�E�����j�X9a�GZ4S��dH��+�O4'O_��tMj��nj����<�&	SX�T��A�� w��1d���"�d����K�9}���Ur...����u[�C<�Ç�FAP�x�w�}wkg#Z��?;�կ~urƖ1Ha�n�c��X�{e4�֐���Z`$K�������hg4�)S���7�7��s��d��6��npmze�wW.����@�L8�2���'>�E����k��~[ �]&���aM�W�
��5bk��GOB'�;+B��t��d�5��'�Emn����ё"Y��x�H�$��*ڠ�H&��LA��6��l�h�O�Z.���U�Ф��W������l{g�%=�<#�0q�2��9˘JP�ueDl� B4���Dv
�'�PUH%_I)S�>��{���g?��G�n	k8����z,Ӗi�=�xE��f�4zU�z�p�@�XK�#*a���dUGe��l	"����26韬��������]y�K���,����z)�����&OMV<z���=��>y�d���u�����=y^�cXaC�+n�؁��<e����Y�BW����y#Uy�F�2cD`4���A)L�w��?��Vq��_��b# ���J�d����K�|�J�Z��В��U~��L���*U�T!�lg �2���V�g� zK�Hs����~��������Q��`��ֿ�Tͩ��~�psx��Y��wo�ph$���&iã"��
B4��ph�����0��Ϊv18g��p���'n�۴�i/$�,vO�8�~�Q������'�C:�?���u������+���(f$ww��kׁ���>D�E��rRnr��g��C��/�P��,F`O��h&�}��ۇ����j�I����\-�}wk�����"�8��`ڞ����A���ILT��ě�W
F�j.��m�F�TY�ȉpN�PP��o�&�=<<ԁ�l���>���ڣRbv���^ͳ_����yEXT-w�#,������F#-�]���S��'N3�2V����u�έ���x��\G�6Co݆[�k<��s���9�2��6�vN�ǂ�Vsbʠg䈵��7���?�-+�D�q��F��gYb%ʀ�=����7q�(!S�:h2��~�H]!旚��4���
,�ńV�����p��y��%�.U9��>DD�JVP�������(�:O�nHH�u�R,��ĩ�^�H}�P���>sevrCG��?��[�!>3o��gI��rk�q:F��,��N��Ȳp&R^�Dsçf��.4�ͮh`sm��qQ��\���}:Ϸ�{��;2����x)H�:G��
���\�P��=�k�/Ͱ��b�x��Z2o�
�V~Spǝ�����$ީ�f\
�=�)P-m�SM��͓�ʅ�I��s�X�𕋐����*YR
�'6l3����W�{U+i>3D��4X��q��J���t��|u%�����?`��7�Z��v|��4�H��V-�j��=�
�Ҳ���^=�������[ho� /��O���Bg:K��娬�녟M�h���e	�[;v��3��/܂C�wvq.	
�l�����*T�-�DT?vMo:aܻ��j��^Ȧ�ł�IE^�!E�]��t �&�!�V�y�oz�ƍ�=z�Ia��n��ϖzu4׳'��d��<x�z!�zC�c�:5��5���+N����D�f;/T���M�5u�"�t����M���/��>v>P�C!��>�0���H�e��?�9�R�t߻�p���il�(>�������x������K\+�9�����6�����c@�;\oAx4�ϣ��X?��N���>]u�����RVm�S�v�i!�+@�� ��&S�?��?K�P��H��8.���x�?�����	�����;ggK����xn����6��i)
�~����^��Q�Vn�4�������/V�h�_MI98i��$��775o�ܥ�t�
�j1����Zh���N��� �C���T�������~�
Z��߄�\�Q��qߨ������,�6	:U}i@^{v�������G?b�k��Y�~]�N�4[�>Q^���E7�i���M�]׃MEa���EGSNB,���Q(���^l��ds;O�z�����A\�$k�i��C¾������v�Ν���
�5�����7Z
��yݯ�̀9(��|���a���t�jj��� ^��z�8�Eis�NJz��+o�5�X�3C�?����ڦ��pXJ�RIq��4+��hhd$�0lڕD8���+Y-S�]6`��?1�^�U�p~�sh��d�IhL?�QB��.�	�T�j==�I�h�@^qȪ��ם�v�,nL��GR$A}�T&#�r4Ɇ7�$~�k�,/���f�%$3۬�+2SJG�#���fh[� �A]��
��t���RE�Eb*P�r^ ��_-����N��_�����/�@	�������\���GzI���0���D,;��y�v��!l�yYHzg�ƛRHLI�.����M����l��>=~�� �+�Q�M�*Q���wi���Ie�1_vT�������*qk�5l�II(�
ㆰ��e�".�U��U=[��5�Y�0��R;u/�<��"^�ܚ$y6��.�2��$;d?��G�Y�p�1��5j�D�Ĥ�=�܋:L4����S��g�j����m&j	���uhǖLn���"p^ꨣ6�^��"6�nZ��kCRҢ-��X"���s���1���mm-}?B�*�b�п'I�UL���@�I��ps���o��_Y]�ڒ�W�ǎ[��w�2�f��H��a��פ�a�q��f�-�$>��W��YZ�J�&�����>Ou!��b����AHk#p�����ڂ��ԭ̅�^3��S(mmA�y���.�l�^U����'׏�$���ٯ���y�kk�_��U�����?��O>�d8�ܻw���ן�f�R�9:8$�	��PTA~�{AXV�����j�A�'9�8���b,�XOqD����3�c�j;�ݓ����aC�'1���ٴ�
��ZJ>tI��y߳qR��J��� �l�(�(�f����ݻw�������1l�ŋ�/���,8]5?Skj [�q�|벒�i��fpP-�@,���r�m�L��$�3SA���N��J���:]%C	��,CV_�D�y�J��-�D|x��w���|~y1eSR"���2>A�4�/}(���,ցcd���O������{�kJ�O.�������}Os���,/�&.��09�0�wh��*8:y������B[��/��R���x�+b��VC�R/�2�?i�1m1B�/8�_�>M�C�C�>��I5MK��Z�a	'�G�Z���T咈��[�g_�ő�|��Y�r���z��x��~�'���~�:�����G��@��c�Kʪ���8\X����.ъx.���l���f=s$��(��u��ui�l<���~�`6}�J�J��HFI����������^G�Lt���Z����E�$J��L��l�M"�*M檒L�4Z3��w�(#�oHО�?��l\(X<�:�W��gǧ� ���e&a&��x�4�,�T'X�y�!E\����yfVڝ-�T55���m�:$֦�������g~���R���\*��ٯ _���r_˟�����C�a���f�[�C�%yM����x0��B|~�����.�����2��ό��*ΦWk��pҪj���/���Χ��[��bb�qm_aA�<����er vU�Q��-��ƘR�	��yC;��p�-�vT��ZIJW��)5�i9�Hu�̭���ʇ����M�52,"���)���Z\a��������?���?z��F+j��eC����;�K���������/�6�ņ핂��w��j�r��Ġ6�
g��0 Bg@섺�WZ��b��[s��A�ޖ�ǐ�:Ɠ!'�x���HDM�X�B|=�X1�����j;tmR�eN���{Wf��A�E ��L�����$bqK�6���hP��u��b��f�UU@r��[qn2��޾�mxl���A����1T"P�-��To"�9=ee(��%qyXj�/lmQ'{�c7pz!gV��gVtԖLr�a���L<(K&,��\e���p=N&v3˄��CG�6Φʢ����q��h�M��K��Z]���3�s��x�6������(.�>}j�"�E`��:�R�=bi)EL*#��4/��Sk�L6��;��^�`r��F�'񱓓R��<�n`dh���@)5|�qE�t)�=�dK�K-		�P�5�S	��,]~����ݒ���E��=�M��a/�Ww�^�W,��'�����v�@�վQJ��%��&8�� �t�aR��f�̼��������w�}{��]Φ9l�u�H���ֶg�-��dsdVHu��_�_F�T��puI��UC�\]�ĥ���vSS!�nG� 4�����E��Ὥ������hї��w� �5��{O��gS�����.���0�<�.��a��ٲ�-��*��l�5��ˮ�����n�RK���ݍs�y�� hC.~e%�^!������z�E;H͖i]��JN�eִw�[��Q�3&�6��� dXN"�~_F�Nvw���7wvX��O]��W+���j�g[�+��e�	����%�e�1��P)5;��n�d�+ �WS~mZ��j�L,qqd�^�Q�A�'�[�p��u������pM���A5������zGL� �q���$�$�k8D���-=߮d���QP
���N���5~������迃����os�+<(G�czM@��[�����$8�����J��aU[v^jrGie��(-���"��o���*�Fx+�_��ן��_���	~K�좝l���5}J/�����PAL!�Y���?��?VV�X����4̖��K�i������i�M�V�Φ��aW-n_�g�i'����	��,����i���WF�����=����~إ�5�z���g�gP��$::��b6Ӝ�@^�$N��M���d�4�qE��v`�Ѳ�H$�j�X=o͑q>W;^V�ۺ
�Aj���Ip'Ir@jͩ�l�0��o��4t�p���<��S7���YV;�7��Pp���n����tҨ��G���fi��g
�$�Eb���|��+M&�~�Y�1gg�=A���-�eC���%re(@]�s^ �-b�h��.�����͛���2���./;��@��Lenoo�O�f$J_om����gC�p-�a���w���6��/�/���ӉTM�����[dSW����RYvO�g6u� �
�ؐ9�]R@�@��C&�6��/�qpD;��'@�l�����t�V��1uk����վ���advT/�l��in���Z�'E�hA^Yl�������N/?�WR�t����̺�$�mH¤"̍����CurY%d�B(&i�YT2��h{�<��,��AbJ�@ݑt[��Dfa�SL`�2T�9}ơ�Pb�ۄO�Wc�ݻw����p�u������_F^�r����U/!�8�U9��T�.�+r��5��;�Ê$�S)f�X��-[�̇��A��$�����j]%Ϋ�i2�ߘ��.y�<����R�y:�j�[�^j
����L9��y���O>��:�_�Z`r�����_����~�|���{����Rjԓɖ�5��%�{�%-�Ӕz�f��?>4J�N����x�u�
�����������F�2��P_l����Z�Cq�~�A0�Zqii�KgW-�!Z!>%�e������C�0�#'���X�[�n)���.j��)ݗe!������Bt@N(����d��#��C2������cz���RǎKS8�-ތ�����R��a-�R��Nx��`�˓ʐ����r�"K~���x�G�i��~�:��bU��g?�ه�wpp��=���ϯ���~�/jb�v�z�l�
�}�Q޿�r��S晃#��
sN"����_̮���!��� tq��"T:<�d:� T�uN�J+^�9 U���� v�9����2ao "�/V4�l���dI㬘�Ƀ�9r���a����A�E��L�՝�[+���)�:O �gzr��jԦ)�o�I�,���'xg"Y�6S���B�Q�-�H� �d��_A͙s��o�=��d�gZ�@d�XΙ�0xX,���Z+��3������z�b���Cز�6������$�"j�4��K,�f ��4! w.x�ʠ�C��ӛǲe6��GG�-��&Ou���*~%�=wazN�|�̉��k$kE��`�f=�����)����Z��9�(A^�Rk�:!Z�ɖ��q���1͙8���Fig 95��<���sыD=j�גX�8K�����[�?���t����;)T)��~�����23���#���9>B���W��o�nZصْ�J��6�'v���F�!�����T}۞��&}��������%CQ,#�OA���K�=Μ�֌�J�j��t�T���rK��)	��~����E݉����x)l�Y|)T�j�2����;� �n��s��kĿ,��x��JQ�U�Z�2�5WĆ&h�e�>��l�:h�x%��7���6?�k*;�0P��wz��xA�Ed���a7�B���M�$p:/��g���'��2:gI��K��$����]���p�T,�-��]�M��M5K^����yԅfOIQ��!��Wt>	�9wA��=5ǥ�0Q�l��:��v�-SBׇ� ���|*\id����S�^3,[�;}�����tJ˂�Ĩ�� 1��p���v�+��߿�;�Xȳ�׃8���w��QjEX�2�ʸ�-�A/#B	)J�,_�+y�Tj]��F��k�K�R�O�Vv3�.��2�(�@Lp���-\�R���I�8�@x��(>�?�QtM\���f�ц3J�#�NZ����̥�J��:9��b#� M^��K��[;De.9�!����"V�q��Xy�d�M�N����� ��Ts���a[^�HFõ��cg���{���V�ڴ�9`I:́hfV��+��K��`�b(�.S���Q{�O���+���Vp�D��ϊ��5�^EC��d�8o@������<K3��j;񯚺UPv�=�8SpBvv��}�^(s����Y��xH��(E�/��Ts�t**A%͠-]�BWv�ܡ��T��}�\ꞁ�h4�V#eS(w�U�%vc��ĉ������I=b��U�W����쒺�)uI�)?M��ETO�����_UJ�ӫO?����o3w']�p@�1-qK�_���_J�&�G2�s�����V�n��;A;sh�����y�X:��Kii������/�	�|�海�~�?��69M��5���<���:����{cc Uh���������?�3@WWR���������_ͯ��˛f'UM�/rh����ZE�:�n7�<-b�K$=\�]�û�R�Yb�{�ږ�Z��u�$�����Tm����	�]�R�x;'�?�>d�믉R�>ʪ�6k�Df؜"I�:�I0\�8T��R�z�۴�iW��ʮڭW�
!�y���p:سB�����
���ZR�샀Mp|uN(��U�m�h�������Z�#��*)�G��/�V�&���\DM����^�w�D6b@(������
@\!i����iǜw0��]m�Րۤ7�`#.B�9D����
�4!V
+��^�hc�ZxY$i�ĕr�m�a4��uӫk�2W�c4�;��&vr��i�4�][l=M����.gp�G��J�RM�%|��	�v�Vtk{�-*؍7^�Xh���ɣ,U���ﾳL;���it2S+B��֟�^u`H���	
��s�-����D1��ӧ� ��׮�^O��_<;���D��Zt]�K����j�\0�ulѲZY�\%9+����,&"">%�Dg��r/E��oI|\��b
�ϟf�l`Z�7�H�i�z�g�Y�NT�+'(W�{-�m�i� &ܷ��<�ٌ�����.���*B��Ї��jN*
�8D�6syz�27 P)P��2d�T��:N��
��m�̱-�_C�*�ݮl۹�a]]���a�A��S�&�G#Wml�Z~�N��>�Η/f���Í	�pԒ�~�'�y��vH�2N�z�Fqe�*�z�`�+l�>;���� 3\*|H*V���cʨ媬|!�Ň�r:�߸��~!��Ԏi�E]�D슏q�V���łi����_?<�?yr|��mS���ٖ���g������������>}v�W��:�y�����հ�Ї�ܿ��9�IfΗ<w�"�Ur�"#Hr��]���YF���4����}�9C����j�@�u�����t������=|���ٔ��%;G-��8��!�J5�	�4)�u�}=dP ���l��:ܺu����([,��u�h�p�`��d�xY���X�"�����T��(qc����l����,���r
O.���$ȀgR�55�)�f�������&VQ��4k$P>~���1<���D�$MU�P�q��g�@X�&	+�u)�����J����	��b1C؏o������,ӷ�� �I���Q���0u2%�`���׊~��wM�NH�D�sIjX�Z����*�q�\ �ǃ��XV®NI7�F�s\��K�i�����8,�2..�$�dE��F�&�0�fS��{���/�X)�eeM��8����`��H�v��k8J�3o����{�w������G�M|p:������Ǽ��G "�)�d�Zʘ� � ½����[*�Fi�ŋ�`�QB� L�8�c7�'g/$�=@�O���,<͠�R���0�ix)�ƅiD��0�oQqfT�@����We���~]�I�<�޽o���'�i"q�Nχ���М�Ɍ��E�94�{rr�՗��O��� ���!�hC7�Q�*��l&H���4�^��y�*�5�~�$f�	w@_I�t��	��_G����3f$�ӟB�`���_���o��6K"1[��1ؒ	B��d������^�g�,�2rڴ� ѵ��*s�XCD�T/.�Yx��g��ƈe��(�W�=�M�/�4F�� �]Õz*iί�khl����85,��+��B_��U�^_g&b霼6l?M��������p�1f�|�IMp���mVy�>}��&Q;�uq�\��ch�;"�x���ҪX6k�i�W�S�?c�t��r�M`�Y��n�ek�"7�X��o(
�����iΧ���g'������/����O!�m��P/�x��S�*�M5^�e��O���X�i�Jp�Ag��`}�K����dxb��;�1�la+�1<G����H���Ǚ��(6�uA�xSf��w'F��t�mW<�� �%N
�zK)�2I�0W5�-��ށGz���.Y��p�~i���O��5�y�����>y��rsdrY�����1æLT�qt�W�L3�#.��>�.om�W�E�7HKN���V��VΟŜ�?�OOH_%|RFe)�\�kr!=%�l6��3���*�7�@�BZ��X��X��(�({�&I��J���XsϬ�z������ �4�wA�H6fz��Q��h2>ц���X�FWWwUu��U����ι��+Bc�`�Q����}����2y�G�v�ƍ[[[;0�����G�.���m8ʚ�'��鐉��!v�?~����-�
\�/z��Yh��0��.B�feO����d��������?�y�6��w5�BI��xi�g)��d���^�|��R%��%�@�1`��vF$-\�2o'�?�Xj�5 �����5|�}'t��ȍN���7����G�5_T�/[�bǷ���!�%>�\eIVս�*+~�i6[*+j,a̴fYҏ9#��sy��5���K5).��#|�W��r5������$�o��&ÿ�����б�<V�pJg������%"Y�CA��W�祥����h�<
Hxv��U�w��3�Y�J.��r�����OX]&�g_|�|��>t����f��������t�g^^DE^_N�h���(���1?��n �������7�e�T��H�����Zs��;Bư2�4-�j�7��#��
��*3�ؼSyk�eE�5�:��w���"��Zi��n��޼��9�}��bG����r9ln��ڻykw�V�}yPn%�%I�[5Y-�
���O�V�F�Ɩ�G=I]k��?�ao��f�2��!f|��A��辨~5ӹ�Q`W��(���y�19�ʯ�_�-9 �_�NB���ɘH���Ƒ���>�����MJ���*'}��I�e`\1�R+�f�Z!g8h��h�`�~��_�����T7+��A�v�0��#�ί%ƚW `�JR6^g���E�������W��k���C8��s�U�����ǸW������o����Z^�JӞ2������-Ogs3��cw��m.�����������v��JfM�YUM�{epG�"e3I��fU�Omc�+ESzsюo7��ʎ�1����{��r����m�v.w�����a�RU���~�\��/���(�����oKf<�n6W����g1�,j�X�m��R�_��R�p_���H�j�@�|���Ӯ�e�h�h��>6W'��j�U��6�]G�Gn\3�k.�fהK%p��ߴ��Y��"fm�?N�d�|v�Wi<���H�[�����#��L��	#i����g�2,5�k< @:=c7���3�n�sNa-��iZ/��)`,O��0��N���X#��H���fԣ�W�F֕'0��2�uv�H�R��-��!�K�҃�^��\��]�z��*���oY��XW�(z��VnU˲-�L����;>>�~�z���E++^�P���ii��e�<���Ɔ-n��pϷnlYU?U�g�`��+�kSA��W�R4vgܰ�~�!�D`�
DV���9ܯ�.k)VY%$�^��$j�����2{���H����(�J���1���0��2I���!Ic��v� �U1*p��I��~���97K�Wo��������/_���y������J#�ȗjl�6���oڙgW�$׶�W�r궺����z����^l�[�iEH#N��廪�A��0�p��"+^x����F���1�`�%e7�p��(�L�v�ՋZ�j�uKj>q�я~�}�����y���p8�,��d<�Tc�{���������E��_��T�ɚ���.�0�1������,w�ܩl*����y��.-����͘>��%a�J�$*���+�ŋo����u;�����|iV)��o�5P���ӆ��������#<������,��U�U��e8�BN-�|�n�5�8��DQ�D�HV��OJf:f��jz,���ɫs��&�ی���1��qfA���}C]���pX�����w.�lx�F�F1�G����T����i��>�J�^���xN�����_#��Ξ����ӏ>��st�@̶w��|WS,I��;;���x@ⶩc�|MaX'Y��m:?�����~Wس)�?�������x�wntu���ȭ'��f���ރ�<=g*m-筲�Yz5b�X�Jb%�5�]nݾ�ͱ���Mg���_�������U:��
ήu�_<��Z�2���t�?�-;��	k�0��vQ�!�v��uAS�ɟ�cU�J]�*)�L�j>�fp4��q�	#T|E�x�wM��I3�
��E���$�VY,6Lg3�	Nɏ���d��m2�����P��:�j�s��0(��sx��e�!4�wE~j]]Y���[�土�,��������}�{{�|��s[�%��d-��{4΄��>-��w�՞���yɶ���,�ʻ���dVx��Ϟ�mc��֐��j��x���u��m7�ځ��O�!�I�b9u�$�0�]�{�e����D���ӜS/��L�6�ui|a�zi���fE�&3��ĥ` 1�(� �PP�|�Y�=�������^�F�"'~�у�_~�e�0���;���C�� B�stx���������#w�cs�Q�=kʑ�����5�9�u��Gdi���qnZ�K�`�
/d[W�)~�o>��U.o��!p%lTLu�e]��4���Փ�F�JRX�UB�\,8�&��ܣ[���z	A0��B~u�_�꯹�$zP��.�8PZC|p2nT�ڶ�3bof��%#��-d>��Zώ�8m
#�[��ә�AryE�6N�x�y*Gbź����y���܅oꍕ�ߵW�΍AF�BD��.�!*5��t�y)�Pr�eJ:��塚�Κ�7�1B�z�ʚ��`*�m˰�Բ�5���[�򻰺n�1ɚ�*�-Ý��|���f��� �&������ץ�����X60yKljSd��*^6hܪ��䗹�����'�:_�������5�_�!8�W�z<�cb'C�rUF���|��ï���L!@����'�R���������|�\o��F현�+���^G)���RWL&Ƣ��:AVV���I)݆�*��*�_�'��x(�J�+�D��3O�mM�O��/��d��_�̎+�_���2��}��X��P������j��vH�,�o$�
�PA]P!ɘ�u�=����6Rf@D��K��'�8mb�����ׯO�Sجyh%y�by�f[�A4͆
:쯞�:�R���-_<`G�J�H�}\I[��`�{�������C�������<��v�w��|v��]�H��=�8zq�����[j
̛�7U� +]�A�>x@w�mr�A�&��k*������>���!���w��$�\�\�׿5��H��Bd^A�!N�Ђ�zHk֠��X1���j-n��	��b�Q���8��Y'�/��~�|�mj�V������jGsr:\N������5����3�f:ē	Εc�����״��̪�_����N�V�pg�?���j�b��0��bx��qIT��yg�x�7#]�p^��`�O(�Z����\u�n_�-�j��sZ�{�ժ�B�z) āp
��{�x!/^�j-D�S�����{de����eU�By}y�Jv���6Bӊ�^Cβ���2V�
�	H���p��TR���]�R��:��7�ɟ�C[֍�=��[|�<Z��!1���õ����<��S�(�K�����'?�����3��7S��g҆�I;��8^�86*z	)%&��*6%������*~D���z� O\����(�/�ͦ�(���qI��rdkEF�z�C����Da%R:�T[�'g�.8������A[mE|�z׾Z������n���A����a�?��y���޽��l8�G�
\� ��}�N\S|s��cd�i�d-/��*�e��.�d�t|�,/�O.�7L�e�6V2�Ǡ�iq�y`�E�KEr�+�n��W2�E�"�f�#SΎB`�"�"��WX~'�8߄�0�v�1q�k���'R�u�n) �UPY��V����!�1��� Ql0�� ��v�o�c��6iD3��¸�C�X�Y�/.g'g�Ua��(�9)D�M�(¡�����y&}�=�˳c�y/g#��;y��`�/���������n�84��
��Ai"�kx��×M�m)(��s6_>}��������{���ˏ~������d�E_��|k���Y���wV_�C��Ӻ�p�%a�~��B�0�rv�y�!\ý��zO�}4�moNv���@(��b��8����q����kmG�����ɫ���z�b�/��VܧO��Īnm�2G���~��˿��?��?�m~���g���������FP��o|�ѣG�糽��x����ڬrl��+�������:��"���-�p\_t��)ŎOu����v!�<yʨQȇA�s���vJA7x~�K..-��6�/�yɬF�>�������朞G\�<-�����/?�l�r��t���`�_�m�"??���u9%eAJZw2���c{�l<���8���prά���^+���ԳǏɉ���������ㄾ��K�DU�&�ֵn����L�us[R�Y?z�>���p^��mPC罱�3�0_�{����>�Q�&0lc%��L��O������o�yqɾ��<��e��`0o�`�/����:}uD��n��ٽf����g�3�U#�n�N6òZ�nVTgB4�эџq�IW{!g������R�8��J�����:!�z5o67�IJfO���7�&5'���༗��hm�>Fq?��jZ���u����]'d��|/��������"�M_Tճw�y���?`nw����+v��R����C�G� ��^@�,D|�^��fe~l�l�l1;|z�����0訳�t��+�n��.���@Zp�}b���O�t!�v0*0�CR�����S������V�kĥiuN��`4VDm�?Z.�w�h�dP�<���1�ڒ� k�A���}���o޼�o<:����?^�r�#-
�$)q̑!\J�"�A��=-T�k^bZ��/^����9Liz��$��d>p̂sp}w�Z����ַ���������O�~���`woo4�\�~����d�e����>�CE��.�&�������S�ED��ӳ��<ǒ;n}=�Y��lmo����P�E`�$���`4�%|(,�C.��5��H4���Le���W��s��1;����f��vrZ��A�}�#��X���`l�~�����i=^�\z�iZ��΅1ʽuf�2^��aIUc�e����=�%���g}�>'%G�����Op֮_��oٲ�Ϟ��v����]�Mq�!��4���@]�����Viq9_�<?趨�H��qm���p�p�.b���G6ւS���x���w|�r@�=c�Qm��E�����y&����S��9!���x�������FO�<v��8W��g�r4����x"*����� ;���(޽}���}���m"�^���Č�ѡ�W	I.�򫨤.�~)h��5�!+�5��3�G6�1����i�)/A�8�Qo���t�"�x4�.��J1���|	��!Z�[L˩y��#�քc�Y��}AhbԮ��Ҝ^l�iW�l��^�<�9{ˌ��:�/Ĵk�4����+"�U6�`���l4����~�����GOO�?�h���/^���O��Bw�)�^��z�󏰖+� ��{�^Y����¨����
�W�(�����lv�g�6��$��k����&V#�����К�e�Sy/�����t��\f��	B�I�i)5ק��s�K�9
�!UF�b(��eƹv����Y���-ʝ��8�	Bs�����ҙ[�������b
my��4�b��_"��t�
Fe~,O���\5��$��=n O_4����bs���q�ɶ��Dj780~�/��{�9�UŲ00I���K��-ȹA8�����%Ro��@����@Cu`sqMX�4�F��:��.���o (���h%���~2���e^�N,R�Ŗ{���TY"�\�]�bm��vьṔ�{�4��]8��,4z=q@�F_Q�W��.�V���
��*3�)�By����W߃>sq�R?$
��8���k�w��]�y�2o��ʪ���2�Wǘ�mn�@sN���>��x�U��"h86G���&!��dn]����vI��=��lE���.��:�\������P0���
f���Q�p�jQ�a���椿Z�y���Z�.c�)8w�;���gON�a&cj?RE+:��(%�7(j���!)_dOJ�>�b������.���Gi�e����V�h
�>�)-����n	��_"���2M��#���9~�7C΄\U���2�1���`��섃/?���0��l�����w��_i#���)��4k;�_GHva�w�U�to����`��f�g@Y�����A�U�R�ׇ~�7�8�'�V�jQ�W9���U9����ڻ�o�'���׿������.�$k��K���ER�Q��K��7Ê9U���ji;�\��7/�tf�S$_�*K9V������b�̡Vq�B��>hݲ�#n���sXe��(�PS��O�N���s̥�(�^,�%�x�R^a����R��I�@LB#�"�ml
���!�"�$�E�!"�k���&c���d��[��qŒ`��*Q�&�$���W�B��=m���qx�Ȫ���׮]+b�l���hol�H[Vѷ�=�L���
*B���X���OGC��:����kfC�d\��s,��7�=�g9��a�u۩XJ2�Z7�X]l�)σ_>~��n�=���Ʊh� ꖊQ"�e�E:���ZÄaҤ�>Z��o�}}\�Z�K�be[��r�?!{�89|n�����V�hi�(�J��>�E���v�RpWl}��6�(���8b��VP���笠��yP���5$V:�4mӇl�	4���v�:�3��u�����lN:��Ig��F6��lK�̅�1.۹�؀�~K�F>�ӝ�����\���F
p�FQ_��#$���F��JC��<d�Dp�\����MF�����H�ur���مA-���*A�u�niU;�)ZT��� .��DF�>�h�_4�F�r���=��o�N�ܵ�u�={��_~�s����~��8����7&�Q���;w~��~�v������'���E &���4&cF)���
<���l���<����+#�����BA����:�0y0jHyD�F�`��X`̖5YŪ��3��a6��5C�����(�_0~��o�9��޽{4񈞢�Ǽ�@�w�3';�88;o �bS�8=��в�����$����lmjD����֪߁��������2.��Ye�9={iylqA�"���i�_�{�Q�H�4W�xi�qݘjlZp�͙�Lr�A�pX\�����8<��{���P�e�B������％�)�l�1E�-&Z�%Zv�{=,~%�y�MB����<'��X̴bX*�e�ͥ�KM!`Ֆr�=:?#���(��YR�p�1ʫ�O���y�=[�FK���a��p��pf66�88pی���>� Ď����ċ9?z���p��.d�a�hi�ᘐ�����WĘ`��ۓ	vǩ�XC<����,�lU��/�������r5^��(�Q���D_ִ��d _�6��~�#N��.;]+M[��^�(+35�9�e�[z���M����{�ۻ���w��q�JUkQ���"eH�N�A��t[�°�����9t8/�(Я��M{���u��N7��@q����N/�Ռ,�g���qͳ�ݽ�@17�°'Q�m�����qk1yl��ǽ����JD%B4�
�o��H�̿��#��GU�0��N�77T�~Vj���P-]��Dd�W<��h�X���|���Tnol/"������^��������SQ"n�\���$�O"Ϭ#��d��_�+p5��y�hL����R�����w8�^���x�w6����*3s�4s<��z����Z�(T�{M����'���Y��%D�s�va�>��7�iׄKuK��0����/�7 d�}�/2�u���恗YչBЬ��Z*R�&���A(A� �gtH�xy��杻����(V�,릋�ʣ�i�Z��̀Z!- ��4�f�Be3Z،X�Ȱ,��,8�o�0R������{�@�گ,SÕ�f��!��lM��ҵ�1]�J[�P$h��(�w�奩)�CX�8Z�A�&�*�y���L��c����\W\��iL&��]�݄:D�Te}z2��"�RH��º�z5G�Mf����mޒ+5��f<FSQI��T�����WIڻ���6��gY�B���f49�t�1�����p1	k��D71�~��:����+�Ҙ�҆������q:dl`����+��4�������7ܠӈ3��?������ݹ}�@���6ǶcRɥ�Mg��ѐ4m�u�9�q�Sb�3�%]�ʀ������������a{��Ltߪ�%bX1��;�=Q6�ɓ'8�F�*�wo,���>����I@��� �]�O���Nt�\��b��_�}�\�M��ԯ�0��T�f�!C�Ek:�1���W^K�{]5�؎TSe��a�����qp�d�a���c��ܖ��C\��'Ӫ��K���A���TP��#�������%�버�ç>���@	 ^pJ�����s�Q(snw����^�ƅ�7n�����yq� �x��?׆�,��
o��S�������elumu ��j}Eg�嬻�����o{��%ݢ^����cc��.&����#�Ky���������)��-��!a��j���;��Ç��u��,�|k{c0$O	�BA�C�u_���ɳ��/�PƤ6p�!���8�����k�P���6��ɇ������[�����QpȴR�`ō�o���-�ՀnO�j����!���J��@�ݹq���k��]�ٹ���WP�����듪��iA%�5����s��wn>~�b	Ã.�5���ƨr&�e������C:�mgƋ4�m56Y0�&��\)8���߶�as��y.Ωy{���wYT�PZ&H�]H`�S�pwy1]�&�;��Be�����bfs`D�=s�qce����:�L(�7�G��^`�>��~���1�����l1@����\��(B�����#���<�����7����q֛U�V���Ѐ����<�i��I��dmq�2��O�S�
�s|ׇ�3�OV�4�ؾ�?��mm���IV���wg�2��ֈ���B�O�r��*����o5�����$�*�;�i����.���t��������8��㩁ю"g��.�,E8C�לM^�'�ߚ�S��ڳ؀��V��,�W�t��`S&9P���q�=����s3V�|������;ҕx�d��n&�R'3��wIN��,��gF&}��GVZ6F�δ�,Ws-fM<U�|A��8�������<W]�3����] "��.��E��Z��G�z�������A{��˘�����8>�F�"��*� ]I�Yj85�ǩ�aêV[�����x�����%"����L����^8��V+���� pd?{�}p���z��<��׈�d��2mnﴈ� g f[�
޶���2���u�ᤫ���^�r�|6�)ݬJ����p4� X�)�ȩ�SYf�z�ν�h8�Ζa��-pI�u/�-���Tq3��bTy$
 E7�N��`�Ƶ_�-���D�ub���?}��9������������+~��ܼy�$A�Y���[�ⳲZd)���PSfp�/N_�+��i1���zg�r�3����ϸz��k-x;ZXt��T�cn��&y|u�;��0�w[$�W�zv���ZY�́�c��$��a	�&L�2�!W׉ ���r@��{��ɦ�s� �v�b��dr獻_��W\?����_������L2v�9���&�gv~��ښp"�D�Z�d,)l�64��������k�x�q��Ϝv��S��W��xq:*�AU
W�Ea܏a;F��)T�s��f�3�6I;x�ߞ��Q��:��s(�e���_��]c�=���Esp���w���wئpzzy�޽�z����-f�ҔCk��`q��ؠ��������/>Ų�$M�c\1%,)�/1�d�t��~���n��]�q��0��g��Eb}�!�t���G0F�9d�z�=��������QZCM�}n�M���Lg��c(��>�`���`��fw����7�waD�����f�����7pYB��Z��l�mn�E����� 0��|�ӟaebˁ��Q%2xX�h*�|�n08>>���ϝ���AQ�h��'?�&QlCVc��zM�@�zyil.e5"1Y�K�d�K��U��)a��=��V��Z�6"�i��UnΞ�5.�-���� Btޛ/��)Q��)^<:���{����*����^\�sح����J�e�f?bǉ�2�V��gz5X���m����L#����->���FC�����߆繹9�1�o�o�Ӏr��F�&+�ںs8�l5?��.��<<|����HT�Պ�O|���K�ե[���jU��j� їi3�Y��k`����#h������v�*�~��,+���\�����A�����ds�ڵ%|�����Ep�6#�|�p�!��!�L.��z'�H��NVi阉t�qxH01��
�b7��|A:���qLg�'�5��Y%9�F����aƞ<9Z.m��:+N�����l�����;;���3�/d!�ab����*h�j�B?�$�5D��/r�E�;�̯����#�|~���q��
&i�$��Q�g�[����?��V%�^�|��� �UY9/b3U{�:���֖u�&�,C��,�Oxmh4�x. x�@&��.ʧ�_|����!�yk�ݹ���裏Nϧ���rzyz6�ַ�����c�nY{�QM#��&��kO��|څ�:�'�ǀ��P�8/�$��^�],uJy�aw<NG8{���w�}�Ν;�>c�Ǐ�Bc<}z4�7��_�v�gYג`S��O=�{5�|cD�ۼ`�;�|���;�0���9��a7�A���l���Ջ���z�F���;?�^s���\�om���s�`6[�{5~����̬Vp�=����@r�x��8g�� )N�EzYi�q�Y��uf�f�^�?���m��#?
� �{����\ex�ɀ~�a�Fv>,Tu�*g��(�Z�`�:�:��|�@8���	�4��K8��p��&*-��&[ۓ�M�OiݶY�5L�����7�ߺ1�����%���e��ا�o���Xs�r:�ŝ]��_ĎF�u�����mԘ���" `��M�1�*��pqA6	�㔰���h�w,�s�QX�19���.ʹ�)�AG���4�Zm����([�&�,�	iwvxfO3�eq�.�ǣ��r��/���M�M�
R�3�JDҬ����x��a�<vկN^:���x1������~���꩕��]��k��=�8�D�<�
�4(*��J���*k؈����z�o 4��� �նw�u����!?��6��d|�����k�j���?@�
$��g�@f<�|�m��� �������*�g�o_�����n�U�TL����$������peVmh(o�V��UP�������_�>}�c8XE�FA�Q�3����嫗gg0��ܡ�>��S�y{X9�ϧf	?�d z�T��8�}��o��v���F��P�=Xj���(1���%�'wY*��:���L��nf3i`�
>:��x����#�"��b�{�Z����q�l��6G��v����q��*���\M�Z��������&mzW����#���=��Q�K�u��,S��>�4p�2��T��-��)�2���Y[�LW���v���5܆U�fJ��A�b�"��6�T5@�[m������T�W��v����:U���S�}qр���Z��1� ��l�JR��r#H
n��-�ϙh��'�C'2y͎_Y9�� 8%���U��ҙ�4X3x3b�!���5����"�E�.ۘ�kgg�ˌ`���G�N�Y[�4L�8~%9���Bu�mt���L���m�������)<��*1�ٓwtM��HB�Mr�FdE�74����2��'��K9{yg��N(t��|rd��k-M?�l����q���7n��!b��p�1�DfK�wvĤn�̪�F��jZ�*�����ƄIK�K]\^�oSNam(("�
)&�ƌ�����)���J8�;;��~�}b��S+�TVH�����$�T�/G�ǋ2s��mNմ��le����PoN6����X�	;���+�Q�KPU���pm�-����w[(%~��� ?�2˫�p Hcs�u�}���ٚ��!*��wBeJ��P_a]�θDEע%UT����[�N����#��a�c2Y��`M ���i	wJ�a��hR50�{�]놖��n����ع�>A[�X�6$�����*�p�C�5��Qϱ�E��k|FBFSjSD�)[	�
��Ë�Eu/�Ʈ�,p�\�/�po����HUcG"������2��԰�x�[o�%�O?y��3+UYY�O8c��R�8I������Ӷ�+�1������M1֞B���ʡq�9�pY�4�׊�u)�QJ���\_�� ��He���:������~�3��`���E��;��`YF���Sa�q>/W��jW��)\v~qj�����]Y0Gf&Q(�p�Uh�����W�q1��˜Z�$�6`M˼���B��Sʣ�d=�&<.n���p'�'�5D|''�DМ8��úag/��&����~������/��R
����{s��|>%�F9:�9��{��k#�r���M����X�6vIյ�㵩Ҷ�����^�qɫ2d٢J�lI}㶐r�N�,��Ѥ؍qzi٢�rmr�G��RU�pw��E��~��*v���2��1+s��P��~���߿���g��קd����V�� f������w�~��S�#�/�=������1��G]�-׊���99"��wPZK
~��t��RSzB�jQ��4�|A�hm(~h(��ÇǓ������d ��I���1~���q`'j��\U����+,�f��1���r��"����'��[�^p��9�Q��f����6F�k���E=S�	��{����Έu�ל��΃�H�e0,�Z���t^d=;�ijym<���YA�!�����^d3���;m�AK)a,��o�uqqq��olwϊ�Dv*_ %r�؂ d�7��cYC߈AM����h�:$x	e�px���W4�~3�V�u���e"��b$͚�U�,���姿�""#�Yt�����<N֜�Y��n�<x������y� ���zv:����huV'����=��{c�rٴ�:��P��M�Z	�#��[5�\��9�KC���|E����ci*b8��r�'I�Ou]T��B�er9oYK2��P��$���ы?��?��4pXYD<�dc�����9�βSJm땫����E--����6;(WKx�[�e�s��1�X_�E�"zн��������}2�F���%�ߏ�^ə��M_�eҩ��uU���3c�2EHHb��\�i})e�{6��{y�Z�̳����0�q�t���!�3O�u��}:<:�$+%}�1���IJ_��2P1E�%d�8��u(�s�A��W�������o��e�vo
�ce��J,��F�h��n��8~3�W���-H��@�㜢��9���7��������	�X��o��xX��A���+뱘��Y�+s����L��j*<=��W"c��t��� �����6���'�P�r�a���U3�����Un�Z�ц9Ej}3_�b�ˋ�i*zVB#v��R7Is*-�o[���y�pv�e�J�^��G��x.Ȱ���v�q�y^�Y[�&�d��`���ē��@?Ш�Nu�N�YD��^��-[�4%�����ȋ�7���)�Yة�a�F�m��Qobn,�rA��Y ���Vɩ�rsݽ��B�~{n'lG�4��2q�Q���v���y�
�`�!1C_���������}�Mm�?����޳�9L����(�f_g�� F�ܚ8�$���,[�.x2~ۏ�Ĺn�lz�ͷ�
�oI�*�i<s*ǭ��n>����3(�I���U��լ�!�N&�<�AӲь��w^��C���~��'��Y=�7E��$�ٝx�v��3B�|��7���n_����-����ݝ]����cx��5���8��3^��7y��6����i6�1���m��NW�n���+z�Hup�Ļ	탯NU�����+�fZ�B��&A�ݺuc��u�,��N�_�z���H�j"���q�?�s\l2��9.�2�n�v*�hcɶ���
�X]E��ӶXv�Za$�J_'\]c:�q|l0�J+fn�cm���w<�Fc:�֔��G$\�4w�0�_�'����m�C4����E�bq�+T͹�hpY��e��ko8@8�s}� ���M��uB-��	���_�_�8w��8�;;[1�zc$�=sY,�Mn O�Y��Z�a�A�P��t���$��ӄ]�*��\�2��]�0h��f�ޗ]��&:�l���Y�~�Rb^6�
om%/\z��"$e��UH���8��	�7�n���֛�ن��ӎ*�Wg:�.Q����nD�זr�p|�1U��,�k��OM(ZZ�g<0l�(���^�w�)mn[ri��aDj.�����|�k����+�K�li�m�N�G�4jeE�I�:�|�u˪���rs���������石��?��}�#��gcs�fd�L��Gɣ�_�H�L������/�C
�m�ӊ��%�g%�=ΈT�,CGf\W���Q�%i�HEd=z;�T���CF�48�Hb�(�ھ.�oþE?�Bq)Mƺ��D���ji�;7��ǃ��|�b���5��ɦex�Uv��M�����϶�Ɩ� �%
=���Î�A/�:'x1_W��%����B� @e��4�L ء�Z4�X��<��t�`ZR!Y�q/�.�`\:[0��Ƽ�ς"�4�V�b���ۢ9+xR��ҥ]�ɹO"���b�r,��'��ɐA{���� O�w�êa�+�����W�_�޻�9|9xc�<�);\�f�H_]N���TԞ�Y�zpZ�9�0��F(4�M�l����x`agsF���\Ng�4�&��
�D��w�)OrN�Z�D �D���������?88��� �ͦuE�����֧Ӌ����V���A��7p1_@��v>�`'�|�X��2!5��jcJ��L�SFQ:��P�ʉ��X'�c��5s	�Z��Q���!��S;��j��%_��jkg��$��IG������~������&�a��ւ�Jh��V��ܾ/<�����Y��ͭݼ����X_����-S5����7v67�ik�C��痗	a������|���#��],��`n�?� �l&��rO��'�D�"�0�b��5Ed0"�bŰ�����q	Zw9�jA�Ӛ��Ω��}
É0�Z�%�Zڗ����{7o]���"b����w�}�'�~���~�db�y���B6b�c0���fƈ�p|�+�Q���t��L����F���ϟ�x���V��	=�����h�����i�L���+�`D�l�%U� z��C��/V���KǦ�s%+7/�Qi�?��4F^�j�X-�!�Y�i��o���J�&�V�un4�畷�G�<�>>~z�0~���T�fj֏B)k����=��NQ�חU��-d:�,�����~*9�3����Q$o4��|r�Ъ;K�V��}]oo#�%���;��ҙ5m+�|��z6[(�Sn�|zv9�[[\�{׮]����/l�Vį���9&{�Zg�9a&[��7����LӨO����;�?|�Jy�HrN3^e�Z^�k�X~�ًWq<���&V�	߂���]�����>�$p�QN8b�)�5]-iC��Aq����F|�g��3�.Ⱥ;���y�s�h��-���}܆:��T���O���+��6b�#g��A�=~z4�$Wu]z��hss��Ǩ!,'X����.{�m���� ���*%�L,F���*�f"��O!nN��ئ������0f����,ӬiUjJ"%8bئ5.vYm������뼙K���#W3�a���h���U���������?���|�;vxx8[f����޵�j6�v����4Ka�p*�6gK�R;�33���>EՁA���g�(�p^b����TY��*���Ν7��٩��4޴�-/�;_�ɉA���a0���Mw�d���`�(���"���1��aoؼ��!i����U���h����¬,.����h߈�?K.������^���Fz��֫����;�qZ�7�l1=��^L^Xf���#`ͨf!:봼�`�����Z$iҳ����A;(����U���J��)W�Q u�\�Ğ"�.#�!�*dR8W�
�8I��Nx�=�$�vTME����d��yb������8"8f�N��b�,���g�˧�.�P�<�}/�!̈W�Ń���e�-pu�h�,�$�����b�&_���q�$���Ճ�a��[���;�ͩ��"�dɌ��ԗ��øy�D���[�<o� p��ͽ���F�\���&�M9��2W�Cl��QB��`Uİ�:&{}��ފ�X�����xy��m����g�A��A���`�F�Vyv~vub����3\UT��<I%��Q+�2D�J�7\�(�ch�=�W+�!L�}G�%|Oq��!�`4�?Y�iC��h˝���`�C��Ƽ�����Q ���>7YB%p��PI�#�3��2��.U�[���#W����l���	ܦ������-��:��6N���7��i�"�ǈ뫋�fB�4H�:�_��xv|�[L8��k�{��œ'O�� �Y��i����j �ږ�W�^ݾ}[�����Jc<�s����+�_�T���C���	_)�����
�������"�)8���S�����կhj��v�;����˼
 �eٵ��nո^�?q$` ^�+*�k���%�~ctSQ�ݶ�� �]�Py�.%�ڸ�c_�mF8��~�O+��&�'�J�{����ٳ�~�����U��_�׫���T`�l���k_]��{��Ȏ�eH��̒ʹ��su�U
PQE9#��K�UtU`���e�U����Ow���ի3�����	&@dv/�_l&�ErjYn�JeL�e8�4
�K�{�PV�c6!��&�W�8A]�^l�D��������h�P[[[�"���.��cK���#lm͔s�wƦ��www��FD��<�S��b�q=�W��	7�&	M��@+3�se�ij�#��T�|Z��ޅ@����Y�u!�w���-8#�R�DV^�t��(V歷�z�����W��z��!��ixF��ǖj8�j�$e�:�e��C�N(����)YQ5]g�$�ެEmt�.��Tb�|LS��7n܀`U_vJ���m1��/6&L����0fVZ$3���J��R-��$8�t�ѧ'B�-�`U5yv�X~_o�
V�7*>QU ��{�z������*sYS|�䂃z/�y4B��O��}=�"�5V4)<�Ut:���p��6hάN�H6e���"%��ӎ���H�,�5��h�V��dUIn����w$W�����$ZaF�&}/�`X����%����7ȇ���]��o���W�<wA�T&�,yQ��ͦv�.2�����2�Vw���$�}nw�*���km�=�Q�#��%9�h�r\B �o>4>::�o+���?�ַ��,���zQXZyv,b!|�*�D��b�a�O���f��F�6<zЏhAV��ˇ��lI}��p���)"��>�ho�;7o޴��d���ev�H̃w%N��X
_��4L���х�Ĉ��w�rA��m;l���E�7�������	��v����7�J��� >۰fŞ�h3�~ci�s��[G��:�2^UYw�Qe*��ꒁMh����)�(�-�n���sܞ:p��e:�	�/c�g���Nz�[��w�AG=�R,3V�7�]�CZ��>���;5�`�(��YZ(�˼C�yx�)���7o��;�8���g�^]j�p�,s�ś�k�i\)(}D�}z���$_*�O[�y�ƸwrBH<��)�_��~���=v���>��s80�7��9#4�����{p1���/��Պ(�O~u�/��/��{�$2�q5ǙV�{��t 9�u�ٔj6���e�x6�Q6�^}eZ��&�c�Z3H�b �޽{��}-���!�xN|+�D&������ѹ����r49⺹MCjX��r&����h?}�t�X��1�n{���8Wb��
3�
�;�s	�+ѵ:Ȩ�Lr�t���t!���=����2y0#�4�	G���\�'�ѧp_�c���"_Eb��t�"I�-��q��{��Oݼu��"YF��=f>� :j�ځF+J�����[��]p�*�|�l�`ZCR$/p��N�=ï�ϧn��X����W<������`�E�r�8v^�^�c������1Ѡ�M����XU�5_��ʖnBE,5H]���A�Nɓ>���N�Tooo��olӃ����(���w�G�6�3��͠�w����0KR��:��_)�L��j#h�M&���Q�\�~܃����0J)��d�J)&+��V�Y��w���7���3F�����i��?�3��Oqz|���3����uq̓�E)O�y�n`J�A�����(����U!��������U�ln�?��?�?anT���38�?��BZ8����G��絍$[��Lx ���SG��C�+����m�R�)����Ԃ1��]�w�Q]$�ϟ?�l!�X W^�6Qd��{�v�3������S!�z��@5��y�	�D��O|�zW+��,����	�?�t	D�,��Ђ��j)��-�Z!Gy��h^���$L�WTWk):x�	h�h�j璼u�%)tH)	�}V��j`wViK�6��9���m��ԔM�vX�S\��닒��o!��q�.��^�t��l(�2{bN��f)̛m��׊�ۖ����L*srN�+�BSx�S�V�I�[?~���
&vNhK�&y���е��Av�i���˵��������Ҹ<t[�.J�Le������@+�y�
���e�����.�W��:SJ8
��6��2Or5"�!�(l�.;�1j��l^�L��_�V0��n[���q2�U���!Ic:��2����~}|p��:H������HY?<����|�.�S�2����j�VwĮ>z��]�}J7�JY��uҨa�=&^z���^���}��ֿ6��И�� ;�%��i;ƕp��ze�	��`��iY�a^�Y-��[.Jb ���~�mD��/�N���e�Ža�~�`k{�Ei�E��4K!d�/?-2r̩t��1cuq4��l B��`���D�h�ͯ����-�-�N���N��ujMOv�L�*��R��DH[�#�[�������|�o��!�11�������`�i������@��"�zu��k{ԥM<���=C��z��1�N/�d\����+(�)�	�Yf=J�y\&8�]�T�L7���4�Y�\��}�SP�"�����Z�)���](�*>��8vۖ��>�} ���H3'�q��_��?~��}��?�l�����oZ�\R/����g�Q�heu�,��X���5��b0X��2׃Aed�n�^�S���5�g���Y==;��/�^����~��!rm�4��(�M�X�n�֩sz��͗�R���,׾6���	��<W��'��1̹���pe�U�Y��٠7']��
3�e滑2/67���M�sɃt��ܲ��+���vR�4`���jÖ�Z�x���-[Lc�l�_)�����Fd�tǃ�ed�<ǌ$<�L��$�S��0`^p�\�����rV� &(,a.t�U�d�,��̣(�e�q��>���o��o�In^�'>'#��^�UK+� X�I�Av(/�$�����E�E��CW�ߜ�D2��4�<s�2�z�f�8��h0\MFJl:�a8�7V�r��ETc[yX.#��E��$5Ìہ����V�f��l:���aB�F�ɬ:�&=5ʚ����F�����0��W��P��K�e�HA�ڵm��׸��XCU˩/���L����N���c�%ab!������l�>�8���3���黌�qԣ���(�$�0�eoo�h�I{�ȍk��!��'-�g�A��"5���mzd�:Ma����[vRi��
&v�qs�Щ�"oBw����"U;�$�m#�R�rڰ��o���ˎ�WBerTt?��_�����Ę��р���|���4yu�"�����ǣ�[TVًz����G��W�^]^N���-�gs?y���˗���e/� SIj���{�q�d����ԮyU����Co��d�xn�WX�~P9M..��O�D~�Jښ'r#
����%�.���C��P9/_2�vʻw��%C�ͭ�h+��LVώ�Y*3��u���h��ƅY���0�!tkk�-)	�����ϟ�f+�d 	_Np4Qcj��=h��,���1x�G&�{j`qJ�r��,���K�˵�u���l7��cɟ{AB�em]-� WuC�eڌ!��r�������7��t�z0�����e��
{�X&��>��̓r}wkk��ޕ�\L/V+��Im�O���7����/?y¾��]�WaDbH�1����oy�2�Mg�%9/,$fao���j��lz��͚a}��f�ƏOO Hwn�-9"�s�\cϝ qǭ[w�}����?��X�}�w��������j� >e�]?R$`MK�g_|n����?���M�tt��ER�A�>�d��N��?���_GH���c"��?<�wi���\+*�q<�����9�P&F��[b���+ Q�������7�,�:c7���G%�6�����z�u�Rnm��gV����Hd�J9�j��֦ks�x��!Y���b6OH`b������~�́E*�A�;9�q[���{��]k6Z͑�x.f�x��j=o8.�a����K�&������4Y[�4S�@�+��Ub���j��0����LUOe������yV]^LE��3�	~����[[[���F�����C�RJ�AfCM牅��1������,��~��z�+p�^���Y7?�������Q/Ej�p�HA��p3��p�#bD��3
�=�~�b��ʹ�����NA
��Ѿ�5�����X�*:�_��,F-,d�8k�U�s���C1���'k�l��`���/D_h�_��|��Bb�c�'54��sr������7��
S!�>"�z�v�F$L��5�O��:����PhK�p�5��z�g�4�(��)�O{���Mת���`W�e�+(6��\D���g�F�j��H3ȍ��O���`j{e�q��c�cv�x�l��Lz������t�[�ϲ6�������ww�{�k7���>��=]�a�^�1���.�QF{=m%�]�(���Ğ��}��dE�Ze��U��	�Q�H�����?���߸��m> M�b��y�������������ۚϗ�א���v��t����f0lݩI�M�YIo0.�X�����M�y�����:A�p����L�Z��$���%��d��C��J2��wp����ނ�!c����#����o��Q�iJ�rbx��h+�3�5�dw�OIX[�h�
.s7�D��#�:��n����l���ʠC5nX�i#H!sOA�,����{2���d�S��@�2ɖ+�}[@	|���R�I�x�q.��K7����Ħ��d�胸?�QAX���q'Kփ�K�A�#P8n9��4,�&����(K�w��Ԃ� c���>�6�e�XVaS"=kf�dI����#[�,$l����pRY)�@D`j�u
��`��p0��޺ygz9j���Y��p�� ��V��\ï��h�~P[�|q�Yުe┑��6���c����;=c�Ɲoo��U��y���4���9�]�XuP����ۖiuR��c����ү�7� ��.픥&���t��OkJ_�5����m�<����G���Z�4���o���q���/m��(Yr5m�r�*�R���ke�,D�@]G���	΅���;��ε�[��.w�^���r2��_͔�n�o�ťQ����۳�t�`�x���7�bz���E�(nLX��M�g���5α���z��;O�U)���+�J�������1C�(4�� �$$��o+������un:�ml�?hOy��g�0"Ln-�n,kS�0�$��;�6}J�������tP- �a�X�VI��c�>z���c�^�ʒ�8��}�k�1y*ꆫ��d0�@[��-3S�Lsۉ�Q�5#�U��l�׶��0�ǯNXd1L�	dd���-��<~�����ˆeO�@U¯.����_ɕ���vw�}ꪘb�V�f���[�����!�2=`'"��t�����$� ��ne��](�<׀�J<a��9���E2,?�0o�"��v-�g�֌V)t��sPAT������Ouȕ��@s&3�n���d�x@|�|97�Nt�v��H�U�1��Xr...�~���R���7R&s*;l��;Y�Z%s|V�XN<��d�l��`G �����(�W��ByMV�|6\���"���%�e{�o�f�J�i���v��:M7^k��ז��XjU���Ç�יIO����!�p���5�oz*0�:�cT��հ�Xp���ia�>X��r�ʞ��u�����]�7W'����k�Tv��!,Q����O?l����W��Y�b�l�+��<�N	
4Q��<ݧ��xj�D��(CD�e/������mn�x����[[�VQ̌�E��ͷ)���V�#d��6�CM�5��(c�6A�_�F�𝑱��f/���фo5ē1��Cp�����-�V�^�-�T�y�QЋ���f6���4��<a #-d���)��aQaP.)i�R�WP	��(6��F3s�._�w�V��r�&p�8��P V})ʢ�DE*�c�iH�,&]J)&9��WqNwww�W�w��G4"64ć�J�����AJ#���H�?hg/��qj�SƁo���dwq��0��B�x�����HA�pX�z�{���'R��+"���Y�4,1 ��U2o̒�^X���5<N���c�V�����A�Q#���T��
U]؊Q+n��X鍢�pl��8NG0��*3
��O��9.�/�v�V$q���������Ul�%Q��6��J.�amL=�?��6԰ksN�,Tu�Z��%۲�~���L(�n������d�%�Ȫ�5,UE']-|�k�^���+�G��v��mf�'��xe&�g?�����K��FBeʲ@���xq�<�D!!`�q/����8 ��{���O"�[I��n�Z�k���3B#��!��6�B��*�N;�\�F��ظsh�i�޼�C�������߯��w�烘QDֱi�Ц�����b��)�5L3�����s�_w�]�"��J`s�R�t��KU���TrO��sEE
s�d(������C��D�A�%b��1D|���&M[���ٲN`Ȭ�j|�tS�����-�/X���;;��@xJ[�U}�V#ÂYU�|c�%e�j#xFVK��%u��*�7�.�q������.��<e�圄�ۻDOx��':���2t��uN�E���R���c���,� H�e.���t��5[����c;��$�������ݢ~�o�y�]���M�@�D!�_�W�����ٳ�WGQ�M`����Avw9K�*׶�K��I��M��#�sK�u�v���Q#���"s(N��s(m2X�WOf35��R�C�2���Y�P ��a/R�Hyk�����U��!�$�uvw��6I�yv��`Lv8�B��6�S^��)��dYISȹ5�;XB�aa��D(�A�M�&�	�qg@�z�%d���&�m���wy�kmYG�F�-�U�$4��M��z�C�Q{���3ƨ`����b�*�m�ԛ�{]iG���1�HĽ����ұL�!Aߐ���|e`�����Cҁ.U2!:�pjp̲'��x<JS<~R���O��Ϲ~}o��΂��m5="ŕ��g�r�읮2����`˖��+/��������ky����lɱ�������>�����ݯC~�5�[Q5`1������Gѓ����EN��خ��I9�t-�;�M�c���,L�h��BdOͱ�n����	Z�ONa�w�����$K�ºI�P���W��.�;}e{��]Q�;^�uk���3Fd\�(F�\�z�aÝ͓�y�T"�0>�J�$�M�-D��`�3�d:��.�i�o��)l�Y\Lɚ5�/�EtF�U��R�����n�hG�-b"�;�:�Yt}O�@��A_�O����.�:��k�*�d&5ItO-�̳�[w�K�P���˵q��ol��G(�ڡ���Sr�Κtcղ�u�����/co�dKz]��y����C���6�@!�(JA�V�z�CV�"��w3���P�E?���
ڒ�0E��%� HP A��F��;ߪ[�9u���k학��[T�Y�[u*O���o�k��hZ�b�+�(N� �}Ӊ��	��Q��t� ܂N㨑��+�AE�e��"&��a��\V�ϙ��|���˥�71ˊ6��Y��>�������h�q�9��/��+������}��q�p?��=���k嗕L�W�A^`5������f5r�\��B�T�����V�����۲%*�@{�`p��T3��Rn
v���vwq��ge�e���G��0G0�6��p`3��g�V��я���e�8���e�ru�ƍ�8�Pf[��t5;����O�̞�Q����.�'ʋtg�l��[��M�s�H4e��Q�K���/�������e:��zr�/á��1�:fz|"�j���"	�P�
VIX�+W�I=�	(�d��;����e��l� ~���i���7��x
�<Ib�!��31z�u	B�?Bp�p������'P�D��+����t�b~���h�aG��3ֆ��.�\�y�M����ӳu�P��+ñ���t���#N��g�Ĥ�sl|sC#�X�����H�j!r>�M�#"��ʃa�nQ�7�ȠmnA9F�)��6�J���u	$�r�ٙuSr��b�8888��"�X���4?<<F���H��A�3R�5]���-�-�����~@:��*���[DT�.��W܄:�f����*��Q�§X*�MF6���^]\L�b{W�!ԧ��ӌ%%)b�e%<4�'�����'��R�W��c�o߾9�����d�_����S��5u�L���x��́��O�%���m�h�2�AwV���h��N���[z-V2vV˵K�>�G�:沓�Ʀq)��)qr)d�ZH��&�`��C��{�'�����68���`Y��������W�>�������$vs, "L����O��^��-�g��������l��3Av!T�[��ң��R+ƫ��>J���5�fe�]��*gy�MG�5�7(O�ą�#f��lt��8��*S�늽�f��&A�B�k������>�Z����,��:�q(�cqRZ��Z�:�I��[s�k�6�z�fi~\v���K�nj�����U�Ni]t�`)��#�g���~�{D��ZS�����"}�fy���C'?�%u���[~��pr~~���c�4l�>;����я����W��W߸w��Mբ��Gu����|��	�����'O�M�l�/R�ƮWi]9���CY�ʦ�{udВVQ�A�(�S��x�\{X
b�������޽u||��N0�u�q�O沎�uw�-���'x�[�n-W$�e:��ٜ<�䓳����_����{W��Q�� �X���6/[b[�䟬����d3
N�]��9��"�����;<::�ɨ��ݺ�=_q�7)LH�;�8&�؎������#m`l��A�sN[�!Zħ�9�@�E2�uN�Can��&��z�h��N	Y\̕%7����Wo\��X\�z�5��3'o��6���}���Jmx�[�Ѳaw�x4"s��)ǒ�.;��ݻ7����0����=2��5=�N���mT���^��*^Q�釧n=�-D=���N-.f'gg���K���߽{7_��hG��L�{�����O����={f<b�O�>�;��/���G��h2�����=���l���_����P�Dr�)�n֐�fF�TZg�{��Y��hh"�V��
���-��
_��eӬk�t���:슦�\:8���PO�Y��	�"8�v�z���U�23�/��YN���A',��g
�D�d>��-jH<���t=k��(�ʺ�}Y+�6�	�Y���"%���2���5�il92���A;�\��һ�^�~��7_��~^,��C�+H��)�0,;�^��*i
��6��5�6,�N�z؝��܄~u�Ӯ�s��U��k)ҭ��/�����=|�|z�<=�_��d��h��//b��h���oY/���(JZ�R�N�s�P������u6m��$�5��XrAƫ�#��s1+92���\��-��fݘ�0F�x{Tu<������&�,�Cy�xXE�P�Nvok�+��0B\C�9>��5�`�U�|4�wa�Y㍭0N��yE���D��
V�9A�%);��)���N�V�������(�+?�Fl��9�!�/�ʰ�0g.;l	��!��#әR2O��6���8	3�$���ѩ� 5� ���q��F���ds+/&���W6��ӧ�t:��M�0����#�E{W�e|��X/�R"�; .X7-��ǭh��y���m��f��f��qh���m��A䊫A�B�A�ܹs�Ƶ=.Q:/����t�A��e�e��U[Ķ�K�(�����ՙ�8��j�3�q�	a�K���>R-�m|�.�:�_�A�����W�?ܾ{_�]��9?����(]��e�L���<�^RW�'�4%��(����I8�4�I4�c��e�L���n^݃�Ĳ�M}���Ѡg���T��N|Z� ���Q��t�h��Obf����� �9�"��O�K����z6��j�N:�ԫ[����5Q���e�*h�a2g׋?Ѽ�9yʘ)\��(��&Ky��<���t�X�L�����~�)�~�N�������nS+-Ȓ���Z�<��p�O|�I�����s|�{̆�Y�Ԏ$��&[��l� 2�j��1A)%nG�S`h��:S�a����V�F��_V�91�nxxx5�Ká��<�,rn�V<�9���>�a�(������+��%.f5�8]rY�D��
Ǽ��YA�f+II�������2U�Y}r��!�8`V���'{��U�a*�#�h8�L���c*�o{l��{�b��ܦDD���q�Ԣ��h����v�6�"(Εő�W���^�%^�_��Eph�#�!9��Pm@f� ���r�y�\O�gSv1'â&w-7����^B;A��[�q�#>�],e�SP�e���d�x���+�
*���ƌ�b��'t�s�@ɇ�BJ�(@�L?~�b=�����&�v�,3��Q6���O��O~��jܪ���s��M�#�+}c��ܘ �2�G��e��)�������}��n^"�^>�8����˳i�>�ݿ������<�?��C���}��9GL� �%�-�(��[JE�n@5һ�)R��MxQ���2)N"d��r���*N:���b#!I��j<�m��"7T�P�� ��r"U��9	t�]������]�B�}�*#���I�=-�R�E�vK�Bg���1"0���O����t������YB6�;�RR�����0�2��2e���Hg�&�V�X�%�4��3���������(�(B�t����|�W�W�ଇ6�-V-N�Qg���R�70k�J��S�X��Fe}p���*�wlg9�ī�"��y��[��E����l_"|�8�[q�*�l������1'�xJ�k�[��9��${�H�=aN��,��xR�۽���+`w~􃿄�X��/L��@a�|��$�u-q�jB��2P8��Ai���_���u�+�5+n 8/�V�y�'O�ܺy����	�k�m�%��a�~�8)8n^_����嚘,̯��ݎ�.#��6�ox"7�N}汯�^�B��#6��n�����NdIa�:t(]�������JbF,�e���vMXMcX?\�c�ի�w��N�ZF�E������n���jn"�b�c��M�n(������2�+�v5��B�2�k����>H�kpp[J����7֚����@:��8�\��0�Av�j'�9�vN�Kj��}(<뼇����2�q<�����۷��e�+m��ᲱJPnZg�=\+����߸ޣ��z8�RU*�����R�r}����I�X�d$_��w�=��1���[�����j\XF,��Ǹ2�ϳY�|&���qd�C��W��l=T�'<��4r�f�&��ug�\�U��W����N���6k����?c������W_��ik��cdՏ��{&��i�Wǁ��QUL�K-;"��?i�V{Ob��Qޔ�?�����aC��ojc��"�!�c-�5��p�6�/5�mey4hh�2G'e���*��&��Xe��&�8a�3�M��W����<�l��s- F;�o�����ʵ[��݃`ʁ�E����*�)��:5Τ���,[a2�]X�o<H�>��L��n��|��s2�-?�Xl�^g�,�u3864Y��&�d��w������=�(Q�,\���Q@��+�W*�����q�ܭ[�?z�+��ǟ|�	�^C8���y�:�y��,D��;>E�0gp��<�G�K���������$�9X8�̆*Z���A��q.����5���E~�$MWX[c#gR�19��+���\��[vsc���_P���ׅ��u�i+'���4��\g�����$p���T�g�/B ��s��6_2�e��2#�ö�g�G�Oa���������S���s]뫝Ѽ޸s�W~�W�c�Ԉp|&�-�B�WMc��4^�N�����P��Ǉ�hGN[TNC������f�8<��3��ӓbǧ�m�aY{���v<]��ܼ	�W�|:bä�wh��&m�^�����N�������Ç4ʩ�����i5�������W:}@]I:�ZG�P��w&eh���.5��("�����p��b�s�՚�s���Bq86��f(��'C�0Q�ΖŪ☈P5�	,���O��!����:���j�j$(4$"}������ݖ��Ƀ�U�'��kqlvA�p]Oj:�O�Bp-�E��x�S�m�IO��MW[�f
��)�Ybs�B��
�#2�кX̷�~�ʵ����<|��Fg0��re���֤`�r�t�P�W�(-��s̑���$�)�Z�R��T��O������,܉�h{s�S|Q�d�c��,ք��Mm�zz�ύ�;Bg{���0Щ�I*1��m4�\+������`U��!���#a��ܽ�<���Mze�F=H���ь������䬖s�jp?W�\��❬2���-���D9��>ѽq�Ư|�8��f�����g8�ԺU-"?՟�#h(��q�l�~���]c�^Ze��W~�(��6ra�W�w�y�?}W�5ܚ�bЊ։�ib��77,oH����5Ff����)�H�ϰ�T����}�J'~EfҘ�^�d8�<�]pX���_�	ٝ��c5L��pu��ߥcBޕ��f�+��Dz���������p	�)^븪�Ѹ��^{��4}�>��6T�t�9�2k+j?���r��n*9+'_�;UW��gD���j�R2Nd�
N� ���nXpi��2y�uW�j��_F�����1�
(�R���۾�"�U��>�b�B�+WP����77�Z��
�����7�R��܎��r]w�=`�7=���Ԛ���}��'J �V���`��O���9���ʶ��{`,�xd��g��줫�AJGm�W�0�����J<�p�UAu�4�RL
i{�=t����uC����]�n�,Q���a�����KM�/_�xc�ٝU�����ݿǕ{_7n��9= �w{w'9x��b�(D�;㝲hkF�� �<x~z�����g'�gN�R+����e]���
<�A����i�Fu�Y-FB��� �&�Q� ���~^��짫6;��k.I���c 9�X=�a�6d��S�#�^6�4���j�gt������߾}
���[~������Ŝ�.��s��c�m�z��W
�K��ei����^�Dǵ�؍�J2�K�f���2��e�&�!��2u���W5Yʲ�G:2�X1\�݈��<�ԸP���j) ���אB�jzQ���ȏ�O�pcY�����<�l�r1��Z֚�7��]�dl�r�O�)�<[����G����)�ZA�kW�զ
"��!���3:I
�A���j挲r{;�;[;A��⬜?}��3�!��
ھ�p��&I')��2��J�G�&w�r��x��k������=~�t�l���E
�MC~0�XR����-��5�{����5�6>�!]s�Z�#1�g�q���P�u��dx����zK^5i�������^�T%V�ɼ��@��NX!L���]�qC`i&h�3u�!���$�[����gL,@�%r����0��X%j����{fu0���o}���pϞ@�`��ƃ����Qg���m#+�C��j�ށ��L�|>
Af(�  ��IDAT��[a��QE&H��9E�����n<���&��_����i88L+��<��`�Ϟ?)8�b��k�TSg�O~����ى��$�^\����1�ۿ����������Ǫ�oz8	�������h�k��������|��'\� @2k�vC�~�[��f��Z)C��U�`$�6��Y��Љ�eB�+��س�8i�<:ZV���Q�{�Kן�~�NW�;ߐ�E�f/H֗�©�Yzx���2j�u���L��5\��\;E����j�AA�@��w���ZB!\�:9e�����H`Ʀ��?^��6aa}����U��� zζ��ƃx�.�
�f�|�}�Da���ph�q֙�<\'IBڎ��V�<7�K�5Duc��e��U�Yn��sa�J��M�(̪|d�f���l*#ڴ-���i�A:׮�T�>��:�k��4��ڻ��$�F�u,�4��0�s�JT�~�ޓ�,�TF��/���4��aQg��i�������僃g����6�*�B�x8P��)���7P�yo<Q��x0��ڵ;���uZ��R�4$W77�="�ac�Xa�nݼW�H�[j�|A/�35����Z8]�����#����BDS�q�(z$���l�L_}��a<ql0Η�z4?=9<<|��v�֐�p��=v��V! 8'���Ƨ3H[�=2A�I+�T�!�C���'9�A�!TLnQ��G�� ��M!ݍW�N	7AvU�D��L�������Z�J��ݽ&/��0�� ވ�'���)>
+^7���K������X d���o���6- 4^��+�u�zY��ԫ�"_�8~?
\�c��%�r��{�^!�Y�lJ�h4P�,�>��02��5�1�̝��������6��W+��Ւ�Y��?f���ֺ(�(.��?���06����~&� � ��ٖ;n�����Ϟ���$0�������p���=�r]-���1�s��c'	Wu4ŋ������0fgU>��y�>�rKY�,�L/�ٟ�-��Ζ��W���u�5�۽Zظ�,+*�נ)k?v�\ٳ�J�$����Y>x���7��o�� �,�l�l�7n�g9D�i���aA�:���Jqxƍ�h{k;�5�ڞ���EE_KVȹ����"�5g��}o4���'���?���o��?]b:�A2(3D����Ln6�_E5_�&#^m:g�)�Gw�޽s�u,�r9��:=9�::����u�-�
���_+$��Y����|z���^�NO�5��!笺P�ԤP4C�n�k�������i(+�+7������d��t?��+�~�r�+V�J�O6&8���<[����YJlg���
ߍSD'��c�5��op�g''�9 q�������"+� 
�����0�n���j���k/L��O���Z�lK��Ӄ��[��Pm��uWs�"&=�I��[ono��� �$,�:���:��օҠXX��9��zqrj�Kd	V�Rc:L���,��k��J&�3h���A�Aʝzyp���Ӈ��8�7�m�������,J*7�=gx��-뗮�Vs*D�LAI�¦���X�O^Ԯ��5(*�-o�����童�0˩g`�E?MԉM�k8�|+�㚗���B���z�-`�B��5� $��ʵk�����V��N3� �$N�*6�_�5%F��f�ἺH�g�wv���rN��US�P��1��b%��֞D���d^۪5��bw�\=}��zAGN�;�b`q�s�ƣ�2s+w�]w m����e�b�R��f0�D��V��1%�z?fx��ʈ�:Atѩo�sv{w��͛�^�E:coro�H���Y����P3aki?�/�l^�s֌��w7G���Nx�✠�E���6���H����m�#�pr8�y�b��g�UB����)N��rX0�:n��K,��G��3u�L�h��p4߾}���ڼ>�rU�?D��� ��ɢ�}Y.2hcz�[�*L��ۦ\s1�$L�EN<�.�"�l�%�c��$���� &��r���I�:���n��z�lU��r~J���,�q�19�������JW'�����$B2x��-~ 	�I�t4��*t� �F/�5׊��b�������@�U�Q�9�d����h�㼚�9��saF��p����h�.-�U �3�#�;��p��ʭ-�{�w#;^�x�؁LuXr�w�.��r��O������xc{C�8�Jbm���L��H�S�0VP	S�<p��Ȍ��rk����щ$ڶao��-QÀ#�l��Yl	� ��!�m��s�@uI:-��0�uY��a���n�K�_�l�dL \K��j�d��wV������ok{È�xx����9E�X���n����_n;��3?q��.��	��@������n��_�uc�$�V�QI�'�uf\V7����q�k��E'A�Bw0r�Y��0A ��0�[H�Z
�_�O�>ŉ����
�mm��XY��i�ٚ�K\�d��rd���Fb����P�Bp��}�<�����Ɩ2����8��ɭ�[ַ/	\*�J��-��c%�X�΀��Q,�R�J���ڰ�7�m��u.%���|�K����~����L��ƀB�Y	�" ����{�̳�Z�r��5����0����9�꓃�]}����W:-�!|�V�}�o�ԕ/�z��{�J��x���*p���H�(4Hx:�%��r�
�l��$�����9=L�  ��"��I�5a��d)��vNN�.��6�2�X9����g"P�/��JMc����X�V��j5Ck�V-W�	��B��ֆS=D6�l����?��w������_�����$DU��4H*%�nډS�Mg��F��G���+��%��*/�V`#L�o�C]V�����WU����_�(�U`M�(��^H�9���	�W��S�DN�*#[|���S�IONN�6w<�����Ϳ�_�q��/��/���/�䏿�(F��ب��	v�eW�Q[o����*9�Bw/ʹR<c����/.��Y���Iw�Z-�S/��%�H�~�n�������]U��Zs-/V	�^� ������]��^�5��۷oܹ��}��V��o��oa���?�g�����Ԃ⎭��
i�X���v���HiiS�G��r��^Y���P)�Lъ�X�@Oڴ�Cm���$�{�uS�e�^h��$��W�~�p?�VNہqN��D�x�#"��p�bP2�:Ox����-Rhv������у�ޮ�gMD3�K}���g`m"��Ȭq��a%�Ŭի�g�Y)E��p��JO,��pJ!�V1_�t��ޗ-LO���s���(Vqcy��ٟ��7��M������a�<쁚MҜvru��/��o�������~�'L�0��>��"w[^�Jb <�q���A��Y34�&�����(l��I�4�&��sݶL����B�{��u4�8y�&����ʸX�p6��)�8���>ZʌIT��{�g������?���g��]Y3s��%1�7��87��s:^W�P#߳�5E�f��Q�+!vUBS��ȶ���5�B��ٓ
Q��D\a��,��J3�O&���` J�m�@��rS��Ν;�.)oݺ��C��9��X"�N9���{��e��9�^�Ԣi.�DP'/h�y�=x�K�Ta����V��u�?� ��o|G����8h3����KCʁ�8��
!�N0�d���Vx��jm�6�Y�V�č�R~RE5��߸q#��ƅ�cq^dPx.R�z��-�Q��̷�	#�P�o,tXv�R�|��n�8��p�6P��
��UwA���nEF������1�=,��WEU�17���E;�Q�u�:�0)����g���/eC��o�9`O��5�(����,�|�U��0�j3�%ï޻G��}�w�O�N�����F�w�R_KiB��jځ��1��+���Ǐ��$�㍖����\�~�M֖p��2I�j��D����NsU$W�R�U��{��D��>���ܹS�1��ZYm��F`}4ީ�(�yI�3�q�u㊨��Z��U������]Sj]UU�1ځ\FJƥ��_��a�897�1B��r:x��Dݏ�G�p��l����<z����n�U
�ղy9�O
��r�H)<\�_S�-lV L�������v���Q�����dkΛ�d�ۆ`j@m$�]����1�j6!�N���_߸S	��[YR����+Wx�Hf� 3�y��K�xݧۡn��1B�6�kf�i=�ѣ���/>�>�8��D~��B�"�=�M��A,+W�ߘ=[�0���p�[���c)Z�c�nh�̦�
3[U��qcS�A�Q��c�`{�	��}��x�Y'�G/^��0<�t�k��Yae��̘��$�r�ᚊ{�1$������ۿ��Z`�˗'�(Գ�Vi紒��ΊbR�V�ftB"�"����B�C�+�,��ZB^�ju�ߐc�V7�i3�f�JQ�"$%]�c#
�Ŧ�	VL�Ň��Y^Ğp��s����1L����q�U"l������I�É���M��U"��si�4]*l�	���\u���N� �gm�D�TI�ɒ�.Z�6�\&�� l��h2$���M}X�NXi����*�	��vA����R�����Փ[�v\d��֦o
ԣɾ(���U��;?� 
ޠ��y������/gBx����s���?W�E�!�xe��}vS)X�����Kg X�ppܿ6{������u�'tcl����p���p�g'�3�>�[+�ú�� ����x�T��~S�R�\)�*�H}��k�wW�"26�m��O�[�	IC��꒫�ɛX�_����?�N�j�ч�`˭\��k*�$��7vl�C��g�"B����kj���l'�[��qV�:fP�k�9]��ӱ`�+�3A�+�e풜�1F�Ϻe*}):n�2���!A����|����4�,T�<���w�Ѐx:�#�9b�(�%��.��K��}����r���O{}�'��N#)�7�ϫ4�>a�߰������I�h�>�F��G�*�Xh���Euψa�6xZ9j�W�Ez��6~.�� ?E����Đ�>�T�3�^Oa����Ѐ��d��x�Gm�4Q2�(�#�9i(w�a4l[����M�y�'�t͔��\�e���^�Y�<;99"u�5[}��k�?���˿�˿�?�/I|h��4-G^(��|�W%WW�t����n�0�ŀ�q�q5^ri�:�غ����GLi�����8 !�U#w�)�0��fd��ԏ���g���u�����*�)�Rl�"�l�HSn�%X�����|g�� (\�ƭ[8~��k���o�R��w)~�2�����Ƒ"7��L�tPye(����@V�#��b)�Yf*�k��&7*�����6_��Z��^B��.AQ
��cdL5rs��(�����D�jT�c=�8����/����?��?��_��7�,Q�_����9��;�=�:��i���b-H�=�Гo�H@��T��ߦ ���~�?V�����dH#g�SU�9�٧�6�ay��PB��|�	��_�Ӝ�'2`�&�Kҭ�wò��&T�#�tc���R�jZV��۷����1��a~��'��űT%b���3�{I�`��]�p���Wr�uZ��� �X;+�&LPh�<�w�������O���l�	���03�%�1����&���)��L�Fz��n���UZb5�����-��,�hP������W���A .	ǃ�ՓG�z���4[=~��֍���-<�?�G������[��9?�
f����IM@�����v�+�V0u���2K���HY5?���鮗D�s���福��S8[-dcm��j`d^��9*F�r|t���&kkv�b����/.����%�o��������X-.F�x��gG�/�}�G���w�-�Zo���f;D���X~��M��Έ+��E6ZC����a;�x�r�i��I+V@��
H�'��&y�S�\���ܫ����E�+�r�f�D�L��鴜rN_�n��d�<G����kvv�MWwT�5~|r��Og�s��,�PİK�q��'GJ����0�Y�V������7��vL\Ө�&\�'g糫�n��� �yyNNNKba&�s���Imfo�Ѧ<�Pf̺�+�;���c��;8|a����<6�ve�U�_o��C���A���!!b����?������!������u���҉O�*�>H�w��e�]b�d���[9��]��y~0�],�퓵���NYejF'����"�
��0b���Q��.�4�LW��^3�j����2E�ۜ��n���m��b�8�(�	1Z-��}��{�n���ٌ\��Jmh8��o���'?����v��t�QH�V(E|�7)q�(t�=}z��~��_��_�6ȥ���r<����C��6�ɺ�n)/�h4��r�*�������5L�{Ԅ��g�lY[�lD�8��e0�Bf��6�p���c��u�:�3������l�C�&q������"Jw�J�K[JDe�ճ�t�cU; �1��������/����>�n������ޮU����o�\{A�ǟ_��n�ٯ�d$�9鈐ź��W��An9?
bT[Ωj�ԨD�C�,�Աe���A�]ێ�>'<Fuv�
|w<*�a_(KXazڬC����C��1�۠F�Z�0~��k@o���>�c�7�����)t��ɱ���x��� �j�q^Z�G����`du���W�������������7dZ��rBzeX�V&	IκNY��ri�2�M��W�{j��0��B>e��9>���;�g�϶^�5DDUf������f�0�7n��}�8:���s&��^=��L��5#V��b:��$�b2�&4˕,��F��j� 6��G�|���}��p���ÍHB(��,��k$ʩ���I���bq~v���=	C��hSM�(�ɝn k�^)��0%�oS9^;��Y��ix��WmPXa[iӓӥ��b{_OӔ��Q�G b0z����<xT&GG'��>����bY 
QE�#+�ñ�N�ú�5�LW�fE7'@�y@'�Q��Y�>�GW�<Ai6��3S�{T��P�p"�9(��H���ڵ�)n����m�^�x�s�^fȤ���x2.��t��x8�<x������x��/��rm�5��ؘ�$O���O~�˸��F��HVi��v��[�{9��MZ������'���i���}oj
���]8!ʜ邝u�qRF9��h�W����)�i�|0K`C�B�(��F��=̓�P��N���[nG$�"��nR�?
��a���dkc��0�K����(����gE��&�0��*�'wDIm�5Ѻ�h���:�,7���Js�������fT\~}.Ec�����K�v�W^�4���!z��s&���cdɃ�[�Nц�q_�n�T5�	e0�E��#<�i���#�#k�"��=sp[d.y�� yVm���y-�������(�ZV@0��C��|�M�{ׯ_��_�(Ε��Xe'�>Q�e��v�{Y�@%��T�7�q�����r�����v�KEXw/[�v.��Y�]}�_��4���P�}z�mI�\9�V(�T@RC���s$	x���s��t��z���x��u��Hy�H�(L���,���.�Oj�#I�px�^�ڥV�k�u��v�n�aE�+[���ߍ�s�U�Dc��
T�?K.��됔u;�����w.���rs-֭az�����z!�(��q�
ӷZ0�H�JY�^��7 ^�E�	U��\�:Qpֺ�p��@(
�5�o�l���^���}m=��C�B�o}�[����K,Y�X���g�t#�Duld�.3�tZ'�%Bn�>��d�n,M����U�N�	Π����LN.(��\�
8�2x],x3�̏���sXT�8mq;�7h���������L�<�?��s�x���~��;7Y�*��1,�`^��T�k�����	�rr/Wc��3� =�b�9�ŹI�T��1�ZY<-���F7�|��g�qY��XM=��D�o@�`ɠ��~�m�����hӥ�s��k���=���B����$^,m�wҖ��z�!9������~m_zo�!�����4e�VƗ��a�#�	}G�ڔ:�s���b���݉�/�8G�����#�>�H�E�Q�z����<A�L�C�ot�p�_��_r֥qi,	�>VlT	ڔ�@�K�$�ο���k�����Ó��`��fIn%J����Ϳ�@�����.��5�g��@� Rm�!I/>�X6��y�(�}����X���6�됭����`�¸|�`� V`������a˟����ǯ|�+������e_��W���@�)�[G@ H�;�y�u��)�J���Mi���s����fѱ*�$��S���7n[��%��I_�Kv�#��b��&9Z"q�����	r\������5�B�(���(�!}��'��ɽ}x���#a��6"/�\IE���M�e��00ɮV%8"���*�����wq8D�c��<�S6����EC�5:��o��<NH�k���ȕ����Ɔ2nP�M����8�́*��c85���)V��blجW�qͶ�$�mzY��[o=x�@c�U'�<l���F�#U��ۮO �V���v
Q5�E��l��������?��6�9����;41��mj a)(il7hUR�=��r��5(
�1�9֕-����B���8�<˘�TiW�!��?}�������?����:\pj�n�1��U�Y�%
m�n`8��gp,7��UT��&&m�@i��:7P!)L�^r"�糾�Y��7|ӓ�d4�ʘ;��czN��C��ou�˶���B�S�Y���2�.�^^��I�ڞJ=�2Mk�����Jj�����L,d+FϸwAY�ҠE;/�"gv����i	ɖ���s��W��%�&�^PO&���w����;�����|�� 0��k���0��sa�U���1[�b�hX��P������&�,`�4�{�����O��
)��S�|ȍ��Vh�͢;P�N�� 	����K9���bW�I	Ý�����ޮd�� �A���c��.XZg�eOI&,���ymC��W�s` y��!�>�-w��9��,�t9��8��"CC���x�CC�3�v�G�����Wy��TH�19˘Ղ���f�#�A8Ĩ?�n\�pO���ڤl���VKc��Vt�����$l{�v�;5�K��Ut=�O���e5�%qf	���S�1�_��{��%\M�����b�a�_�u�S�J�1=�+��ؙvlw�_��x�Da������@����ڗKC~��J�j��%#R;�l����U�x��ŻA�Mk.%��1�rˎ�Z��=:�򖵱�l�R3��4�0����o�[W�"P�:�v�6Kѫ�`���Ip1Ϡ���/[t�vi(�򺄵�D���w9�W����<}~_���|����r����n��d2P�"���J;R��%��B?���e�����U���`>�)y�2��J��mp�h4�CM���^Z����W��Ԩ�+�����ɓ'�d��u�h������};�q����Y�Ly���25���M����������X�9v�Z�y_��͐| ��\���ӭG��+�qۜA��]t�e����je q��&���G�vS�Wv]t±JN�nȆy���by��	?!�9k�dXgpsLe�cu5,�Ne����e����ۿ�j���>0T�G`[��]�-���[�>�����vEյ^�g��M7������;A���.�e�"H���v�V�D��ٔ�m�9X��z[����U.��������t��מ�n�6n6�3Y� Ur#���D.=��6�`�f��!k#n���#b��ݻz�ڿv�Ϋ���}�z�د���76�5�i-�>c�5�1��f��r�lUF��:���N���^a�xغ��g���g����\ޡ�C~jN����4\^�G��9�X�E����,]�C��x��w($0vm�������;�;��ϊ�g�����]���\zXu��ٕc��FU^uWh��7Ewo�t0D�˃jh���t�@�%$��M&M�M�V����$m���Km�2-JC��tA��Kx �5�,��0�ބ���У�nòp���q�o�	�gWt�6�r�+�Vb�6+�2��@0U[ۛ��=�'�X�G_q�ݲ�S��$�`݈;8�0�����B�{�^���j��D�6����f�l��ws0�KS����!,�ȌN��u���Y�S�iW�Jt�1u����s�﯎�]3��n�~lCB�^�<�H�xI2��A|p}x�����&t=�>|� ���}���Z.h���E�/����s��3�w+�ĸ�iC�Mg�5S{6�,h\�_�֙�փ٫��2�,=ڎ<�Y%pB�t����C�g�b���T�T5���￯��h��,v�2�_��eTzxv�ǿ�����O��ß��|�>9�<|��[�C�q���v�}�G�������@@
��?u�L�e�PMU�Y�c���A�~���I�Hu�[j�X!�1���t=��A��8�w5h�l�à�lSVnݸݬ'9=X���}<3�^�BX���l��_,]�W>q��LlT�o���l��P���onN
k�������;�����9�Z�K2���l�|`9ӣ�?ƥ�NR�
''K@�b7)1l�Lu~�kе*�U�2˺֜�>�.C#O��
)m�F�Y��F��(�W?��͍ѷ�^-��_����L-�4ŋç�~z�/?��|���[���A�*�C��u�[�� ���Y�1����)v�� G�Co���M&wn�"Sϓ�Y^��_��T�Ч��lVc��y� �����^dIғ�цcu,uK�#�g�7GGG�b�( A�xc& ��$�tYkt���p�#ߋ\�v�Z{1=+��~y�-/f���H"�kT9��3��҅�U���;�/��l�6�E��5|zE�E]���+�bs�e�X��\�S��),M�C�� �Fx�b���Č���4vp���5H	�8�5V
Ңo��I��z}��fTWl�T���8r޺����^��~�������x��^৤�<^1W�L@�Ei�<q�nB5�fp�۷o���Zxpj����?~�\[-�t��M�
���_l%�+&$�/,�������7;6Ԓ�X�����?y��k����}���>��|vA>Ǎ\*%�mt����[׽����dkNb�����O�<���TkSP;���0���J��GX��۠��#�M��C�C>9��e��#Zj��O�Eb��t���y~x���[ׯs�ʚ���y�b��H-�}�U2�?a�:�j�{���yY��	�����*�%o�,�'��������'��u^1��V���������YNG~����^{}f���ׯ��m���`%��q����D�A��ĘX�E4J����c���g�XohF3���l��6靝�YL���b�6��D�N�h�E�S��8���9����X�nI��sfv��Y7��M�q6_֮��r�������!�+����Y�.W���eV���Q��U�)����"m�J�-��H����_�u}4��7n��j��ds�=]�Xr�H���l��Wiu�V��h�Td��#?l���ǖ�)î��c��,��a�Yd��p�Q�|��cuܜ�z']�������&�Uʖ��7쉑{N �@��߂ɀ2�\��{ЍΈ��^����d��ݻ��������y��l:��Q��_gV����Aۊ�ϸ9k�)�Ö����+^�N�9��^U���
ڲbE��j�������7��^�/��X',S]fySN�O���+=��dzT����߆�S���Xg�ѐM$��wra���1��w�["�#&���Ղ���ղ�
y�)Y�k��,���N�(s����
�߅�ӰS����m�j����X.�:K	��4
ܲ��#�M��h���)�&�2�f���#�'(�ᜯ�K���q�-�w�Vy�'r���|�~�"���%�Dlo�*�`gu���o4�㓃�EĳSf�f��Ñ�0��&|ҀӶxx�fezq@��g�ܵ��zaU{����O�X��2���Òf��ƉE�~��g�^�h%"��/��@:��p�A�z%��N��T|JX�m3C,&�!RR�ڬ�m��"$L��#cz��.�HB�h�0�݅fB�38o�ڕ���C7`gk;�y����v"�&���U�P��^mu����c����0O�s�O!D�Fő��$U���d����SHԆ�~6�
�tqb$Wuf^7���(��x�)��L����%��oeG��Fd�zَd!k��GC�dww�e��*N�N��T��X���?���3n}��|���?��Cr'���+��Mqĭ"ԃ�x!0E�u�M�k�$D���}"���s�����6�q�9�����u�򝗳���jm��ޕ��ݝ�x�ǒ�"�����8�{���P6(���в�~,��|��<a�-���Ku ��X�Me�،%
9�Pk6�����'�|��U�GR
��篼�|&x0�	桲
J�
zj�`C�'�n�in�yQ�NuH�p����H�}�}C{�~���Jy٦��4G������	�eۄ�� s2�'κ�*�v'�?��p���wȼ�XW5ͦQ\�-u:d��d��7_�U��>!�s���^+�.�h[�����n:fЖI�˴�\!��J*`ְ?<��iH�;!��
$ú�0R�PFK�����OuiADW�t M:��✗#mH�U	3����$����X�,�F�!NE�7n�{ATp�|�BwMڲ	��^�q/*��l�/l�&�>|��T�6#��ӧ��.~��o���|8����7�GQ�Y~Ĉ�+n�z�Ӽ����ɿ�E"�Z%�N���%��4K����.2�x�h3(�T#�J�W���_7��GD:���M���3�P& iK7���||,T�j��q�sͼ�ͧF�2�����Rz[��#W�Y�v��$�����{��rU�ܴ� �p0Po ����,�y/��v�B=b�����
��oh�Yh4vJE��<�yqlQ{"���e�͠�H`��j�Xd���/�$����������~�̩���^��ݻG��"���Lf)*iq�b�X^([*�~�'
q'�O���Xw"�IԪ/!�м�ROTv��6����3�b'Cs�����?�Q�c�D�P�S���k3Y�ـ�����s�E|��'J����ѣG�� q҂a���Ϟ=�GO��������_�e���������#8�kemi�>��E���bo<�u_�9;�a��}u���U���|���k7�鸥�j:���yGB�(r���>����7/p�b'����H9SD&�u�8 ����p�O��y4*�=����n�Eů�$���VI�+��#A/;A*�nB\aC*�x���/�����G}tu�7��<9@���P����&A��߿�<uc�)E6q�����c�|k�?\������G?�n#�Ys���1.��\�k�7lӧUNͿ6iY�[zL�\�p�%����a5�-[+6P	��t����/y�������L�D�O���=�0G����y�N�)�U��KW碬��<;�W�EX�c�;����w�֭� ���N�-��!#�j;��)$��m8�@V��B�X0�0�Z�-Bhzx���ҦO�<�b���]�V��/~����n2�q$���+({X4��;��y~Ks�:6ܣ�P�`J�R�� �oCC�B1`�8��[Zg�\BM������g8�8���������1G�,��m�t����,�ֳ?��E���q7_��������H��&��p붭��(J��G^'���62�*�ͯEv������N�[tC���P˩��
j��{�>���[��������ų��G$�'� wH�ö��/����-�ͩ�������g�a�>I$T���@=S��;�[�\k�iuK�1����dBzu72>D����>|�NH)��X�!^������3
�u˾5�6ِ� �ln�^#GN�iiD��%8�<"�,c�g"~���z��׿��ML8��b��IふD�b�����i]u�k�BO<�m��K�=�V>�N��|2���)"evl1��1����=8�'��R���U�J����cp��87.`r��}
a�Kќe��j�8�'��>��i,�;���9������P���1y�h�Wp�,U�!��o��k�)�SJ�M^�<�gG�[���] P��Zv�Q�S��]�JT��l[�j�IY��`ʇ�92��K���s���_�ͫ�B����K&#����CUDI�J��d���ۧHz�#
!˅�Q]3�F�ʚ��B��2�v��]f,s8�Ґ"Ih��"�v�e�s�5gU�|i,��V�5F�	nƇ�@O!B(�j�&ݴ�����Ui{�~K�t��k-�0HHS8,�y }d�t��%������y��H����Κr��|ƪ�Q��-�K���%M-O�G�������T��+	:����׵�ri7�W��?��AC�bFհ�Y�U[tקs���� ����2_�vS,�}�NH4�>��Yq�	�/R@E�}ZfiӺ����墔QvEb���¤��	��������$�c��	ܵ�
��K����J}�������K��q
yw�8-�c�m�Д3Ї���_̐������([n�nR���x|��h6;W�c^�X��� ��!7��x?ژ �}.Y���s�E`N���}�0*{#��0΢���[�W�f�Y0p"�}�1&�+3�T���-I�>U\W���=�yZ�J�z���ʲ��-l��������zNh�B\
;��W���z�޼qZ�֢v�x��x`�TJ�������P -!�:��.ع�X'�!UiC9��2s�L�o� N	������Z�a5/g��	w�֖��T)�K�^eM+I��
���{m1�.눃&�����L�S2z�{ׯ���mK�K!Z�N�Y�VF{q�3t����)>K�|6u�E�ҡ�RK����sieZl��(	���V(������Ԑ�_���ln�[�
�nҐ"s�Zc{]�=B[���1���l}�0����d�㇑�(���p��I6Ū|��޹s�����q�=ܒn�ro�騤�,*��(=kH6���HV�·I���=>��c�	�9�����������Yc�̓�zkck��ݰ�U��q%��Y��+���IE�􂗤6�.�;��ۼ�h����_���
2��}�
O$�٩��$]�z!%?G���T$4�����5�Ɏ�Vy9��8�������Fc�x9d��ViT�L�6�ONO�qx׺�ŐW�)�V�܊�����\K�L.V�A��CG�e�;h�^��D^8'g��:B�vņŨ;� ��� ��z��믿.�>���-H���j󬬇��Ճg%cta��<j5���	����E?�3\�xtӤ�ǁ�L6��6������Q(
������Wfi��IQ��F�Ș!�s,ҙJ���5Þph�&��7ur�]��bQ�ȭ/�\�*�7œ2���������%�g�ΰqJ�_��^�3����FE�P]�F����߾��{���u~�޽(��O9+ ��k�q#�ӏ?�:�l���1)N�0a#��[������+hwxჄ�X�ILs�S�asb�uuE� M5]� ������7�u�a���:�o����KY�_
v�P]JNC����*�*WR�������7o�U�n�.��{߅�<?�|��Q�����O�^<z��'�r����g��8s��(l~���d<���tݗI���Ī�ȏ�ѓ#��g[%�Ҭ��ivw ��e��gsF�n��L���$��B�m>}�B��y�{Y�R�����L<�E�r��n����������������H��ѓ��NqXF������3�ml�`�+��7#�L�>�C\�'�0���&�A�я��X����(37�,�%�P�~i���G���曎��TY�ɐ4���	���G��\?�C�1�;��ȷ��.�q
�Ϸڻ(��dnUzN���ZFmwo{3Y^���6�66�4P"볽��ݿ�����l8�3K+e�%�X����W�@�)�M?��k�߃s߄��������͛7�� P�>BcL��[}�ʍ�T�6n��b���,>)��{���U��\-<�z��o�P���~��7&#</qT������|�OY�D��Y���شur*@D��Wi��X��0�PY�36t�\[���R1�⫲��6/^�F4�f���\��mJ1u�y+��J�)ʒ�ӹ��7�.g�ۃ��]ݣ6���L��m�� ��0t<{�����ˋ����ty��~q���W�b{q�U��gL;nl�.��k22m4�K	�`{���h�{��wY�R�E4&�_�O����� �μh��Ǳ+�`�����W�99���k�LO�!fm�r`�!vҸN`Vf����P*�i�4�xd���kd,�S��0�5 KX������O?<:<����UCԪ���[�J�@%�ҵ,��ܾ� Uv�憪*X(;2k���P�2�¢��ҹ~�6l	>��űZ�kX3�ђ���qj2Yg�*fa�q"wWϝ�gp�2Y�h���9̦��_�*��;̋y^�uu1?=x��ӏ>��&`������#�T�;�|jB@b#̻�\��V���XʎX�����w����Bߣ2l��5d�C��\W�0q�$�����d�Z<�XF�m�e���	�sa���[#͘��&�91�&4�*o|7��S�;��b���Y
�*9���1���J=i���T���֍�����z��]��p����G�f�w��Fq�Fk��,�B��:���JM�<q�qk/(獲�&��W]@Ҧ�P�� �Y��zt�;9��~�E���2}Qr�n#Mwv��[�p���*�B1�����&Qe1?;>x����Ȥ��VP$��r��'v`�6�lr��X���K���xܠ�Pv09rv����XFR�?��XLV�	�������
��t�*]<��z��b�`g&�AM��ڸ�˼/�$~���e���V�C��u^����Xh�e�nR��-��&�XP���&�����S���t	dt{Z�������kڑ
��*֓qG��,n��$�X��4��fdk��|�@ b���8{����k�=��Xt,�V
Ǡ��F��&腎z~x�㶿���s]�[j��T�*K{8^a�J��Ŝ�̐��1S��O�u1�P��G����$�.�fA��hd��H��ɨ$&������ﰣ.��*{Al����t���H����D*��7����`8f��&p��M׵TbD����b���Q�Ӱ�]�4tr4���pbÌ�,<�t�J|El�󒽌���E翔�/�Z��T*��BY��1x��}1��+�[��Ѡ6"����޻e6�����t�[����i+�p���S<�T�j	"��1�l�e�q=5�^;Q��x��D��u4?l�Rt������W�1�S;���>��C����#�1�[�6ae��Xn�:��1�0���w;,hٍ�:.�C�5-����{��5mf͢ٺ��j��ꏗ��ˎ�[\�Bv�EYv{��*(�t=���zJ�9�/޹�E<����dQ�bȊR�v�U�]�����^Ѧ<�ڰ�bE<����v�ٳg��s��D1����0��@�#�c4sa�e�:����"��S�^��ϱl7�"7�8D������7T��;��ׯom�����K/�7�(q��|e��'�ܺuK{+��'2��l�jD��m�t`�dE�����ZN,-�	�-$Ks��������*�*훹R�=N;X�w��2Yu���H�֢�h�.<Wض� ��u8?=#B��/N�^<<<�{�կ~��x
����&���#��t����;F����8::��b��"T�3p��h"k�O�GIyxҸ2�3K7�ԕ_z��9��4lFؠc�����'�X�P��8f��6���^�d����-DI�JI��PuQѫ9-�k��?99Ad.V#��?nIgGU1k�;8<tE�lđ8�Q̮��9W����*�W����'�?��������^��!
��[����Dݦ;J:N7 �V���ӵ��p:�GL�߭�o��.�7װj���~;,[+�u����s��M�S+�I�6̺�S�����2
�҈�.�(1���فސ<���{��>�p�c-�sk�Nm�.���x뭷��{��=����G?�>�w����_������h�k��D�|Dp�v0|e:�����Q[Y��R�<�'��z��[�6�TIV^�pǊ�t��?�uL�����a�����(9�"�Y$6���'?���77YkzK�P�m@�ҙ�JX0�{�0wf�)S���[�xa�����D
���9�Ϯ�̂ű�����7k�뼮�|� @� @�����@�,�e+Tv�.��������ⷎ?t����pt���B��l�$Q�I� @	�x�{��k����$H��::��Ld�{�9߷�=��v�ٯ�eoe�T4�ƍ_���qa;r��<�AgL,ڗe��F��3#Ĵ]�[�p|����[o����g���'bc�{�b�������qW����Bj)�2����z2/`����4�,���UKb�;\̙��l�?��VU�t��>�+_�Ja.����HKXge�)����MF��G���w[�R#<5���m_�&�c[c,P\y����V��A��Am�����^?��Q��Vg��e��hݼySΕ����F�� �_�ƈ�6�^�O���y&�]
R��F�xVJ��`��#�\�5�^O�l.s&���ԕ+W�c�� ^��-�j�y��C�Ir����%鷨d�R��T��ޥy�mh��Ѕ�)�C�-F��,��X)n�`4�_~�-�sh)������y�� \����]S���{��
��Nh���K�T���L���9;=e�rq"w󻬵͆��5�}/f�Tu�ٜ��Xv���;w������*����t��l ����������5b��&+����͈3��"�=e~v�`�z�x���x��%�c}�.��;����Ĺ�4�P�m��Q�Hk)V�]w*}��:��,*�S����=����aܔ�����������+�C���sq��E�lǇ~xb<9�+)��Ô��$���ܪ���D]��~b0'�c_�������J�����ӑ���]�������K!��Rw*lpUKw)���|v�Y�=�B�\�8_�|�'r�7c����ɷ��>��2џ�:WR�mw+�ʣϖt%^ܳ˒�����BBI��ed�$���K��YXǅ7X"af��b=����ļL�&�a�#�m@D_x���ql��&����h�&��9�A�%H����ȧv|����{�g֙��;;c���6빴nzѠ{�c2�!�ZJ��m@;Uծ?�^eo��6�����8@�C �,�AƱ�qW���㇜8��M������X42"���_����7G�S��h�u���M&� >=���4�=�C$&e��U)W������5�2q���ڍ#"��0�Ii�6��&��r����v��Zv�΂0��<��1�[$z��05�L��m���� ��Ɗ�
�h��ʲ��gvSН�1K�"��mΘ1|{+_�i�p.��K6���/I)4:Q�����#I�\�%���&��X�դ��b�,D�r�Y�;Ufo��	�w^Q�c;�5�2"Af����5��ݒv�h�^�U��I	�g_�Tx �E��j�GP�O���*��F�Q�N�c��Sԅ�l,�ھ��M�dΤK�G=�:$����~5-�+���T{ⷭ]]��	s�;W�d�Ni��N;��-���4����a����ɫT60�]��q��j��v�>��M�qc�(,2�d�m,ǖ��=<>#%y�����ꏖ]@��dh��G�M¶)M�1�6vZt���+��(m!�m��2iI¢}YT$5�F�{5�I?a��.�l���jI�*%u||:'[Ȧ)E'O;�B�_��jx�뮧�6�|vc����l�����r�w����_��cO,3n �6�(|HG����X��C��;���i�.��͎h�q9g����0�>�~�� im)��� ω��۰�Uҋc]���Q�����K�ɯ���"���
�f�����><�ΰ:�1�3=Ԛ�����ܥ��}�P%OIpXb;r6a�A,���OcC6QNҤ_�h��W��s�;W�K�&DPDz!�1qF��t���c��;V�o�����/Um�%^��럍%��*2b�G[�	<)�*>ZI.c��u]��6�Ŋxatb����ՙ�wM�1"K{eL����j�89�9����
n���|�d�pp���_�~��5+�;�	�k��ϭગ&����3��|	�=4D�r�i�(�y� �择RxD�l��*!ʳٜ�8	!]���q��}��+#)Y�N�X@8���/� �<6Fnp�r�Ash�r�،F�����j�#�G.͇7���4�Y*ۨ����M��4�/1y�E��I���i�O���ӿ�s�S�W��/}Ŧ�x����;�ܻo4�i�p<ƟBeW�A` ��&j@�ϝ�[@>�p�em��h]�b��}�%��F��"D�*�f�������]�X{���!�Q�l�"�^/��g*����4����.�S�WJ�4�������+���|�3#�4ǲ|r��z�)UѴ�_����~O=�\y/���V[�Yk�֭{J�~�����W��_���q;� q�D8PG�$L��E����xe]Є���ax^@����I�pW7n|$R��/p���.n	&�ב^W�06-���d�j�D̟�6������:��,�w>�,! 7?��1"]�|!��`w�R]�/����>�5��Q��r=j���B-i�K2�E^,�u����aS&��۸�+׮�#>��AU���D��r��ڋ��ҁ�R]����+�w�9�_e1��|X���ýd6�C��L�l�14e��,�S���d�st��m�v���~qz�0�c׎QTN�r�;zn�H����e95��-a�O��I|A;b�Z.��`�D
Ð<{��+W�2�E6FX1�9C��>�+�H�Q� �SѨMV#2��&"�Ta9�&��@������4��,�Mz�A:��_��G�.���QPm7y9�N��j9�m�ȩ��a2��d�U[���?׃a�|�2��%��&;hgH�����֌�����B��[�GCCR�I�����KD����Y�E��٫�A؛Mb���p�B!$<�t9��ȭ�n�@�y`1��~��|��������򚊣�m�Ν��DK٨�9A��ah#��=�b�_!Z�M�%��)F�ZA�s{=n'ׄ���<�ȷ��pݲ9��W�O�z��D���p@�zǪf"�ٚ�Fq�^��(���ï����=��zƻ�&�P�P�D�'cu�Ǉ�����3���f���$��9���&��N�x`�F��^^0��wa�g�$�ݟ-Vr,���Z�lm�<��u��Ϙ�0�e�����W��l���O^�'/�{7IW��֭[*o��7o��� �� 	c�Q��$��`�k+�e�dϔp�><,E��� �v���C�K�2��N�S'L��^���]8o�f�цZ�М��)[s�`�f)��z���䎪��R�hO\R�&m�Y/�յ���?�w������w�I�dEy����hl.�L�
�Xy#w�Y몘��0��ǥ9�tr���œ�����]"\��-ӝ-&��0(�
�`19}x����i�a���s�4�d��4�к��ڕH�<Rv̳4ߖ}ِ�� �������3��ٟ��ŋa_~4���{aD*K��7,��4�.Qv^H�u�M�ξ�����r@g8��\6�⮱	�MA������	m%I�����l���n�<~�O��a%�"+��o���ȋ����X�0�����ɻO7�? _`��� 
���K�C�o��?�u�i�Gܑ��s_�ƹ�bS�G7>��汝)u[�f����0@(�Ы�}�	�(Σp�Z��c�����'KK;��p"9�wSMgʲ���ñ�Vg�E�Zd����wn�����M�r�~'�y�̥hp�8Ҋ6��O	q��?G.)5V�S���g��������"c�z�ײ���bS��rm�wI�6� =UX`6��ȸ�W��`�e:gG�bϺ)�$T�
?WuZ�9lsd���7{{�RJ�u�����Eξ�8x	�ŴnRǺ�,WP�����K�s�qj��'�r(Jj/�lol8�%e�	Q��p{c�(�h�!9yAf,�lj�7ua��r��8�/_O�
0��|�V�!P-d��۶	#j��W.?��]�>B��˯<��[��HCo�И��T ���AtU���Ӗ*"Ga�� �̥2}BB�,�����(���F�.�k
f�R����X[���f�E��f�`-�Q*�H�����ơol�I��\h�hߥ���I��-?lK�O?G 3x����{JG*���*�D�'7�I��V@�lVD���ޥ��W�~���E
� �>�M��ɜM�Z��t����GB7�I�B�?~)w��`��Ko��ԓ��34&�N\8�أ�����C<m�vO����fAU��b�KRú��ꌩ������tSԡU�J�|tO��F5����8�|pł�޾}��ɳ���h���R�M� ��J�����5z�2�gb��ְ�ru�Ų��ڶ��R{mof�+�kr7�ְHg��m6�S9��M��M��ݙ4p���: ^'
�����g?�s_���vO�#亖+��q�Ww�j��vV�ʪ�J��2Do��$Aspp�Ԓ4�u�U�g��ta91��J5�-��������9.��d��+��u��6�z6
�M�>5MT���2>�8�H�/x�u;5��ȉ�:͛LGehl$]�i�Y��P���ɚ����X�>I}�R�zUըO+�h�c���W0[o�Jv�x0u��v�m��6ީ��m�z{��L:���	�
�C�I�;6� ��oN&,�뗈p9��*���
�c��(�@�:�e��v���W�p�xXx~�4'ltlr���k��P<���N��H��=JU-&ߴsa������+�jl��g������E)���cR���%QT�Z��!z���}�R}��H]p�<�R�K�X\�%�]�����_��a�!�o��6e��.CLpoO?�4.~��m���Tu�8I�_�x{q�ƍ�z#��kQ��fj��y��,Xt����Q}���#Yǌ�W��!���C��#F�ɜHY��tǈob��Uq���.��3R�3�$�y,�љ�ڡR!Q�����/������BD�1�N7�����_y��-nLC]f�%|H�i�4�7Ac����je��������s!��|�<UJ=:r�A(7IN�0�U��|+�P�ϗ���\3I�t��ʗKG>ί\�%�[l��?#D��<�l����!E�u~~o$D�9���Ņ�vtD<�A_Ze<������姰n���q����}�Ifpi'�+�L��g��L�O��xog3�&���`[�_e�u:9��	#C�2�Q���! m¢�#W[�1�Bj��p�~ӷ��n����rͩ�Zf���JP�d�FB�t~�%|CMj��̿����L�A����n�>�m��E�"������k����ɳ���y��ʋ��4k"×�Y���]mV�I^�
��Y|y�e���ڼ�ɩ������������b����6�%���tjmA��j���ۃ3��}��@�~g3�u��I��R-D�02��SR[l�Ǳ��3�H��,�u�C�;;�$ݺ�� ��7�7��#�`�RhN�T
.�59=��z!T���f�sn�� K+�P��|��D�	)ʲ�x��	17JՉY�])�5Y�7�+�"u���]cؖ�G<�I�bŤ�2P���z�Jx�+W�m����9��8�0�SQ��ܷ/��$%`�X0��^,`�oݼyzZF�h+L�tQ�J��Il��t�HV�Z�ql���)(��Zz����EW��])�	6⩧�b���ub������dյۋ)i`�P�83w.?3��u~�XӴu�&Wb�Ѡ���Uƨ2��2�%����	'eK�)���t&�nXa���
��A<�t	�޴�
�$G~�BS�ǕY.Y��k_�ګ��*v���������7�����s��M�Ƽ�p3��I�U��;2)��le���ogU���a��.�h��*���J�3˖�tӈB˴:2,)
eU7��1H>0���|@���+��%��5�:���7�߿��`vp0�p�Z4N{Q;%�������D�ft꼬��D��qM�Kuu�u$��V�β,i�1X]��B 2M7�~����D��mJ��LM4�����bJ�yV�|�.'�%b�����a�yU琄����m	j_�����v�S��芓�&C�PZ��g��5���,Dh���g�K��������+d!�8g���D�
���폠+��c�f>5�>/��dt�f]-�0�jI��F�V��h&�,�U��m*Q>�QK6�T�O�{�^�vj��o����	�֭�����v��2(D��A��1���F[�I��4y�6�
(b
!�6+:*�����N�M%��vCZb�u9X�U|�]�Y�ܲ\?�N�_����j?���;[�&�����v���Z�D��J�m�(I�r�g�t	�����˗eX�vB�z
c�GU-MR����){mǞ�� �m��㥗^��W]7#&t:�y�՞&����x�JR&��)�y�s��5��G������1	��y�dq��Y�Ʌ�뷶�@"1���Hx����o<��ٜi���䭼6���D�gJ̑���+O�.N[��Ҵ����Zѫa�[���_]@�B���a\gW�ˢ�ٸZ��2�_F�ܤܺ}/�
�j�0O�kB��-�t�p�W�G���M�B��]YT��v��t����"@��!��^ ��#��k�
�ꥴ��v#���gݔ���ˆ坼�N戡�r����s���v���YmU��B��М��LV�l�C�n7g���P{�@]3��{5��k��U����.M�I|4����>��<���ޣ�����a�'�i^�{�	Ya���-��\���a�;�zd�;4)�	��R�>�}�V^���`��S$�ge��!jt���-�".Ɇ�F�i7�)�T��M#������r�����<6R�'����d���t;5��t�ݖ�� 
��Z�D�"J�˨^ד���J�x�|�J�=��"�6[�Ϋ*����u�&ݏJ�]ۙ!]��q��Oɳȸ��ijD�̻�� ~��_��իWq�,�8��o����pa��TX�� GYU�.	N5ن���r�Xʹ/9���>ڐs#3�F$Z(,~�,v��̕��J� 8a�c���bhL"g�)��s��:�R��̦�i�w4���HX����y1[T��>x��'w������r[x�mC$�7�u�_��ѩ���lNK��5"�������ӑ�ssRٖ�1���ߐ������3L�����8_������zo�n���L��0rk���z�aԖ(�D�a���FAK���M��=��-Qq�/i%g3���YQ>�ԓ	l�Kҍ��r5�[����%�X������T�&oa`�]�p�vHn��i\�&T��1�[��뼉�R|=�>_�G{����>�,��{���_�(��8�w�����x��^x�x�J@�j�q��陋�Ǚ�|XFG�:Z���H]/
S�F�N�R��)QU��v�>@8���&��x��S5z�v0��(NI6�.��*ʌ��ݹ�^z��gG��G��+O-5�y�����Rr������?�o�5���_�źu;�'1��"n������^�I��w�����}MT���r��㲃$&���kO���X�Ħ��R�9�	�RM*����&qo4�­������r��3e�cC�k��L�:��9�Z�'�?��d:1<�\�(���1?��8Qv���r�O�h�E+�'�}��� *���>�n�5�A=�^�����I����	}x/���q�0$p)�Y��cM^$k'$�\.f��=�`>?9�Y��+˳�ŀVl<��br,�B ��S%��Nt��r���7&�Kϵ��D�a��l�Rov�M��>7��?��$���G?�M�]͌�.����8�~�XeM;��l�$ե�Z9
����U
�``�e\:A�M\���y��0X̧�QWo����o��E���3���Ύr���d�F�[��x�2_gx@g|����h�{1"��5�×�Z�2�OVg4�kTK���d�X��k<2��&�NN�bC�+	�t5�EƧ	��:��¥��X
1A i��O���"[/�Z��X����՚�¢�Y����A�-X.W<����s���/�?x�÷�z��`@�5:�!'&��Pj�w���DA%���PL��u�s:����x��;zF����l�2;_��p�ĥ�x޻w?��b����a�G��nH4A�P��3�J�m�u������8�W����P��2��#E�,x(�ܚ�������:Ri� }��^�%��D�b殹L-x�i0�k�-&=�e�l`Skj�;8:��v$���C�	5|	�kB�q�V `8V�J@98c��ZW������LBj��K{�Ȇ��A�CWl�V��jg����}�֜��,��|��w���fJz5�0Ë �e��9q���\%=vq�ᕍk�y5��m�:U�B��( �4N���,�����^}���������y��t)G~�*�y�<ܔ�:oS�A���?ʋM�m��7�U!�!׵.�7Q(B=���|ʊ5�8(כ�������Ѱ����(���YzaQ�@e��ަP�������άSM�2�`ź��Ԃ���@�mD�Ր�D�K�]{�+_~��a>�M}����~�[�����O~�"�ś�ye���M �98Wl���]!���������f)^���3c��'k�b�C�%��W�fu|��ID�{�{�&s�9˓�-k�ͬ�&����iO���$v��8zG_8��3����������}Gud�6W$�x�y�M��֤�6lmU�9ˁ~���LV+��F6B&+J��	
��F���Y7�-�h�>�!m�gi�^�Zf�,�%O�I��G��A�3�G}(�"_㿺̒ȇh@-6E�� ��=���v7j���8��a�D�;;,�޹�r=�@V���A�]+�An-щS���K_��!�X���|�ͬ̎�r<3�u~:9�$(G���7|� ;��v�O�{g�U�N�b�KŶN�4��n�X0����｜џ��~�+_�վ��/`sśm�[�VlQ�<7</�we->Z��"�I�� j#o�.�p�򼮱cgG�2A��Lو{���p�\��䎎Ƽ�rg����}7���l��2�cRz���U�*ê�Y�;����vIUn�]Y°Mle��/-+Z5�c��[�Ǹ���:�h��t�ߢ9,��W^�Cz����}&˷w�����!b (JYsHx�(�6���d�����������:�
�X�&�u	3wng�ޣ�_t�qv"��%Cc�֌a�;��4Qg}�X�C�ym"��.׳������[o����6~�})��GIuI��Z��������z�m��9����a�6s '�L�Η��(��?�G�d�l��f������ٷ��3�Ԓ.�ٲ���t?���{�i,����ٟ�ܛ��)�7='p��I��2Mf[���ɂ*�,ͨ]֤ؒ�>��Q�BY���oZ�i�6KQ�R0w��
��^UulC7�b���ɣ�5X58U�M1ܰ2��.]�&���J9��t� �*>�>��S�<S��^I�(��ᇂ�M&����3-�05*�]O���S�lI$�΅�Җ�9:�ݬ�W�^�q �J��eg�[A���7��L%\������_��I7�5�6%�Y,���Ƹ�!PZ"=㙁�������p��"\o��^��W���\�)!l�+��4fV=���t��]��R,0S��a�y+�܉�������mȧjǁ��t
���6&�d��;t���vY�5�X�^�ɞ��L�Cx��6�5� ^v��]�gV䚉fˇ���;9!s�/~���Ә�O�9�l0lg��?cm>��`~`�iS�X�-��F̒��/��\�Y��שT�	<�F�ǩ��}�^/�A0�?��/�
�THҤ�-���Iy0�̒�e`m������7M�2�������gX:���:.������tS8�\������;��'e�Bz|�J^��Z;�Z@��v�x���,�-�i�φ"�q�������zT�2�|�5U:�%b�ק�ظ�<��
UnP�j����-�޹O-�r�oU���*J�����e�������ҡ���<
c:�0Î�Cڃ	�,�w�m�`=���ZZrvG��"�	�����|�]�����<�7~����}Ϙ���������۷oܸA��O:e҂��I��R�F�1�l ���-�Q�)Y�#�U�R���HO0��ל9�J2[���^qF<�l�f�h�Y�,�k�M��e�$JE�C���x�:fOv���;N�͔a6b�l�vd�a0*a'R���������G�Վ��E��kqث�%�Y��w�I\ue�e<��v[��UB2��C�Ů#\�B��� k�_�j�;��
�*��À�5�&x&1E�Ν;z
|�{���pJ��gIe#��x@G�5�(�n(`�bO���h�\A�:�H�f��- �^$?�"�_a��X�cn�j�2�,O>���Z�C�*�Q�Q���ӫ�e�nG )D��6��z�֭[x>��D�~��}��f���;�L<엾�%\����������SLG���\ w��d�P�s��7����z�!��yVI������W.^����_��xn�B�M�KO\P�YYW�؋��Pxh�V)JWb��� x�J��*d1C�x��C�������V3��KƴA�FM� i�v��L�E�.�dr6���i@'�&�BV�æ��VvP5Q����_T�[�E�qyʰ{�$�(����8��)j-�E?n����	�=����@��y�s� �=�,^�ѝ��=ό�s=��U��ѓ�y�ƪ�jY���É�!m{��hF�᝜����������{�{�9������Y�o��v�
=8���Rl��J�?�q�w|AR��⴩�Ӆ������V7�i���O���}�nmȆ#�W@l ~�u��ض���e�67�G� �s.�!u�R���L҂���V����o����!���������X�A�X�M����Gs���mX^�Uî�F*ʰ#�)��<5�D~X��k�ϰ?��|f���0+��F�y3C�+���@���@Z�F}D�<���y��ՠ�lw�q6�i�D��w���օy��.��e��<�.?�k¹7XY���������pбOJ�S���~������w���ょl��VE���ym�a�N]˭/�le ��r��9��tf������|�&b��9T��(2�9����W�\	����?���0	Y��Ɣò��[m�NB�U�ƒ�f�vv�NI[z��(��5�]�<=#n ״��B��[�i��d.n�<8�J�:8/���}�a�:�dն�*l����[�=��J������86>nu�룥4��B��"�;�P���G�r��� 𿂋r��6T�b����f�M$xm�ϑ��#���e��hm�h��)[./&O?�����<���΃v����|�Lk� h��L�.O���i<�p�ri��,]g+����}�����&Nj�nƫ?�&#��v��i��
u����t�x�hxߣ�X��~�ﲢTdk;�h�Z� �˵��Ʒ�K��4⑮K��
{L#��l����h	�b���^K��X����h�n{ξ���hKT�=��4n>�#2A3"��>Φ�~�������o�SIqe܃F_%������q$�	'��eI�_n�q�v�s
[
'U�!FB2�4�C��U�E��+�"ޱ=�]St!�J�lA�c]�ũw,�!n�A�\u���z�Yh���f�˹��S����
ԡRxiAi u�:o������u]����m[?
����C��tn�f
9|r�m����n�:@o�GI�I��$�λ�G+N��Uт&\�6���EXbVݽ�z� �����p��4N�?��֘1��
K�7�<���g�ܷ��1Ds�>�2��ڜr6���n�6pIk�9�:�L�z���P)	����J;t�R��R��ι�Wa��c�S�B1�b<Jl�oJ�#ù�aS�����XA<b3N��j"��(Og��6I�*�Ѕ��MJ��F�k2F�#�FkT��z.kK����!�n�7ƥ�6n�����媀��q�X��k���ѯ^�Wx+��/�K�a9*������{���O?�ù�ߐ�<C �(�sc=���$�0�9W�C���^c����v�SW+x��_���F�t����`xngWק%(�J�E��G�>RzQ��k��'a���"bx�ưu��b�L[')�1��
��U}��:��z����
|�_�����h�HLP����Y�����q�i���T O"�;H�� ����N����K�?����<-R�-�X��馽�yu
5Lu!�]`�q*R��n�QUO泪	n��8/��+�,U'�h� ���-W��7��7�xC�dx0�M�y�T:�W�{�fn�{���6o*|���E̺��@>#&��c��qi�܆�9ǭ�΋[P�<f��6��-/�r�x�/}�K������y��F�m�z�Y�So�b�K�b���2���x�%��w�ygrJ��A4���]6P�*�VKlW��/����ONJk	�Fe�Te���p�*�(��7�<882�F�	'U�A-��^��lqW�#n]o'�I)q�3��eS[y�W��v�2�0��g���Xe�h���^?��?=�O>Y�Op�89qek��G"�?<|�@��k6�5tm>9��B�ץq�1��i�C�A,#���NR�����-NO��z���`�$Φ0�Ũ�����ӗ/x�/VTώ�v\���x�ڑ���N��Xȁ�aB�0���������?<�9�w��A/1t琭�[ۢ ��ޭ��~�W~C��XϫW��C�=�Le��J2�,`����R��q2��1"����B>E�)V�1�]��?RrAl�,W����(�:�9H]*�I#�hz)s��k�J�M�9'���������0�q���M䞑�i��ǧ�Ӻ	��媬�����'.��m=��FI/�s�n�v��ѱ��eEwe�Ԧ�P�'�QY��JS;�[�4���~����rS�4y�-�/IePf��4�ޞO�%��R�&e@h��~�Rm�|%Ӵ��)�և'�6ʕ�,�}j�S�=�d�i�(ɨ`�н��=��i�3v�\X�Sy�:�}?eK���KQ�0��
��X��~�ގ׿��KPk�y'�^h������+?�䓓�c+�p�+�oq+肁aa�F:�'f+��	��
�<(�!�>44��R����a�H�<_f��(����\��G����;�Vy�XRg�8��Q��r��H��/7~���s�e┲?88P׷�&�k�"dGb,�^�'?�9����鿃nľ�����[ڠ�t�o2�	�����%53b�?f�4���t���(��Y̧��.r��^�h8k��Y��,:87߳�30	�r�a
�^���jr<��̖˂��]o�����R4n!e���#��8�� U�u���J�](�^��2k����n߼��o}����2�%��	�O>�ZG���T�!,��6�7�f����[��k�Q�-�7�O�MSrf|-VjmL\�G^5�eS����[����`����W�|F��bh*�e�k�E_ q��K�u�A0�u�~��Gʶx����QW���Sԡ4�# ���|s�bd�SO=}�
�5�w�<��q���T�`_���Y:Jz����g������zЋ��?:�'�8�b��\����CC��<��ra{�����㓃_|��K���1>q�q��#��~cL���Eᑉu�[ůq�e�&9�=�x���	e���rO��@e��ׯ����A�\�x��v|t×�t� K}��P������;;��O��[ou�~9c��p����GR���nn�|+�>t����G%����V��D_k縍G`��-Ȼj�"�EA`;�Q?��3� ��eJR76��+سb̿���|iu��d��)�9Ɨ�K�J��CS�RQ��GM�}����.�x�8�v��h��-r���Q:�#��%�&�4��O��{<is6�q6=�@#�B����í^��������Gm�\PC$�?����Y�H�،U��N�=N!������������_��LС��Z޼�Ơ�^�r��-Db���/�-V���a">�|�6f�v�
0��5f�=
�F�:Sk�
ފ��6�K��go�k���C6-)�^���^#��A�������`�ܧ�wZ�-C���k�tY���a��M+c5&jn�F�Fb�9|���:���!~�1���+9�Ǿ�WVg�t�A�H���s|���6���l�d�V�Ǽ�"�f��-)t(,�L� ���������ה��Xm���{we':J�w�MW��:�a`��6�U�3�ϴ�+��PA/cсM՜O�#��f?P����{���A�Q0��;�0�H}����RiWU;ϲ$�k���ϳ�|�,˩�j/˽~?*����L/�V��������ͨhi"�UDg!8C�g��m�nԆ��f3g�����F�1�Ĥ�n�<�y������x��p}5qk˴k<���z�b�P�I������YL7<'��B��Lew�ލ�@ѵV�cߦ3��n�,?�̚-4�ބ�F<�r��s�*����o�-kb����m��j��ْE���^��U^��X�ܫb��m������FYnX���a�L	}Y�~��V�E3S��)�$����yƷ���iXP�*A'�lB4�{�X�y_�)E�]ۦPT�	��y��[�W��g½4�nG�K��Vk�-��5�Xi�$JO�A����V֑kjgW�\�uM�:��1��8R�٨���A��B�*�����=���/�6�o�`��g�}��ի���w�����_�"�������uy!ݝH�,�KˠWaP���6��}��	-�p�^�?��B�*m�z=&ʛ��1�$�OG���E���6�T�M��=jÎ�^"���8�vc��V�����ch����~�!�x�S�V��m���(�D��W՗.>�לL��D1."M2��� � hX��ݻ;�NS��Z��mK��j,�_���0_���c[&�i���Nq��Ka��/����p��w9颮nS�ԕ�b�	�����Po��ߪ��Y�5U�6�`�$�����t�2Y��L�8}��7��y<�fk;�Y�'&eH�.!��6�N�&&�78`��C�-�����3��������5���&-��y��5)���|ٚ�r���ը����8r>�5�X�Mn�jo~K�T{����@�u����N-���f^�%�~���#����m}	 $AT���5��)��l�w<�8;���0D�UW���Hh�S1�ЈX���GHDcT��B�B�LH���L�҃F%&��RK�:��B$i�!��b����W���o⃠��CN��<�6ո#$�s�y�:�������з�Qp9��uJ	o�W�@Zk�����¸��v<N�)-��+UI�����awn޼���/�{y�ʖ�� �E�(��rn3g̲@;4�)�N��V2��w���b@lm��].����'cO�Ԯ�YEMW��?��sǍ�IT��T�	WHӾ�<M��~/'sc3�qĮ\�۩6��ɩ��H���mr7�TV�ݩ���|��<�*?�Ɖ.�/_�-5�C'dV ��繹
{{{��믿��k�	��8�2V�UJ'),������Ic˦m���hqj��vqx���w���M
���W��[A-�XX~�9K��S�!���My8J<�Һu�����F	r2������b������ŋ��O�tgk������/~1�N�d[���:�s��x��T�6�P��_�y<-�q�z^e��q;�/ӪB���� 4�)�
�	��T��U�e��7Ʋ~�t��~�Y+�����{�x�ڎ��W^yE�2����o��o��g�������TZ��2L�Ԇ
Tƌ���AӜ5�I��sj4ʊk�{�͢j�<��҅	�S=
M�C��y��M����U:���ʵ�5�Bn<�̮!*�e� �} ��[bt�ajV�l:�FL%<0.���X(Ǟ^z{d	��0�p�2��D x�B�B�M'Ư��t})��|��F}2�b����ج|c���^ߐC\���P�6� �p�G�.��9�`;�1"3)ʱ����/��oh�sn|���������{�~�Ν;��+����It¸�".�(�����ާ�	<.�b��S[5��%������fv�o�}�lAn#��I�+��Y�?����]�M����H q�^�IK=Dg2���ry�^��s�	�(���A�v�_�r��[,n!D�l�vh�n]D/��$�ʺ����ɱ~�7�}%�?�xx��~�e;���g�
�|�8��<����H��ɚ x�x1M��w���ˬ�n�B���
�%�dh�3C&K���~5-�/�>����&WD��sM�ҕI��V҈Ym�F�ȕ�J���|I��F��iQ��"�����Z]�o��XA���I.A�V� �L)��0�+GNi��3�yC$X��`F�ܸe+֭l8?���uC�C��"�ev�%�����%�MZN��d��>���|jw��m�C']2TĊg~i8��<��y�����ĳ?����Ƴ�����3p(���\��K�I=,�w�M;=S���fע���o�Ž3(K�K(f�^� B��[8�v�ft,;��<����d��NҠ��⟰���������Y>��,!�O�el\���"�ɬs�]WTI�݆ޔ��G�����$�B�6��EQ��u����.�J�R=2u����+��	.l��e�??���c���)���`ʔTA�t�>��{���s��#&�z+���r���`8ڪţ��<gJ}v2��^+te}���0�`8);#N�<[	Ƽ��;�[U��	Zp8��o2��4�,�[��[C<\m@I"���m�V�q�e���
߲q �w[kjs�`ã79�P��w�;IL�>�+���:�:Q"�br�	�]�L��lW��̶���M拜j�>��*G1q�]�pHSG4»��J�!|�F�G8)�<¥/�A�s�\*Y��j Oj�+�mNuT5Ǖ��q)eP65Kӓ�t2Oy�f0L��t�w(u���6��C�O��;0ʿ�P�Q�X��+�}���92j�@�\$�Ʇ/���-A���0At'?��x��-�\x�����[Q�s"�SY�q8a�g���!<!�[��N���	����\˃ӎU��1��iS��4Ƒ��4Ջ����RiW��A�� ���97�p�����r}�=ط��2�<�ٻy���K`iT�	�
�׹V*�pIg��w��}��&��U:@B��Sz�eŞ�u^�$�Ԍ�~�O$W�����Ã��W�z�a��_�l���QB�s� [�zQ�b6������Y��G�M�D�����M᥽7�E�e=�X���i�E)��l�>2%�d���<�\~�*�]����6�fhbI���6�%�V̭l�.	���^6yuj��������"�HZ�;@��]_3dA���*��hQ�M���"�X� �lF�:9Z(~V�^N\���|U��;|x���;Ji�wƜ���7e?�Ī2�eʦ��.KOv�S��d����<_��R*��<uQ'6�R�~��G7a4ONfa����K��K8���܅=<�u7���������J�q�b�A�}�2�\l�K|zi�l�o��K@��ᇟ�
'�i���e{�l�Ѩ�8���f���B�����*^ʋ�;9~��ųW���c��lv��*I�@X��"g6�Q�/vms�$c~ຶ#N�T��{>��Zf?�����3� �%3�"����dRm�,f`��_��K�ן{���)��t��������z�����
`��m~�&q����fx||b���@�����ܣ1���K������T�f�6GGd<�cDnJʛ�������\�fݨ�Ç�£u�=Ú�R�F�j�a��8��56����(4�A(a(U��^�~ڨ����µ����[�����L)E�D+���������֯����?���Pn,���{��-���W�����u2�̬�r�Y��S�Ly6Ov�_aUu�4MQ�
HyFOf:c��o#�!�e��zIߒ2�}�C�v6	ƌ3%��8L����V|��m�au��q�h��@��O�2�]8lG%(��d�r���l���?�#N�_��_���_z��o���I��?��'��R��ȱL0��Oj�M�>`/9��m�En4g���M��k#�J)�0��KEg$�[��d�g�0f.C�m ��Kb�������<���x���(�%�{{{b+�[�5���U����WOl3�'��L�����/��/���� 4~H�:�/\|�����9���K/]�����������kV��Z̧�G�(��m�B��CGf����î+v��� �+<��h��KҰ�9ٛ7n�'�l)3����6�#P����ܪ���ߐ���zju����	����~��5_�㪣����GO>��MI��H�{1#�A��=�mR�+:�	��Jfl+妉e�LuW�x��m �C���x{�G� U)ww��s��l^���礼�k_�"���4���GjS���B%ϧ�x%6�i0�j���3���ɝ�
^*zM��5w�����t6yp�p:�=����}�2�m�+)}�K!,�|��{�����E����������i��xj����7Щ��
�ױޤ�AG0��3�U�P-����
J'�XB���5��I�dn���j�
�׹�Stlk2P"XD���H�5�2���w�3�h����wy@�S���Q��f&4=�Rn���6�:U~TWm����_��	���oFCL@?��mܬ���5��ȳ�׺q��ZVϰ�4�C��麤�ܿ��L=���-!�]���vSyS[�Y�%C�Q̍���Z��^��7|q�Ge;�Uك���,'w�� )6�[�I���y�]Տn��ɨӘ��)����̴ϣ��b� ���G?��=�3�]hݹ^�Ru1�e�߉�e\���J�f���bh���L\$����R��VK�K95���z�?o�G]Ə����n����Ɔ|�7��������� znq6�����`}]b؎kQk��cu*�P���xa/�56�[����^��
��#n�t��������ƺ;�2ٺ���.����{*d~���pnO�&Ł[��:/�M�EG�:�/�L���n�m9���f���8��a)���4�Yk��Kzl�ќtQh-�,�(�Z���?4��H�TxQ3�S� 叔��۩��e�(����:�kx������sx���{��+��p����)`��2���l��c�ef�ZP՞���Ň_��_#+��|��h��g��t������a#��a��76T	k�-�q��#��0��\��%�^�ԙ�^��bR���jJ&�.�bXt�0�[�k�5�l���>��*��U��J���Oe�%�*�+��%d%�ʏ+y!v�u����嗯����9Ea��{�eڇ
Lj*W����E���<��x{�U�y�:�))�Ư�<W-�e��L�ff�a��0mZ�����t�����G�y'yJ��U�DZ�\u��X�PVJΫ������-a�+{�
{�ء�-�1��;88<wnW�m����IQ��v`Lv�IB$ᓲ�������9ƒ�.TgB ��ZiSBB-�G��^B�t���	�K�-�����UV�!�������"��Z���60��&h�l�_S9�tz�`��ha����� �kCPK���s]��4�/�o���/��׮]{��Q5-(;<3��sGiG�}�������|7��y��%���R��x���g�����{oܸ�vZ����>W��ሣ~�w�Qr��}�����R=>��P0.��$Ѝ����ٗj��C������N</�Y���n�W"&�]�#�{�a�`n�:����vy��y�ݡV���=c�S"!w�.��T�7m-������l�D��g�)m�R��v:T������8C��^嵩�Z�߀�.4�*��r"z�*i����?M'Dg�{[g+�X=l"�W_}ꓒ���P$P�Tj2 �B��&��ğTݑ��RY&��~�D������o��u���$�,����]}/��$QZv�܌�E%�~#����x��i��rekιVr�c�ÁĒ��H��)\��o�Ϣ�Ǫ����P��'��Ԕ����&iT��3��T�&Ʉ����$ck�#�P6M9�wv<�0/c�Y!���g����ҥK?��Of��K/�$\A����i�	
���@-Sq��g4)jF#�6hSj��C��'TY�����iz�����u�瀞�2zQ۱�e����xI;LF;�cUX�^��(��8�K=<��ϭ+<���f���B_���Dn"�G:;.�w�t��j�^q)��7��im�Ա�>�u�&V�+C�Z�)����0��'������z8f�R�>��BdLtqs�қ���}*|�u%��&VJ�������kV���J;�;�F�(HL�:�T�9gcr���v�	y�9�qܝ�/L��/��2�W���H��4�'��˛Uj��t뭓���U�i���8^0G2�҅�6u*#�.Hz��{�lq�X����Ko�#Ϯ�4}��'�* ���݀Ow"o�oA�F�@$ �Zf�s,�1����=�ɹ������*K&b�6�Dd�=8<��|����4ѫIv�}Ѿ��7���(՜�����E�أ���K�6�{�E^��V�r8LU��w������S!�X�.�w�E�C�M��6-��g��������?��uE��^q^D�E�n\�%� ^��M�N�έ�|:�2'�}F6��p{��3�u~���96���xf�^����[�"RP5H�k�F���;���>�ԣ4$���1EX8����9��e���-��r�$k��ۀ���o~�k_�m6�G��3b�qe�p�2mL�|�K�/�#��qK�A��g���c�e�	i1q��j��E�/���s�=� œ�R`���LS�ͪh�'�?��چ������3޻����*g�X��BP�FW8Q��n�Ց�X���BjȢ> ���y�QU�f�5cZ��"���r�d|���8F��B-i����o1@f�Bi��0��0ͧS��͋�M�tI��f�|�$�D7��o�}����>B��!��(�#;bԠ�G��m����"h����<Oax5���믿Łe�K�jsy��Jd
�d�y�KjѺ�1�x��0��Ǫʈ�k�V%i�)F����fM�63�I�V?J����<�i@���FSv-���u��)�	ߵ%5��W���U͆�NXܐ a/�ԆZ;��'Ӭ�p�J��0����Of�nR|����h#�3�-����F9J+��p�3��cJ����$R��}��{n���`�d�j�:hW&p8��Gr|�� �RN��4�Fw�|��g��ZZ�L�TYN��g2�fK�Dzp_�*��;v?���"[�:0�9�5�A�"������o���Cg��r�'��4��7"pr��̦�X��&��bM*�&Hl�f����I����t��vS���z��m�L�2^�$"mPx�$�Ga����}
^;�a�M��d=�*9�3o�aVų�
n��`[mVf�#�cns�g-�):�*��#�ʼ�&[����;[�e^�!���qb���H8#�Bӎ�q��Qx&[ބ$	*N�2������}�����s��?��I��T������{�8�C^��f��[��^?�K�\�?��.]z� �K(|7:f@�^���zPL�d���Q�B7��Zc�2f^z^S/�z6[XX�-��
Gk�����C��[/�J�Q�Ppf��0���Z��Mb�BWY����[&�N1�'���Oks�l���)}͍�~/��xL������r�fA`1=�g�:<Ƌ���뛯_O�G
e�6	
��O<A���Û79S���že�v�-7�P�?���`H��H�&�oQ"�:T��������.�$P��d� ܮ�2�+^V��!'�:�IA�L�c��H��i��l�d�UxWFKೇ��r�� !���,O.ϝ[LOF	��m���o�^������ݫ'�����ߏ��J�'rΚ_�ͺ�����x���,�G�!�t��k�9S���b�ɽ�f�|��NO���ɟ����?���~W�u�0YZ�����	�:�䛣lÌ.W�����ٺ��$k�����Y�4�O�QL尘����nIOk�"g?� sABh�4�8�\��}&˭Y,���L�)N'0s~�5Id�����K´�W�bHWH���
�V�$�vz)�o���p��������?ȫ��'����sNaSFOYi��$(��Z+A���1-2��FF�����B��,�'e�|�\l�؈��w>��J7�sP��ǿ���'?��2���BmPX6x���-��~�Vy5ϖPT��\ ٝ�v�Y�y"_�K�M��S��y�H ���9���pd� ���̦<qC�,���	��ײ}��׈��5n�(N�n������}r���q���e��)a��~O�FF�Aߥ�
?9�v]K���MU��Cb��g��a��/(�YLL�S��R@�fo{����������RF�����;��J�#f[��-�oІ�a7�⾞�DX�1���ڱ��Ǉ@�y.��rgCrU��Ap���������ȉ`�#+-p"jt�ֽ��O.�/���������=e%>�῭-GG���-�[$=M��x4V����� �mL�4�
�<Kd�|ᅗ<�w!��%�j�%2���~s�f_r~NQ=�8��x�L�]1R�OϺk�q`1Q!����S$͹w��j��x��ә���H�V�q.�V���$^��l��a�m�^$u(���l��XzIc�Ek�͵Nb�	�ev���q�V�}�b��ģXxxx|���!Q�mPms�I놐�����w����wE�X�b��7m�l���LY.��xaD�F�~dn������u�� t��$�<��u1�B�~�X�<��l]�אυ��iڠ��9�ɔH��8�B�Z/���}��5�㡱d4��g��r~�=�=s��h������z�0f:eqh�/H]l(�v^��b������"l]*�߲^���z.��Ofe@�G+��@h��=��,���>����o߾=�*���H5�����@�hA��_b�j6Wi91�C��������g4l���,����j	��22+Z��|��1��$�Ʀ%綶%Ջ��U_fu�g`�)����3��!���=+Թ�!�AȂ3Oz�;�^��/�����������q�Xj(���?������\j��.�c
ř��͢ET]�%b���"G܆?�FF5�MJ�"qDÊ�-�B���R�V�8ۄ�#��^��b����>Ϩ$�d ;j-��ۻ�>�V��bx�C����<:Ɇ*@Vd!�N>�h��O=�ɳ��~뷾�u�'@ �����ܾs�?���k�W��Z����g��_X��!	k�2��S^�z=W��\����ӈ���M���c�O�p~�=�6�իW�k6b�����P�@v��p�m�ӽ�x�ڵW_}r����?����x���>ˤ�j}z|�T���׃����j�>�-�4{�͕�r���_��g���n|\�5ⴱ���Cl,g;B����d�d��<_Lp�b�x �b����_|��.ۃmxa�8dӭW�Y}��������}��+�Nf�[�pr��zl̪ӈ�F��Ǟ��ո$v���
��P�e�ܔ�N�����3�/N�a�t`�/J�����k�xM�i�?~��������o�	�w���a���L�10�݇����Nn�)�I�fv�<rkqo��?��?��_�j0��r�BP8�5́p�*6*�B�üy i,ΐ"e�~�_@���7�Q'�����(��M[M�7/Eϗ3?�2e�C�t2�?��@�4>N�v�"
�Ⱦا`0�i�X)ˌb���'����j����T&��Z&{:��gDu���Oc�I��u1VD�&U�Oݸ���R�Py,Ub�o4���Rg������#�M�Ee��0����Y�����Y3B���Fc��j7���=߾7�'ND�(��u��v���}9���K�s�]53��u@�Ѻ��^��hXj(����Ñ4Mj�xd3�/��'�(Y�b�{A�Yͯv]���D6n5�"���QY8ʾƧ[U�XSw�X����u}n��{�����,��͛75 ϳҙ��^���hU�q� �� ߧS�n4�����sM�*y��dT�g�����ߩ���OOq�tSGun����ܳ�y��g�{���j�叭�ٵ�؏��s?��e�3_^����{�Z*<K� Еt��W�&)*�%�3u����<�ޫD�ޢ�wxf�DT�tY*u����)�
�Ҍ2�ꢢ��
���9B���b엤;���nl���3%�W��#�T�v
���A�B�h$�� Cۮ�����Vp��Id	��ʰx
_�Fi1�j����C�Ѱ2W�>cII�d�pFVNm�]I�vdgXUO���:���5�͟Lp'x�[o�ew	~sXFؓ~��א�GZT���߿-��rY/���Z���x��$�z|Yd�dN�*U���^�p�p,,�$סk�VE�M%�ca���կ~��ŋ?���I�nSI�F����c�B5da�$�ⶓ��Z�q���-�;OHU+� ^-�%c�Ƒ�m60���-�Hl�h!�CeI���C�0�q�UЭ[�tRA;�;7��jxƅ��g�:��N���s���kf��<�-!��1����\��~f���3����*�H����A����Pk��i�yJ��� /���	NOW��*�2܅��RXi����6� �τO�q�N0 3�#�
���=�|6[�@��0SI�Ƅ.���.�� .�0�K��pX���������ɉM�X��6M8I�e�>'qp��E���.��3��}����1˖)��'�eW�y �v�9�4x��/�d�ؤ�"�ka��wpL�YO?���{rr'�5`%E8|Ǥ�g�u�蘒�Ѵh��hsoC�.UuD����r+HP�4���_��7�y�����{�k&RY*WZ,��E0S)�E`�҈���*үB��#4�Uoq�v���1�+&��wx�a,s���4M�����͊�ͷ�P��LmGY���/gW�n�{p՘�wVH<\Xg�obQ}��������=Y�՜��:s��_��%8��Z{IE��'���w.V�g�y�i�;X-�F�������W�d�u&x]�,��Tu��o�A���3���2���F�Q1�oz��V1��P�*�����$Z�!�{���ޕ��������wvU�dTTdeݼ�7�?�;�,�l�6ݴ�0�JvK���U��Ι'O���>Tv��G��~J6����(6�jVwN��4*��SY��db5%�|#S�NtSgAd�e/��H9��)�$� �(`"�嗏?~�ȑw�}Ww3M>��b	.�
ca�`�Z���Q,���M�sV�S%m�oWy��4��
S �����"K��w��>3v(��4�����kKe��Uo����kN@"�Qi+��כ���jĺ�Y-JېN]���֭[� ��D 3��gP��x)Vk��1>B���Rմ�B��"�[,3�
�C����OMM	BJ���z���	.FD$��M�p�Ȅ1�7�)jkj	,�҇�Wu��3��x�"�M: ҲPKKU}��ݷ	�(>��PX!�v��(TK���h"}ZZ�[I��u�&<V%v�D�&٦!S�d<��MS�-�'�V���/a����Z������*"���8�F�AMќmi�Y���ihC�(��2��6�u�D�.M�@�����
����1�G�j]3�q��Dr�Ƌ;�O<)UhLb���[�\[�b��O�>-=�2Y�}_O��M��('P���%�l��2���9d�G��t�[/$�]1z�0�k׮��m��!��o=�������j�KZ���R�$r�� H�56\T����L��w�w ���?�aC\�aՆFG'''�y��_����O�E�̎�sl�����
v��NiiARk�e0
���C6�A�#�s����V?����5��������,��u�]��x��da�Zo�cSA,65�E󤞠�~l�-�s�q��\��5�t�qFSnyx��B�[�- -m�Ǜ�0��0I��Q��I���� �1Y�=�&�)�Ꝕ���,`o�hz0"�{~j��i !��Cs��i^_�n�T{$8�0�.м�)�+0�1y[É'���7��'�|�T.���7�]��.^�x��)��Ue��LFx2M!�fPUNL�x�ZB+��D�S ��uր_���j������d�AQ[�L�6ށP�lĨ ���>��!��q޸q#(ߚ�̕�6��D�g:��:� 1H�K��N�L��)�����hV�Nq���3֭���'Y�����N����u~�x��o�]��{%��W����Y�-;�N��c�h:'�*��A���&���L�>�K��y��f�7���C��i���r�B��+�}w�5ss�9��˛���5�0UI�T��Q����NR�DLD7W9�T�%�UpeE�Ը�A��H�D)��N{&M��Ν�k"f
k��ި5s��z�����~_���Y��9v>�<|.%�(�g�X{{� �4eXB��ӌ��L�w�6��Md�_��Q����T��z3��騴q.��Iy�����XG��a:^�m^�I����a����tu'N���իWmAC���5La>�MMw-E}�s��mjW2z3�kP8Id,L
��J�"�R�J_���OݞP�����E��B�"J����P�2��(=���lD�n8("W/_��_�������}NJyK�BNSJ�X�c�{z�d"�����J��b'æ�v�B��#�{W8QZ�3��Gl�Q�<�5�<�&%��2w�m�; d�Gy��x:u��?�N|��B��G�b��`_on���[0�hH�,�1�rښ�z`Ӄj�Ծ���g<��X��F=�H����"�I�e����Ue����5��'5񾠪9�q�)YZrX�bb��&�|E^P�R��*ơ�v5������*��Jc�Q�k���6���m��pH!���ZF�bH��lN���U�vh'˒��<�(l-..Em'8PH$�-nl��Ev�l^[���l�5�����,-���פ�e
S�ܶц.�����h0Zm3�Z�j�q
�Ol:?���2�)N�}w�������~�!>d��MQ�6*վRO6����.5j��gŧp�Ƶ[�n,�-*M���h��S�s�D]O�lHk>qh�4����gS�Y�\&*�}w��UVڊ�����X����)��b��4A/W����bZ�����"�7IZ?2�l&}CLf��S�^Ң԰=0q�J��a6W��W*u�llP0;i�Ɖ�:��m���MrYw��8}{jffI�g�qە�9�S�ߚ��RQ���f���4�Ђ��"4�j_��l^k8
����7�7��x	�E��t$�Tjjw%���TB)lL�)���@S]J�=,w��[�7�������P��V�v*��d0"����\ϙ尠��'�ntܖ����r��q�!�c��h�!x��2wR2軻V���,BV�luIPQ(�7s��|��f4�R����ns��U�UBR׿b
T��iR�V��3(��I�%MVF����ҖҎ���VV+�@K'튞�6�����+���N|�y	��]/ܼyk||���(�����4ԞԌ������`��KX�#fLW��6Q;d����ePEV�G_�*ss3�V�b��jDa��l�u�h,�ff7V��ރ���ѾI0��M��qCZ��>���D���ݙ�y�<5p1lQP}�e�Sv҈�>�G���aV#�,m %��V[<�%�L����b���=���!�AB�+�3ԡT�1�)a�*\D�,/���mЗ�Ú�"��>�N۰J�M�IW�Tp�%&��*�b6�KdZ8�l����%'���[����{�����V�g3y�ڪ#+R%�i�r��H�
�7e5 ������*Hkpp��]��0av|��_A��I�U1�K�j��0d�`�C%��<��e�j\�P��M0Zj_��y��9�+̅�I9�e(i,0���<ܣF�9NAFϔu	�4��Fz�|��-AL�lP�:��k��B���h��S���Ҫ�\Ij�LPeT��0/*i��u��ћ�(J��VN}r���3���� z||\�{zv������'��*RT�Ȳx���Z5���,�k�Z΅�+H�vv������ ��fn�i��u��	��	�<�e���E�7mLx.AS� ��� Q���Je����8s�́�~��D}܊������$֬��mxxJ��aI�a�޵��@���n�$T��hC����Z�r������>�H�[��*�rafz�J�:�؂��(���I�B-�|���P����Q4�2wPNS(ҁ~�8l�� +8vaY������+dm)$�f�e[h�q���6�����%���H6*I��pn�fA�|m7
!�æ�6����Q�*6k���m[��av;wls����Oժ�颥���1��I]�3oK[u1C�1�T7�*@���m���P9�T�6��u��'NHn~�'@��"�^���|���{��ܹ3��L�,"]H���ŀbD�(���-V,�����5�(�$��3�A>U�J���l�?�Ҋv�O��柁�@��Pɗ��c����ӳd��m���Hʐ6���{q:Q�����x-oK��Z�����x�o��{:I�{�Y����/��ZW�Xj��w�Ys�5w��;�u�5kq`�O߶QR!@��=EW�h�'[�١�a�ȴ��r�4��3�j�g�z|��3ۦid�9�׿�\Q_0�����6b��W�ƦҶ8��6@�NW9GV�(㶎Ov��|5]朆�X+h�=�p�u���Є�ޙ��N�w�Iw��v�����D�w��:κ�8������y���>�-L�Q��&�IkE�Z�H�v�����!$MZ2�$���6�D�%��J��3�4|�)���LK/�+TO�Ō�����C�a������.�C��5��E J�5U��ԃ���o�I��7V�i��(�qzI�gW ��8��)5h�6!]�EmZq��a�RU�2�p̦��S�HƢ#��N�.�zC�Kd��<�ޭ[Ss33� ]���,�r"�9�)!D1�]V`rr���K?T�|/��ªO�"����)��QĦ;C����}X4�Q*����� ��0w_�~	^v��VY�"_�>�}��\[��"�[((�T�v�!��PN�Ƣ��i��*BC��E���S�����a	�ԇȂ�R�2��0p�@ߏ��IJ�g���R*pֱ�.ޠ��t��H�ޅy��J4ب{���][������W��crҢ�z�A`Z�833}[�&"�������~։�?���������ݖ�0v�m�0�Ōd�,DY�P��5E!���1�h���VT�$}y�$�#�5v����D�	�cq\�4)�$Ǣ�Jr��ݶm>���:�s��gq[g����ImV�I����ub���u�Y��ھk�`4n�G�������)�Zoێ������I��v��U� A�#�
+�&�M.+� 8�z#��\�h���6=��]K�a��Re+O�\�J�$�o� X�����ںe�ȑ#�Z�ə��Q��i;�O=�����Re��>+dsL��]��>}�ӳg�h�j��N�ᾛr�t��2������`�9.ZA*2<���Ix��O�7���������|������GZ�S�Y�=�>���j%�����%���m�)+n�w	�&x��AF,/-/K�E��~���m�'E�����#	�IO�����j�5gy�,�zK$NSܦ��FՒ�߮Յ_َ%H�������@5q[�%���3kA����W��ڗz��]�A2'm������3k�[ZQ�v�8��Ӗ�}KŶ�_%��!>��ڻw/����z��+��m��������ʘ���� ��#��h����=
/ϔ&�gf�2-.k�;�K�ߢ�;>/��i�S��"P���⏴kD��R/�Y��}��J��Lb'��rc������@��A����v�� ��%G�8�Mj������z^�/7��1J�3`\�����fzF8x�p����!�c�[,NDŁ��;=[�L��G�A%�ij�-.,3V*��;V��d��Qoq΃m�A�����dM��:G�%��][ ���M_�K�.]�v�K�&�+)�ߤ/|����,-B�L��*���vg盂�p�L��#�L�ݛ$�M{�p�SF�^u��:��d�a��rK�<�.�))��=4q�q�[�TZ-�:¨̐ �\R/B�w�3��5_������~�T��,1�x![��ZnOI�5B��q�b�*�)#����C�7���������e�øu�v���nBа1��2E��ߴ�x��&�V���X=9�a:���k���l�t��qs�98Z�!ks񀇚T�0�=5�wfs�q���i�B5����H�`��6m�<}��~��_���?~��1H�k_���cO`%�|���n��sGF���a�>v��ٷS���#�-W�SR�X�F�ҁ�h�v�㰺R厳v!��A�~�{�ÊAɁz�����o߹�U�>��������H�8k�;O4�h[�v8�J{�ɉd�UW����.,�s�3Zx�|X%K��j9Z�
�z�Lc��@k�bs���U^��.��@eS�'�c�;`�9mv�:UI�4�h�m"��$ҭ���r�RՖ����A�G�-PYu]�	u/_��سg��� ���a?����ⱝ���B{�nz��޲�Qң�+������<������j`���z��t��f%�&����	.sG���rI8Km:>����q0�F�e��5�-s�@`R��5���^���V�K��|!�d� �.S��z�ĭ�t8��[rϯ;_�OL~k'�������tx��co�01@��M�'Gu�;�U�����:��*���E*^}��9��.���UHCJ"��6Gw!���>�	��R�Q��:�b&�9�3q����#�����oޞ��{����\*�Y�#Wwyi��ܣ��;>5�{���%cB��VV=,���Y�i���J%7'��;d�;d���N/��ڿ;�����5�z�O֬ҝ��ce������_D��{��6��Y���%/�ǂ�7�`2�X8�j�� ���$X����I�����&�JLb�E%��$&1<uG��.��w`�����t- ^j2D�y��=���%[pxhH,� w��>iu�
���E��� ������z�" �a����[+��J$Y�d�;Q�^����튥�J���(N"_��9:N2t,���ۡE�S�0@�h��CH.�=�����ZQ ��ԝ*, ܼ�#����&l�B�Sؿ � �hq��K�C�0�j��R�l��>9>�"ATt<W̿8�@�`��i��K����,�"�P$��65��n��Q���0s�ڍ�`�^4q'Rvgxx��+�D�Ei;-!��o֛�����R�L��� �s���:�lJ�iT��HIF�����i0DKafLR<���Ae��X q�;vE��������B^�2 �\�(�VَH-�iR׌M��=׌���cMq��6���-Te����}�k'GJ����@�Z���Ć��>����ٳ�z���F�o�V�P.TZW/^�X*��|�����x��A��S��2��_���ؕU��|j��.X��P5�g������՛�L�M M�J�(6��p �Ѵc��r�1��h�Q+�Cّ��3L6��nݺ���b6רU�v3l)"�M��=�������o�n6Bh�=�	�v������y��ǡ�ҕ�������"��ڵ[�l��~��W^yeqa��kii\y�Zo�M����x�Jy��c�=6�y���{����̈́�>��&;���ɱ�O2�����҆g��a��b�~=&-Z��t�z��+*��C��?��}�G&�v[�vg8|�����Ξ=���R��+)��&n����:t���O>���yI�/�|� �����u9Š�Ǟx�رc�\YƷ��ئ��U�|�GyD,�$C޺}�5�oܸF�c�\��矿��˷oݐ��e{z��W�<��FK��S/ Q۴�"���k�֭łx�w��#vrMPd>
r��G�J��@�s�϶x��-,�����6�XiI.��)�J^���=��L��xC�"6�Ps�c�������06LH6�����KA�R��Q���Ŧ����܎�4"��������C�u��<�٤�^ƍ��3H �H�!�c����;v�x:w��\WW�j���..=>B�cu�+�����v�E�bʇ> �_�~D���&sA�1���LFXk6�Q�0��aA�`�Q��s	����g�"4����0����pA�K%���[i�j+��Po��bD�Ֆ�ԥ�O��077O�*�˾�N��HV%]l�l�RY�1m�V%9��%��R��n'�N�l6��D���>�+6���3���+�K{���hW34�E���"Z��"���*�m1���
��8,]��N4W.��k�v�����#�W=����s�<�w5܅!�0%� �����)���F�S�>�<4�l �#a�\�B��Y�e=0#07�HE�D
�\�M����VBivJO�Ɔs�E.-EՊdF/��$&��I�y�Õ�N��#/�Rݢ�N炫0�Bx�W o�u�"�s��:r��VrL�5j�v��QS��j�K�1�C	�Uk�D�T�gq�<�:u
���^�J �P,�2y�3�뤾>��CB�p4fgg��s����M>�?�C�QҨ7��a�f(;霜u���Τ�i^�E���	�4��όv�`6:7���ra�tL�L� ��i	�L�b��K��]�T$��õk� 77m��裏>��C��ѣG�x}۶mP N�8����J�J�h���\m��D�ކC�	�{	[>��r`�[`N�ל��A9�X��L���>}���ݻ�wW�X�\�/_��`�A^�MR����[�J�Ψ��$��S6��O�gS�US}{z�vQ���
�͙��.��7 ��>�p�̙W_}u��&�kbXU�844t���|����ƿ iZ�$a;#��d�Ԫ8��Ź�W.M]�J�\����gD߃�ƀG`��-,�F����ڼy�uw2d�؛���6�C��n����7��OwY�Λ7n*����6�J]���̕k�^{�5zl�?�L#�N�`dd�S�ޒ�hdb��D[?�ұN�*��0��pB�B�F��lD�s![�7��f_�|^e��b��=��0@B�����6���|bM*���
�i��!&l��pITּ�Du�Wf�Τ��tzZ7�=\1�.��!�E�/�Ir�U���(Ǘ�����/��d2;��7��� ��Ml��By���qRFj��tԕ3����>ؚss3�c㨿j&z���`��I��A.ll���_������t~�{a�Լ���d*���:�)�O�~Q�X�������gʤ
�X�#�#T�Q:��W�U���I��O<T�٥4���sL��K_��h��N��Ư������?�R�Z�La�*�"�����\�� /.抝���
���_�KC�Zm[�<4��<����"Ca�k��)���
)��i��BY�4�T&5�i�3�<��/�~zz$�֋�]��,];&X�^Ez0���Ѓ�����U�+�w��]��ǆ����oA.K͆i��/߄|��JWxp��(��.�����M�YsT��+�qCWa�lu�g�;'-�)�X	�aJ��77Po&U@ؖ,�X���j$ttb������Oh����*�nE���K�J�h�L��L�d(`��V���d�0*���!�cN ��r�S*�s�A^�;c�P�(��������Z����밓����7]�蚴"�����T"q�d�/�&���*��n�4�X=�iO}���Dd:r��R#��r*����F�Ӓնn��6T�֟�C���P��uR.,m|�U�aI;'����֭[��
�~O��fLQ���+�s6�+��`�k[Q�Q�9���19���x�-[��ꯖg���ڪ� �YEc��/^�~ݺ9�l�q"e�@��V�1L#�2"CQ₭����E�a������c<P(ϟ?��WΓ�7�����v��	��z_��n6D���E�s����W��(�����>��v����?������W���÷�x�\Ш�d��c/9��І�0�����g<�@W��_�����|饗ɊCmcg�c��t��O>�����^
W!s���X݌�c{
�ݳ��
,�Lp||�Ǜv�I�	uA�5��W]Y=p� ������g/`ה�e�Z��СC '�����Pd�\�x�f�"ݴ>W^1����;v����_��G}dA|�}(��ظ��
$��9���胃������pxPL8��'�RC��G��]Sb�,�����w����UbCI��JhZ.j����9%�.]8ϣ�&���=�ց
������t�Ʈ`�B�I��e|��������s��'C�ٵ}������ ZH���lҧCxi�Yc@�^<bF�6�+0��Iٽ�Z���0�6�z��;��Y=-C2dr�0->K�VKJ�Wȑ���1F�>w��sޙ��	�����|6��O}s��E%��!fjj�d�8�3}@�*t�dL�@G�g�s�|'{���X��<��W�|a�tV��-��(�}S7⪈~�S[̤�������]�5O�I>_��+8G *Jv�s�&���&���j���[�H��r�Ի!P;������-2
v����\��B�:S+�A�r]?�wr�)�t��������F�A����Y1S�&4��쇌i��K��jPa���k��1�
��mO�	�A�@�}�v�(}����E;2߈tn��#��b$	,��H"N��J"t4F����NQ%#�v���J���US��&51��'�6�%T.�E�dM�t:�R���V �9ƶ����%�	N�B�z�DrN>:0Y��m���-��<�\��f�/-w�%ȶ�_�x� <�� �i�XlӇ)�!��'!9#F��M�5ztK�F��=ii3:��E��0���΁L޷��N۬���0���L�q,���xui�/���i
?�.�Ul����O?��D	��ӫ���a�������u{����g'�M��>�)��p�Х���њU� ၷnMAv��[��&���g=q��3����<5Y��@h-N"��K���Vb]��b��=O7q��W#�md1y^��ה�bw���{r����-/WWW?={�S�
�L47��,���pJl ����!�ft��I]�x��{�(�*�J������DKi�-�t镶�r�����9�N�ny^\N͟8q����xQ�����7���� ���C&��R���:�I�(��I6i�����|��H#:4i���ԳB^�]�#���>��̆�``�z��T�6�.�r��)���=���Id`�<�E�_Z�zaq���h������t�|�k�e�}[�:d��o��'fJmt<��'���uu�I��M����Ɖ(�\aҤ奎. u<��E�G)�����AN����+x�(����B��H��J�Z��+��
v�g��i���7oe�E�O:��)Y��vj�R����*�$͜��]YnZ���I�:؟��1�S�s�z���ӷ�޼��ŀG��UOא��S��o�۹�=׏��[n����'�!�O���XA�V��U/g_ߚ��6׋Mbcb���ɷ���/�ܱI����j��N��Z�,�{囲�T�l|��7ډ���XҰၣ�=��1�É-E� �ID�;Z��Q&
o-n��Kvu�����/) �fSb��B����c���(�Z�l�l0�~�8=�ȅ?���OM|����v��7[͆8Z��|92���؉Y��[�1�3���3�q��1CnA.�XxH���Q�2A��"t���	��8̗ݵ�������n�!������L��w)�7�KT̻s3����d"�`Ka�����W�V��RR��� Ԧ]���F�o��� @s�Zl����{�N�C��m\le�f�+A�~����Fz���>C�&�ZD��Gg�	�"�{��a���e��X"'�bHM��Z�����S"��ga��;�B�<U��V���A�P���"����^�O��-�\�5	�<>t8^�r�ف��Ĳ�n%髮��K����#�M��y?_C�P��6�=��O�4P�����GF���K~���?��?hrec�R.l�۱c�ѣGڿyb|hd��Ud@805�좛
�B)�}��9r��g��r���H�Ph���4��J��T�k�jQA��s���|�(9�+�T��'���⩩)P�������?���\"���� ��h�䖧�zr��}�]�֑��3Z���������P�@��zKKbsb��F�>����x���|�xЅ�8�S�"^��|��I�ި5%�n�<���"����8S6��F1�������|�Z���h�E���x>��������&o��/*|�Y��!PZ �Ⱦ�ݙ��᧟~����`���Ǵ�L֏#�J� �>�j�)�Ƹ�Y�ެT[���=�gxt��_<�կ>��c����?�aQ�����{|Ϟ]�V���zFG�aU��ܺ��e�8�X�4�����c���LdooϱcOtu���_��ר1���&�N�X�+j��݌�[��{�7���4C<t�N�$}�ݴo#S���������['O�����B+U� �wm>��1�ҵo�����cU�9�������/>���������D�b�w�yo��C�� ���,N���vLႉ��rY��j��˗/��CL��~��Z\Z"8�ڛh��XK.Z�W`�\��^G%Jk�PU��A~^�Up���4k���îA��r�f���K���4V���I[��i�&a$�2����u5J���y.m9�G�D��B&��7G�m�L�Q,L�n;� ��x -Yg]	QZ�!���|��$e�mD�n)�`�F�VUwT�RH'z�c�:\���j�M�U�Tf��*�]�֒��\���/䥼$Mn0��r�O:δU=$m)*NȘ�HO� ��n���,:&�㈭(�b�K�ꪸ�6�7��/U�ȨHKtV�P�p� q���Օ:�4
�Pס�V��M�Y�q�
EO�Jb����&���YO��Ao�Ҟ�y�*uE{4�M�Ɇؐ}�����n���>i�<�*S	�"b/ب�oJ���y�⛂k�Vb͘�x4x�h��ܾU��"�놋�{mġ��j6=���I����K)�(l���l�S�|_%�r�5�E�)�:V v"��%^�okOG�W�M�&s^�$�i�h�;�<|O�
��ƍl�X�c��y�;�h;��Q�%� ~M�a6M���o����s>w��!(�쵅7`�L�%��ܹs|�ۅQ�%�F?l�Җ,��;�i(�\��i��:0ՑG��>�5�8��+פ��\S�l��O�˶��suiYQ���˫+K��ݽ�!x��ԁ}�w���o=���[�l�!I�^0�={���8u�{�blDWeL�Kz��B�5���g.�֗��jҍ��u��U�-���ΠN3�"^�e�@+�$�I��l��\��.�<�_�pqh��4R���Ȓ�$G�U�P
j���#c�O��"��҂u���3���h��a�Wp>�VsN�
����Y�Y\���9���0S�!T�(��f��8���K*��AiXhm���v1�(\=���LwA�MfH�ܛ��|�������Y��S����(�0���n�Ԃ��U�W	g��N l�Abfd�������b�b�\NCG����m�tz᩽D���)��W�� Zй�Z�b960�m����=$�g3���f��L�P�*��/e��
�zr����[ׇ���f��zTґ%��uYse��n�������kq������]f?���3��E��_��|��6�}��Y�.���C7�� �!'!��� �	B;�ɠ�p�1��_��w���Y�5�A�c/�06��q�ԣ�\T�|���blt�W��6O��}�pzk�۴H�D��"e�f����u�����Zw��v�$�p���;S�=�P@��k�u׮߽D�ı���bW���8&�4�;+Yt����i�I�րˆq�iف���<V� �Ѕ\��E�'0Ep	$G�Nw�1�������ǮA��Z�	F~�FGG!t�%��"�gAÕ�S,|�P�N���������]?��ψ�&�}��۷o�GpO��8N0h�'ӂ�U�OC����̓�''�nܸ�U��#����ڮ�*��SdR>y&�$2$Z2��hD�Z�忶�O~*��%O�z+�`�⋘���-,��ǴtZ���dliU ��j)�]%h\�A�~��ǯ��z=�fҖ~Ӵ�e50�|prr�	���[�O�%���M�0�u�M��PjFZ����1�~�l�(�B�$H����3�!�p��ƅZ-��%k[o�`𚝝�	48�+:M֏L�T*+�p4�V�>�RQ�c�6�IX�s��$��[�������/�k��<I-0?-Wʲ��2�g��玱٨�s�h	�L;���b暬|�!����?�ך���~�k�$Lר�FFFr�n�^��Or�x�	6���H��ϫ�_�9��P�A����7v���/��/��կn�Z�";v�駟�R>4<��,2��\d𔗂<�x≁��������w���#��'@s��j��B�H�1uK}�H�Q�� `�A"�@�0B�ן�:��]O!' ���w��/T�&���fJ$����T_��z&&&F�G���S������	������r��j��-2�:r�N�>,c`P��9F�ȠŲ���Ķ��b�u@$�4�Ҥ9�7��	ҭ��w���#�3�M{�ke���4�LL�}���Ų�0�4'�KmY�X��89v�O��OϜ9s�ԩ��y����`��hM����ЧƢ
���)U�F;���!�n}�#�{�nV��M������FU9��H�c������$T�3�X@�䴲a�D��}�bj+�$�^��hm�$Ap.�>~cx'N�x���w��aF-Ԭv���8&����L#������g`Zb�8�X\F'T��N�r��q�D6:�#���ݻ��Y�+���i���X��~�R�LX�q u��\��(�i��V<���C
!4I��)�N-�~+�}ͷH�+����}E�594K9E���j4k�Y����S+Ma�L�i�^�"�I;���p�}��	�7:��E|[�����b���q�d5A�0�2�hb�f<k��Ҝ���o�&�wcU|�O�nG����c�A�s��X�����#E�M��P�kF�l'�Ϣ��F�U*h�ۆ6`�	k���U��e��>��	�\K�[��t.�c,�X�Br:� �>�"�,f�&W��U�7ֺ�'��%�[�:�9r�0�v�[o�if�5��A㹦8�T>��Sۤ��&hF�j���l���g���j+��&
�:\y�*�K�ǸM��&R��ap:6xxgn
�K��E���T�~�d�Lk%����*���D�|d����k�L�nj>tv�,���{�Q����ӎ�]n\Ӳ�k��k�<�E0�_o���;���c��?3a	���@�&���م� Mf�(�]�f�b֐
Rk�&��Y@�����3nĶ3�8G<d��/�]<|WŐ�wdp(P�<�ǖV������m�C�VX�\x�����{�1�'�%p:��{��#F��@�1��i���Ӎ:P<,���\�V(	"]�@����|^q-^b2ӭώ5-�����'����k�Bljer���޽��?�4$ X�տ��K�6�B_:N�<���x�z�HK̀��Ҍ(jw�)s�#�E`|�t��%�V��O��igQb��/:څ�+�Gc+1�z����s�����Rx�$U,�\�&O�:��;�#��5�w��Z3��;����Ң�u������X��D�R�AK$c������Y�|&B�ȡ�2��)�1��)�@v��_`�pK�C},\72g���`�k�#F�4o�
nu~�9VضQ#.������C,9���~֜��݋�S�)�Pk���:����R_�:6��t��/~����W�8�����%��扝���+�Avw���$�4;Z��姈�BBe��i*��V�Q�(H�hS�(�Oٵuj��Il��=��ǯߡĄרRpX �v$����=)���*��m�_ɂp�E(����H�"���
�n���\��\&��V|�Y_���VZaT̲k;��,<zU�r0�&<����;��wH��HJ�\��ŝ�!�k�q�Y��%�5tyO�O:�����w��ҐL�I�0�72ż�x]��Z�^J[�SĦ_�Fћ�S�e
o�T�l4�8���zX���6���y[ѷB��h��M�Z�F݉#/ж8/#�n\%�����C�i���V�rq�����S�����årV.�f�ϰ给�a�<ǰ��K*a���˛�7~v�,\���R]Y������`��@8�� �rXG�'�e��O��-(�r�'�+��d;�[X�`C�">��s\uld�����o���}��6l�$���B��S;�r.���Z����fW+a ߒ��Ҿ>|�ZN� �������O~�92�Ez��@�P��(�[�3%�5]���.׊�]x�I����ưV<�P�Iue���iN��%%��Q$��9}�]G��r�0_�%ڮ���$b�73��o�-���ׯ߀�W�W`G
���QH��nߍ�:P��|��!ݳZo��	D������܅��TJ�C�w��$������ĉ覭&�B�$����6$��c��0��~ࡇ~������	�hA���}�7��n�8��[jEMe8��>|gE�&<q0T��s����x#��J�]ӳS�n|��C=t��Q6T%��ę�9 �<>h?m�	�m۶����7ofs�S�N]�t�Q豥p��L&e,���*�㌧��T��%����H����˸�رc{����O:?;��58ԧ���~��GX��J�f3N�@�l��5�R��0����=|�{���'%�8�d��~6v�˫�������>��ߵ{{Ww1�sk�e-R��D.\��*�λ%i�,��hǞ�/E'�xn7�Zk�E�k����m��%k��~ZNN�Rָ�I�21�X{>n�B����v �M�F�h�m0pEf�Ν�����֭�;vL������hV��[,�K��������(��g!��!(���{��o���0�����C�Q����$�A��U"��6��Qb^�(�P1a�m޼qӦ�l�����Vʩj��`ǲZ!�>��֐�r�Z��)��B�۷oǊ��\�R�]�7��7鎡+�~�[����K�A�:�t*�
���h�&�N~�w��-�~��?b<�e�ax0�G6�`6�V��`M�}d��h=����D��Z�������UDt��	�w�}W>ݩJ%|��݃����&&���c%F����>��j�E2M*���W�$R�J�i�]+h�t�n�#�(�G&��DOPhZaq�yu�����������eO���j��:���y`X,mG�l&�?~��o@�T޼�3�4��b��.=�m 	��\.i+'-�D;g||ro�9ي$0��<��P�d�wtl;x�����L������Ɖ�ųΞ=;�a�>u�v�Yk�S����]���:�z�r+q7��Nc<`�ҳUm�D��,��?��Π4�� v�#�uG!R�,9�5\9;�\�`�g�)T����+��f�Py]�c����/���oƽÔ����cd1���8ڞ��t�_<��{��aR'N��V�JL@�V+�Db�B��-�,4b��2:��i���`U)�]��ƚ3+
��b��4|�-����Q��C�e7m�҈=���i���	�>�U�BQsl1��&*
�Ċ�XZ��Hd�{V���R s'�$�2�u���d8��B�T��'ӵAo/����;Ku˥!�9��t�S?'d��N�BQ��)��P~�����C�+dee��z�]�a0�����Ν���>0 �� �0-�AS���O�����|�
���8�K+{�zp��бH�fp��R$8�w�jp��{ұJ�G�V.�{��f����Ü�ؤF���K+�m&�vځ��gđ�u��0��ET�hPL����W/I���=�ϥ�KG�B�<B�@~�a�	�Z4!��'^�v���r`L!ʙ�F���1\߳�Ǥ��m����Q�g�.|Vv��Ÿ�#|2Mo�Ҧ��vT�GF�U��Hk�1	����g  k��0L���~����i�괕v�޵c���|JXP}R���6�F7�I�K�J:�gg�v��al�m�����=�� k|�8�ݙ���P��E��K�1H�o��ƥK�0xڕ���K5dᱞx!�z6�o�e�7n�x��]i�4@Ό/6Z�ZC(?v�r�462
��" �E���c�a�Dt�_iK��D`�\�˦ܛgН�oZ8'�!k����q���69����ㆲgz��d�{[����x(�֫��K:���/��+��*�F���M��"�k�7�o,V���jÁ��N_�����=28;?Y�Ȳn�{zT�����������y��};�&�o��p��@���!~�3��Y��=	ՑBji�A ���������N5�V��T�>y��U��4J+#2p.3f���i�s��E��MSϤc���b���JF�G���^I[�\�f���)�+GU�@��U��p�D<d��i"�rK�.դL�f_;�$}�t:ɢ�kv������Wv\w��ܻ�fs�ew�'���%��ļHXT��5�⭴Zb�.|�˦+:���X^��KP�P�3$���3̠�Z�/Z�`�R�/-U�h���J�4J�R�K��ȳbS�%0�mM�3��@+��\���Yb�VL��_��;�����G��ɭ:Ń�ei��I��p.���͛���oc�SS�0}W+u��K�qW��P=�%j�-SF�Z8C�ԡ�tX/����˝ Jǰb,��d�҄�v�mah/��D�(�D�S�}��+�J1�5$N�� ����CGw��oϵ��K���`���k�?���믿>=���a��$���tsC�c�y*YSնdLWj�B���P�ǣ�������h�+%�ڴI<��?�����%��31�N��j�<�;c�'N�x饗�',�ٲy��SO=�}�v�����b�B��	����̱��{�_���7nܴl:0���z[֫�����9Sۖr�4�rL���"�{����jׯ�Y������	5��Я$��}��B���A���:�g�֭��@?<)��`��	�8)�|�[j�WV��iEZ3�+�(�d�A�6O��p�f�BNgZS��x�����7o���o��aF�Ǐ��׿��O"�� �����X��@³wP
���&w�Q����>�ǎS��_C}�Ca���.���5��O<������qp���gcV�h��M�Ě�ܴ�*y���,wk��d��8��g s��L�e����Q):�]. "�ee�;(a�_�t�-�̍L�$�˅�q��|�Mlbδ��&B�U�9s����1���x&���1"�>|��*sI��fL4VD�
*�%u�hY�3q ��"����� p�<�;cl�:.���v���ps=
(�<S�>w:G&&&�������߇���6�RG�]0�Ԟ_�*���o�j� �
>V�"��v��~�v+ʙ➱Xș3Z�R��� �@���ū�1u�d��у�ì.�6E�xpl�.2}�y � c#�MU�f��|<'��@���)rK4Yb��� U�7=��Q�S�O�\���b��b�U'l�Y�:�W���W�\����yeEIh* N�E�[�2��lD��
�L��!)��5�i�T*��ޮg��>�[6o
L)�$]Z�D�`��=�?w��;o�K��2sdo\Xn`��CTcގj�X"�/ĮU�J��=y�$v�pq�,.�2Z�a������,�:U�8��$G��hQ��*h%4H䂨Ř���\�b&1`~r`�OH�GҀă��)�XY��4
���s?�0]��3���+�����t2��4��$�, y�͑W.�[8�ܵM�*z1��N"Is�چ1Rvd�K�:n�t�Թ��	�P��J�b�:�V�Iߤ�x�p6��l���?�̆$Ԣ���2f���*�r�J)Y4�~��X����YY�3F�Q�X�H�L�n!��y�M!|E�Q=]���t�(w��x344�����|���m�/-5�Pp7\@6h���c8�ͩ��9m�y���+�1FlC�bL�5.r�@1��Ȩy[�_,f���,�q�\4���$�B<V����W� K�����?�BWW�>�r���T��k�%~GQ{�#x0�\�[֣�F���=d�P�������(���A�P;�0/���A/�a<؎�F�46�hL�/ް�m|܌�V,#�t�U#��PR7��N\�������l;>���(E����͉V���_aL�	����~<����G���G���}Zb���qŵ
�j�S��M;������(Q-Oԋ
z�z�*��HRމ�xFȗpg����p� �acW�%�͆qn� q�Pñ>&������I����T�'{���¬iq�.�0�u�V�g��҇r�Ui!�#�0���/�_n��3dL}:�З��l�β�)�.�Q(�-X������T�Vn )J���U��b���Ꙫ�κח����e,k\4ָ�'4�
f�{t�+Fk������N�O������``
��=�ʎ0L��3��`�^�FԬ���8�Z����_��l	|	�沙T���f/���(I���|�ܙ�Y\<����7n����`-P����+�yg�\�	*�Ԅ�� ã#u5��
�qs�@�,mB�cĉN��ĝ��NoZ��뤕ι�s!:�g=Y$�mǗ��΃:�'����5#��$w��wy�퇝�J���$�ߙ�o�ڭ����cV�I��c��V	#���ה\�1J��d�X�S��_�d"mS���f�Y��/
�F��#n�Pk��H����X!7��i����$ހ���]�~�Ѩ���۷gll#k3����K�CHr�#�[�F��*ƻy��?������tJ�+�������@�C�{Y�I�&(ю�]%Z���w@  ��IDATH�f�d1\<77O�{���)�!�N?��D�O�?aWlݺ8ku��?X�HA%���FԠ��MC����~����u!�BI��9��޽?�0����!���Ǝ=��d��X�BI|u�G������
��L���)E�mK�U禨p�q;H@vj'�;�I��c��7��v�0���k�u�ҿ|(%ܶ퓓['�z��o���W(o��N��w��Ç������1�2<(
V��mBGe�����]�����ZX���?n*$���kO�M�F�%��zƩS�xʨ[Gy�Q���~���۳��g�����?��c���B�D�"tt_�hZ=ʏe���f��fQ,����^�@�����8<R��H&�����X�rw�@;���pNC�CB�Ť�z���nM��'L�#�a�生H�e�uE��T�Ȕ��q�z���Bh��n�Z[��%Ź����%��O?�a��矇����'_z饕9I�f���KF�׍��\��U��h]KW�w�Ƒ��R5�W�+Q[�n��?x���_{~�����+�RyqaE*QF����r��;r�!�#ż��S|P��E}}=�|nxp�Yk+�_T"�9>Д���R+��M�:�v�N�U {�2RaJaJ�":����O}�k_۱u���ԥ$�����3g*+��(xO��E�ڹg���ZQ��D!��DA.H�D��YǊ��6�J�d\������� �-���� ���/W�K�e���<]?�Vj�,Mp�x�_^����� d�D���{��޽{'�=�!�t��L5�%�R[̃�R�KJ�����m%NP��� ����.-Γ�4�+���U���ڱ�ԉ��f����-@�U���2'L�bqt�&[MNN��׭jk�P�,/�1b��eW+��� �Dj�n<(�H>�藿���<�X�R�P��k��U�4̥�2E-Ҋ�s˥�yƒN�%��]���?�w�Nj���/�[���3��!f�|��ɏ?�xqYj�
��M��/H�={�l�8�4&�ק�~��g�=}�I���V�|�I�:����ƛo3��s�Rc��cv4��]	Փ;IӝR��������u�����Q BX�O��x���b�d�fԸ��2Bo�'�y��d��-�����OϝΦ�@:|At7oޮV�0�u������R�1����l�СC��Υ=��ŅeE����r�I)���0���̤({�݈�(�/[��7���Jzـ���?���DLJ� ��զ���+8̋���Qu:��i^����	�T�(�b1\�>	IT<-_.�$"�����]�{�I>ۇ�����^Z���]�#��R]�Ÿ��Y�|w� �#�nЃk��&��jD��&���u��U-V��"؞)�@�'�����ե#�3��m�|�Rš6̦֓���(��,:�/�Y�>i��@�d��n z��7�NQ��3��:����2x&u!�
�N�@i�"e�ԫ9)�d�7A��6?�'�pV���e�j��DlW���L.�g���*�8��=evVQ'��u��<~���3��1�~I�<4�ď-n�A,ߔ��W�K�׎�$#a�z�eT�B���)��%�E8��Dr	N��� ��[�P9���A�咅�g'�Z���o~J{F��r�
,i�3U'W���j��RYm�B��)jz2a4��qM�K�A��*ɸ'�~�� C}�����;w�B%󮤳����sƔ�qL��F"'4J�;22���������~�;���ʖ�>N"�a��B
,S-h�ۍ����eI�.{�������цgg����Q*	[h��?�����[S��M���#�S*�A�#�s��p{�%�*5q4[m6)�$�L
�'aG3\�� ��=�*�l��6m�](����iN ~,�?��Ĵeӣ�jcH{5�v+�\���[HQ������x)~88�CGm�1�����S��%�U����.n61��)�& b�������1/�;�é+
�͚�gگѕ��(���D����j�I�?�L�v�4hͨ�tw��$�ДS(R}��M�/�M�q�uzQ�'�v�^sg����_��ٗl�_h�{�9�yw0���k�>�L;UZ��YB陵S���5��Z�6�wU��<#���,a�=.yBT������,�;S��6`�K���v
�X�8��(f�
��蠣tb��3rH��[Ŧ�w���S䶅@G�1A���S�+N�3��v�If�K\l�b�ĝS�t�u.b�~ߛ�^����Ϛ;���9	���d�:u����r� ���r��\�aw.��3S�$&`Fm[t���է=�Nn��g�P�k
�[���/Ue�;����8^�PPh'��$��W���6`e�*��� �R�QnR�q�F\666F���v�u�*IA��e&�0��n��C��a	�V��TP��IC�X��b��B���:�
�������y�8[h
ْ�RW��wL1u�C����w���h@[+
y�Z*d�l��.�:�N	/�6p���͛���G?�V樾�϶�Òk�)��`�\�t
L���xg�1o���qRݱg���2]�BS���K\�ss��T��*���ܤ��^p���ҏ@���D��S�#��[�Z��d��� s襗^b�Ig�G7�Y�� �|���͂�XQ���@�����{��G�z�?<����v�r	f������1�4:�/�4L2cG���Ċ&\_����z�*T�@l_�x�5M{�9��8�aa2#�ɤ�IcY<H"�����?�tC����U�T�w��K�.��J+L�@�ӗW�'''�n8pӢ��� ��̌�K4��*�Sl��#�6����)��jM
j�bw5��:zNS
�Đ~��_}��_5�ڵ�L���ZY�7��'3ŀO�8���>����X���K�vU�V4]�3�D< ��"1Pn��1	���Yd�1�c��sE�L��	�J�n=���`���r�fG�e�*��T�&+1v��<�k���88�̿%�pAO����̜<y�ʕ�0�0�͛7�Qh�[�%��x�۷���&,#�T�;1���gϞ�����=���dA� m ��5%V����o�rjgΜ�|���<�~��k�����>��Wl�M|�^XX��	e���B�0}���cZ\��,{݀?����;`�b�,��Ԙ���=���?�1E���𕮮��.`HNMMad����m��f}�ڵ�{��UA����b��c�+1d�
�[��n�G��hL7WM��b���#�?�r��;%�b������|W>����=�ܡ���M��Q�=�a�T|�\@]X�۷o{i�<m��>~�8�plÈ�J�Gy����ADb��O<
�J��#G�<�̳�������ɓ��$�J4��R1Cb�0�qr�1�vM�G��M�hMb�t�O84�U�h��JR	,2��嘢�T�$aml�n���b� �gnn�ʕ+�)VHD*����Ķ-`� 	\�f�~�Q��!������JV��Ҡ�d��=c�Ih;_J����<
k�-�hd)&�
GB��7��F�y-l��F̔bE�^O��¾lQ��}�]	q��w#>�1ur�1XB��Z\� �-�(�b����QZ3:kgM���eܱ�]Nf7����4��:�P30�M1� g6l��"��k��$��y����ǐ�5I�J��3ݛ�$r�� �)ȢqtN~�B�edը������=�G�:�h�[�r�ŬU�Љ'%��jˢF�,k`�8�H���#+�7/�Ԝ�X(w�v����@�%�Dً ��9�?U���F��c��>l�c�a�vZee���=ǯ�>�x=��h�2�hQ?L�PQ� ���v�V岨�诤gD�M����R>WP)_�چS@`;��L��^0�r@��
�ڸ�T}E�%q�B��� q7p!:\�j�#��3�H� L���Ȁ+���꯰V`��˗�Q���f��6���U
�0�|اvJ[mO�6����%�w���w�& ��\M��A�0�و�c��t�Fü�Pl]�'O�(�I��ԹǮ��tgcGl�U��If�d,H��Py�-~�=��Q���V�~�)� `�R�>�'�U��VWx�xءo��-[�������&"cbS��e��c�_[_��]�S>F��.9�#2-��[��z�ԙ�s�lב�T��ݤ�8��y����TH�aV2�����g���(�Z.�K���Uڏ���&�	���?b)��~�+�R��_���Y������t��܎Vuk����?��)k�E�O��[�Ƞ�oZe�tT���eP|J�y���ʭ�=�TT(��w#Sp����.l�]���[�F3_,�_^�;岏s���I�[ub��� ���j��^ǲ�a��5���)����ҁm���0RA���3rb�kVܵ��5<QN�X�~Ǐ���s_O4k�;��]+����I|k���:wΚmZ���{Z�-��1���tu���^+6$k��o�������y+M�H�Q��'&p��厺���"����Oue��i��2iI>����X9�Q������_"]a��$;9��\�V@JZZ����QSc&��7n��4���C��eBݷ���ԩS��!۫�.�}k��ڊ��v�%�㛏`jp>-��X�����BO��ȼ2�(ui�;4�����ե�ze5�)^��B�a���=ɚ�Y��4�M�)��,�.�/��n�8��m��288��l۶u߾��� q"q'��q'���)J�a�u���J��u���	f� +��N�u`Z��E�"l��c��'v]E�k����33*9<J�)S��8�Vr�N���w�s�f60�m[w|��s��s����W��!� ���"Zi]Li���rii�0�Ii���{������N���9�Պf�V�UY1�*����-e$�����/,@��Y̖�B�qr�U�#��6??7��w�葁>B&g�\�6�A2���zҾ#�����Y¡<�L���2u{�R�9��,�������z�Ъ����e�.�S� R�9���;�JM��M<k��� � ��P�����
=�ٳG\0�+P�a�TV[a[��`7Y�6�l��`���P	\�tW��x+a�[����O����򅋟���K�=��=��8lhd8_,�9G 6��l���kҨjq���'�@O>���-�Z>�q�TeUu�W��	;�ξ���Ã>������}�a2�]72Y��?��(�N�ܾ���)ɯl	��-�gj�\6�%u�9�D�P3�n]!�����t;i��m�p��+��ݺ9�y�f�kX�=&POO��:��񉅚��[�i"s�#��+��K��o�Ol���|.ϣJN�T!����~�Rw���s�h�X>	��M��W���~������܌ 47��3c�p�c�-��D~���}�����gа�x�Ӿ�ύ�.]���_$�L�֬���!x]�9e�D�s'il�U\\���:ˀM��ori[�J��BT�R0Yh��|�g?���a��2M�_�j]H���r����k�d�5�=�\��'O������Ѡ7��4�ϗ��|�H]���H�6
�Iâ�(
:��Zo����z���j��J}p�g���x9rd���0R�L��'�U<��{5)�8{�l�
rꡇ:�/X5ٜ�5M?�5��I�|���L�@?m~vNp����J�}v���S��	�T���5b���8�QRw*�9��g�3��9#ө/�#;G<x0���7V��W��-W�,�*KЕ��x�`�aW����Ο?��M�s`hX����� ����Z���?��W�2(�Y�N*��k$�A�qRRSX��*	̺<���ռQ~�6%����;N��1pl耣%�IA��4���ťz�JeCj$���S���х�Fq6�JeI��"��-@����sS|�6�UƖpj�9?��[5�
b?�eo4ø.�b[��a~���z&�{-XI��]-��7�*u*1tA�\"(����ͽ���T��t�fMg��˅P#��,���:����7��$��o,/�J>�d���}�=kQUIV�ՖKr۲����������4�����a4�e�fZ*IU���ʬ�3�3���o���Ž�̲5�~R,2^č{�=�,������j�c%�9�$��Bs�����]Y��N��@�� 9;B񇕺-�Vdff��8��4����i�r62K'�2O4���S*�-�߶��	�4G��`�v���I]{��x���	,�=W�����Rj��m�a�������r2����mALj0N�2�ą�]+�����ohh�-b�� �[#Ĥ9�C�p@���IWys���ֺ`9a�F����7�F5V5EH��8��˛��8���������g�}��Ǹ-�˃��ˌ6t)�82eom���؁���C���J�9���'����h�Q�)\il��)��큅^%��b�����O�-7���v�O>I��蹧�	,��Z8����Ji��G*����h�-�6j��gF�T��iw:u���D�%��9�[!=i6��r9���,:?�EI���:�z��í-A+<3`lS
��h��ƕ4�X��Z��)B�#`�=�zp��ZŎ&����<H��x�f�7�nܸ���q���NKK1&�h/�f�D6��~Y�mii��9�*ys�@�����N�Pz9fT�A��p�n3l$N��֊�$�-}E�zJ��FCκ��p&7o����F@� ����9�ls}C��Q�t�mt��J��|C��&�ZA�ʭ��on�w��7�|���{�ɧ�����O�������8�͇�n�.��=��0�w���K}[�u�?�Y��G7��Ӿ�c�s4�{��A4��6��[r�>.{���CQ.&�OZ���r��-�\�;è[�����-�g��vP�l
�DbH%Z({���5��ݮ�U��tq�+{�d�z�E�h���������o��{J�7��y9�s*�0}�tq̉��d�b]Md[7pn�.���2��*+�Z�M�[��K=��8��~g������Y{�m)�*��qW�|��B���5�ܡ7�3�֭[��׸�48^�1����)���N�?�������CkCK*!Z緌�ψ�r|A..ֺ	�a�)!(.OV��h�'04q���q*ql��X	b ��ڮ�i�Ή$�a�\�zU��#��5&l{J�S�)x�R�YŘ~`g��1�c�vZ�.(އ��[���hDxY�F��B5C���[�~�lD$�6�[�*.�����w�݈aG�L74�ݻw1�����qە3'+�OX���ŗ]Ƹ�����j.O��ӧ����_��R�1�n��RYM�HP�Q����]�(c{���덱7�x�wޕ+�#�ǳ F�����^�|YS�]¼	�#�Vs�u>T�zb�AԱ�O�:�V't*(!?�V��ė!�_���KW��Đ����0�~�$����Zjg�Z������q7X-Z�|"��z}�D���O<}���T�CIq���y����1*1<��1l*JL�H�N�[[-��,W���0���"�o����Ç�;I�<�1=�T����/�l�o.��*>�㯏V��|��H��r��D�)+�ɿ�����SO�"O:%��r	�I��1Qe&�w�ޗп2L������CU����lC-Zr�������������6R"��[oI�\	���u8��ܼs�/�p'�����<��s���*br	���fg�)z|�X�:]E���,�d�N�����_�v��͛�M�>�C,!0���;��3D�>0�1 6 6Y^��!I����x��Z���;�p�q��X�Px���@G���I�|��/=�Cl�!̱cl҄ZO��P����O�HT���LN�i��8����%�P�O�/�בF�ssssJ��eX
���֨.5���p��F�c��Mp@)����7*�\� kj�,sIJ�)�w����f�hx��~����~�;��N���bي�,�KY�=M�/��捝s�]�1�X8��3I�L{H�3*kqJ�g
K������e_�x*|}����C��,�D�Zc�ch	p,�U d�Ck0}����Y�zM;n�s��S�1�OX�AN#�F+�I��P��!T����[����Z�r���_y�מ~�ILڴ�#��+���èp*�U���|T���������Ж�z�[��>R���:Ac����FY�m��ٷo���(ɁK�.x����F����  �p<a1Չ'p^{�H��@3�aK.'obÛ�9v=�	n�/"��x��p����a�_]"+"��Ҽa���m��sw�,�cC4&���ߑ��rFF��v8`ђ��)�����'��lw`�����%��\	��o9�)r4`T�e� ���(��.2N����)AX`y<�����|7N#tb9a r��e�I�a��7�1�)l,�eQ�@�Dk��U���J�Y1��fg'����2��ח.��`��!��?u�����T3>B����}����a�7PK;oY�)����a����W��Hc����R+r�Ԓ�j�L��ěB�����ڝ���yBm�B��c�<�����7;��.\�����Z濙Z((�;w�p�<[���=F��9�^w4_������o9x�[��%&(0uЈ/��՗C�BBr߾}8)px�0Bp��v�xj����h�$��n,H[�_������M>��sL��lU�IAλ*G��]lz�P2Pu��7n`�n�3l}[8��r��N�R��:-0�X���3>H�f"��X6O��D�m�88p��Q���/�O�|���+�V���a��w��5f[�+�?bt�jw��4����:��s1�\,��D�;9�N���p
PC�̃2���l�
մ��'��A_��<a��nwy��@?��P��O�,.)�v�⡃l��$=�ki�Z��$w[[�Ī)a��f$�MX�����y\@mϟ�[��|4b���á7 e
���0��������F���{=��Q�Ĩ]G;����v��m����@b�+�א[��T�;)M��|�J06�o
=��^t�]�ߴ� �7%�D���7�^R��;�)��b�w�l֜A?�����4��Q�����]�n���%��4u	��`����8�X�rQ0]��G����+Lb�a��,��{8�ߍ��R|e7�u�4��� �םz̨g�#a�$���C�F�NG��'�AvEM9h�9?*�%9F�Jfe�"���o\���3N�����<������V���i�������N��\kNL�O�����I1���R�<�8��8�'��ڑ
�4/�IW��ٳ�Q(	s��ɉ�	��;�����6��da� 4&�d�
U��i��v�-"31�����X�����z�4(L��B��ӢM��4U��1'Owq��m8���Fp�a�^����X�8>��H�Oe�г�q05!=��'��~�V��@���C݀��8#q�� ��M�"�@���I��M��cCW$��Ch���щz��q@B=}���l�E�T�DG,�39�q�	�~��
GT�65�R����0�L7ط��������"L�0F��I�VέFy���ކ����Q�{�M�G��S����dd�0�K��ܸ�o�s�n�yy�R��\n�"�!����
��n�R�rBp�Ò��]�&ݖ[[���8�X���[�J偄)a�6�����no���fm}}{v~�ĉS�J6�O��،�'���ǟD���O<����_��m�ľ_���R.��$����c�6g4��B^��t.&�����ɖBq�c��<󗡥�+������
sT<�m����Ri�ۋ/�*=rd��o����������rjxa�/m�m^�xee�v-*�V��%W.\�� {���a���Rƺ�x�]�x����8�|@�ܾ�}�g�8>ڄE,ZD�'�
��Υj4��&��3�ǧ'XO���6&�Q�I�~�C��8/goG$З JM�`�zc�a��k��NĈb�x�r����������kk5�����S�ƾ�9���СC��-!;䄂�TQw������vQ	=���V/pu��8v��?��?�?��d���4��?�~>t�c�,xӝ�mL���rĄ�^�h����_��ؙ8���I�������?m������~��SO1����T4FI)�1ԯ����^�������X+�&�����&�1�
(�c��0<x��{��ի��I�eume{goU�-���>���:1��(�x��ҥK�_�?w��]:rׯ_ǋ�qЁ��l��ԋ��Wݓ{+Z��Z�VnբR��� ����S��N��ږ���d<g�e�6\��tĎ�a ��'�y��l���H�PhoL;)/|Ix���$�{8�K4�E�e���I�����3P�DT��;�D����7�>H��!���fl�&�o�$�Y>u�`uU�FF�!g��甯��)�p��:��QB�9b��u�f�H���0I�H �� ��gi0�6%)�><���r���,WJ��-����g��8��q�P[-s2}e�&���1H����ҕp�p+tS���ν��K��ַ���2a,�ж���~�H�_��׫�v���K���4������N�z����q�?�(��)̲�5����A1�T�P���6�p�>�I2.������Բdꮁ&�HʕJ����^���)�of����cN���O�iY�h�$�ݭ��=����a����<0cı1څ���zqqQ�U q�v��Y��9�.���Va�A+*,��$���m��Rl��ۂ>��N\3��a���R���C�?�o��KO�C�p۹�)�}t#���2'd	�q�*����.�Ҥ�z�O<AJ,(�l�<1.�SL��k���������}�{�
q�H���̶�aܹHC���0nBÒ� ������煚e�����ijG����ѳr��>����5&%�������������S�5��Q���>4�GǄ��\���<S�W�4���=~�������Ơ7p^D���t~^P�ɁA*[�!ň?KD��Č�$ZM�rKCfR����d� ���ɓ�����8Z���9"��ƍB滹�q"m�g�g�}g��W��.U���o�[^�.V�������`��eB3o5剙��Oe��a4НV��A��ރ&4��w��.[-�;2W<�Yj��MF7aX9����Z�k<���l�?���O�s����QfR6ޕ���8���߶f����{xlB�)�s�&́[� �I�����_�y��C͒F �̙3�\MU�w�y�طq_�dr|b ����-�vC?`F�e�`���n8��a;��l/`�e����q��(�.�����΅��a��,E����
i���j��ۺ�����e�c��y�t�c�� ,#�B� ���E	m�,�s���
4a�TYf1�{F��1CL��\r`C<�@uYa�Vk�\k*����$3K7���G���@Q�#W����@So=��K2NdM:A�@�c��J~b�˼��TŁ�W7���ܬJyBE���4j������@�J�Q'�ة�Z�T���o��{�h{.~w+�~$`��*>����~�W����D��Å���IOM˴�F��P퀙��i���`@*.�U�7�Z
�g�F�9��u
��T�{��a��V�;�ʠ��Y��zt�u��
���l� ��L�j6X A�n���ff�BL>.é��V���b��a��+R'⠽v��8��/��
�x�����tI��&''Kj���y{�M�Cp�p
v:�/��r}mC�nd�ۖ4й�yx�鮌�SMs$��a^P���]շ c�Z�������s�_�52�즙��	g6����Z�4R>уp[�Ѹ�)���������Ղ%aB��,�s�El2ۯ�dU����f���3�<��s�!ߺ����[�i�>Ɯ4謊���Iɬ8Lӡy�O���n8q�}uG&d�)�F���%�����t[�c/�͈�r�q����_�V�ቓ669�}��4FU�T�$�������B��R��X���>���d:'�8P��͉hptWS����ŋ���r�5ś�$p�i���f�HK!������Oǣq���z6�/~�>�fʵ�W�}����E����zblnLc��2�NiI�1-*�ad��0QRq�>�����}:�D���zCF��y.e�����Vvڍ������=v��\:ɞeT�ᅱ����ߏ��_�;&T��Tk�Ea�oA���x��^�-^A���H}��K���~��+ƻ3j_��z�ByY_�.�Z�-.P�\e=�'�!�%�
�b�|ۓK�w�ۿ�[�,����&C�ҩ�	���>� 3C�̲�A��H"M-ǈ���a^���c�#a�Z��o:.3�� ϟ?�ӟ��h/�PПx��~�3���\\�Ϸ��ȑ#�'0������$�d��~��Y �&��C�7�3���,i�VEy��>�&��)o0��_��b����z��\�|��?��G����~r_)����Nr&�
��+\|�'?�gH5��*��xe�#��qQ ,�;���>[]_�ȹ���A 0X�����+?��:��)~����#�MWbW�ZB%��.&�:���t����4)&��Q�گ��J�iT�51 ��C��?��?�Jl�������7�G"��s�L
�hW[X$/[�R��2��9S�������"��b���;&\Kǖ�Ʃ���s|�'T�82U��`з��4Oƨ�e�	+u��u�ҫ4&�K�9g��ӻp��e��P@����/� ��E=��B�$����J�P&
?~�1��u��hmRr�K9�Z�p�+7fh�V�w(�����\��㕹���s�~�,�_�v�G}���~��d������!8��Iȕ�C�*���T-dU(M�L�ذF�?�+��F\�̖M9s�X</#�81X��kxOwe���m%�ok<��p�_�~���ݨ2�(^��.c� �;���/��*�
�C����Ѵ&�祗$ފM�-056!%�[��S�I���U�M�μu��lI�.�H�[>�>Y�90�����0m�3Q�����1�4�#�ј����~+ߍ�z,�J���s�KIe�),L;�u�1�ލ�뒣U��c�BT�
���� �-�P��C�b�qD�R饅��k�6|1��JH
�D��Y�	�����Ϟ=�&~īR����U��|��3OP��X�͓�V��g�z�6��}���t^Oh�u�T���.���:	���3��Q��8yVWםbd��o�;���R�%,�d��i�j��Ιe�y����G�yls,1�J}ň�JÇ�xh
����&U(��蜏�t�����_|�9��>�i6��!xG��|�k݋��ŏ?ۀ��8�?ѪB�x�p� �v%f��gm�	iu<���X��&�� ���(�1�P�T#�"�4a��(ξr��&s�M�ǳ��+�q������%v��h�E�|�/�p��nP��.n=��!�UɣcM6yh�X�DKA1-�-�N�x_Y/�E��t�㘰.آZ嗿��T�Ѓ��"��d>�&�h�}
��f']��⊌%����"�i����^�+�#F�ʚ��ǎ��0����2h������4�Ҩ������=ћ�L[�J;r�*�q��Pa��>�}pvWR(#��T#�f����4�_#P�Z�����+"��]�Q�C�)LՑ�:�-��<|S40�Q��6�i7� ��0��P�:�d(�^WB�ڑb���4-�]���m�ZH0����Ν�+���Z��j���z�R2�j�ݏ���Q�1ќ��ހ��a �L�m�`�!-ڽ]�ۨ���[ڇ��`]QbL!z�0���d8Y����n�B��yL}���U�fk��Pf���\�9���w�ݫחV�6������Ĉ,�����(���}8�B�es�m�hγl �%P�"c��5�4y6��Q3Z~�vgtt�*U�	�a����#�Y�S�{P��_�����J8� �pc�/^�7��k�w[��R��LT:��r���-7���X�8H�o,��$��d��8K��[��7����w%!���,�\�����n��F=����;�N:���gB��&e�&&ƞ|�p]�6�4��Bm��Y�.f�+@C�V�!qX�aE�a?�� �Dm��d��DJ��cMLWNϬ)�h�QE�_HÄ/\��.�ʏ��������{����x�ݑZ ��1R�#"����7�_5�h���Ǧ:Rńy%�t�l1K0c��JAd�NT
�����\}��^�����tBB�AS�a���&���[�N�JkR/*�vK՞�)�?N4^6AJGj�z�?�pE��r�%��_YY���lm���1խ6�	��
�	̆;�-��&|� 
�^g
	󼹱u���wn�ּ�Ԙwv[p�9z��	��4��`��!�3f��KҊ ���wqN�д0̈�;� zN�M�����Q�w��}��jd���fcD9��eVd�߾}��?��{��W+��>^��6����+ǽ�W�ǂR@�X?^�������+���j$ȅ �g�F������䱓R;66�����w�Y��p��կ��(�5y���&�ml���h��;���Z ��TSA� �����fU�gɽ�!�P��آIgCK���~Ha���(�T(����$�0�y��v<�����$������?�<)W��'%^��?h:�S2q�TF+~�c.O�:z����Iz�ԓ���6�O,&娞@�(=&0�f$�����o�[��_<��o�����􃾘�,���ږ���P�~�n^Ms$�r��:6�)��LC��&7Jb�O7����OSh0����ͭ��?�/���չ��I�cO=��d��斅nL;c�f�Y)+�ys����h3�,��f�ۏ��Z)�ps	c9cs++����2�AUØ�T���6������������ܼy���w���F�Β:���%ucJ���/�n���?�O�|�g�'x�r�'����-�~�6�aكGQ��R,��A��|�:�� ^&j߾���	��brb�ᚷ�z������O��bu�5�9P�L?����W.�?��!�q��AU�8+�sX�¼��a���_���=�i����h�j�������C%�f���'���-?�l�_�����
�^��s%�R�=ݠ44�"^��^��C�����!{M��P���k�r��$�q������J�ܜh�����! �pl\����2h�۝;�5�_��gֶ�٢��B�>��|n��.ON���tV��Nq%��7T�l�8|���K�R�Q�T�����Ѣ��F�ԓ`���ˈW�cc��k�n`/|��p�&�g��U�R�{���Zŧ̓�[�?�'&�5���\��_�௿�;�:|�\�ϴ�P{�mU&��8�3�|����!^d�)��`<[[;���G�t�lN�3��������kY)���C�%C� U����zW�k���q�V$��/�+���X �R�Hm����T����K�xOo���7��lo^�t�W�:�JX����Fk���f�څW�6�Y:��?�w�3��F��`�����s=ڄFwZ�+kky L�-�� ?�mV�7`M_����x%�p&�'�p՞Q������M�C9sa�����_�K�A�_C���/<���GJ���I26ZgA�<�4���hE�nO�ӳ�c{�jQ!+(_��ː�Ń�qP$�����j���7:�8��a(�7n���_B�_�$Z�6ʲ�Aγk��SS<������f�N�NV5���v ��w����Q�f.E��Ѻ�C�Y`T���U��cS���z����VY�ojl�⥯WWWǧ&����O�}����c�/^T*�+�Ĳ��ۿ��!�8����¾�m�[i��&%�����g��	��С%��D�Z��l��l� r(�� �����/�~�i���՞l���7�&g��� �d+d�u�ծİ��Y��vwC�9[R�
D"ݑ�R�*�/n�F�Q.�U���MLu}�1�ov���SO?y��5<q�1���|o��"lh/�l���R�[���H�ASoby#ͼ���u�$r��n_�@Bn�lgg��,�W���06��)~����$D0�����6���$;]	t��A}�>�0W�G���������۷�o�d	P:93����k �sC��嫺v�ܾ���;vd߾Y(I�i��&��c�cb�����d�R��@9$���Z:��n3Y���d�8_� �sn�V?u��[o��E��^�ȱ�l����(�L�\�v��Y���P��n7����	��-�)���;�Jp8C@4 Ib� �O��S�+8��c�z、�
���>ai�@��a)���4�L�&�����}��	+��HھI&����ɱ���i��,��G�J�[E��9>1�fJZ��V�6lQܡ܈�c��/����ڞ���~�������b�E�ק��O�<%�,�v�׆����5i��w��]x����as�:�S�{�n/���KY������[�*!�^+��Iq�U+ؿX�Jct|k�]*����jzC���w��<��O���$�&�!�a8��8>��q�=�0���ۥ�ښ8���1)��a*��B�ݓ�r��Ԟ�8O`���/����y�����m���}��ʕ��x�ӡ�t�`�F�^"��H�:�:Ct��Z�bN�Ԫ�m�&�C���oTэ؞B,�H��ǗњV��,���Ґ!s7.V��h2ϭV��1v?��
]��u���w�nK9d����
����q�K�da��Vͮ5j�&p'h��VL��`�>(��
W��eK��=�,� ���Nm���M�|���d��0���}��Ɋ{ʣ�
[=m��,�0���pO���R^y�F�\G�h�ѿu�K��cT��>��$��a$�3�̞ƹRW��q�[�_���E���_2���Uo�g:�����c�J������]P2��
,��P��j�V"�,��!$糸Ͻ�n(�!1�8�χs?S���0m����T�hx&6����=�ٱ���b��-VbZ�ei��$��ab$9ED�ዿ�կ.]�����խ]��;���lD�'[��<g~ 9�~�߽>33�G���ܲƌ:��IjJ\@`Bli˙�̭J�	&N}KF&��r��}�Bƈ�C���-��p2�F��T)��Y"t�g��O>�a���B��$���SO=E�,n�������,�������/��R��`�xLON@/��4?���cgN��E�v"��3��Է��Y����Tjb�X$>���C�}<Ma���FR�P�m8�D(x
'���&!�jI��v��<Y��0�h[߿�P&)HDϰ��ԕ�p�g����kN&ɉ��������w�ɜ>qZ<"��q�Z%�_����u����o�MM�Ʉ1AժpN�I���t>mjk���� S��Qќ*�/�/�S�`�=ՎQ8�Z~����GL�0�t}�3������`9���b�ا��t(���ĝ�-22�{���cGO�|lw�_����!<(Y��I��FqGqd�Q�;0QT�DXHg��~�i�	�q�(�$N&���?�sX��p�P+)�A�G��j��]2�r�O����;=,��B9 ����=O�60懪X������6~h�VT��.����������(��2�b��m�g���onH5}6vg���H�v	3�D���|���n�S��т������;|��!��^s3a?��C�+��ˀol'�<2���X��<y��{��mh~�$��d΢����,.5�O<��k�-d��`W�G4��}��**���G�_��� "�����O����@a���3���AH 8����e2�i-�M���)E�����Û�[C��mPe���0� @*�� ��P�N�(������KKK�o���PK%��ϋ������潪��.�iFs܁b,���;���rA[J����xz��\bK��K�h�kW�����}%��TCN��N�>��*3Vmзd ����܄���ݼ���t��<w{C05R����P��kK����O�ڨ�x8���O�ĜgM���s*�B�X�Y�L)���Ohk�d;��#k����СC�(��"�֤ �?ԯWC��A�ey��o��З_~��|��gy�ҥO>���0��z>����P�a;�F6a!�k�e�y�����J�������r���(0w�o�yH1ɺc�)�a���I�B�8��'ʩT����0��Ը��8�ؐ�t�"-my�:�ˮ]���tXx�g�~�i��$'L�Hk�jE�b�mQ\�Nh6�z�β��__�Zή�� 읅#��i'��JN�o�Ce��:�ųD��Єd"d���cae�m�F,IWϲj��/.,,���-ςM�ן[���@����G��~�s疜�bz�����gN��}sd�w�7R�H���YbG�������1��+ɘ���a#�(�Ւ��n�̳J)��,����/�%�^�Q%S����[i�W��k�uujw2�[��.���D����ž��E(��,�@V�0�N#�%2E��e)���� �����2fR��	�;3�|��g�P���Q�LA,�W����3Ȁ�rzNMM���ǥL#������1{�V��6ۑ2 �F�Z�" �M��g��Z�myx���P�Á֜V��<2
�;?3'��ļ���Йu�0�OZ &�~���a�нPl8��Lb�I⌈��Ԓ�6��X	�I��LC�%��A��8J<Srv�^!�}h�Ai���H���G9i
I��:8+bW�y����.�B�0��~��M��'���G��������ԸAh�sKj�X�:wC��#*�2>�]� E!�-�Xf��:�=�"�M���s�)x��l/Z�x��g�{n�Z�`1j�����s�0���h��?C:��h�CMMHL��Ɔg��< �bC=�]�Q�<��E���)��)A`��'��(��eŁ�8����R/$,w�`�_��22�ھ
��pV�KL�+��k^3�B�6G�d���.oB�"��i�y������h���\*�{�Ɖ�_@�>�K�B���~.�����ME�G:���S��	:IU�D�!S��A�/Q���z�a�pB�7i���^̃��;�:��������K��l�'�@�r��|�J�ȯ˄�z@��)9d;�a���YJC���>��C� �h�w2�?/.��������S�S/1��x�b+`g���x�j$�?�&>N}z&�S��(��.������R��Z�w��>��8\qe)�>�]����`���@�ĉ�LO>B%d�p�^���$���=4��ob\����;w������2<.\NEl<s��z��%'"d��!�L�0����?W�|��@I�꩐�ŋS?���Hŕ�x���/	!�%��{\�vE�Ȭ��/]���+�4F�<����Z�*��������j��7��y|R\�+W�a`�rn���g����]p_~��8'A6*�M�|�Z����Κ4ۂ��R��G�Myw.��A|]XBs�pQ���
�{w�?�F�0c��U��c�SʵZ��z�B1���l�H�zlr��x�v��K$�iq.�28w���웝;��s�~��#���x`��̸���%{j�z�޽�q܏�P�~�;k9� �1,]��X�%c
�Wp�A�)G;�9c�Χ�d�d>�MZ�L���y�ssS�iU`�_�����r𼦖�s���{���@?�������w��8c���xV,�>�g_<��A�i'���\��D]=����d����]�r�Ν���w�0����Ԟm���2cx��'�L�n�s�����m�|�V��n&i� 
a���a��ח =��/Q�T+b��꫍B����ѥ�$�	U���[�%*YJ~���#E�u�/I�ԏaR��<������ �c��X=����&�a���?Ɛ�xa�v��d�8�e��_���o(��t�*e΍���������P���y��i�����K/�	?v��r�	���6����b��*���by��x��G��P������7� ��$���,h+���1w|C&	�͠oHZ.�uv�7P��E�S\y�,��Xkã��OZu�uc2���-Sz�*.T*4<�\N�U�J)n�k�Ν��N[����ٳ����*�P�5+��!}�=@��5���F�LX��n݂}���_�����ǐ.^���ё����Y�Y��"�3�@��<��1��Z����2<���3�$y�$������	N�{��椙�î����=�x+t,��w�^���a���~6L�V�bqq�����N��G}��LQ��4����Op�a�\�p���Y���n��i��{˘��Z����LϜ:2+[�g`��Ԣ�o��Op��\�V�U0Z����R{�w 򥯁 �X���ߴ:
�	���O?�c���|�;єN_}���x숺�}�y�����kHbҖ��\������eM��g��<F��E3��ijۭ�v������W�Z��A��4cI|.�TX�h4 7����HK�O�A<l�7+�Z�6��yRk�$[_ۘ��o^x�C�����>+j�$VCWCW�Jba� 4�@L$|v~���4[]QӾ�,�bj��Q�1��-��m$��Pe��D;K�ei|O�"Q�µ��(�H��es'FO�>Z���>�,^���mH�v�(+,�>���{�a����mz2�S�j�-�-�b�΂����"�i�CA
-� %ĳ|^<�K�l�]��Ai}����p��pr����?^J��W�ƷpXh�sL�� ���b���ue��^�˞��=���&.-��;~��\{v}c��\+3.Yo@r0�A��8q��L��L<����t�/�]�t�K��"7Ef���Bɚ)T��`��y�	v(#eXh�ӧO�L�i�o�#�;q�v�#�$MҀV�>^5������ ��ţM\�Z��T���J�@�gҞ^�9�(��0��^'��X��Չ�y��t�U�J�'�2I�2!���.�
� F�e��� ���
ih���!����xڒ�3������dsu�l%�Zx��F��V"��m���H��cK�Ë�����T���*Q��V]��J���~����bD?�]z�U��2K׀�@�D̒�uǭ�.�d��H������8I����w�9�H���Mf1��క�3o���T�0ImA��;��,=���f�|����=���_]���U؋�_��?Ř�{�o����-n��
��?�̷�FcU�v��qVi�p�J��L<%V�T��8��&�G���A�����u�aVh�Y�I� �gJ�U�n��hcl��i�,o��_"<�kث�wѷU 9��Fw��!iǣ��<hp���?C�2��_�+ч>����p�c���*>lv�uB�}C9������<�<�\������I�M��X�"2r�H��n�U�(*Փ�~;MI1� �����*)p��	Pq�@�:�[c3~N���϶��Y%-�0����ck���}��g0tɬ��s:��4����P��dN:R}Cc��t F��qŕ�j+O$��)D��5�|�{rh��Qc�툧��U���d�3a�B-�H�x�Δ7������\�6��, ���LO�}e��~�����:�yrz"���8?���F���>�L����a�Vz��� ��V�wQ?3�s���[N>�Ė�3�`��. ��mR���6t���T��Ј��:Y��G�Q��K����]�@��F�o����s��~�
�̙��%�짟~jb��?��Y�j��}��S-�Q�`������������u�Ϥ��3���rd��pay�Y��� S��f���4�WVV�mI�Hn>LX�jY�J�������C����Qҥw�"NcG�X��A�z�b�4D8v��v횓[�G4��Ȼ���n�~b�d�Tj�����D�0���{⽌4ǜ~�����=�>'H��"C3�pjR6����Y7����ak�G��������Z����] #/�����Hʶ�bb;`Je�˥�^_�/�[�$;ȴ�N��`���ؐ���
��DO,R��^G��;�KE�໰8 ����64���ӝ���.A������Y��v1`}��˗7��昱�0"�Å�ݻG����zFln��CzT\�1.4�)\�=By(	��&=1�@/%�Y�i�b�TUf"w�7HL�]�s��y�|�<>�l��G�{v��Y��ۢv�A;~�R&�D���7��2<ҞD61O�b����I
-|'�]���:;��af#t�`�JIL4�]O�.rԤ��C�P����DXw�6
`4P6��h�M�9�en�W⿬`��T��1�裏>�䳏?�xc}+��H����8V��у�2�3ш�Ci`u��	Z7GB<�A��zF�ϳ�>K���������}��2���]�Q��e����u�R����Ƨ~�f�`𽸠��lVƷ�Jc!���S�Nq�9���9�&� +��qkk��a�&�s<Ǎv*`U������J���.�lɚ86I�#��V�x�"N(%hcf��!�� �'䁮m���˿$�E���uN�6yCw�:s�W�+t$Č�|C����gS*h��٤�"��5h��%093�
�px	VE9������ѣb�KrP�Ş)Kr�S4��J�2��\�
�/S�`e�|N?S�Vj�v\D��ga|ejBA�t�i�Ɍ���;d��C�W3d�PK���Hb;8SB:�ѱ��g)���hE���􃕕���O
�R�%梨�?e���"f|��Up�8>�?~��T��v��"1�.��Z<"F9��&DB�r[�Wx�P?p�3%O��Z��Bb(���u���Q9#�'�xH�੧���Z���._��0� �� ���`�������9��c.���)@���r.�z�q�)����e�;��)Q��DI�lrM%�Ut�x���N��몔\D���H�؅�Cε-�"��Ѻf������-�!nH	X#'�{O1h�,h�&��F�b����i\ilKk��a��[o���縠,�(FN]0,tY�_3�s�`x������/� X�yC�'|�]F���X�*�Q�Rv
�~��������������Ë�^DN�� �����Jiol$�^�6���kQQK&��<���$���w��uK,0�H�H���g�����u:)�>]n�l97��B�Z�A�
����2���aנ���{��+�
Gmh�p����23(��e���ɸal�;D��ku��>�E���am���$��,��?O--6gP�A+2��iw��2��(�Əv�p��w$�9L]��R�97։Yf��j;3��쀺}KWJ�P`��aWՋ�H���_�F�g�Q�L���G?��3GQ�GP���W�^{o뜔Ǆ���+���6g��a���+P`���a�%�l%.���T��t����~j5�E���7K��tɗ�c���_��Ϟ."ZB-j4%�-�
� H�?�O��.��Q���r��$��o���v���8|����Vk{nNؚ��+�7�������b�C��s��'�e�P�!6p���(
Y���=��{�^p���I��=���垩/�����yT�����)VV�n�ı��iަ�
{��+�cNJ��Zo��O1��{�j#R�y��0�T�<t��#��Ev\eT۵+X�}�ա�������Z3;�]h�R���Z��4(#)�S3ӥJ9�م��b���A<�ޯ{����Q���R��N�(���C�&eS*N}�7�(����줰})�?oH� Wĥ%�9��/�}��?y%��Dy��?�6���qI]������2ڂ΂��I���	�"���d�X^Af��[֓�7l��ҏ�V��q[̒�#��[D��rn�ὅoB��)e�&�Ҍ��>�������,�s��c���5����ϳ�S�O����8�E�x�X}�����#ﭯ��Rye��:z>�|�[������?���V�������󢛭]�8�{�n�t�>�ę3g^z�SOH��Z��ɲ/�fкÔ�#yq
2�%���$��R1~�xML��� �
W+*�JO�q�����M*�SHTʥ@�q��⼑q���Q�V��v�c�#o�J��R47#��.]"�gnߔ㓆=���v��J�,u��gR��<�$�#h�8�l�
O<�$&���?���2��ʰϨ������lC 2�pb�jD�M�3tU_hj�8�#���5^���jvd�V��խ5�`��G�-���K7Ե���)�ru�f�Vq0׌n�|S39-�W�e��l�I��t��^C��tڙx����N��mv�6���p�����m����X�-�w�,����~���k��6�(v_`�l)C[f9��V�U�F��"y���񳐙b�s���/}�W�\���} �{ڴ����{8�!E���&�J��E�	.��?�C����6�/��b��K}{i"���8[[[��E��HC3���}gfGG�%K����ע9�D}�cǎmlo�]��\��
7Q�xem�7G�����*��C�D����3�E%8p VY��_�Zm��1�gl��݄��Y7+������(��D��+Π��%��T�_�"�G�ܭo[�p���b��W.}a����j��VY]�������=��s�����k ��i����M�oG��XB�4�~lb������o�=+ �))�Ƥ�h�믿�;
:�&c�oo}Bz)�Fq蹸&�nk'�JR�����$��4�s�aD���g�A�ʁ��#X�ν��C�R���,��Y�H{���[���j����>|pffJ���(C�����L^�z��٨� ��̨ �b�E�{�3u`b�ь���,��I�\��~8]4B��r��Ӟ6�M��g�߸q�W�Տ{�D�!�� ��a�~�n��"��m<��`�����	�O�KwBh����������O��OZ�6�E�6քPeJ�#�j�1�Q���4����/��9ș"jp�h9����w`{�d&�\)-:�C�r��Pc�{�B����Jl���}����i5��;��rq�`�;-�k�T��$Y�0���P�	��;�����BN*ڒ#�хZ��i�)�&ȹ���`���NU�!	�c�nr�d�nf���44��9l����-��h�c/�q���Un�i���FX2	*����C�R�fqqQ:�_��F�x���,�i��_HD�JU����7w��!��Ҕ�K�a̅+�1�xv@*4��S:���L�3^OpiC�a­=��S؁���B�pOȹ\�l``��=+e�,; aH;��3�Νe���wV�#>Q:Ԏ
�օ�H�F7�qMR�@�JZV77?;539�L!}� sh��ل	�����]�tcW������A�,�,)T��|ý�Y0c�,N��Ǐ���+�y"�ܝ�xC�ۡ�F&�Wt.:�<�7�mV�W����4�"�u��c�?޴߅��p����ۊ`j9B���>B�m�1����"R3$㞘@�Ɩ� Q(��U{>���Vs�����ݻv����*W?���cΰ*��fJ�Uf��շ_~%�	��t�U���w>�]i�>>��S07Lݹ lj`�}��]��ug�f6;h������n^�	�YZh��J�hW��W� fxGqba���������
˦�'��ƃ�L�덛2���ӄ ��:K�;�}�[�������;a]J�ꂾ<Km�\f��"u���a�P=��첻@V���~�8e�z+��7�2��-�{L��ѨȞPI1����RM����o��|�=R�lf�{���a W��Lq{^�{���f$
 ΃#�<W�.�D�Hu�T�TPq�ك�9ࡧ�S�i�[M�}���@�
0�B�ţ�`���QJ^��l+w�6i�XޥD���3��Z�y�<{������@(�6mk�p'J~M}��������<񋡴�JLq��$�uv���=7/~E*T���T��>.{�Z'��
����1!�9�(�!!�^��juV�E�b:1�J[���l�1��"���	�'q6L[�"��/�\फ���4��ag�Q�P�BD=��ٝ��$���,��@��VmH�O�a8��F�e��aس�9�J%�
L��0�V� ��`5\h�Ji}bw9s���
��nB�66	ƈ��Bjm��s��ab���;�>�F�79Qz�&GFB���ċk�f\L5��*y�g_��C��:�櫏��F�ȗ���}�B��aOPi�_
�d�6f��&��%�8	�ۣJa�T*��DN����x�������]��V�Q�0���fQ��T�YK2M~"Xk�����y�����򹷼�>y��O<��o���ӣ�c2H]��ve�`�CA=+	���m�)wz���pqU���=\��$h�8�7�ؑj�P}��h�%�;K�<��#aYa�|��q�F�"��Fn�%��#G�}�]%Q�nm��6����/���sg�>r�XY�Vw*Fu�����������ꫯh��;�O�9���_��7��Ay����f���͜V�gre
r�9H�
O١���yk-��r���}+�����	������ƹs�.]���Obᮓfl\ډ�:m�nk�`
+� ��Q�Zb#���n�Hc��n�k	S��fk'�zR�b�Z�yzL���@��Xom�\���}��A��h:�\)f˸���$�\ ."�&�۔{yv=�>�쳐m���tl���|�˚�*3�1��N��Ǐ㞘y����& �1�
'��
T����s��������?�#"�bs"b�(�F+�	�氮�٬�Y[��uW.^�XBl`�R%��xb[�k�R��{�%g�⡐^�����t!^��&f�y�,��3D���Ļ0�C��Z��##�+5=��G(ǁg4W�sֹ��D��]Ԋ�t�y*ѝ`*H}��Qv��"hx�2�V�U�#R�+e�S[ ��KJ_�����NJ��%t)����/��/�Y?8����m�т�^�y��r��a���eV`Pa��r�2f�ع�z<�i�`S�6g��Z�Jɧ�l/N���-����"��e��A��4L���@�*���$;~T����}���Ю��L5�����%Z%���LĒ��
��Ӵ"a lK�Z,e�9��
m钆���K��r���ڎ$2��ӟ�tgG���R
|�A�׍��,�`��^O<[�QVW7�������O��U6{*�¨��J�A����zIl�<'�1;Zy�Vw
O+�L�τ�wx7O��m��("��"j�#�Z<+�{�xU1c��X�LiX�8���OD��ц�m�c������x�	��B������o�{޻���i
��@,�s�B���7�ff�z�ĉd�*�$]]]�[�h:ޜLJC��ӊp���*�,XEy�Nc	 �/���}U%_6��Ӈi+IH��h�a�	��L�:�Ծ	FT�5�{$��nc$��]ե�O��KR�P��܆�9��5�d��еa0#�_�]_�s	�����j���O'9�0]j���b�ζ��gA\�r������!6Ԋ����~��_�c����PK����S�؛Ĳ�WVV�F���[l�4����7��^�b�<[x�ٜ+e���=�d' ��=L�gߡ`�L��ê-..rA����f/��]@���B.`��8 ��A�P��y:}�0Pѷ5��������u=�މ�Sb������^����"'564*<(Ff��A��.���u����'��R:,--���BNtg���4e��'_�
9��c{�B4툇5�@}.�7�q9�*DJ	_D�/��U��sM�[B�w���g�yv��~�V~�j^w��������*tlL�G�WX �O<1�~�Z@��4��E�y�B#���|:�?iM��2u�'r����%dMu �������S��p�b����E#���
U�n]�B��<�=�y������8l��zs��lL����h�C�Kx0��l�2�a�
!+���R}�l>Hb�y��Nɂ�?b@�����qv��^��b.�֋��O�m��?k a�ψ�/y~x�ʵ}��ibjj�Ν���Me��m����v:�vsl����(n�������l�S���$�*h����d�������
�@�@�o���C�i+ʨ��P�yD��;{i��/�!!Xlm��V�[;��ְ����xrBț3?+�ou���ёQ�S�P1���[y�>5�l�� Є��D���(J���O��H�n��� '�K��X1�`�z�J�@�$f��Vr��t!\
t���?C	��4����>v��̨��3xh�Pd��E%2gQ3�ڦy���~��$�嗝X�Nk}q3������Fc�\Q&����<h�1<G���ċAk�.Q��4�~e��H-�Hf����j�L��|��O��M�^.<JC^���A*RÊ��Q.gCKM�����Fc�0og¶Z��Z����bE)�wc�DG�"�4'67@=S�>)��NC3�;�A���$'P�Y^����Gz2Iw��s	� 3O>}�^8{�쩓g�F�TQM�&���͛��nܼs���u�,j': �Kn��@�v�#P�q���RO"H!�����PȩT�H�bw��ŋ0�2����"$��f��s֝;N��"lzL��V�����a����7ۭ�/������Y�#+���0�V�yz�a�ӏ����=M2L$��%Q�;��F.���A7nܠ�6�f�B*�k?�A��Y�X���0N{݁t�b���X0Cՙ��|A�e����Z����n�z���>~E���)�R�:pb�C(�ߎ����ת�����݉��n���ay�ı���$%ڢ��T
��J/�G^),eiw{KzG\�r�ܹso������e�����?>6ʭZ�	=���Á���R},Y�2Vwg[0��J9��y��00�O��0�vn�VV���/GG��d�j��	�$�6z!q%���#aTa��U�qZX���s�|�ٗ��w%�����8�G!q�Ml�/��ի׏;1�h���W��x��_��&PD��{����k�p�^�4��31>���ϯ��^�x�Vk`��u�a��JW�Lr��S�g���t�H��nm�r��`بU�,�ɇ��@�D��b�2zVQ��A-0�K��Q#6w�����o�va��̸xZ�9����ʙ��<��t�dj�����?4�l�^<���'������dݥ��&w�#�[{�ArX�yo��b�ؔ���;�v�y�&���@e,]����ƽ~��G5��vz&Nj�rk{{r|<�����*k��iw�"5��-Z'��O��x��#��������n�-�������j����:��܍y�.je(�#�^<zR�3H��k��.`.D��j{`��s��i�/P=,�d�G�#A��hÛ�����9虃���r5R�&D��,X)�ә��m
�"�������o��ǵ��E*�J��`���Om���ù.��+q=�:�7a�L����
������A�ڹ�%}'��bl��:u���Mh��/IϓM�Z���3\y��n�J��;`,�^��Q'b���?�R�bIy�=����'���b�bor�奰��)�Y��cd�+�'0ZvU	� ���u�cI�/��RK��P����6��!m\���J�f��nt�%�[Rj��:����U�+kljz�91&}i�-���$�Ƨ&���Z5cY��qWmH�o���R��3���jY�?�1u p�R019y�ĉ�9���i?x� �
�S�����������TĖ���b:��}\�|yjfvbbr~�<YA�̅��}Gz�m���"15��P9�p��^i�;a���˴�Fr��r�12Zot��D�|#V{`�����(!H�$����n_�q��
��ڕ�k�҄�U$R�z�&zbk�=�1Y��]�i�l��'O25U�S��0ͳ��%vp�u+Qe���QGȠ8��PP�fȡ�Gcr�+%�W������0`�A��v����S��H�%���^��Vg������}�չׯ{yܼ������|t
�!Ηb?�ܮ�+Nc[��)'Q9�mm3����-���72�XXX��zP?�l��F׳{��,�B4O��ɉCG�on�Y����7�˖�U��� r�'�6{�Z�̋�ﴗ��ݻ-���{�O�>"ٸ��zm�����1�v�n������������+�v�N���jb�C�j}�wpw�~�akW��<m��s�4f&�4H�P����i~��#;��qC5�ӟ-�]�W�RTK�,Y#^:f���V֠nݽ# _����Vk���\�Dn;YǁK�,�7Bѕ�zH���j[1�q�h{���g�>��;�_ֆWf6�}J��.[�ì�Xb�5�j�L������>	�aؓ~x{*s<y�B(�^��5�#&}�7po��c9i��q�C�00��R4{{�o�٠!QhTXn8,���s��X^�b��Sy �����'`��1`��G'��7��vI�����<�U8��4���ay��.�K����ٺu��իӇ�k`�t{}�u�Mv���`�U���m(z��M��c�ǹ'<d��1 ��٣�/�{�?��?�aI��E7�H���'f�P��p�9��jV�c�2�W� ��5�$�*UJ��ИB(�VO�8�n�R�<CKI����L�c%�g�sH���!�.�6�(�F9$\999�a�&+��m�F��*�.1�عuV��x˲p��*��`��ͦb2ĻL��%j�N��A6��*�擋SZ��C�<�y 3��."T1�t��ΐܽ�[���0�$n+`�!�m9��Ә��p}1!#��xy�˷<#<�hLӔ���I�ml�4鷇##u�6q��$�zO&�i��Ve�B��dp�h!�'�C�����8�)�|&�(�CK}�YeА�_)�<�̕�	���zs�/\A�dCdÜ˒�e
h�ay�>��k����s���ec��VQ�����g�}�����V���y�>�"�O�����e`��	>Ml!$Cu�ދ�)"�ٛF�!r�95!+]`�Ӫ��'�ĺT��������L�_|������ï�~�6kT	�7�|�g�b�7hf�{���5���.���ls��;�0����cXRp�n��2$
�mUn��v�b0��2u��g�}�QO���Ӑe�'���0��7M����&��ѣG�s�ν���-o,..�H�[����U-ȯ�Ǐ*]\G�`�Z���W_���G|���6<3:Zmu���(Q����$ZJ��6AJ������ժ�EC��j��̨��UI��O?Wv�tZ���*;{�,7���Đ��M��CaP/�3g��ٟ��3O>����:��ԩ��[�u�g03,|cT�3��\�t	�4�ML�;wI����ge������Ly�X��R����v���lm�2R��i��1D����\�`���[�!1*U �F��S �͆�����	�L-]^�2-�čF�Q��!rw0/z0�!r��1Τ�bH�#`��N�:������q�/eo�d�u����9U�Cee��*L�AR�ZpK�(7Ö���=*Bᇖ���zQ��r�TP
Q"[�6	� U(��y����f޼ә�����T �3�dV�瞳��k�ַ�ø�_�k�oƸ����Q%�b�~�M]���6���F$W�$T�ꥰ-؎w&�-����F�[�鮞�dhz�Vq�ȭ�805#���SD��Sp8�o���ך?��/^�Dt��(c�������r�>$U���|�QA��}|zM?�V��2���"D��G���d�ӂ�Q�s��Y�y��߉N�8�Qx/�����ſ���{���/���"Ӧ�$�։w�>>/Ɵ��9����>�v0���ݦ��(���Ǆ'�|bn[�T�r(߾}����p�%ŭ[��/?~<��;����r�����v`X��Z���_�k+����o��֛o�I�;�c�.\�p����q�#%��:0d�l�@���P��p�7�Ϣ4�2��7�����N$2K�η���~��>N��[���}QwU���S>5<B ��O-�� n�3*��@�c��Z���.�A�Cgf<��"�-c'��ÇGX졫F��Ѭ�ˉ������m�2�݉`ֆ|#�|es���ԥ�傃��;�oj��ϑŃ�Rm:�Bϓw��u�rb�������x���8�&�����~�� xJ�\M-� ϣ��4O����l~ W��p���M�GC9�g(�G�XZ£��[h|:s��,��ŕ��Rd�ZͥD��OQ�s�xZ�F��t�%x`�z#�øN �Z	�ๅt��;��K��7!��~�=F�k`��ٕ�Y�"w��6>-;�[_�UK2�Kڈ%�� ��5��:K����֨2?%�?��Hn�^�[ΚoE���-�;����P1,<���H�U�q���~m�S5�gg��D���u�@��Y���RM��r����~!�k���.Ѐ��/�텙��(�Ao6��t=Y!��΀��%�S����5�j�~\�/��D��ZYJ�z\yu}M<RaQ�f����91F����L/٪�ؠ��#��!*sss33s��N����iC�,'�E�UFku�QDE�f4㲄`��8��M*\m���� h�&;�5HX���h�1��HeS��ʁ8��z~�a9E���
��<'�26�Oq��T��_��(o�T·���hԮXs�x���4�Ɇ_\=�-t4�BU�.�����뤄f=�3����/��lZ��ԭ�[&��b��R����P�vʕs�
�D�
ۀ_�����77;����//?[�O��zV�eE���V���٧�d�oߺ3=�gb|R�2/7�'��xϤ2�ژ�6�8�󔸸��/�l�P���-�]=0vw�J^�qW��[̌���b�a"�=~�r��)B;=���,"��>�d��my�6��:1�1h�\��nx�okM�8RHx�3.,i��L�X7�O�Y�E֡"���ɉI6�Ҟ�hJ�ەZG��}���BDoB�P��B��{	,x�ϮJGڐ�[(���#Zp�?�КK!K��ݎ�]X�'@��i'���\�D�:�Pj=3W�&qtywM{Ef@�2-��pɖ��������\R��+n�$��5OcWb�n�"a{	<3��d��Q�YTz��K�R ���������:m�1��1sE�D�.�Q.a�tjq�lUl�Lu�LWU,1-�]X*�$�(�e�BN앯�-[핕U���
n�Գ���:'��l���lK7�z�2֜31�}ȼ8�Х~�X�}���ϝy���S0urp�`���v��p�����K+�{E�4���㓓�M��S��HT6�Xt(;���$?���|1��l���zO�$zKLmG�_��jW}Or��(��gb=�)�Dx̯������߽���?��?�r�&�+��E�j����~�����F,�?|�h�[��Ԥ/#Pso�����ޑ�{��iG�\X��Pu��$]K,�K�2Ҭ��6��W�
?W��|��\B'_@rXW�a�S}����� �����#���c��T�C����[�
En%�D�[�&b{�PH��LL�K��Fa\a�Ɠ�'�}�?��QY�F�_i��G��Ǳ���r��#bl��F�$;5ln�Kӡ%����Mavóme��*H��z%�Y�z=n�wZ[� W�q�9r�S�k�����4p��\�|��-�������o~�иJ�$��,�B��'N��8D�&�������&��[<���k��/�5�N'!IZ�+���j�%�W���������!.�駟B��={��L�8t�4j�j��3��,���x � ������sIv�"h��θ����޽{����I���{�N��,�?�Ň���� Ͻ�ڬ�٨i�YO0�}c{6ܢW �>� 5�/��XϣG��jK���bH/P���mn�C��HݿW0���oqqqϞ=2�0��[B���m���]��e�Eh�C�Q�BM�D��޾�3gΐv��HX���1����[w5�i�[x�f���pA�V��'����a�%�ۗX���a
8�$V��T: O7)Y�q�͛7/]�* �����;O���s5�)�l���X�E���-X&(�����Ri@Muzg`�y����(�eOLà�f�$B��9Ӿ�2��HV#�+�옙l&	�{.�G��+<��X��Ǐc�]�M������BI�hG����S�5LC�)ʴs¡��e1��-�4�<ல�r��#( �xj�]`�M�7o�~�W��� F���u
���ے��'x牱{��ž�S�VCb�m�w�>�ʫ_��7�Ȉ�u�f���V��������-�MA�3[$D�3�=t,t˷�Z�Vx<��:'$��w�r/շ��8ع�L��"|/g7�7BJ��J����piI��[�zS�<�N����j5��F�5�J�8%	KJ�ZB��7�S=�AW���u���n����ys���V[����I!��m(�Y����.�-����
Yлv�ߒF�j'Zh-��ti�\[�v�ڭ7�M�.�z�#�|N�gZ�"�H�8�Jryp���T��761��U�LHUۭ�����YL��p��˰��61��[�I�+.��ǡ%���QQ2�D��f�g8�+����x�t�P}�
�e�F<џ�k�B6g��wv��=�MgQTc��>�{����Y���3?��4馢?�1Tw!�{I���E�{�.6'R�)������~��0���tq%3\�/N5����",��g�}!�޾�[�g�Wő�{�2����xw͡:��B�+̯q��y�-G�h�8�kձ�	��؂��t��f�����z3��N 8��*���Қ�VJ�6� ��^�G�ǘ1���`T.8��DYi@��<�)�������y��N�I_�p�Ν;dka�K�կ~��_���/�L«��G$����!��Zoq�˺\pjx!E�$=|��(Q��B��hF�8�2y �$3�s��-�gW�=FFe�Y-�v1DO.)|��i���::�cq5z�s����OU�kT�N�<����%�a����b7S��P�灄K�0�vx.U���Ϛ�+�M!�&��l�S5�T�%x�#��_�Jɾ"���eW����/Ͼ�����{{9���N.p�L�� F��"�('�%l�#a�2c���b=[�����v25W/�S(�R��,�-��c��gq�w��3�5��x�\�'RR�}����O��3�<�|d%8�B1�8~�4��C.=,�ΊV�\���Y�I�Y�w���v�잭�e<Vǌ|��Ns�`��~6!��>+œY?�6�?u�������^���"�`Y���Ϣ�1,�ĥ�ȉ��ع��Ĺw�v�T$ـ�A�{%ɕz�v�7��h](���9�E#�����1���������{&y��Ѥv�]qA"%-bƀ��eɞ�m2�ѻ�r�v쵓���[ ��O����3�/$�T7&��hЄJ�
_�ޞ&%+�}^�$���_Y��'��u��b�2?8W�i//\o@�ۥB߿�?�������X]]���+�ik7O�W�LeO�a`%�t�N���4�t��Ȱy,36��Yj'���$�7/ͥ�8�v
���hq��W^�k(D��gz�����4�i���©k�x��h!�[�[_o��ڬ�;���gϞ=x���Ç�"��"�{��ŋ�\�Z�N1!�i��� C��L ����t�Y��w&@��k:�Z�8h(��Q�K +�.~Oq��B��C	
�-�m��6!���'�P�/�;Χ�q���d���Ӱ蜥ۨ��������˿��V���2�	b���L�����QցU�+W��Y�'�4Ï��)�4N�A_�|o/�y���!+���v��-�/W(~Q5cF\���c����$�FS�W���X�cǎ�u�9,��z���<u�����}^�

O��&z3�_��_��̼��+��1�oS~�P�V����1= �Tݝ��$ЕL<��-]tX��CʸE�zʍk4�o����s�p?p^������~��y��n�x���t>|�L�ŗ��1�_�zujz+@���*��#G�����~���X��{��� tap/_�������p"�߾���8p�?���ee�ğ��...h0-,,PgR9p�U\�?*1���c�_�j��ݧ �_^��m�I_z�������oܸ1??���faq�n��:*9��]�*X��#MLnq�0b�zV�&��Lo'��@u�X��G#��Ut�>���p�''Gqp������Uq���_t������z��.�x.O��릿UP qhh������`��:��4�MN������f+Z@�t2�QcW���-��P伻�q)*H1�X,���5�X�`',[��b���[yFj3N�v�*�d"7�i����F����yJrϙY�H�bHz��+_z��Q�2I�,u�Hw0�hb͕��gV���g�X"[��	���=��ЕB�h�'N�XZY�5��w�adx��J���G�ɕ�,蕋��FB���� H�3Ǒ���Al�p)���FF��\�i4��Fv�n���!�ś�F�ס��7OM?M���_}	� �3<:�'����V{@�۷oGq��c�

�T�6ݔ+LCC�ƅM͸͢�ǅJ-y��c h��g߷�#������pG�޷���S����7���~P8Sŏ`Z�5��g"6t��Z�Xd���B��#+˫�N8�=*����T:�ڑ�|^�ňh��r,\�	�u&Y�z��nO@C<VJ�[�M����#����
�����	� M���J�F~I�k�|o9�%Q b7/�^���1W);��)��aͨ�)<\��qnN�P0���.�,u�%N�N���T �n�K���� Ok�{��S�t�)C�<r�M	�������w˨�~*��uFMc�q�L��ҋ�I6���C 8u=%�Bu��"����UK���������1?z�(ܡ��)2��M�y�-�*	����f���N.�m�#SK�md��a���sf�m���2D�%�u�#��3h��
VN	C7��J����:Xmh!~
�ـF:�<!oD"�O<t� ��4�8��Z���U�9��1�|��sp���ڪ{79���e���|�qA(��Ñ	T�I]���Q���ʙ�tb[E�<qE�g�K����,�ޔ8B	��-o�ۗ�g^!�j	�3.N���+�sE�2w�l�J8�3T�Tj�r���G4���[�v��p��{�^�̗�O�]��n2�{&!S���d������S���'S��^�_�*�If熥��+�IT�3XZg���d�v>�[d���H��)��b�e��f��!'Q�[ܻH�M�<yÑ��
���&S��M��F8����,�␛����Y�7̳%VBF� �h�ҼXZ^����/�yA ���J���q>�4�O��Uu1����v��5��qT	|	�������ݲ<=�}�:����Zw��<���U�L2
�������K�iH����2��>Z__q�$�N�R�Ԙ�pg�Y�R�O����j@�*l�'?�'�]<���ɔ����G���H�F��-v��Zf��\��/'w	���"�י&)6V����Bb�G%x���QdiS<�T�2��Y�Gf��q����6��{�e����M�cL_/���.��)��<"�D}�;�E5�ib��٩�t��Ůf4�!��(+b^���]f�2��+���2pc22��OJ�hj<K_F�L*�(d/����d�Lw��� ��e�G�Бo�85�Ü�+�z�aЇp�L_��J֎��$�C�)��䦗��iN�|brltl�ëUFtbkk����=������-�*'7�^��L+���3@ �a���X���W�����^�ׁ����3�eR�kZ�� ����������p�.x-�,X���3D1���y��z���Oͽs���d��sIiu��5� ��C��;y�������`n���Ga�q(\�I��fj!�!Щ;����s��OH�EW<v���cG����ɟ����N��k;991<4��^�?�o���^�{�@�N=\���ɭM3+|bl4��zUx���sR�e̲�����Q-����d�۩�rEK���-�`W�o�M�\|&p��+�祕��N�"��ƺ�+ڳo/�;����e�Qn6���?p��mf%&Ƨv:�.���v{w�<�ػ��\�?b�j2�T����qp>qQ�'��$�S���_�5���+�d��<zH�31�wx�����D�:jX+�w��o�{㵷��X�㧏}����H����ߴ��7:����lm&&d.�=���Ё���2��}���a������<1=�k�����2C`h��4򲴀$��t������?�ɪ����8�0�V�ί������_�ş#�PV�U=??�}���4U&��%�e�p��m���ӱ��5�m�$�� .�p�������R��j�ر#�ӓ�7ѹr���kסE��?~,g��0l(<�FEX ��d��&'�A���������*��2��d�PA<���z�ezr}���6>>�����L�^�~�I�n��76�x饗^}�զ?�����۷���>���h2�O��%�7���K�sI@Zd�h��m�,M/����^01:V�c"��#q1+Z�q"�-扦��JmS�Ox��eD�ؗӧO�-��k|dgg�֨�l�ۅ2�5b����QE�*%6��Y^�&�Y��-����P�F_z܆j̱�m&@B�Z�L3���q���,l�'���ý���@ք�� [���QH�M�\V)F����z�M7�H	��ӏ�kNHv��A�T��k�IKda��\Яp~e��n]z��z�i�W�9�ĬԪ�>�����#���� +I*���D�7�g�p���PN������ {�����o�y�����OB`��LBE������wn�y����G}��g��
0)�8�|`��eW䦜8`����T`�vD�|�(0��]�j�����A$u���b�Q"���������^�X��w�y�d?�m͕�ƚP�������f%���j���<I��������.� ʇ�o��`VO<3q���I�x�&x�x~��2'	yO�T%}�-�A��%�l���⑻�~
��$[c;px�W~�Օ�7o�ƎG�z�Ɔi�ߢ�|ۘO�k��=Z�\���If�Ȣ5�g&2;A�G�yእ"�������7n�����}�@���!����W6�WaH9$����"��q��0y��$���ӳn�Th3@����Y[o�{�$�"����^w�Б�R�#�Ҋ75��wJ��)m���^�rucm��:b
�3|��d���e�K�N,�w�f��C\pv~�E5�����J�~��҇>���B����E�>�skj�	�k׮]<A�7�SO5��)�aF4F��8���[:])�ap�%�$�>H-�;�ַ~���A 5<��#?�����T��>�4��C�O�Z�����u\�1Ԥ��0ܺu?8p��^`�Ky�˖��3{l��b>���*������v�����l���';(<˸�Qjf��,0��6���K[���0�#e8�x=1O�^�ͼХ����C�$��+��4�Q�Y��H �&�	Z�tD4x�I
����R%mow�����w�L7T��G7�,f�'XE{�h \}�.�]6Cl}`jު����m�(���8B��aHr!�.6Um2Nn�M��j� _	|���=w5w?�J��q�r'�)�r����?q�'/��7��.b�᰷T�FH�L�{$�">��L3�@V�f��(�G_B(���H=����JU�����_@)9����R���w�kI���.�U�	q����P��<x����C��޽�xeӸ��k]�"������Ŭ4e)I{.�$���9���8���$���'2��Y.}{	'�?�[��h-ܺ�K����*�,2v�e�8u��R*���a�3K�@O����X�����r|�bI��K�#m�*��+�l�tJ|[#M-T�b����3Y�Y���n��9R����e����U\��Ɓ�	Ss���3��#���E�e"�,�cǎ��a�oAL{��ѽ{�V�l)�:��;د�+ ł�+PS9���δ�\@f=ܺ���^�*��*�U��514r����y�#��HBY�	-�?P��Ċ��-W#}J~���6#:,c]>�B��ٚ�e*!\�<P.$k4�mu��%����6<��k���ns�/.���I�5tp�g�:�����5'.����00-Ɂt�6�������k����T����M{��+�PiR��U��o���BG=*�~�o���<x�����w'w:R��G���L�
Գ.`ݝ�oG��:Rbe�twEh	w���Qβ�vSn���6�)�kN�[��x㍥2wtH�����:��ŗϞ<y����u]�X�-%�>�Y�U���D5*~���o����G?�\�����fp��J\��DsO������\�7�+++�����ҋ�T��)Pc�k�m;���%��-΅�`I�fMa�ډe�V��q�؂.������$炧��x饗��@i�u�j�Y�����xYh1єX��a�mE���a�j�
�n|nj�a��?x$�3"?���d�V>,�$(��ա4x߲}����Z����&�q4|x�H%��ַ�u���}�=q7�_{�)W���?Z�b8�I�Gh��<.��s���f[��V�e�x�"$�y��|�+x)4�k=ƻΞ}����?}�?c��݉8⣰Eul�gk�bC�Ș:<���Ζ�(���?�>�A=��8(ى'�������Eq����ÇϞ=;77��W"��.3�G�G�9u�.�]�=�]��`�Z�Ρ�ڏ�Z.�W ���:u��5�?a����X(�n	W}X��^��i�ȩJ�B[ij0�Ѯ� ���D��Ĳ*3���s��ȲP�Ii���X�P�+�[2��xa:��y�gq��J� ex�~��=¦��	%�vA8~�3jcl��h���I�8`u���*��B�C;U��Z�c9�dR�n����:�����S!SP)�zj�Y���R�<[��-��©�D��Z9����U�8VL�9z�Y	#~���A6�_���ǿBD�p�\u,ذc`�|p����(Z�}��*�8�l�v�m��"�"��HY؁3Ue��f�z�ĕ_��Z]8D��1��iЁQfހĚ��r"��R��vz��+\kjϴ���&M�v�L���C��O0+Tz^:8(�+Ϡ_�/,�U�����3�t	w\�ƱA���w��a���2O�$~NS���ޠ�C����-�d�2÷T�Úe��@|��^Xhge�%v�p��*�fa��vt Z��r����gY����CJf�C�#cZ���rS0e�/Ib���q�q�@����KZ� ���=��+�a�@,�IE�^	��4&��b�ȋǩ����Y���Iw���j FPXH�˰("a���o�GaO��ȡ��7 �J��=������-�����NL�J^�oЗc��@ ��)kĪ'M��,�/z����ȶ�j�P��v��Q� �U�?T�
�(+TB���Ȧ\j�8��T E��$"_�z��s;����R�@n�/F��Վ��`/�_�V��������Z#�B��%�PVPO{x\̝h^��� ���e�M� T�ƶ+��9c�|Yl<�0�R�6����~۱���A^�N��g�,�*n�S 9.�4�iN��+�;��-�����*ϯs�\��q.�nQ�Y�H0i�ԻU���}!�u`���ʩ�M���WKm�I��:w��}��D~�ȱ(t$O�K�"ό���45c?��%L,⹑��O�#����G&��������9J��������u�6Q��t{�A���N�k��_O%g�,������
3��ɱ�.-V��g?���	,��g��Xoܸ���Gh�<�"�.3"��\�R
��PMg�"؞�k����	�p�G�W�f�Mr�p���<����a���<#V��.k��m7���a��8�5���-D�x�⡃P��g��Ile�m��6��O��}�xyttN�n�h���������,g �[�I�=U-��S�쇖���$c�[����d �f��`��?�yZ���`@ѻ�ms���1!�@�ރCp�dX����A��E���N�E;��k�p��8�m���z8Q*\
9 �s���IՃP�ҥ+.b	`����>;?��~��(���n���<M���_�Z���ߕ�xcm29=5��xT��z��)�OU�:2[�T��-�ڢW�+�����R5vF3v�̲\=��.���C� �f;Ta��˙lr�V.�*���Պ��ޅF�u��݃��v�-dmrI�K��f���9`�9.yJ������=?�}��z�a$ST:Դrs[���6}0����x����HuZ�nH�dX������Df�9��Dw���͍��4���l���w� �io����ў����������CCմ��,����7�:y����^��El*���:������Ï���&�F-߫��T�9e�4��kh�3����2�~pQ.�>Φ����ȩ'�Po�._����ʂ���}�MP��0qϿ���ꫯ����oݺ�<��Y\!�;��C� 'U���1M�İ���6�=O�����z睅���Ua����QCR�Ӆ�x{����
�u0茌�m��P����CݬK�W\��J=�)-��Nk�� ȼ4�ˁ��E�� 1D�dc���2���&3Y��z����3)QxP�La�ٳohd� ͻ��'�룏>��"��aQDg����m7��	����L���,�(ID��2q�4�$�Z�����I�ό�(�*x?3��aIx� ��_�s\���Gvmk{sy�Q�Qݷo�ֳ!��ر#���M8*��G��N�ŝHt��9�b�u���.߼q����8sss�6���zr���r�d �������=`�
��"Á�w����Aϝ;w���#G}��'pZ X�3ɧ2��S�%
O]\�4��BMK�S&.%V����� N�R��!�8z���������>.{���݆��ouZ��߆�.,��sPۧ����7��'�$=���_{��S�NA3�׉B�HO]���K�j̖"�dJ��N���������Y��<��C�L����>Q�<K�D3���2ob�O��>��N�S���pg�ij�,�k(Α�>^!���G�e����
��&<|�έ�JH"�����gH��jaO;�6n{{k�^�ݺy�СC�A��B`	���ʂ�ȀHE �qTL#�g�Y�k�U٬�xw05�b�^jyWU�:{]h�l���S�g
�O(Zb.i�4�N�Pn�̫WkYa�q|*l^����gch������k�iOirl��.ˁ[6e���{�W��C��T�c��|Ph,����w[X�+^q[n�l���=j����κȚo*�2�ls:����x�ҥ��N�Qa�������䅚�m:r},r���^��=������,,.���CMg�
�+
�4/-�l�o^���k�n@0a\�\���F��-�L=E"(��sa9�فe\e
�y���_C�Hi��T���4����ZM�"����8"� uK�#Ń������jX�E�g�����]�hA�} ��QYP26i6�����eb�b8�ú<ED�t��{w�\��R�3�\��j���lϚ��Lb�g�/3�!4��i�vmB���5<�:�=^9|�������iX%�e��$C�aR�H��R��P዇�	�w�t�#�p��� "K{���}�x�|����M<���]*�?SԹ��p��|]��ѣ���Uh���HhǪx6;�`�,��D�a�*�=7L���#uT@�aӤ/s����X*�Xmn����T�#��g�K�' o\�2�AU�Z����dk���� ��葉IVs�ѸU, 1,Ƕ�P2�Y��\,����oܸ�3��sd�|���+| ��
g)�S�8Ϗ�Ǖ�)�a�bDqj�@B/qc�iÑ,xzZ�Z�����{��r@�^�:26V�:�TM��;FC�&�@i�;m����0RuG�?��$xƝn�Up�����&��_8�^���n�E�`}��`��L��>b3�i����0C�p�$�H-@�9��d��'?P� D������m3r��<��f�o�h� ty$���#@�@��~��[[��Ε���y�#N;�2��#Bӎ�Ʀ#���-̋�H�Jid�G�~�X��X�#������H��N��Z�2"���.J*�]v?W�3��̚W�ÔS(.��B���]�J?��儕�B~)�۽+lq����I�/�-��� RX2���P���#���H�]����*�X	�����p�W��9a������8���q�����373�=�;���L��*-r��Q(,ћ���(>����j0Yv� �nIz�,�������8���ʄ���M7��o�u�r�ݳ;��6ե�$����>A~���gS��E�=%�8�>�s�I�ۡNn��E`�zT�&�:�v�}.kF �ˉ���*���P��Bb5��DG#�<�rA��xaQ���m�\m�:Λcv����.�lP<x�;�������`�Gǥ������z�,�X-�����p�+�R{k[�M�VŊ�	؜��&���� ��+�t{���JK�g��r����<[��iՔ���^5�@������$�����D���p��P���x�j�<���1AA�>��i��|.]%��J%bDUtb�ťq=㇉~��X���*�$��r1�����,l�	h'�AeӾ^
���dl���"e�����]̈�x}8�8;;,$Q�r<�f���fQQ$y'I�W^y�_��_y.�Ш,l���(��\Y^�����^�r-Ԑ�V3t$��j]��B�U�vD�g{E� T6\Cz�A7���+u�@��gPjt���0���%2����2]4��	x��F��'2�� xp��zx��v��v�v>\�vE؉��կ~����8Ȝ1��"|�/���?aBi!�K��>��#��{O�ޅ
�966J��휨��z0�0�o:�Sb�6p��v�YKq�5Q��2i�t�g�E���޽{�Pxv��N��ѣ��`�n�h֞��q5�$��P\������t�;ԥ��4���y<x�[��[��4!�GԂ�4V��]�|۴E�*3Ş{Ԋt�L� 6�Ľj�+Q\[l.P� Yd<#�d��~��,4&!a<������?��?}�ᇸ����'G��y�%����+�A��쫇�`?�x	'r��)'#�������@��������:{����W�^\���Ҫ�a�P�n0�g'�� d��³��>�81}&�V7J���sss�Ν;p� �>����Pc��AD$���4�|�V,�4M����6@�ņ{�ia��� ��h&�?~�����D���[6[Ag�����n���U�s�Xf�'�"J�7���
�W�#R�]�Ǌ4&��kv�pj6C�\҅��9�\����:���P�u�]��yag��$P*�+_���/uL�\�8����yK�GC	C��HҎ��?��ۜ&��X{aR�Q�cGMK�����Z�h�.�X[�DJY��� �gN�1d �$J�����EdJ��ɿ/\�����ѣG�N[2bӓ���"�ώ��H���U�l���b*[%���M�ey�7ҔФ�Ü���s���F;FT|�S�$C_�N��]��^y?��f�"���E����БC�:P����������>��s���AtV�Nh�R>����f��?g_V�cdc;���2���)�Zb�n3;��v�o&#f�k���	���FYk���'��0�
�o�k��`,�B4��!�����X*����k$,����ܺu��ŋ[�m�5��+��Xf��|�ut)	�=)lcJn�yt]3J`�q�(�����#x������!<��H����B��ֳQ�ޖI�3��q�<K��+����vc��$-&A�j�r�����ȲǸ ѩP���.�	,*X��<2�5��ϡ6xp�uH.�;�7R6�,�>�O�e�O�ۗ�6y38�ł�$�����'�	-���$J�K�R�%h��W.	[h�VdF[��x�e�(f���ȏBg���@�Y7Z1��2��v�/�7�9~�"�\分J�A^�fZv� �Ŭg^����"H���g�ve���̽v�Z]���:σ��c�����Ş�$��a��]J#�|K��Y"EZ�K��k5�'���fMy�[`J������tm��b�9��{��n*����R�8#���l�傤)����#I�EA���J-[:�D��:٩�)��[�m�֯V$ܗap��#͜`dGq��2�Dc1jT��E	�[X|nb&|�&����F:	���59��,���d\ٟq�n�;OC�\�PN7�ѳVϳm������(��,6��O��[-�s���BT,+���Ӊ1���-�7ŀ	,I�ٓ�۴,��b�$5�rnwe�Ȑ�2�yɥ�u)K�YN�V��'��d�~I�<��Ffŕ�;��4�e�]��*�ZD�,Qq*wЬw;�N��lt{�0�/}~G�ȑ#Q=���'nvn��\����2$}��+K���xtl$�!���HQJ�����������Ey/��]�(%���w�yꋿ}j)ܟ�LS�#��/s_���Z���x񳥥e<k��?_��R�<��d ����H����)����+�=L��$�-ZH�^,5(�$�}� �s���<Z\��U�Q�Ğq��ː����������f��4�`�n�7��˝p<�<uun,��dHNQU	#2;#I|V�1���/�ȑ��N�F�¬��'�|"Ϯ�
ݾش�ӥ�L��%�-�D�]]�ƨs�fw�-02�w�$Npn���H��e!}Ŗ#z9u�^��0���������S�O��;�o~a,�LL����{�dG��ta�@։4��T���e�
����X[�:O�%�����+�3��c2�a��yUn�/O�q��oR�*������D��}��O��R��+SаS�y��p�A�G�.���'���Ư���[o�������� M�K�����������\����h�����7�T�������G�*V���>;�LotISm\��*g���g?�t��pS�wn�D�g& ���Ө�-�ِ��J�:37�ېP_.������\�t	w��ʵ����QؔB��0$$�פSy�(t�q.��E�,_8��?����������\��Ll��`�Ӿ{oA��.�4���.���'��{��wmXb��ހD��ސ���m�0�W��l����W�ZI�o2���"ͥ�<4�����{p��� b��M6\L[�6�A0 E .���a��H�߱;uM���>s�~nI}�e�U�>=�v�LZbOwU�m��A���}���-��@2ޑK����z)��E�/ˌ�[Qh�������}�]Qbq� d�J�_�u��2�]���D���P|��X?�h\�O����|��Pښ�-�@y�⊀k��$:��Xg\Z�֘��GW�^ź�j���/UN$��aH���v�s^$����?'��rVi>B�ev`����T��K$qK\!�R���ν����ʣ���ٙ��n�pU�r	y��/�����F�G�ٳg�����nm�3gh�~X��'&�Tq��Z52�,�W��$l�Y� ��XHD�������nd���d1�~m�m;��1e���b\��<>c 4�rK� �ʼ0%�~"N��N�*VQ���ʪ��|ޛ7o�*8��`�=��?=�	�c�/B��~�z����NgbT�"��I�sQ5�V/0�!�L��O юB���3�?��ft]�ѡ)���"�Ğؓ���V{;�C��0d��w4k:����ƾ3k����Z@�]9�e�'�dff�y�J���)��/~!�ݐВВb;8R�پ�~�b�eޟ�
���g;�2;�ӳ)QV�b�!�4�y�lb�UP�E���4�ؒ�:��Z�{�g�sW[��A�O*�X��M�B�s��_?��sX����&i�W���FԐ�˗�^�|�����N(�\%�s���Đ&����ƪ
L�6W�X9��I�aʥ�S55�\pm};IVr
�]��Uf���d��)B������vj����.lmAl�'ٓ���yk����ƛ�LJѽ��[<oųR������/ =���An�o{�)v�ϩ�ih(�e��ӱ)�&���~�޽8�;����:tH�*��,��u=�e����N�;h�##Bŉ=����#c��v톫L�5�D� ��=��ay��=w�I�*������Ҡduy���X���E$�ѫX*4{��0k(�������D�$�8�ԉ�Lm6;;AR��166����:���u�fM�s=���V���I/\�=��;�E𹜑�̈�s��caY�b%�j!�L'5�J�����\N�"9�`�ޖ�ҕ�ؑ.Y�ێ$��c"��I��\A�D�8/�N ���(�P�1!�a��>my�d�p\�U��b2�)VÍaփ2 �I1��6�	_y�UK=oBc�5�JMӤ��`��L�/�r�!�pU�cx�wM��'!�2�s��ԁT�B�Af�t"$�JY��#z�l�x
B˅G�H��+�(,H0����Z�GȘm,lњ�h���-�gM��#�CdR�z]��a����s��BaQ��e÷��d+s�Q�4¦C��~�u������ҋSœ�3o7��D6�%����?鷧�q�ˉ��u�M�;_�ٿ>��SW(����D��ao߾���Ӻ�}���,�&������l �?�;k<d��8���|; MS1�nw'�V��Q��n#�p뙱�����/*�\�(Z��u(sy	B�L~�Ygf���3qm+�����Ǐ���W-J'��,���=��9A���s�	��"*3K����-=�,��)��-6���*��������������F{��n��+��%��ں�>:&����I_T� ���\��ʚjQ����44[�+^ݩ��r�9�Fw�#;������k�� ������.S�p���X|Ml[\�Ϛ�q2ZU3�2y��1�(����tߍ��$;vP&��ő��R�670T�8p��	)��ɥ��5^.w����j ֈ�;������K�����y��}�Uz�D�n��̃0Z l��\�z�
q�������Y�j0\sg�Z �TY�[��9{����|��#Z%����i:"��D�L��D(��7?7��/,,�%��3+��رc��ۿ�����{d��X��~�e8���#F�Yi�(<��6���(li��~��5āڶ�v�:�]��/;�/���#M)�cN�<��/>|xna���c��i*GP-��r��~�׾��sp��x�ʔЭ[�.\��ń �~�d	O�@�^\UZ7��	wW&��ѿ�@g���¢�������I�~����σ�?�U�t�$��8�?&5�n��I�3��z	�._&vV�����J]��8$z5�"�Be�ƥ��߹s{q��:�CQJ�,'���n���i|'I�� �1��C�`Dp��V_!ZRUªGQ�^Ear�w�=�F+f
vn�����h�5���l��a���h5�"ց�\c0�Nm#K�4���l29�t6~^^^~�����<qS��N��$���t��$��U���w�풍��2�b�;ӯ�W
���]`�Z`f�K�Ti��,3�p��33sSSS͆��I|��j�4L�6�_��Oc�>��{����ĉ$�׷ne_#�*�,A���z��KW`�ۭ��2B�L^@��
8��C������
o����$��K�5D��r؛�!���XG[�D,��o��,��៯�����n�sY�w_�����-N�����s���_��8�m�+�\�l�?��O������
+++��_�A�2�gc�)Q��a^�����K�@�"MLX�aZ�3??ϓ>33#�MP\B#�ڹF�zCv�Z����	�恱��nܸ���H{�0J$Y�sʹ}��@�\9��8D�@�V��dV��6oJ߽�u0�IS� �f�T0�#لA߹1���8-�.$�l��p*�Vƙ����v����; ���5����r$f
�KR;����#G���jt�}ŗ��B���|=v�s6�rqi�=;���)b�
���`�)��������	�������:1���n$>�߂�=�i�t�'����f��N�~!��nﭢ3Xh�p����;�av)���,����a!�X�7n��?�3a�#]/Ә���[R���ʹt�d�m--���L���J���僜jez�7��.���_�2˯�x$�G\1-��yr"-?˜�='G���2E@��(ݹsɓ�J콀 �~�|FrZ��v$��an[�!�3�('U;>8��p�:��6�/a�z��K���i���1��Ze�I�f�	D���Tp�N�>}��AFMs7���&=�5�8�jNK�Vh�pd���"$�!|(M`	��ؐ8�gtW�S�\ӳJ,�bn9%e�BӤB_�J��}��Nh$"�'?�����zC�V��]��L�l
��4�WH�n�������cqY�i!�����ԣ��J�+�ec^<sӧ�~*�2�/v��ӈ#t��|��3-�@�^z2`~
���q&�g9
�r"��瑻lU�Iy�-����xv�@���hlhR<�q�͔���=�ʲ ��lw�v ������1uy	���௰J~P��A���AMN�a�abF��1o�C<>�ʕ+8�S�&��
���FS���gJ,�����B;eX�2�����r`9�紼�N�܈L�_��D���fT0��3����J9>1�] u�vb;d����#�eIG<�e�ǲ;��
��VI�]�20dQ��f"R !�2�:�����=�!m}�x��O�/���:����C��8,E{ZΜ�c�w�0N���=�E1��/I�=��/��s�ʯ)߆�T����dFȺ�>����k��0>�*4F�d��G�٩J��au�:�oؐs;b��r�o��R�~B�П7>�D"��W�=
MD��
���P���4v����G0���jK�QӴ����HLw��V?�,`)�Z���<�q����7��;�왙����������2y���%lB/D<j6�����<���8It �(�Wڝ������s��~��~fϗʟ�A���G������q�5�EDK���v?gb]���VSB7��M	5�ʂ~���t�;��� �C',Sn�1�.����ju��д�f��x.����_0����ܒBV��.���omo�m�K>h���N�WO���y�ofѽ�5�q窰���,p�ȡ9�f���&a\M�J1�9̋��K$�}��t�-�6�_��m�m��n����>�탾�ñ�Gj͉���<>��׾H����Y��M7�5�Ժg�1 l�����Kk�N0	��z����a*6���X:іj����'%�\*-2F�5�F8~�װ1p�)��b�-Ƶ^����7�Z�n�/�������+o���������
+o��'�T[T��lg{���wn޾q�枽{ff�y����J�.��{�!<�|��^|��̋������G�VC����d�ǹQ�pK06EN�E�KFܳ�O�#�:���yg
���k�F�gߕ��tV����P}h�5G��K�����������s'~���I:�G�g^>{�ԩ��9���w�Eui�8�Z?��7�kg^z��_{��W�.Zo;��.�S�~�Z�0�q�ko~�s_a������W��T}�%��
����8��+=8��x���ڞ/p	�1h��`'=����ue�14a��z2^ُkw�=���������A�R�6miVf�󫵸����'NgG��۷n_�z��(����v^t�Nr��uh�={�*'O����lg��W
35b��;�B�7o^e����2N���:�KZ읙�`�7��у�����Q���=ac����J����C$���qP�V�&&��ܸ��	X�O)d��㍕�Oqڶ���}9� �"��i����-��|.bT��ի����S*U-�ki��S��@�s�w�g��[x�������l�v�����7n�꣏ka�W�g{�%c��d����br���#��"��Ƈ��;����	f
������ɚ5K�U���n��������;pRϜ9s��Q�/��T����5�
1o�IE��no��?r���W�_�_D�8b�Ƚ�����v���No~~?-Q�+n���k�/���d�������������6����D��R��i�k[��X����n_�D�����[w?��/��?�����@B�ѫ͑fR􅻯A�K�H����0h-�R����v�J���4� ��@I�j�A������������Ã��Qh�����(�Z�[3f���jnK��`��4c|������,�t%!W������8bK�O�R}eI2{>(��!�G<屢�����K�8rxu}C=�M%�_
�F�y�K��'�^�4ȱj��eס�[����4<U9��φ�j���ku}q����ŋ�����Wu�.h!9������ǉ>�ܙ�O=/S/6�ۛ����>��CA� Z�~�6g��\�.�_X����vv�A�U�M/��/�J��⪔U�<����*�8����z�LK�;�ՀW)�a02&��'Xȕ��lm2.y1~�����8��+kb��'Y���^{M���͛7�=���˹d:|fX��х�n�PO��������F�}�L�P�O��f��'�
_��BƈÑk	���r5��_�:�{;�4�T2f7��㍎��� *h���U��8, ����̋�*߂��jI��5��zĊEQ[Z� l�S�3{�6�8��>��We�V{��;����g�,�3/���`g�YY_�5al��;�<���OK��2ŅI*pu}m��xe�ڵk}��D)A\o�{3GK��d[o��#(������:Tӑ���c�&C��ؒ��H����M�s��`p>��P.e�=_�C!��l�������Nw�����*b����i�8@�c����{�KI����LOOׇ��C������~��&~��H��ś���*�LS<��/����t>����'S�U.c�g\t���֮j%�MU�%d�*u�"b)�{'��b4�nG��i4��Q���,A)KwI��-�b�m�.lm�!�̯���;v���H�q�z��UM��s�E+�x�Ӓ�_X\�t��p8�������-���ȧðʱWʼ�����E�J��$:�1W$i�j�&dQ۱����3;��ӔsU��E��>6*	�-�׬�dP�;59=1/a�Դ������R��Z�
/�!�����~��
6V7�9��s'�;469&<�q�+K ��������JATNV��������[�O��.o
j̋���s3�b���^���T��dJzT����.�(F��h�\ŤׅF��]�wj�^������\OF[Baͬɺ�C��jU����eǖu{��v��lC<F�����~�@�sM!,�m����t89icks{��*� �ć]���A�+1�A,��6zC�U���vg�%�q:��1����hkK�O�Q�I��/����d�~�*�C��?���߮�"7���Ǹ���ɜm(X�E���S�%ڑ�7Ҩ`�v:>"���eT�޾}[���V�#�F}�Ү��l����$�ɩQ�M�P�CCظ����{x�ν;���[�e�_�9v�X-�@3gQ����ɱ���VO�V�٫�Ff��`[%�'B�z"��6u�[��Aļsn�]J�+�ᘲ�V̸¢��@&Eh�W�F.̰�FS�Q,PǝN���%���qd���<�` ie5����̔���2�����$Y�R(�F�A���̥0�cz4/h �O@�Y<&C���5a���������(��̥���Ǔ���?I*�"H�4Y~��������A�O ��K~Vr@!�1�s!��(��w�e�x5|dO+҂��tY�/U�N�U	+��`��lP�9"�
J/p������j�K�G68�/��M���T�n�\x�j~����9!�6��D�5�Ă1�4�Tb
���un�^����2���LF�=����s"�|�Kr�Q�w�l�c��`�C�xO�~w�_D �_�U�ڮ�,2tq�qU�|�3�$T�ݻ�nݺ�����4����o�pYG�������g�������4��kG::d_nAvtSD�i�Y�	1�N�r;g�����^seLB-��TU5�N�y�*DD,��<f�R�JQ��Ç�����U)�������R����A�Z��jtQʿ��"Tʧ ��:߸~��?���E[p�B3�8Qg��i�v��O	,щ�U2[ 7���oq�N�����R(���ܲK�P��Q��L�q�WNHϱ-_B��U����+"z~�_�k��{gg�Ibib䣉��{��tBE�����?S���Ŕ�g��͐\
�_�ع���9[�D�K�˳W�S.^Bj���W�gL*��:0;�n�<~��ŋ32^`faa����\,J�	a�믿~�ܹ�'Oҡ�G�/SS]K=�&� �gO�u����w!Z[[��)QͰy�tZD%�	�p�)�\�����}�-A;듞p�&��#�UM�?�W�u~1(ZYZ�lCz�����?�޽�O���ť�^�����7����)x���H٣_~�E�e��@����<�S��\}����+¡y�ܙ��I|������C<��b0�=9=�┬�nnm��A\�K����7��ɖ||A�c����tg���NJ
�}ó�*]N����]����ޛ�^Y[^^���@fp�	_����q$v�1��E��
b���`����?�O$�.S\���T�T"l����x���R΅�...�F�c�
r�[C%� �A��[lL��t�}//+W�>I4���7�hԅ��+�7	���531��2VE�aw�$��C�._����t"3i1Y�_ZZ�������o;��i��YJ�IvA��p� {�cB
|��=��R4IER*�AWU��_�9�<��-��>
O�����wG���>��i�K�,��G8͒`���l��2�`�C5��NEv�&�Ϥrc�����Ȯ`��3nY
�$Îm?���:,�\^�v�iYЌi�˴��ũ��s"�B�!l�ю�+�ӝmEr5�	�D�4I5�����2B8B$����螺b�����������{�t��ZU��^~�eNz�x��`��3�������ygc�7��S'��9r��ڕ�{����,t�ipA<�BBv[�|g%� �̎�(;'�0xJMO<��J�r2�b����a�`�ݻ�dlbT9��z�=<�}{��@Byv�%��ʕ+�@�
�I�7�7��%Z<pJR�g�aաC:�j0E���j{�y�	��{R���Di�I,%J@+����"K����eI�"�ٱ~�퍐�Y��T6�xd>�cE��x��R������<x��3/�^�&Z��ҎP�mnn�TNz���"R�з�ZfAL���d�А3�(4x���l��e��Y�0�͡��F��B�G��)�qU�\^�>2�/"�=9k5مb1��lJ��(�,2GU'�:'P,�̌�q�)���56��>M ~��X=��	rC;d�b)�
�1,.R���%�WU=1a=Vo�7��o����+k�6�9�c���>�.���S����"�60�V����]�>��K����2��pd�kZa:����C��4Ldۜ���k�Z�@�Ghg�U
7�^�R�;u-=gC�3��\�۸}O�m�o�p���1���K/.�#&�B�������Ն�y.��������/+�����%�1��>fe�Թ%�+ӲT� �/��:��@����P<�h�ac�ݾZ��R�8�c��k8���}��$��&!ddW���f���I۸4�MJ�e�2�;ө�
=k�O�nV8�Rtq�����կ�o��H�fX���%8?�.]�>�1��/h�}�fd槰=�5�
c.�i�����)��#����ڱ��[�/\�Xfp���	!�N�R(j}�#�q���cǎ��{jj��ą�ȵ[]
�(�̤�Y!0�g��V	�eX��%"�G�҈[�Ms4�������kɾ2�ӒR�u,�I}xL�:�n˰�g�m�L������L��e����'���1g%�ot�U��{�or�_zew�<�%|X]Y�g��9��$K��x%���=��[hhȁF����V�m�oq��O��=Ԉ+�ӟ��%��<���������͑.�N�m��
�r�� k�g��L��L�g�%��:wĳ��$5��(ӊ���[:��2S����0-�{gK�$�.�\�Ν;8���q���d�&�,����#T�C^i]v'X���9".��ϊ˿ 
^)=�4��6>)��2�����Jx��J'���
�"�9�xA����-�W��g�}l��9�T���D*��E�w��*�`�C|1���m�Ʃ�I=��Z�b$�t����<�£m�+[�
ý��xh��	�[915e,z,,�[���ޡ\�3PP����;Вc�������Z^e)��v������Q�͵Z�x\����	���Jl�ѻ�8T�E��7n������j��4.�o���W3��x���Ɩ�I8��R�rb�r�D�
��/�4�'U���͉�8�g�R9l����;�[ �Dh���N�3B"���m(���������ɩW^y�ĉǏ�BM]	���gy�{8�����=��G�������CN�lE,A)�8�n�]c���4DW�х�=�c�o�m�W̴�t��$���B'<��5�i�/��'N��`���P<�,}0<�������ރ�|����=w�y�\��d�i_�����舴��Y��[��޻���o����~���?�����������O������|�J���%&X�`#\q��|�-��/_�z��u�盉�����667Z[����}���~�̙��O>��>��jG�8��F%�
�Y�T޿�*D׋�CAq�.n��W_�WA���ϟǻHڂe���m.`���I�Q�@���L��|��D�X͖.//�d
<$�w B@<u��a\� 1 �#R9 �`>�O�!X.!H��s�~�I!܁���|���Xz��Ua���7���H���g1cx����'O�x��㥟���7�]W��5C�Z������J���6X񙙙�����)A �,���bv,&�$���j�)���`}��x1��LX�6ٶ�W�
�qk�hWx����t1�zt	]/�мbrZ��!�T�M�����������7k�뺮�cU֌y�� B)Y�'K�n��r[~������_�7�(ڡ�dɖl�"�	b
E�&�\��sީ���S�Z��e(�bU��{��g�k��9Qp@�׶W4鬋|�!$��/~�����e���Li�A��{��	v��~!�LKR��;Bw+�����?�������
�]�ZƉ�BO�X��q���S0~��Ĕ�Z��O3eK�"���FWG�ԉ���akk\"�BAcl�����kct��p�\�b�*.�nؔ����Z�jnoc��t/�����~��Oq� 9�;���g1r`hA=FߚF�H@f�ۻ-C��v6�3F ����Ul�P�0+8׃�HC�/�v;��}�_�����������7���o��w������J7ɣeK�1��J�����g�����"_�|��ᣰ{�͝v�x��L�⚄7��a��IL��<L�K\��TL�\z��%�cf?��Xcg�3$P��leV��7ߐ�(4�K8:򄔣ͦ=>y����Bh�K�����R	YK0�pJ�'�V{�Β Xͼ?x��\�G�,--De��5KU���b[:{�X�%/D1�
���V���@{?+:������]�ha�f���r���Bl�n2U��'�:�J��������y���w�}��ɓ��ժ`�RY��Ip����ڔq�8n��+U�d/#�^�Σ(���t��^a����[�U��RKI�:�aKT_칡����u�̨!�ј����`�R����3o�e�"e
��/����k�B�Ϊ�s8�U�;[M���7$׋�	W�+f���`Ly�qq{|48����@��T0DKQ�����^Ϛi�`�M��d%��a`�v�=|Ӣ�+!�|װ���������g��:<�¹t�䤺7Z�͓�P��X�a��ɀ�jN�8������K�r�̈�"�'uA�U���,� 7��&�q�?.ɠ[�ş��עˍ�/Z=�!����$2רו/��{��g�# �p�kB S&AΔ`nW4fl�p7o�-�`���?C�$��H��&��<�뭝�jc�{�,$/˚Mb�F��m�{d�6I�v�Hhi�<ۑF�@�d\VGFHY���+�|��=/.\9>�-����n��oMf<��	��{Bs��w�!�=@�B���d��H�dLܪ]�/��5x㶘=���J�G�:5���իW����NNM0ۂطo����ss�0�@W/U�E	���&�'<\�$��M|����N��;c���`[�p�x����I���	9B�dB�4���)Ө�7���'OAغw��Q�'Z^.w�.����֬U˕r4����8����@�"_{�X������^D�{MÝ����<5d��� �P׋�D߾h�)iJ�V�|d~�l�65�9��f��Լ�%J8�.�k�E�rn�}93��k_�����^�ü��q�5��)�k�b~�{����Q�{�׿���-S�^�x�U�� $2��b�6�����Gtr*�i�Z�P���r�,�����i5=ˈ�,�92�Å��ؠ sV�����!4l�����δ���o���-Id)<�̳�tB4�� ���%!�D ��n��Ɋ�[�۰�d6��z�hM�����
Sct�_���P�NV���a1��$�򟹍Thɜ���`�e(����"t��p(Ex,'�,�'�>s^��S�%5���ʞ&f�Ӑ8l�{s\��&&��rOS;)�l�mQ|�1r~��X��;g�;R�v�fy���_>y�dnn���:!	(o�Ge%%l�dB�=��\a��'�g?~��GK�Y�������YX|�?66
1�tI��W��}��a.�؞$��o~��G��}�K,��� qF�SR�5=]I����}1ID�I�ӉP`�Թ�0�6I�.��gΔ;E]I��`#�t�D��0���&,��|;p��T���~ǡ䘿�E2�jw�+>^�����Dݳ^Ċ�*���>Z�W;�ط%A��'�[fb?05a���1��3)C�G�7"�(C��N�д�q��O �'B
v�(��Z3�!z��8�2�M�B~��3��ߏ�	���{��ܹÃ��EO�ݝ|���y(����&C�Վlӊ3��#���bf%���������M8n^J�J���PCj��LO�Y��G��ި��gh]i$������Y�����g?|@ߋ$�X<�_��_����`1���"��[	�����T�=�<7�K�-M���E������BK[@�.Md�	��|̃��� �������j��w�˅�{���u]%SS\��P����ѐ���"�=N�P�h/p)�xdBV.;V��7�ĳ���x̉I)P��ђ�QAX�8�S��p��G�;�[�ղ���q$���Ԣq��5�(��=S�w�7V<;�SiC�'[�(i��n�3�� C|��m&gsQUgS�ST�?��?;v�;��ε�W��t{6��-���,t��r�<�̠�u���5%}�����s�vF�,^Q�V&VQ�ьfJ.tL՚D#��%��^�)�G:ɡl�%�q|:�����Ѩ\R���$����~�YZ���L��i�u���@j4�2��J�׿�5bi�2"�Oy.\D�a`��
�b�o/Rn���,��[��N�kvv������X'� �79Z���o��:<
?*]�z���S�?ՐY�%��~qoP���(�ZY��^������ݰO�(C�����]�maaf�0b�����	�e�Z��b��yv�0i��\�B���m*�?�jM��t�ґ#G�K�RfIH&>���Ю[�7�W���H������M�GXj��Ŗ���Pc�0��̼������|����˾��b����5vL��9l�A�X�	-11k�]B�J���GB�YDqsT�f0��r%?C� ���h�N�Ks�\Rw�)}�ש��/��zh%������:ԭ3�4�b�<����UH�[j*��~5p�xlHrL�lZ$ޱ0(�iy�2 �*n����g8�®C�8.^�=�y��Yf��-ăܾMOhn�l�4"X,#VC=O�$NOO,�B�JE�;�<�
�6]L�����]�-���w��k��\q�[�rnG0sxq�*�q�5�w��Vd�BV��(B��֑�����PG1�}��i!���,r��W�ВM��l�[D�g�
�s"Q�S>x�����4^"a��W�ZJ5�rn)V�H�Bbg7�*�>�e$��/cx��.\����u*.���^���&� �JP��
5�k���i��ѩ7n<|0Kv6�q`��0.f�by�y�]���8�?u-<� ظn���#�q��}�fx �R�H&~53h�6fW{?E6T���e*s�N,y(��p�l+�;���? ���Q�u�#�b1��5K<;B�p)�7���n���<����jS���8�X��`
���S���]���z
Y���
�4��8��L�P�Bf��ϣ5Q�|zt(vև0E���.��Ѹ����h-�O	�<�5.�Q�$�O7���)gŖ��l)�V� |5�3r
-��w�Ƈ�R�2�%�t������x9p�9��2���I��
U�;Ȧ(�B� ���|���r۞\�T��0��Y�W���Mqi�b&����+�/瑊/wW"ќ�vɴ����9���C!.��e�GLl����"L����2$j��ø��\����X�n�֧�p6������
)/�!�|��cg�r5��T������:g��o�6����G��5꾭:��m��/P䖢�u�'O���]�Ċ�ypz��!"�a,�}cs}�>J���ejƟQE���sr�y����\�B�qo�4?�Ģ(�EyzEP�ȫ�^aβ[}�I����8���dm}snO��)�0�H	�ND-,���j��06c`�i�l��KD��ʄ�N$k�L��$ J�_y���[S�,EKP(�����.0Ez�B��X�̲��M�V�T�6��m�K���!ɗ3'K�jX�����@]b�G�VV�B;	��?�"Q)�$�%�X�FR���³�ě��'|�h����~����l7��cY;w��+d��G7o��jsKa!�"���$�Qw�t�v|ۆX���:��=��0��2�>���J��۴����c�!�Is����デ�ĉ(Y�rff
��e�E�k7=�&�x��Z_�x�����\ks��믮o|���<�dvnbf��Lsw�~n'�)i��������Tltw୹t��ƒ�/ZFfPV��<M��Y�J�b��S3IVV)Ϊ��fy�fsw{{��폎Ml7�34��>Iq#�����cwDv�$#4<��Ͽ��'��ꘞ�����k��=���*/��^ܡP�E|�OF���	t��TC}ms�|F��L^��Tz	���V0����"�Ղ�Uj:bq��5ͼ��vg���ْxr��v��r��u�x��*{���I���B��5� ����.)(J�O�[��=ś<~�G���ҝB�7�&}2I]�x���>{��Tx����Z�6e3Ð��?�<M��B�%��'���S��7��� �.�p<P����`ЃS
g�<T��{�2�A_����\*����?�xqq�v��&���	4�+o:KI?�����tdD��R�� ��0xL��!W��;�\����w�ڵ��N��|V�RD�ۆj/��d8��VJш���n��C�e�(�؁�m�X<j]�A�k���5J%�bh�xR%�3@���#�)���%b�Ǐg�_���%��[��n�a3�ڑ�<q?��Ϸ���Wuyi�Ν;S�ӧN��*�{���Ws�4�$��'o��ֻ����{ڌs�表�ʴԐ�0V��H���5w���c�/1J����suf���d�_?NR���D���^E��ӱ�X_�84��	JH���Q�z6E�Jtv���8Gx$:��UH����}�l�~����Ç��~��G��9���[�6�ƜL3#,����μ�5��Λ&ҊZ���"���K�La3ݖ��&��p.��$�8v�4���4�8�-���3U�0v���7�`�e��k.�Sø��C?7UޫW�r���u�j��q�������e�KG��O1f*V%2�3i�bN�Psap`Ә��Μ2��Y@,嶛��C�v��� ɽ���,r��a�p����k����nsc����
<�j���)Eյ������MbȻ�j��n_�u*�Q�Փ�����oݺ?�w������mVj�\ &����!��oɼ����9��z8=���&L�0Q
x\��4Fc������o}��Ƣ��$|;|�}3�S�Ă�`*ˍ��}���Wm�D�
���	��l"��=x���,-�
��j-I��)�h�k�� �6!�>��t�'F̜r��u�-��e��_�Կg{b8|	O���啓<cT�������fkWX"�AGe�%��ȑ#�})�JSS3�Z@�/�4V�B�tiI 7#�3H l���>~��H��!�l �7nb^ �a�',̾c��x,��DT��D˪��3mG�Dr�
o�[K��+�˸[<,M����\W��J��h��;vdgs���.�8v��ٳ�uXX�B=���]"���,��BϯWk��p�S�F��~�:Kmc4��I �T�Xy�QS9����9��1�����e�j��ˆ�L[׉�b���OI��e,�2��|��V}�m�/�β�������33�'&�ȳ/�)"ꠊ E����u��)ŦȱӼ�s��[Y�>x��n[B'xG̞ck8Z��Ą�s`Xk����X4BVK�E��f� Lc#&L�����x\��*+�!��9�.��ħC��%-���rn��������*�VtDDǧ�#��/��O�L��/_惘<5���:l���x߾}�\��i6[���*7�o����B�Z�~�>s�fW�kD�IC?��נ�� #8:�@�InL7�jmu]jוZk�]�8S���כ%�"�B�a\�\y��w[k+�K��OR��>��F���L�^��)v�N_S�RV!<�*�~�z�k�<�{�����\�s�����8y,C�=Cg3���r^���	7v�+���� ��u
]�>1��h�<���Ր�&b�2ה�ou�����?<T䕔\n����y!��"z�'�W�͙,�˯�$�ο0/�M�[!���C��в�i��I�@#�_��[V��T��X�W��V�u�c���?{��m�5�  ��IDAT�� ��gϟ�D𼵞
Q�X��Q�����:�e/XLޥ���@��/�����	4����hC;�8�-�������zg��̡3�k[�k�c>5P�RM��&��xݺs�ߣ��l�4����p�Xp~QVl�$��G_E��m���u�cj{�k�,G�ѣG/^�KIƛ0-I�xN�>}��6��J�#b�yW������mW�Dv~��c^����:��1|�^���؎���A�gy5W�tV?��|7_=Й���XJy�ˬ?�Z��i�70l"qz�hF�(U�!�tǖ~����lmm�-��ir�޽�S��ۆ�����L-d%e;���5)vgӗ;��b��>��t�4Q~(�Uݭ���X	t��L�B�X�Dh�.$�0�+;;3���R�lnnV��+��FX�����
��"<;s�̠8rT�}Wj�=i��v;�+t:�7n &�_��u�S�:(h���Y�5/rYB'�.�����R��7A�̈́�Uukb�� ���?��Ok�S�4�;���(VZn�]A�'��O~��,..��p=��1��ϫ���Κ�LN������4�m�rB�u���7Yt7O�S���Uw�i���qu�d��� }>���d�7���:5a�1��Ǥ��5�OH�t�X9_Y�4 y<y�ʊ%Q�BGsF%��1^
�ޙ3��u�ڑC��+P�`�1|8Af�U�����L����9�
Xd[������pZ�Ȧ��,���X_=��T�v��W��h��w+�C&���=��<X��L�����$~�p'n�x�R�B��T���ae�F���Ϝ=�������7/^�X�8!�ς^f��*������(���+��g�·3�tx������@AKh���w��/3�nʘ���p���"popy��VE�)&�x���.��DfkP!�Eٸ��RA7j�
.Ns��b�66�S�'�����/]�t���'N'E/G��`f9��A��Y��M����N�ń��L�S;����,��:��ug�;�.'ݗ��S(<8����h`���������/	U�ϐC���qg%
U^?_�+�a�t˨,+@H�i
-���*j�~T�M֪lY;��M*nDQ��Ɣ!���3Hse��,<��p<���qa�=��̗H��v�(�*�����Pjȿ$K����6I.��e�\�H����ڒ����g��(/4���B /ů��@=�hDD=cAŲ� �m�q��8T!������,��_~�^1�B��q$Ss��-�׫���,N\���JU\�n�UFE��2޾u6���8;�� �R)���"�����K7�\؁�����B��jx�X��A�o�=��3E�H{s}*kyq�ٳggΜ�^��&�zcD�ek���Z{���dy�&>�o��|RD5xL�Q�,fL����ְԶ���I���r���A���g�+��1p`�R�y��o�A���@�U�:��aa��G�Ĕ��=r��_��_ݾ}�R2�,�{8v�X��~L�j�oq��o�Լ�(2�0B���0qq�ތs�� LN�$�L�k�1蛡%w#Gd	y�ix!�Ri��_�K]��8_k�Ȫ������ Y/H��:�NT`���MOeR�D=BJ:�j�qn��� ���7#}���S�E���H�믿�Z8'�&�hW���b���3;&�m���*� ��e���3��Y4^�ک�z��e,K�:Me�c�ٳ\��e{����z?O.^G�ǂ��A~&�&ue;:���zv�3�o����2�?~{[��@ǚuea�"]fG��n���ָ M�����B�u���g�G�8�
�M,��f��y砚4:Vƛ�Z�Z�`d����cB�|�RJ�!|d6P<�D��X\�ʕ+���d�O�� ߢRp�x����q���DD�ǜ������r�>5Rn�4Q���R����:uJcI�-�6q��[jh<�����j�yI�:W^�Q��@��Cy�^��C�;[�L-��Qq�B��Ђ��������s,�����/tV��R%�4ą	�m�w04gv�y�
I�<���]:�J�������¾�c��Tj!�ǽvbOs̰����!��3�R(^����^y�����z4�S|�����?��j����M�������I��TY/+��6T�(���[������Ĳ}��(���Y�}2��^���N�/{p7�1��:X��v
�5|&�M�Lg�y�z`�?�����z*:����8Nf����x��VK͝V<� �FG�j=M2�٣G�%��#��U˰���d
�,.Ֆ/]HY2u�H�h���;�/�����$`񯯼�W�ڤ�Hr<L* JmIVvqe0��lK�K,�)§�����啝��A*%M&{ �%/N8����ɁL|uFE���LMh&��%y�8���t�E���ާ
���g�rk�u04�,��څRL^��[�� �J~86V�S%�Ɔa�߸y����yUf�DyXH�K$��7n�������g��!��j��L������n��݇8�
��\[\X�fD�7�`�h>66A��@�U"�m�/�&紉�^ ^tg޳���y��;Y_���vh��T�]�)�-�d�^�UʇI������T1\}�7-�k܆Ei7w/\�@�O��������� �qF��0�ן��k�cS��x���24��ӧ8���#��җ������My�2��h�UǓaO ��{hB����"y[�;�VV,�~ƚ�IJr�v��Ꝼ�ϝ� 9��3D`���iۿ����YIh���F��{��������N������?����3N�;w��^�숞�gO�D��]�?!��~�lK���+�i��G}����t��L�B���S����e�,Ϧ��x|�W���N(�u�
>"(<-%��ғ������NO(x�}�����m�>��A�G7p�{��/�
������P�}�[jj=�ʶۻ<�8��ӍӧO^�t��7�����X=hc-$ؖh�-�w���'mȌ�q6;9Hߐ�@���bJ�NsKN�,3��8��z�҅�*8�^�j ѣo1h]K �U�9���U����If�jay����.�4��p��?��v�+9��-�Bx��j
�^w~��x���^��CX�ё���ܒ2�wr�� ��7�<|���鉝��)�����E�IƟA_j����3����x����`Y�eс�_��b��/�s������~�k�Ͱ��iy�{��Q�����sq�5��k�����G
���R���Ͼc�然�*���J_�ʚ �G��h�ڥ~�����{�]S���V��_�	��r.�t��<�3I�0�N�(��W��Y*I:Lt����|֪���5��^�q(�񠹽#��f��%��יڻ��=Թ����jYGd�5�߁}���$���?���G�|ˑ�jK+Cns��Wg:�>��h;���J?��7��=Zg0�]rm�B�",����Qw?g	��%���k��*X I�C��!o����JbVʜ���O��U�y�ؗ�`ei�Ν;�����-�X�u~��i;�^��=��ֶ�P���.���IEdbbD���ajcs{�ՙ�K��o]�8����\�bл�,���r�%�̆�<~����0���#���<�~�.��V�4��Ib��/����k��::������X�?���n�ɟ���H���AP[̰
���C|)BJ�n��뿖�^�{G��X�7����q��H�UM.w�IRHWO%Z���\���+:�"�l��F��ٶ�V�R$5�� �v���Q�����n�vW�V.\���,�k�ɾ&':*׹�ϟͷvw�WW�\y��T�>������7n�|p�S��T/b���$�=�ȔA�VF=;~!����]bԥ'��r�ܢ�29��g-�$�RC�E������qI�7������h�Z+�$/p���r���쳙}��y������I?9�ɋ�VB�<����<źd�G<��+�YQ:l��y�7�6��	߫�E�#� ��hC����Fv��00-��њ���I�S�a��l��O�����ҡBGFG��dħ���0m�v��&�`Ǚ��/�n���Sp;`��D��7361>1=U�Yb2l����*�"���:�ˋ�S�o��0�RR�5r!�3�%I`�ҷLԁ%K�Y�9����%�F�2�N�ɪ+#�����|�Fd�{�D쓓�������>�����9s����/N�GhŠ���6[�����J��_�vz�[;"]5f�:�����	�k<�p@ny$2˺� 7�!%����LL�ˊ�K�u�b�S�k<rԛ:{)��3K�4jY�-�*JVϦ���T����azb
�
�6��5O�e�_�m]X
�����������((� 7��
ЧV�j@��D۬w2���H��PY���Ν�d46�����RQ�
'�g��%�-ߨL/N��@��kV���\�YO�l�� ��M��N��s�_	�����c��~�J��ɤ..HU/�`y������H��R/�e��;�[ܒ^�ިC�T��Gml?0USm�(k���@AI*ͧ�b\�]t:�_�˞�7�ь��y�ERj`�bw\��`<�.��:�����8�[�s@�-�ƺb�nYe��F�1V�����h �J�%#ͫ��z%E��>�/_����?���\��C�,�g�9_��{�k�T�[P�A.�Q��%�>�\S�>�'&�KH�����Q�3��u|v>E�Wq�ӧ_]�x��i�ӭ�@2����NRR'n������!��eN����3g_]�����ڵx�Զѥ;H����a�ѯ-�55\f�T�'��B!$Y's<~�M��o[���-֐'��+ս9\|�a�ɰ�a�-�$/$w_������{����;q���F�LQ0�Q���&&�:Z��4��%����{������3�Z>G���-��g�`wA(5������l�o��H��Ky�Ru�=m��Z��=;A��;���h��%�E=ɬ����-���X%����L1M�`��7�}��6�'��>�)	|��r%�	`0��<~L��i�R�s��ǌ3�HA��";�/�44C;Ñ�R�L[Zݛ^Y&��ϟ?O_[/�C�<��T;N�2 Y.��?��Ea�@��Rq�1t|�):p�V� �~���3ϐj���o�}�KzW�WAO�j��.�RU\����<��:����J{��@b9]zcl؉,�S�FQ�<����<y���Cu݉��L�M�,X+z�0�_~�%��w�y1�O~�&V8�o�r�"���oߖ��J�RR�v��)H�࠙Zh(9G�N�<y`f��=@������B��l�a�N\�;��3A�F7U��Ө���v8#���D��;�M���ﳐ[u��Z-� ����E�(Ԓj���'{�o�ۀ�U�37h_9��+y<��ď9��|�;�y��w��Da}p}X�a_�onܸ����Y�u����(��$5@@y-�ƥ�~�m�:}2T�֢���ff���]Kn%X6/q�(xwۦ��%�r;	J���1�$�1d�)�[o��v�Ѩmnv��/^lNL���]�-�Qy���e� ���F���Rmz�t��_�� �L�@T�uˋKئ��uj<,1��+DS�N:�^�ԐO� ��N��YU�So����N�u��Q%/�C��z+����[�)����W��կ8-jF��̤Ql\m\S���ҫ�m�O�>vL⸙�w��]�v�o���BTth#q���C��S���ؤ��C�tF��U7@���o���u����gౄ������tZ��;�d؄˩NHB�*��欖l!���"���YЦ[B�(����� �f�Œnnn��R�x�'F�D-G �W�-��<)�Ujd �r�Ľ��8
� y�4��3� �U	_��3:W���H�1B;�*�&�V�	���%v����;+�h��\(����&���j@�vZm�hND\�1�g&�}��v.p���q���yl>|����YP"i 5�F�W']h�R�a.�Oň���~��� ��<����~��<��O�.<��K�i������B�{R���J�q*��x��&���p�jIe�
�;=Jk�|'~�����{	 b4�BE���2��b_��j��5��>n��Qb����[
ހ�w�7毠*y
�[���։�_x��!�4��]*"I�T���� ��߇f趺��ַد06Yg;0�Kqv�p�G ᮕޢ"7��+�Ξd33�#ﰶ�"n�m�(S9�"kl.����B�8&j�b���[�V��(~���q����d����7�N��l���ѓ"@%qJG'����#�L��kk��+#��䘔�t�,EI�DP�u(�]ކ@pÁ�;�-��Y SK�G�:���B�RV�ѩ�ӈ(����(&��ۀ��N��2�*Kű߿��J�tLhcV��gl��# �^��j�.�3�����PrG��E�2AyXI��y�WD'�r�0l0��͙ųu��� Q-;�p��O�G���ֳq_���2i��{�Fd1N;��Y{�Yjiά`r��xl����jфO������
v���T	I��W�J�2�ub19N3Ǘ�S���p>2��1��)�09u��C��s��;v�}uE�c����M,�����#eB���7(
�o_��y�eer� V����>V>�V�Wנ�Fk�x=�~�Wo&t�.��33STԺD1�Od5��NN�svJf�ݮ(��7"�%|�㌽�^�r��x�����7%�$�k#����S�#�_���؋K8p�����DU"2���������J��C')n	��̞���bg�9�C@�X`&����Ef�a̷D{����.o�"�����Ƌ��XL�A����c�l�"xJ�t�¼i��i�����Y�.�l�o��E9|%K�����^�I�(x:ƛ����m��I�L��i�X@TA���Pm2���������������0�I�o&�<�8����%��R�dY�$3oE7�0�m�n�����׳�>����5Z�4A`z@`Kz��[|O��^^��3-�O���A�����|���>�� �˥J*$P�@�bJ�"�3gΜ;wN�J�:�h3p�U~J'.����z!����\�8�+ 3���)�u���?E�*T���,��y���!�9��J�(4LfZ,�j�Lc mނa�Q|]|���ϩEM6�rJJ�˼�<�2�:�ɓ�Cx3��&˦~	�*��#�N�7�ȅ%m����Ļ�%]H^�V���������v��f�K�ё���i8������? a`��hX�xO�+��BDɌtp�}Ne���������~qb�J=A�rһ�0զ���(��J3��L��sY6'!�g�r�ye6P�h�I֓�ӟ½�5=��¹��C�rʫx��j�F�8 �ng~ib?Cl�@\�RJꇴR��wv[pG[��8%�k��7����G���$��ӡ%����^�`\��$��)G%�t|d,6a8��Ħ!v��Ahu�X��ߕ&\<�T��N���T�Q�3�ӈI�C�{b�qWD٬�X{���å�j�/�^G�:RoLNL�v�1S�ס�ճy�/�ⴕ�i�%k<�Wޏ��9���ׯ�IJw�(<,��AdH����ێ{�3�mvn���J�To϶Y�҇%N��J���amd4����5J6�	#LY4IWg�d~�^�A)��<��h7#�\d	��K3��B�,�k5iB�������	eS���m���s��".�lg##�Z]6���ɉ��[���¶9�FG�'�����v�̥Ko��&�dya���L��͋��0��R,��ٳgl��!�rҢdӖ����W0k������,;ۦ������ENt�Pjn�N��jώ�K���Ȏ�v^�������K��	),Z�?��w���p�_����6no�ܺuk|�����n����ac���<��aY��jr��裏b%pĒ�8qJpL�掌� ��nl��p��+�����S�~���������P�8� ��7���O��:q��{���������M�$�CNl6'hM�'�Q�~�99���e�[���AP��o\������o_�r�Ќ�v%o?k��qA�={�}18�M}Q���/��)��k#u�ŋq� �7n܀��#��F{��'�Q*<_X���>9�X�/��{'����$4g����y�����G�8���Y����g�p��Ո��n���d"7Ӑ2Z_��M�e�̄2�[	g-#Lf[�@d`�K�,�!	�:��hE��3;.�~mm�z�k�Ih�� :��/0�~T�U0D6��?޼���_ޝ}�D� J�D0�'�|"��㇩*Y�rzQ��Ǐ�����ts�����������ƨ'5
��0S��jt��Y>_�$�U���QZNz��:Qgz���3�V���ǯoܸ�+|�߀O��w���;���rԶ��wRPZ���Y
�o"���A�`S����	�-��ƍ[Q$�?�.�0/���M�w�4
+��
k;�s�?�^�"�E��&ĉ*��&�J��P���Ci���-���Ԣ��Vtq���hYd�2�R���Qv~�9����Hc_p���~��qK�10T����,�K�r�z��$���������rss[��a)�YVG7a�K�o 2 �Jz>E���Z
Mk!CJ&����SA��ܲ�Dڮ�̠�~f�����u���e�J�ʢJ��>>t��t�i�MFJ��)�{Y��4S�����-� ��_XX�lÛ�@���ut�p.J���B�AAB��1�� (%����Y���a
�uf���Ϯ�(�Z��H���s�34���z6�m����>~�;(^z [�;�B�v�� _#���Z�V���Z�Sk�߻�����q��}<�d��(4�N��u��ZR���A^`������>p��X*7�@��p��2xa���"��拹Jt��!�7-� ��l�lu
��%&";�y��2 a��o����Պ�ӗ\'(U��a�?q��?>Щ2in��p�����Ү��w���8��Q,�A�Ղ��W�ѣG���4|�����ǥW�
\����'�e&A�s��T�m]$�.��mļD�I�ľ&�D�j2Tx��i�����{��Iq��]�*�ې����͵�޿����e����HPb�@I#�N�붺�M�O%���{�H]�he����о�L݀\�d}��W����HC|����+s��2�����he¯86��&���e�|3��AE��1������ϟ?�XcJ !$�V����GGǡ��lJ�ɩR$��f3����VST��Ǐww���7�1����W�@T o��A;�Qd��D�9�oo&;@I\�@����%1L����67�Lj�o�� T���E���=�R|˯�Y�����g��nXb��L F�_�� _��y�h�x�UK���T;�Y�g�vU_<_8��K�.���0�X*a9�6
�zB���q.D�O/�2+� �\7�{ND;j�YCO��'��_}�?����7e�u��+�Z_]�\1�xC^��՜���"�W��BX�0�ԃ,����ea������>�L�8�x����TK,�a��ǚ��~f�����S-}cT����po�p^����7������.gO,�L�"�W��evЭk�rΆ�!����&�m2e��7��\�z~Fg�T�i��xz��t+�O�=�<yr|b�N��pfzcy�y��$x�qس}�~�a�+dU�B��+���NM���z�A!*z!�������`$y��:�o�,+�I��^���K�eI��f�bˬ�w:��Nv��,-Zf1���XF�̶ë��ų��=���y�8�ܖ��KJ,�7%��&)!-�{��x���+y�R��V>�9��>�@�v��י�QQ�hU!�I��{��T��8��</n���-҈��"H'*֞g��Ȏ�ʘL޻̯[:.~b�+��ш0uUQ�����.�$[cG�v`j�r(�\���s]�:�EP��J�EԒ:R��EB�ͼ�B����/��ɳʷl��y�*B���+���vxfE�G:ό2�\RKx̬1������I��j��b JF�3��?*Yw9WJ�5��p�o@$��8q��iԒ�\���׿���hPe(
y�j50ӓB�G1��B�Bfv�h�)��b�|�C��uG{L��hRۧ�s~KY��%�I,��ӲL$30�X���r�Sг�)�VA}���&��u�֣Gd�\{��&�;u��_��_��� �>�%B�r��]|�9�e��cU�NM�Q\�9��[\[Y?<vl�|ay�?~����گ~��K��3���Rlm�`��ܺu��O?%�c�8j -��$�s�&��; ��ʧ#����=NĨ䚕������8������������ ���ɿ�ۿ}��u
�S�t�]��������w�ɳ���{�����k�߿Zh~~��ӧ��O~6>^��V�p�%; p��_�СC��w���o�"����\`z����p�-;qcW�\f?^;�-&��S���:,�J�-KLԪ���
��Ѷ*�.i4:�2,�޽��1�#�/_����я~�����~��m0s�w�i\<��a�m�}�#D�9���ӧ��/�����k����_��W�;��3FM{B_��*e|�ڵkx���]L��{�._��������$R#R-A-Ęb�E#���۴���"�1��M4�j'�\[��O�>D���o�Zw ���{�	���L�|u.�hr;�8��2v�-r�5��"?��v(��U�̰���T>��@���$��O���ө�0��!�M�p�e{2��&�8�P8Z�����̀k�;�������؊�r���g	����Wp����ѣG˖���]f��d������m�K~9��uޗ#`�Jճ�zv5�#�0x@��	u�ޔ������=�EV1���j��+�j5VWW��G!���6��ѐ,�f����Н�)�@�OL�b�g�Ce��"�C�4�N��<~hh�&�|D�mlI����/�V�y��T���|ۮ��)��
��>q�K�1�@�q�����/ Jx'[:���S�tX�B���0
]�zt\�-&�r&����n�*e:��F;��T|�c�H���m���Xs��A�**+^����~ÃC ��>z���S���.�9sv�,�b�����k�� kpc8P��N)��8�߉m�s�ۉt�J�!?�^�~ϭ?�L���=�Νa�H$$1X*l�ڷ}��3$�+���j�Ն��@ ���!Ԙh�у�w�|�0�E��rs&,�t��Q
?ׄ��,f��m`'��s��v�x�f��A�.�t��Ȏ9�]����O`���h�kٞPv�r�ϱcǘ>�6�_<{�ء5Pe�D��G�r�
N�0�!&iqI&��}��A,����[��V�I�� F��旰KK�#T-ʌq�eÁ<�{�#��8=�+&�x�e"�~jz"+@\�G�G�ebA��ސ=���x(\���l�ugs�g���v�P�g#�73$�!��/�2�kP�}M:��i�v����x,���S>{�@&���LO�kv�1M�JKH�HI`��d��87i���g6������U�hܾ}~(2�-n�G<��4��(�t��,
���O�����3:>6��z����0�\����q�I[3�+��B���F-���pF���63Xc��b1f�K��R<�.Fv!*� ��VXv�X&�;gB�1#;�X	P��8�x<������Sh��3������6��{��20�,qo�|N��j��'���ů�(���Sė�`�qX��α�S�AK�%������d�f�|S���|#C66)8�z}�D���^�R�{����,μ4.�����2���=o/�ZLx�\�)5�۞�f��K8`����W�5T���A[�J��v��,eF�P����ٳb	���ٖU�%�~��cF�V?�8y��^dQ�Ra�BkZ!��T�˔}]��>�Fb0,�a�K����A��f� ����0�ٹ�v�;��/s=q.3
���#�,�|�H�gb 0	~������g_��Z�
&Fs[`��7Z_mF��6����2Es"�?ݳ'��,��u�~jY�EEf�oa�U���?y$sS*ò eHn쥦E]
j�J�?9!(�����ו�a�7�R-Vhbf���=O�.ʳ3�uG#��*�48Ŀg'(�9Ї���ZA5H���,��5������	�TD�C�ff�E��8��;w�������y�%����H��l~����Z"�e�Q���XS�BZ Z���lʘY?:����-�A��T�dC��F�n��E+g �j�2����̰q�_L�(�!-�q��MU���"F!T���T�ˈ)���y&�W�2�"aX*
�ZUiX=%�uh���O�9E,9�¥:3����b�!�T]��(�f�@���U��ri��қ��a�왅 �=�hL��ʜS;ΕP�?Юq�|���?2^E�V�*��Dz}��wT�=B�GK���o������,?s�} Y�,�H���T������� ��/��h
q��;�^���Q���WB��#�z�
y��ҁi�����/"ؖ�X�g�V�v�����'�?Y
��8�D��:#A������Ǐ�o>��c�7N?�����p|�߻�;��ޅ@ћ�����������'�5�
�w�~������.���0Q�ql��83B�p��������{G����)�����c���_�!]���d����>���]�@�ط_�Y5'7n���G���4_�z�|���e�Z�Ǳ��k��n�Z[}Ap��y
�ݻw	ѭU�B����Z�`��C&J��wT�����K�7g�5��Xa��,$�u������=\���o�:�h{N��<M�L��
8k��.�v��'�����{���-d�F?������\C ��V��v�KQ_����\s�I������CE@A��[�teq�?��שT�:;;�P'��d�B�iG��X7�ۉ�g�9�߿oMv0֘��`��hl��S�7�;^��B�|��GG�ӧO=z��jW�¼N-~�v�-|)�}n�<�ZR�^?�!2�VC�T�1���i.�� dcL���V�1K����2Fe:V5�^l��XB}���^I����w��& �[ۛ8��Σ�������3O������0޻�@(��[*��
ZF�&|���ӱ[�W���뤤q��w�aŔU]�������)�B%��Y�
���0���=[TN�˷c�(ɮ���u�m�Zf��m�u���k���v��
��!R��3
�߉OiGpY/��C�~�V�H��N?������(¾*y)	�$��j�\q~yj�f����YEh�K��<�6��p�!��V�U�iO�at+��W�o߾s��a�w�J�狻5L9M�����:2�BX��f*�����ln^klMlt�-����	p��2���+��>憎����8'!PС0���w���ΊQ��8J�Vw�"�"-�;'S�nX�y5�`
�0��F��v[mu���I˓��S��⮢L��HBT]�����vZ;���M���?�$Ώ�c-!��uY��l\���)�wN:��V7^,��V6�-g}\�,���2��������:^);0�i	.d`�^���i7w�^��s,Q�ju�\����'O⼰9	?�v����+�$��3	�+/6�׶w��z����{�&'�E��>!���	�
��L�r��z���R�l�k��ȑ�b?���<��e![[sX�fDY�l32�V�«r�:$�+��0�0�,�-.��Wj����a��d����I�2;;���C�x<e�Ĥ��.,,%���ݮ��:�T�0���O#>��Lo1�cw�oO�bՄ���<x� 7������ʴI����ꉇ-%�4^\�;_ޣό�a5���P�� �'����ܓY�ݠs��<|���I�Î=�~~޷!���rj��R�х˲A�asg[��^��{��I`�Ls��f���uȾ˪M-��R@�q<�y` �L;v��ۦ��͍��L
,��Y]]��) o��T���B�K�+x���f��Ǩנ�w���4*:I��X}����W"Ò\B;�����A?�v|��`�\U��~2dIޡ3�X[�\X�65����:��CY!IN�Ԩ~hE�ۡs.9CLU%K�εc	��cB��gN��{X�C��t��95�X"eL-�K������
�w���ĉXOz�X;�đE<�5��T������l��=t��@T��_
W�g)�R�T����,=B��𿍵u�o6�R�&�����D�ݞ��29@�+�d�d���`�~��Ԃ���4�$P<%����xllf��J���������0�e]]�,
X��,3�g2A{�6/�|�J���l�,�]˻zӡ�{����g�����YfɀEG�1?�ṹ9�j����I(=}�$EI�h�`H)էn<�lr{Y����c<����N8�¸a�'W`q�o����Z�ev��hҢK��Ѭ���R��6�PR8���庚£2;C����{:�x�,�8} �f����증!�X�d�(�~"�{}K!�TdBwa}u�3#C'0Λw�W�2�#pU��"��S�A�;F�+ז*���í!�B�<�̔�����
ե�]@�۶e�t�,I*���LQ	ŐZ*k���ӄ�ȭ�{v�/�Da��r��SPҕ#��X�-S�a�W,���E��7��͙�Yx��N�Ƕ_�bI,�g)3K#�@1�N�C�8���d��Yތ���28���R\dl+�i�)M�0`�e"@�ӭg��iQ,iO:�6��m���q;�����bF5��]��N1�rej�Ԩ����`;	��|[��,#xf�Ԑt�-��H��\y�dQ!��R�"K��"�qm
 O-�W|\���܅��E�©��c	k<x�ɣH�(��٦3�Z'?̰�Mj��6�9��/���'"�Yhf� !�I�+��j�+6�ƍ�����$eY�~���}��^�t��hdBL����'r�.�/����w�Eh�?��>}*dX�Cn�3��p�Br�����H���vb#,�g��Dj�P����W�\9}N��<� l�S�N��wo��duvs�^�}�&�ih�5\Y]�������~��|@H�ӧ_�N��������o�&��ϗ+��T�6V@Bӵm�k5����D�?���b�	؍�=�$��\i�1���~�Pǎ���iA���s�b��		<��m	��~�m��o}�
�V6hq��W����gI<���� �_���G�B,�����#�x�bu|�g?�	�V��Kt��-�2�'
R�S|�ܹ��Clހ�C���G�$�p@V�:˞a�a�S�ND����2n�<��^��ի� V�1х��Wha����U'���(�x��p�����b�9;�f�>Z�=Ķi�S��C��s�&hn`i��2��C���\$�������E-t��f��[<�g3k�Ki�ڥJonmK�mfL���?��x��9� ��t�PE
r��q6�8$����&&�M�Gu`nX�wia��o�n.�H,��s�yH���-�w��K�G:u�e�(A^���lwp����]�5�f#�~d(⥥eh�H�γ8�f�G��NقCw�d7n{�t4^��B۽�i��fι�DT,�.���uHZ+b+�.�_���o�^R��jE��O9��Ӓ(�\��*�WGHQ����p���K���2c����L�m7O�/SC��M
/����)�V1�/���Ɩe{S�B��
���K�m�+R���e��������0D���,㩩vŨ"����cHx�z�)�T��q�9�4�(�jubl��	�'/)9F I%2ƭ!Ө�v��=�!�ut
6���Z��J�q�s�8�@<l+�gR���B�_���kLz����fZ����n�U���<�@�?Q�g�����Z��1 0���.H����Z.SB�\F.��Y셍L3w2[�v���d�	t����K��]c6�R�~@�	o	�caa��L2b���C�q����5�Հ���pS���~볺*�P�X�J�D�,����Q���I4�RE]t`.#hޏ}���(O
�����!���z��
Bh���@i<���xe
	��8;;KG�Qd��m|>E��{�����8>��YYY��!�t{X֥"�=M���q�7�)����(���5�Y�*{i�&��RW�Z�uR���Yr0U�%��2��D�ƔU+�BzrkR76�8���o���K�e�S/-/��9��$9G(��Y�0���"M�&��0���*5-���z�;��UpM%lmAi�t}>{�X��A͙�6PXq���1\!��J����<��{P��;E�UQ���F'�0���H>"l7� `����r�'#"�/Pz_{Rx/��?���b�W���6v���})��R� f!&�g!�c�s;�k{TV�6��bJ��.ԧb)4+���J=F
���-&vu�h�x8؆�Ȓ�7�]b�ʑb�3"�DD�
��!�1S���BK�����M�|PV8���V)w�D�@)���<���*n��Y��tvI1���(�v�wkՍA��>�d��;��9���ʕR�uqL+ү���>{V��LC{Y� ���Y�K	�D�sJ�Sx�t�˟rM2�����>��w<9�/@�� �\�q�/�od$�BI\c)<�O�87��teBb��r��+�lu1��d=]���Ebie���6�%Ș��p0����\�!SO=)�/v+��'zcl0�@�l�Q�*5~T.�%�|W�K���m,A�:�	o�Kt[�%b��^��0``����Vw�qP&=���ib|/
�o+��5f���27K�]�)q��gss�A���T:���i�}�t�8+���Բ����-K1�%�'o����=ZATt.���|*��v��3H��e�����\��Y ��O��jRcT�d:�K��B��dA <A����,s��Y�M�3hg�晫�<�Kd�P��p��-�K���[�/�YvĐ�V~*U黳��k��Ezl_����ٌ9#g�2�@��)k��Oj�PH`����G8����M}e���$�W�>P�Y~�Ԅ����:�����������3g:�LhC_R�������`�bW��X��I���x{W��K垶?�m0��fR�+ժ"���G%���L� ò����+���v��c#2u��g���V7�����UG�<a���wtRS�8�e��<�58d������?��d����6	�����>��l���+��'�x`YH�ٸv�ڑ#��y�Z"�?���d�v������&.U799K��j�C�_���f��LC�<y4?���Сl���`��zf�+����`-��~�ԅ�'Ob���:
SS����u0�֖��~ �kM_Xax	��ƣa����[
��rS��N�8�p�%5 !ô �K'���g����#x����'��q��ѣx��/�ߙ�m5w�ݞ�{B�f�`ٱ���ӈ?�]{���qa8��;�O���#�,o���7>������|��"����%��ĭ'v �dF���og�F��`5Μ>ɪ�ݻw?����a6�l�g�~���;��eΆClp�����:z��_����Ě�"-���o�S�b*���I$/�Ԩ�R?�;R6�~rux ���PSп���&Q{$��%�#7�b������B�q�%ހN��l�[T#�LGG��=XO9�Y��tc���jt�d���j�����s�]�T�Ղ�ɩvwicc;SOORZ�C�&�U>��R⾒,W��"��YȘ�Ö*���sV��Dڭ6� �.�/�2c���͚W������i��2о�'�}����¤�i��%`'����<A����.{�76�2��)y,Y�Q���b'J;���܂#�qD`Y���L�:U|�
�$Q�b7==%[��j��L���`N31I�=���=<�кg�7wZ8_�=�p����p�yһS�G�٣��B�$���Է�g��p�`	jC^�-:60�xn���"+��Ʋ�Yƒ$33�R�	J�e�e�S��%��c;"���SS�A%�ǒVld����l~A~�Օ��g���
ok����lX��$m�$k�m(.�	���I҂����0J�%mu���Y�L��Ҝ�X�wֶ�26�ʜ75Hb�V�V�.a���{�/��p���gss�������-�.�,�}~8����(:��<K/�X�*�%ނ��[�V^�^�t�=}���{�sN<��w]x��SM�e����.HO��Xiv�����D���,L��[��SK5@G�
w)�*�`���	� wMW�]^^�m1/��,�6>�� JJ�BU�����S�9whI_G�Ȁ����r��A`�R�kKg�S�?O}mC�Dg��=�q�A��h*|>�M��	vނ��Qo?�F§������Kt
���,�/~��w�}υ�?}�R�O��tܪ`�uv����_~������b��Ɔ�0�z�޽/���ҩS�Μ9�u����'�o�;���5��ř��#߹so텐�uZmBC�:�����n��Ī95@nA5�,{���5ƅ=9�u��ӹ�+�ZX\?�#��c�Ǐ��{t�vw۪F����jȄ)[�q�/++kp؇�}���8��M둌���0���(�PV״���}[KK��5?�^|�L�Sㅳ���}�{iw�Qɤ�K���IS�1,9�R�bR�ǥ��c�K:6�D<�.E�b��� S���rѓT��!#;*1~#���)��.û��u���R������<ϭY,v�:������L՝��^.��W1��D|���ټ*�x�~��@��G��gs/^,�@���/.︾4��/��d���H��#�F����R�R]�ŋ׉G�w��~������+)�L:�S���ذ�O����i6��oc����kut�2�IrD��*:n���9jδ)��+J\v:�XgԹ����y��	Q!H'C��?����ٸ���;651)�e���(.i�k��p��y*}�y/'�bo��
M/C!�ZP�4'�:���7oބ�GP�T�&
�[x.+W)�Qb�a�.��M�ԑ+�&�I��=��e9��|.m� ��U�$=Q�\�=��Y_�lM���)2	f�$���.����D�O?�%��{gP�˗/���7o8_ߘ^�T�����e��
�����x��Q�27=�<�e�&�f\/Rb)�\��_R͹�v��E��F��%��x���a~�������Ms��^��ju��Ţ%��"�gIi��w�S�HeM09�vh�.����iO�tiA��c;�ȳl�����K��j��5��֌C�1��<[Kѐ�]�D��D�1[thT��13��텓j.2���_�j��e�M��W0�_��*]Pe�r�v� ����K�q+5�0�
��Ì�g����oy70��p}��XJMҋ�����3*ԽYa��_ ��5�$se�-��L�7��v����R��ݾ}�֭[t���SPC���u�_,��B��?��?�;wNFO(��knN�P񛙙�Hym����
��[��I����h/9�%	,|�ÇC��ڠ� ��B��b��\��������!7�#!X�x�v������Ϟ=#���܁e�γ��?l�Y�e�Q.��x�2#2#�2k�IW���F-C�5/������	`��x�3a\�
DIHj!��������!"c:��s��{�,�c�TT�9�콖/>w�\'�bU�A��Ƴ�?�<�>OXj'�0��֭[C�˖�G���מ}�a�xT�.1b\Klo�E�'�	'i�^�β�Y�#7q���7�Z�>}���_|Q:�4Z`>����޹s�g�2rh��д�����oÌ޺u��ꯪ��p{�c��V#j�Z�T;���ƛ�X��H�\ ��'[c��ų�,0��>����Z�H�u94����u���l٣�x�;w�;w.�q���/�KB~�����iB3(��x�%}�"���!K���/�\k�<�������w�����l�E�s-����&�U��y������y�Ua�7N���y�����:�%pAx �e�1&��!�bm� |_6�߹w��i8Ds2���(�ʁXZ����IZ��`ܗTw���Q�6�(|�����&�֥���o<�ǃ�X�?�oò`�7Y����O��瘟�UKH.�1b����4ai�@�+l��{VWS�Kĺ�Z��B�z}yy�s�r�,5 k�(N�Hf6ȏƨ����BJ���yǎ۠����UmPk��E�
�� d��o�3��=ă�T�BgN��in^�aQ�ѭ�{��e	an�TS��S�{�3Ku�~�lk�/���'O��,�\����bdx��1�>��Hzfy���U\��/�,�t}��$�M�Ͽ���&�О�x��-:�xz{j�Uw�䊴���<o�]9i�ad�t��#�c����ӅK��"��0�m��O�4��N.^|zxuU�VU�^|�����Y��>�:�.�KY4VFT�����?� 2�~��Ϋ/��3����j�4����}SS��욄i��8�+SR����J��NN��y��\��,���XK#ſxX��x��Q���/~�͗/1��w�(�П�ڕy���.,�B�v���˗n=�P*�բ�{�'ݟ.�=<Ԫ���)VKM4��-���8�r<�୲�(����Z��Awh��扯�o%1W͋�g~���L�A.i��u(�� ��� �3̦<s�*U�ڀ3 y}����"C����S�γ>�7Ձ���aa�!v|���4�hVPp뙴h:c4�������=���W��Vڥ8���;kk!j�Z����~E��9�"��cGM��3֢�B��9g>�G�	7#��W��R��%��$��
7��a.����]��M��1����>�i:���BK�.�xo�裏�Ee͂k�V��a�fyy���R'�qF����8Dd�ܓ<��h��楟@��c�6:�E�n �?��3�b�p�J�����Z��Հ@�K�u��ilm����qL����xi�(��V-t4OJ�ui����j�s�KR�D�U����ӛkZ��׬�fD���F��t[�n��-:��S'������
�
������8��������[wn#�eU���g��#�c�����&N����`e�i�d��^��*��f�����V��\?��n�T������d*>�P'h-�*܊���,����6�li]��N��(Gg���^���7FZ)w�J�k�9�F*"�KY�,n�B{~�a�h�d�@"�Z��ڴ�qqz v

euEZW�z���)���u�N�H�lZ���}&XwsdTz>����4�:m����a�q�?��Cx[��y¢���p �-Vؤ2G�;�z&@Њ��B������ZH��u�Dv�Y�kxc��"'��܃A��^��b�8=n
ֿ�:j��E=_�p3 �¤I��&77S�'�%�nSnF�і��*������ڹ7����r-��W���Q�wpQ��D�00�QA|QO�DK�%���v�����^��^8=��X�9�ʕF�uȏx�R�ǡ�`q('��9G���LF�:����Fi��Q�!�����J�fօ�T�	��Zz�D�+cu��,�k&3�?^-��\�[�Ț�c�$�;�7��IJ�PX�FP�?�oyY{��M��}��U<}��JuE�����d���Gbþe�v~��gqeXz��Y֦S�[[㕎������,�6��{΀K�Qu{F\�C�ـ� :��ܦ8��-ϔ��W�+YU�wU�$�ic����.!>�5�b��V@Tr��Ʒ�}Τ	��K/<��o���_��A'8�ZE\���덍���m��/� }��K����p$�u�����{���?��\-����f�D�6���l�FՉ�58fL;y�v���������<~b4rR�A�>}ze����īZ_���z��������U_�ռ��xv|��s��vx��LWҲ���������Ν�H2lNg�`�76��Y'�={��o���k�aq�ձ�>��N�K/	�`_J�ox�hSZ��K���� �0u:���nk�fM����x��\L\y���J:�Ϗ<���/��⅋���/����o~�=�w�;��;�Ϟ��)R��<sfD��:mQ;���&?�h�d��4�m�c���w���Ō��9��($?y�?~��yM�&\���Ν];z$Ҏ�D���JuK�����x:��A�Bj��/��j�7�D�4]_�O��Z��Τ?� ��'Μ=���N�<v���(��ώ;�����<�p�a�q֤�N�4X����������k5�������߸z�Q�t"�*6��xK���q����Cҫt���F�!�� ���uC2,��\�R��l9_L9Q�]$�/f9�@*���+K���1c�������ރ(HW�c2QЧT}����BPv�����9�3	���?�;���~��ؗ��67�[���9�,:��v�UN�CRT>8�[lB�f�䖿.t�ǑN��m�C�B��P�1��t:Qcݦ��� o2�\p���fx��С�S�Ψ��Ǆ��/ ����.��&5�0��E�`j��nIN��'���%�h+S�롡'���h,uMǡC6+�j�v%e�������_9tx��!X�7��mܐ0�÷����2�ϡ.D.�Ը�4��1�(��ٜ�a�^�0�[T�[v�Q\bc��F`�C�p۷8X�e�0h��6UOX�Q�3��@-�TV�%��9_\�����zR|k-��d�mѮ@	z<ܺr�
�,5ٕ�񇗖DɄ�z���xAW�}��{���oH����R��*�4I�1��ln>��eY��~�ՠ�'fa[o{���5�;�$�q��]�5ҷ{�ꗚډ9��ݻ��򮦍&t�����^�����s�q�O>��Ν;����?~�Ï?�}ai�x{�~��J�����0n��V��t�0j�h%?5k�2?ȞU-۹�m�E��BCat%)3(��9��S�t��eQ<UX-ў�������W���L����ӗ(356����� <�y���b��d9DW��p L�tG��"��)V2&6B�/��</�B�������������*��D�J��a��~02���@���M��|��W"}S��2*��rh8\��^�?T�)?ĉ T�
_vS�����h�]��e��Q��6hi0�FS�x�����hX@{4Z���Q-���w�s������M��}8T��4�``{F}��K�>OӯY��t��L����O��{aX�Σ���45Ҋ~���뿊B��T��q=:�Xc%��?�x���RQa�M�m<KQ�[[�T��Tv�Ԟ���`�[�¨Ѝ�o�������$�?)<]�Uk�DP�/H�(a���l֢DjUI �R�K��i���?cR�/=�RXG�W�G�!p�&���=r�������!	�z�wj	ck��¾\�v�֭[д-��N'��\���.�-���W�R�hU<�~��pι���?���X1
��'{�N���7�$�:���j�uN*�+WVb���^J ����@��v��e���}�R�
�t�m��:���"4Lj�##���6�q�Q۔�`�o�է�T/'k�z�B@�Q���3���/OAM��T��`?��4��ϟWG��j��L��cv�)y`��_�y����1�x�,n����o�p�qWP��ۻe��aa&����=p4��c�G"2N:	V5ۏ�[�x�,��5@��-�}b�OB�v�i�>߷�kB]Pqdp���}s�1U��cog���b�(�RAgg$/��ECA�7�c#b��,,�:ʒ����>(�PZY�{?!n�*�dj�>+j� ]�qwJ�H�];��L�H�ߤ-��.��;�0HËi&	�0x�(�d�����Q����I9�'K<R��&�G��?��e��32�l&�x��9eil5A�:zi�5�Hhd�u��o�g�6�+�
<V�b�]`��-\ig5�K��G����#,���#TMe��vm��Ќ�QPVv7t[�i
6Kx2����>��#O:��Kˀ�:'��c��'��*5�L�re֏�.�$��F��K�����$�(�ՀD��uܑV��!�J�,�pk��+K�%��nbb=�.�Z�ؚ:z3u�766^՗��̻�M�d�������XjD��ܹsx�hg�T,�Sh��ǎ�5z���\�hޤ0jwL�G�B��c�������<���/�8}:���B�V�n��g���7�ރ��͛7�y��y��x��*�����ַ���/���|�OZ�&�\��=�aX����|^e���"��m�<��n"�ca/�d�'<�!�9��?a�Y�h)-�v1��7��������o�>��{c7��̹�쎿~���kWq�O?��$����8�?�1��X�<)%o�"�0c��
�g�}��믿��K�O�[N?����+�K���I(���6�r� ���rh�'3y��r#�Z�Q�|1��N,��8���7u�̡|����*#�� >������L�^�'?��;�b$Z|<8����ۂ8������?~�����'O���14�,B��o� ���X�?��?y���h�����Գ�
��s�޽{8)R�S�d��)��������ى��҈�b�M!�(\�����A����Ƹ����H) �;�Ne4dޚl�2���gj�>%��CE�ܦ��QE��`�B8�δb�H�b��ɬ�)��� ܨE��W�0G��a���Yb��t���6�uYj�J;�J+�u�����dXi�'_D�\�|5��z��2K�5C|/��������7�|Gy������������c ��+x0��au��2zӼ�� �����|Ї�L�y�;�ꌶ#l!�r_m"OY��mݶf�=���u�,��ip�r�"���6��2���%��f��C��祐��h�Җ�76���d�J�ޖYg<���d�]?zLN�T�%?.5�%�i���6�`;�@��YZ���cq���뿴�|$�Վ��חoo�PgSba�.���j>ZJ����c�ά;#>-��D>=Vm�"�zO��,�f��<��,+R�D�^�鄄GEt6~�ӟ����k>�����6Ц��ʂ8��V.*��������`� =}z�xi�É��I�ˋx�Gx��P��>�#  �뛣'6��<N�(2Vr'?3nS����*�Y�E�TG��6 �є��+���)����mm���/�e^|C�L�����/�Wk�����۰G^����y��"/��:r�����Vz�Z�z��q!���*�:$3��`D�yxc���
�MdL�tL�Y�@�|W�Ux�/�>r�e�b����(��2<��Iü/�6C-�F���������1s4�ق%'�]�Q���ő�?O�-�k�	/�,�ϭ7�`���N��\�ޠOX��@m�F"���F�U�H}�t�kez��{t[�*�t�����3��Һ��K)�t�c��I�lĜ{�����0��s�ɟ��E ^�EEړ�N,�/�ެ؍; �8�9�6l.t���$+�Uա��gݝ�*,ش�2��*Bb��~�`�U���T�����ыv�����̭��W��fd%��C���|xh���r� �z&Z������M��.W��Bk2lR|S=/�YWq���(�:�O�v�̋&7άJ�l%74��\p��H�W�z0���!g^)�T�����$0/�h��"|)�
!����#��=��dg<ϸ	��;�Y�����Y�b_��M�`� �d"m���<��r�����_^���/�B/+|�f[����Y}]5kk��UQ����;�^�[�EK�\�wMD�|���W^IN�=���\���ϵ��D�m���3F �z:�
N�F-�B��'�b�%�㌫�ʩ4I򖑱k�r�JR��+eq�B#v4dY~�$�f�*�ȇ��cGp��:��?{vI�YN%�j"�e��H..�3�E�,I���d㤚OgحP7��L��H�������Bp���3��\To���8�x�PKu�Oe���э�w��q��@j=c�54�Hs���B�RI-���TgES�<�Y#r�R*�B��EŐ��#É$�j�Fؖ�&̧���3k#-���p~�udp��U[ڿ�a�,!(fvN���z*�otv=  :�h#d}��f�9�*!�[­��J���n��9�4�������ज�����G\+�],)~+1������%F���.Tֹz���{]$F�IH�8��¤���i=��&�v
�|��z�k�����Q�����I���ӬH�����6ʛH�<g��++K���Ov���Ǐ��/^ğ>����D�̵�2#����`�����j������%=|�%}gG�@`g�����L+����|o&r[�p5�M�B��B��C�!,��W��ԠkkGhű�k�G2��<���L<�َ@��|��tu���Ұ�ϳA�$u?�3�f��ݻw?��s��*Ĭ��,�-�1b��2b���q����{׮^�t�W^y��7�8thu��	���+��/~r�����`i�D�d. w�m�|�/*����֘HOKԛ밫7o
���ã�%h�DZ6�i���i�y����g��G\�B��7��Z�/7Ex��g�PeyTV�1�F>.���x��3g?��3�F�0s$�Ȫr���ɺ���a�J�8�1�jkU�=�E��=�w�A9��]_�/���!"��to{{���4!<��������=��Cqf��c�X���4i��e;h/D������	�}�e�]H&�YCQ�k�WN?J!a��U������
��y��`>u�ر���b���OO�z�����TC/�(��h��,�}O67-/���CD��-kn߹���5Z�a��x�����^~����wN�>��+$���y�=ޛ�z��d_�`�Ţ�E�Ѱ
���4�_�����k6+����\K����i�V>Q7�GRؔd��s9��n�I�����׿���&�������D�A��KV?�e�'��� (� H��nK0�۷�l>��8u��aVO�AȇQ�_|��W^~�ҥK��;����o}���?���J�OJz <5C5V��dE�D�Y���ƃP)yQiO�b1P�L�X�t���m:��YKĖ��K��C��io<4W]-!΃Z	7�J/���K)1Y<׾č�G-�$�G���D<z�D�������/~){��\�����PXy�o^̒LZM���x1"إ����]hc5{�1q:d�#vЛ�RJ�̨Ĩ+r�X0&j�bF��T0�A�W���i��yߕ��w�,R���ǫ���:�ί=��{�r劎]�ɜ��r�?�ܔ�Ќd�N-gZ���3��7s�f�(�
Tz�3c_*#FP�:���Zg��W�3���ٱ��_$^b#!B�I<���G+�<���P�B�C��uAG�6u��{�iQ��T�d�YvP�d-[��BG��5�js��,y��{�bY&3	��LF֎C7��I2b�1��ZH�����a`�ZĄ\�PV硅�4F����8�c6'&ٖ���� ���T�E\�(u��O
�+�oi���[���E=.�8�x�;�M�i$��|�HJ��͇�M���������L��e3V�a֣�@d�?O��V5����*4˨���ʭæ"��B:l���Q-\�K$���	YC���7J�Z��X��}[S�W�Gp���6�+*w_CA�vvb���h󠚞�W�QwW��Qxq�v�Q/]��2`!�rwz�DM���9t|
�a�j���o��?�@���>�L�  sZ�H!M���/=���dF�H�n6���lK����MM�/�X���+��҈������;��Ҝq�
��m"�\�`�+��j4JH�?7�x
-4f�ݹ���NX��E���Wm�(�D�ٯ��w� /�Y��3�;���*�X�)!B�m$���YFe
�L�`�&
�ò�Eg��"�^����=<1��X��*�D�fQ�EA�Q�3O.�2�2N�?)�H*�?�YB��BU
~Ϥ1J��@�*������]�S5�|a�x���>�������[���ݺu�ڍ�u��$F���}���`4����T�9����p4%/�0؈s���d㥮���iy���G�;!tN	d,���#P^�l�y0&����"��������*x�;��R�8�H-�h�<^9����&U��Xs�w�8��ƉI��m�.��q.�E�~�>�#�=<j�*�NjR�)�T$���V5�<c�,7�)K8�$n�B�T� 9�B����ݻs��͛7�^�%#�"3y�Kmhİ/v�F�Gu��fok��J��K�4a�0,em:���Jx�u���.���!�S��vf,�j^VP5�C����;��Rۤ=�o:��&�qĲ|��:����+^�L�n
R"�EK��j���^�4��`M-�C#��lVlԙ��-�7j���_�i��1&[0� ��u�Ȥ�r�=x{����}͓FO�H1��� �<y	= f3j��:c�y�<5�y�����8�,h��CI������ߨYd
��kU���D���z�l8��u��Y�<ok6�p�%K69� ��I�qK$8�F�.�?���EtA�6��6Fp��*�~jw_��8�3f���*~���������YtzT}A�k��6�p�:�k�2#YsP?��+��~e*�@ţ+��r��%�l�5#%����I���nD��q�*�t:�s����؆��ۂq:PI�ì�Jln�����ȂM��ә,W��Y�;��xwyӡ��[��F�\�4fI!�߸�f�
^ORUFV����KeT����o��~���nֶ�'�Ν;�O��������\C��9���!���}z]�Ս�V9���+����f�F���Zz?��Yaε"�-:���"s��P������9�xrwr��F�f��q�(�D�D=~Oٴ�.ۣt������կ~��=��ی��!�!FԬs��?���JIC�x��7�z�\�'O�z��s�ҥFK�y�)3t権X�Yk��r�ӿT�fa�y��k- ?u�y�L۷'2���t��ҫ?��nݼ=��*��*` �׉��%⨗X��-�Il��"��X1�I�|���[�|l�NG�L1\	��ݻw��YؗJ���;2n
�9B%��J��&,"�Z���46}�Ƞ �*��)�[s����c�6����1��-hq���O(��z���ȑ#��#��` �yF���&O�Y�mO��?��������~���s/^�����cǎ�����t�1"���{�z饗8��E��X"([�l>�N��`<#Y��	�W�]��5�>ʁ 9͌��C��tJ��/ϟ?�M�2ҀL#�3���+7�Qi�U��"��jl7�s?�N��5qF.\��}��uA� $������E�!�����K*��6ר�2g/�w�� 5��x��gV_��*/�`��c��O*c>�l��[p��E�&��ѣG������S$��h#Z�`��
���m���P��Vt��!�G�5V��!�;^�@��o���쾉��!_<��+�����������q�A�Ъ��M�l�4-��ũ����j���Y�� &����0	7�'�5�`�y�5�V;���f.����E��=w����Ƌ643��LS�����R*���q���;�X�����^��&KΦ�h��-�W�N�7�ı,�sV�Z��0i>/���Q2)Eb%�/�z���`3(���9��]�ol�s��Ŕd���ݝC� �e0dg���>x[I(�����h{e�W�y��^\ ���J������;�v4h=�w�◅M�p��bT$��U!v � -cl��M�y1��J�p2
?�E�!4��}X2Ez0�z�D�L|O#@�̌ ��:���v�Eia�������.�ё�p���'�jtj ��y�($�ոFP3�L�d��>���񶃵�Lf��&�1���J:������?tU���!�V>[m#O(ɂIAN���g���'%��ϫ��i~)��`v �`f���7����~����<�|�Ly�K�ݬ�W�Z`���S+]u�xR]�c#����Sm�J��WV3�]0x�uܸ,i�Ԉ)fJD֎s]X��i�x�F��؇W+�<a<���ޖ�k��w�s�!�l��Y)ٳ��~p�a՚s���7I��"XEe4�T6����F��ף����;���1�CD�)�RV֑�{���u�#��>��Q^�~�����������{�e����]��Ս�'M6���,RBGn���E� ���P��Y�ZUu�s��[e��&{����v�ٿ(�����dw�l1'�N.��pu`cA`An*��&A���a�|��\ӨQɆ<9\�������E�^�Xѷ�/�}l�Yw_}u�V䄤Ya5������u㞁����꩑��g�k��w���J:҄Q���4�%͉�n�hg�J�Wh�B�7C�V�eu�B��z��u8�ء�l��pI"�����>��@a=���pd'�S7ե0&.�f�R����rI�,KrĆ�r!���߶_���,Y;G�'[�
N���-^�������d�a���L���cB!��c�v%��L��+�/żYl���$\#G`L�X��Z�v�k�UҺKA�F�����u�.���s��X�x�Y&��%F��Q1�s?��Cw�i��#[i%�("�������f6����R���WDF�^Kfi��5�mRcEj^ZA��F1��i���f}ĝj���:^4x�(u_�]u"[��`�E|RFP��i��%���<��p�,n˕3w�Pq{ ��rm���7)�(r�D�V/$WK+�ֽҚD:�I�\/��9�Ǆ,#)��`��F�p��6N�D�;w� ��q���Y�[���ܾ'N<z�xt0��V��*{����,QF�ɑ���	l%Su�,L��4&�xa���z�^L��8�0� w��[���g6eE�)=�&g%�v�5�y���_]J�p��a��U��"��5w��$͜�~X�/l�p4�x��h0D�zA[��ʃ�x�����4�8M�B� �t���~��ɓ'��믿>ѦZ!��:�͵V�����GeCJ�:���ǻ{�|�2�F��1V�ҳ����)�]�ȝd�[��B@C|X��o޼�/*1��d�g��w��]>WB����Z9`ʖ�nb��G	�^�����k�MՄ,4�Ɯ_Zi��D������x�OkKv0����.},���X��^T�Ϣ�O1���P��;׀
O�����E=��o~s�葷�z븾�u��h��U����~[�B�{`�/�VD@xD��J�T?]pn�o�(��k�C<uC���Q�>f��Nv瘪�Ir�����?��֖t~��Mh�o�H���'�����M���+�+�	�4�8���?��׿�?A���G?J�%��S^6���,����ep�q���gV<)B����g2�Ne�c�h,��?�E�:�ݡ$qc<&Tk,TT�9w��N��o�&p�J�ٳg�8Z:���8Ԯ�e{��G�^(*]����1l�~����|F"z�^x`�+m��؆Yw^��>���L|��d�<���������u2�"Dw�d8��Lz��	�FF����C��!}y���Q�ĦFĖ[��?�csԄݠ"�֧��_�w\�(<��`�^�iT�X���$��X��(�u"g�ѽ�?�'�z�M�~Nړ�(���a?����G���b�t�ݗ�*E6,� Q�a�c���o/��V�7�t�<�4�.]�˛�w�R���?N��>�2�7Y�#E�1Fow�\��p��iǖv蟫��J>jY]a�At�u���!����"�^./�XWտ�=��|½}m��e���c����5�Y�ӽ�>�7-*��M��vdV�Y���i&zjƴ�Kl�/?�s-��n%\��BJ1��Ζ��P�j°�	g�s�3��~7�4F�B�Wƫ��/*��"EGEU�j�T���b�=ʪL��4��;x���mj�A����	��"{Q��^�2v�8�)=�k3���7n�7@^?��I��P��k5)��pLw|�(�D��9|x�8�O����	�+�l$ �%��Z�D�2�PZ:�6xjx�	g�>I��sxb�&�bR�p��P����	r#�c����KE���O�G�֩%���orex�q��a:i��H:��+�����U����$ƥ���Z��=�:��)8���U\��2��7<�v%@UL?�%��!c��c+��_�/���mQ����pd�oܽ'�cN��{����7���5�P8�/��,f� |M5_���v��;O>�qE���Vu�dr/�+K�Ъ�x6�ѠЙ���#kt�6Յ�T�i���/���T�v��
�۷o3ÝX�~�sEʌ�Ԡ(����Mɯ��/�U��G��
��z�Z+��;=e�?��UP�>��4��q�H]Q(;Yܩ\�>����WD�4����2�?��^��h�X��oCql� ��:t�T�lq���m���B!n\W��j)��6��R,�G>��h�"/���p�8�������wgOgY�E�H�1؛Ʀ��s�F�
9ݨ��}��_|���{��)���+W�((.�<�--��!l���l�rQ�=�r�����h����F!�6֋�hM��J�F���O�����B�DbDy"kdp35
��F��� ;u��C�ژ�Iȏ4^i��ڵk��T��a����R��_�ˠ��QBD���Xi"L;T�~~hC	y�"��旺k[>VU�œt���ŧc-�4ҚL}C��m=���'��E��-���f�C�vp����]QTj-J�8<h��7�w}��J��D�Xޖ���1���/B+�8O��v��zώH����$\�(��VdP#�Z��hqv��?��Y
9�t�͉T X.����[- 5�ΊP�'l�������2�ÇmZֆ�/凬��cU�+��3���	���� ;(�&q.���#�Ӻ3�E(������o	���Xy?O5#԰0���7ך�e�p@T<����Rd��<s�öE�Қ�,��K;6��O�v
�ҥ[�w�$��LO:U���(�j��Y�C���4]g��Ё҅*U�ѥK�����:$?���F�,��AF��@� �=���dp��'7����q��@�oỠ�����!֓7���*�~�wC++s�P��"���d��˼�̦�Ueխ�=�E�'NLu���g�)7�nܸA(J���=�]j.�\��!�|��ɓ'7��V�@%:/�t�R!�0�,�����9<���5��7�`�*\7V:F�w�!>E� �&��#� ����h*�`c�*����֏�|X����?�4vא����U!��W�]�~I��N��W���=/mg��+Έ�Zkw���(i�8�������������Ck�Ν�r��G}D$�V��qo0t��	��H��Q��f�z��}O�{�
�%��3�qc�Ǉ�`�Y;� 9�W7 kl�B�)��qc��w�֟��
6��Ȭ���`_
?�̕�KW����Ǐ/��rf�~��<�Y6�!:*,��>=S%5��+,��R�j��CZ=��:�����ۿ��?��?�S���կ~E]A����M�3D�{�X�d�8��Hz�d��\��-��ڳ�=s���Ti����LV)K���-��VKK��u
��2��ߨ���rm�j��y�2+j#f���C���QlE �q5�kY�̗c��̫{��q�8DEy�Vn���V��^��(�=
s�4���jU��խ�SOA�Lyis}�X�!�g�q)Љ�j�7���,�Z�]�Qr�ׯ��%�a2�(;%�<��9�ޅ���a�g�G;m��\swC��?C��N+Fdui��M�N�2G�^�H�Z�sl�%�r��J��V�[[
�YMWi��ե!fM����%I�i�+C��X��
tg,(�����[�=n��6vY�J�J���處�sM>Đ�f��2�d� oX��g#�h�%Zvʤ���u��3G�y�����!ӈP��F��95Lcu���b��'���q�3X��Re�h�hf�Ur�J�>L$'���vm%x~(�:D�����$�N:��L�pݸ��0�X��m�tu�;	K�Ŏ�˭1����sC'l�l�$qI&�f�x��׹z׿�LM��I`��^ET�	�\�8�9�TZ�@d�:�R\rx�^2➀C��7;x�,�:��ݓ��޳����^	�G��Jze��#E��v1�>�=)�����o666`�����>�B�ꫯ�:��&��)���(�3}���BJUzʅ�k���Dq�2"t�������<By0]6��0}G��;r��TA�π+lo�+��u��F}a�&u{4=2�e��FH:�7V�G�]2=��:�����J��W��K�H B��X����ڒ�8��U��iE�u��RWh<�!J�.El�+?2��]rm%K-�=�&j���)Yb�	N��x�uw&��3����x?V���a��GgFK��R�)kْ$�Υ�1I�u�Tu�!��$.���ިnҼ�^?���x�,�Wa�vv�[[�������7��*���`��aQ�G�2��,�n�yD��+\��ѕ��T��L��3��+��w�<�֦�
�X;�wfC���=��#ʭ_ؤ���Dk�p�>/u��ı3��T��A`�v+�=�:{{c��<++˞�I�����Md%�4��ٮBgCV��v�4�R:�Z�;��%eҿяhdw؁�z{y
��q�&(�����A��r��MZ�	�E;˵��Ȱ�� �N��pq�i6�1\��HoqK��*7��m�{v����(7<�oSe�}~���b<,""\ zp{k����mUd�8L��c�*� W���X��am��Ϭ��%�ݾ}���I8��,ɂOד���-��<�*7�~�;%��|����=���%lO�l�����j1Ԅ��l�M��fnM�Bjj,��G��`��ґ�w�Vja�e�w�wN8�#�-�k��AoЇV-ꪞ���e�
k2��:9Y�r�d�gΜ�O#��DP�8I����ż�z����ĉd��VL;�}�s��v:\r���l$6�=�Xd&�v�R򤳩�s�F�����|@"|h��)
d$�Y��y��;i�*��:��]�mgְ?�����<�ҫ�;qb�%���۪5}�9�AebLV���+���� Xu�9K�jT�Vd��l��Eۇ�V���$��b�!�P��ʦ�L�?�im,��¯��� �M�����lɗ $OtǪ{����>�܅g��qeuY��9"&|�bV�)=Š ��*�nkuܧ��mZN������� ���������mi�	�S�jT�C��R�O��5]ZZ	M\.)<)�DQ�d��|Gzx}�*}�pE���L�����
q���?}Z�ww���)LҮ�P,��<�o��]�-��t7�*�f�����s/�+�ܹC���<���Um�3�(��ۡ�̘���Ny ��2��S�e�V��z��I�2TU�B�ޥ6�ka���|||��jRXs�/�T��1i�[����=D�F��nd�����,�����{x�n�9�t�9�Xϗ�
u`���_�����[0,� �т��-�_�.
.��_�����������Ç�z5:u8��67�k��{����g���H��U��F���r����������ӳ#�#(����f���{���s�8�g��?7n�nR$1b���6���ɱ'R��F�Ɛ5�+�Y(__L|I�f���Ӌٜ����;;8�'1�f�} �d��R��%��l��sa>�e�+��{�E�a�Iw�	�:j�%�Cӈx��Pc��;O~ǆuV�O�]��Z61��S`���;�:��O�[�>��z\��Z{�J���4�v1Z��j��QCP�L�N��#�M���=��%�A"�A=H�rw.�UQ����F�DWb�q�Z~��w|3�b%���=��zh���u����*N#����:�R��=Fsr�4x+�Nab,��(���]��@�1v�61,:����Ȭ������c+�h�;#Q�l��zqx低2�urj=������FN�X�9�jN��m�	�"�A���x�g��;���!����(%o����%V&�a���;�|(�l��-,-ڎ�q���p�#��Ҳ�hlYv S4F� /�Ö<K�_�(g�T=�Ѫ��5x?�x��<J��.���ٗW����Uw⤑/�j�˪�'���Be
F3 �WT�8���v.����Q��Zz��ھ��qD)�r�սT�c�ʆ�����D��gX��?�X�G�xÑ���k��ܧ�:yv7�lv�W�Ɍ�Bb�CK#a�[L�I8<���+G���̙͚b1��K��h��|ڇO�O�@�̧H{��J�L99s��X`�ؚ4���U���ׯ?�����&�	n�4����	R��k{wgk��x*�[t�A_����*�+��Zc�4�31R�R]���ôa��x�ߙ�.x���]3!���DR�2n׽�A0��Aj��43�8��0���r��h�\�gJ���w�sVB:=4�Uy0��4�j�O�N�Z�����"���"�������:�R��E���5:����D	�P���a!�1��O$��+����w��O��}�3ayyP�TY�I�J�a�V��;E|���h��Hm��ŝ�`���J�"˟g����8ZY~aw�b��Y�c�B$T�,=@@}
EFe�ֽ.�_Sk?,m���2����سg�ѽ��dz}O�0<p�#�$7r� ����YH�칶߸3O=X��(��F��r����(o#�b��
�#a�g�5y'���r�yeG�<l6)�=Q"t���[���R�oљ#�;�L���,�'���ۉڦ[m	����d��l�3��?����[���!=P�<qƓ�-;,��B�1�;f���K!��Z-#z�xM��E���r+�3����u؃�:m0��*�+m7�p���(�Zz.`j���Ό�x��\�[R�ҁpW'@�@�e�V�#�Hp�nqe5 �&��(��\�C�)2����pL��]S��%Q�Y������mS8����,��-�h��)ri�h����G=��y��$8_�d���L��e���~6s#���Wej\���Z�I\#�ƥO�RG�H��ٳ��E?���{�\��\�r�Ν�gN�T�*D�c�|�p0��a��w+UWV^{�^z���s��D��oݺu��-8�[����[�Z�ڳ/�[f�k׮=��s�հlo�1u�BYp:E,�Գg9�@��n�ʔ�ejIB�~��c�-c�_c�<wn�yq�_|�Q<�8Џ�b_y�u��Qc��:
��s:�N�/�,��q�n't�w��guT�䁡����'�,z�=�QΩ<����s*wb}��)���d�깶����5����h*�ܚ^�P�e����ƍ�(Z�d��ۦ3��������+�ƍGO=��By�RMA��򗿄19�d7W�^�t�4>uE��`y}���P��n|.7@~B�CH��h���x�i#��Q��K�^ZdnGl�v�b���	�\ƺ�+�$^v�nzf�3j��-��X.�<�\��8����չa�m�j�'☾^y問?��VSFz����4�Zw�<�ƥƧ>��؅�'OrtR�zzz�*�"뾤�P�+��f/h2 i�LPY��@��Y#��o��l
�l֪�3�.%��l��7�z���5&�1*���-o�ꋭh�O��T�}6�j���ﳄӃC~E�h�C.nY���y}����jO\]ǝ�%�Č{�v�5��A�����PZ�fc�t����΍`'5�J��V��V��t��ga-M����:+�r��v�R�ڰ����5K��)"#�ԫ�Hӝ�P�aJH����r0�m���W&g��xM�:<�ܬ�S�:l<<����%�$�SY:�=^�v^pD�*����C�kCo��reH�������ŕI�,$���C���]_+}��,=���m����S��l�	�I�91�ڻ�zƃ5$y\PvJ�tU�*
�p���r�p����x^9�:w��W���#t�U������B%��'0��x4�~�b-qJ�ƙ���GF�S;�ګ1���ɿz�*2���n$莜�~pa�Cc�r�h���{��x��G%�.��R�bk�ʹ�e��G��/�w��_�x�Q�QjS#\S��3G2uҌ�)>��
�OPڈ�@��KZ������@JKm՗~��C?��~�/�Q'���b);C#ʯ�z���� e6ޝa�7#�Oɨ��C��m,7�ӟ�1ac/��-CgS,f�U����)��r�TLS��+W�z�o�	��	4�1zX������-N���/Dl]
�hij���f�����H�i���qG�@��'7đ#o��G�����p(cǼ�V�V�稚�`�AR��	́}���o,`Q_�Z$�K%|C�/ZK,�c��������Tf�Fk���ԕ���.ʮ���D@僱����e�⑫U�-�Xw*�F'|h�0]���d_Ɠ���Dʶ�zs{���4$�0���Y�+�h1]�K��&j&S8j����w��	7U2�u��D%���U-��!,����
m�gn�x*�}�Ј(8�C��/d��$ :IZD�ǎ�W�\�G��%Z�:�u=㪨��Ž
o����١�1�������;lw9���A���H�YcG��&:�	�?,--�S�
�n�|Q��u'-�Y�`��`0��x�)��q+�;o���&����A����wwbcz����]s�[B�~��?����KVv������:}������k���{��P�9��tKa_��(h�B�:7$ŢL�8u�vADO��I<�>���n����h��%��ͳN���ř>f�Ix���{���3����J�˶z�����y�9�~0>�C�]�x����Īe��Pd	$v�kR�M)��*�S�^Z�'��v���N�	�%�3!xR|���TY��a��w:4���oX���F��N7��{�������,�lV�j�+�U�NU�q�x��e��ʗ�Hq������F���<Ɵ��[�@ �K������O��lo�>~�E'
k���~��7��罿��Ʋ��xêS������v��ܺ���{��^�*U[M4��׎&qV@�6"ò�R�̈́Y�A�A�m��~~P�~����˝�$R����w�F'N��J?s������{ｦ�ga1�[��M����Ν���勪��^���Ԯ�זss���.���1�#��y��>�������8r�v�>������;ۻǎo0��T5�8��-%t�3gN�:����iY��jͪ�mcd��f��n��H��Ubџ�S��́�@Q�sւ�R_V�WW�^�{��/>��+�	�9����xA�K�	���x0p��|Y��7|������߼y�'�Qˠ���L�0,���Ҕ3{��?p��� ���o=�.+�#�An\Q��gp�A��fq�h�Teղ.�9ɦS���˳�b	�ba���A�C\3���=Dm���F��˗/���V�������������g��.�1Ӽ��	�AE��#.~d�q���dY��f��L x��:� zn����/��0%O����+J�t����ɓ�NA���1R��e2R��FӢ N�m����,���ƍ4|��u�:��??�]��Wd}[
���w���������8J�Mi���3�x��F��+;�����3���w�%��G0P���7R2{��l�c�A����-������p��q����0�ѕ�+�P'V��t�s��j�x�_�G��wZ�(Օ�]��~���JG6�2�,�dwUL�����x�A�v�8��=�扅YF2���-j ���׹�6RV��D�4����XY�i�NR*�q�˔-V��A���,� I��@"� ��O��i�@3U��;B$����n���Y��íT�g�
uP
@�Vj���$�j���<��2<�z:iKDs#����J��!�6mt&7�6����ʉ�Ep>c���$��&�
X@:c^JVXS6�|	S����%2�߳�t#�suQ�.se0D��h:B�rE�Hޛ�Gp[�+��v8��H�]���&�ߊ5O��m�O�*g"���9_�}��������x}��F�6���P�L�N��D���W�pi��N�r"&�I��> ����!6z����S+�h�~���Fkz\�v&$Z#�1�#��U�9�����#Y��b��ɭn$�g�QNˤ3�a�k��Z&y����|D3��Um�ݸ1*l("��ΘB�$��<|��aQʺ}���l�81�{�1/�;ޏ����T��)��&�C���8Z����FdE��/���Sx��5��Q���� �E*�(x���4e�{@I(�چ�>$O}Դ�)��V�<�zU����>���i"	��`���q�jh���]9ԛ�w�P�oo�� . ;�a:���`mp�4��x4�r�G�w��.��h���4ˡ�Jh��.���d� <�U��b����m�tʝ]�g��x��!�����}�.H3�k�����r�L�5�7��L��+�#W-*ׄ�c�w2�����gj�<67\<��p���b�<5����n�U,�����a�W��G�/� ch�N]=9L�s�:2�C�܂Җ01�r���U�Of:Tޏk��)�k���LB,�_M�?SZ4(gJ-$��/"	ſ������`#���y�g�L0�-=�=B�0{�`�&��zt�����>n:�6rx��s�\�y�W�5���#Xy�c�����LR�a降o,�F܄y��8�D��uvk3�/=i�\���k�;�W�k�s�bV�U��ț�,tV���7zK�7�����kt���N��1�6�b4M'U�!�m*�CbC�ee���\f�}���<��h��Cj+�t��� B�YIٙg��Wקuj�Im�\��:����ͻ*p��gݑ��J)�7E����߮��h�:����m��6�(�h���&�3S��"�2>�g_�#��`8u��V<x�jA��.\���/Y ��.���+k����Ch���3���a��;e�=@�\%鯆Á���v-���*c�Q���<�j��x�w�w���"�Rg��&c/:K���˱��݃�����U9���������_��_���;Pt�d1<|�0%meeUKџN˷�~,�+<��>k
\��
�ظC����j���g��>c{Kfa��gw��������l�����Ш�=����:3����_|Q��.S��� �+���K/�aq*�4�^x����g�/I�ߓF�FRǸa�҇�� ���q����r��Y:\^=}�4+pcC�r�'�`b�vĴ��T�mQ�h�U\�	��#�|��(�I�!��6�2�!ܕB{"q�k��X�/��B�p%냍;~�8�O��������qeb^�w�U��+W�I*��D��X*�
_{�[O�r.@�2x��b��]�������:�eY�t�Nzc��p��~�#E=ωr��$%ׯ_�𦨰_�Ib�˹�i����j�oss��O>�{�.�j��Q�¸�����{߻v��5y�ĳ���oS���x��؋�0i|���搔S�<����y���/��[��)�
�KٌF9t��=�ԉ'^y��'�c	A!�J��g(��6��1*Tz{eg'z�/��2(��1gϦ��'Sڨ+F�ВrY3��v�m3��}|��e��цP�h�y6�P��i2M3�|�n8�����vWm�w�᥈,�ӂ�%�zbUZ����ܫ�:�P�@�{�*rh 3.�m�����}Nb:0�:w[L4�N���~)K-�T�L���I��Ĳ��BT-v�ӌU҄9���X��̱U��Ѡ���Pi6M����="�r)�\h:i���9�c���
2�ċ�:�hq|}�6O��B��~Vo5V��r����ӵ��o�1��j�~�:���'3��fŢ�&�v{���[v���Sm�9i���y$g�E�I$���ϔ�S\Y�Cl�%M@d`�.b�&�#J�_���B��)���z��J�:.��N��6v##�\?�q�k��s/���I��Z�� �R��$�q�A�8�����X���"�\�u����l�eZv��r�jE'yH+�&\� �Ż����z{=���~q�"cp�_-@j=L����u��m�cc��U��E\�k�n�˫h�JmLSl/�xez,M�K �B6��z(���k-X�\�mf�Z�ڨܼ���z�v��J�~M<� � ���٘e:��s�*�߫��H��N2��Ԙ"\Q�F�E�f�ʹ�e����F���a��Z����@Pl��Ce��2	����̚Z���v{/yi�����lq%"�N삔[I-���^�����|��dG��I'D\�]x��zh)�JXJ��ÇJ	5$M�)��F5�Jɗ��*��l�k/8��F!o�(8�H4_.F���<^�7����)?nR���e:\���rٴmI�t�:S86�7ѽ�^vP�wJ�Τ��8����A��d�"2�6u��
�?T�k؆C���G��"�㡻���A���-ia�Y���v(gm���W�ʑ����+�i�a���J�u��ݽ�
k�O�{��j��1��������d�	�e<�s?I��9�XmYh�&DjM��#�C�gQ����)�P��4��C�v��:p��n���<xP���E{Yu�]wK����!��_�	�\F�\�ƌ1gkcc�(�8��h��ߢ�|���U[�iV|ãT͙Q*��v"2��g��|���R�m\b}+u�j�Yc3�M�V M��j)�K~�¦0;wFm]ϕ��:2���z:�>�!t�v����w�K�-��m���L�K���O�[��X�nȸ_e�����l��q	 �;n
��EpϾ��u��q[>�Sb��U�MQ�{Y���'��<,l���=�u(c��
_�gPZ�$]�ں�*�=��_R�1��s���I���ʣ�g�m]*a��tD7d���p~/_����~���.��?�s�`O���Sk��Yj3|ԫh5x���'O�|��9^�Mp^f�z�b�`@��s��8�4X�Ej\��}�`,O鋎��[��߿O�J��默�g�E�g�>�\�Or��Z���?��=.���݇_|��{����}�Β���M<��겺���ˢ�^o0���i]�~���c�+W/\��/Ub�HI��S��,3�'��c�݀�g��>��� 0�v��n޸-MIQ�<\ae�T��VkL	��|����7����?����<~�8\�<I�&�l�=�n�'�	݁���q|�ڋ�]��ލ���^{��~�����C�V��B�(�T���e�p�����9	x�իW��'��(o��R�ОR��{�8(�������H���>�nN���m�}�p&m�o�ll�_xa�(!��A_���A/_��U��O?�DR_b���D���vMb\Z4d���!ZLD����
�l����!�B:���TS3S�5cҚ9��e}}7��B,mq^����s���B-��@B��./��bB�S�+#l������G��<uN���]M���L6l^�yT)Z<�{�.��S��Ν;���/q�VVW�]H�����b=�,�.]:z��4�A��Im��6$'���X��ZY�O�5���5������Gd�A�ecz �vn(*~�4U���m�S�����F�M������G��Z�Z%�������LJϡ��n����pk����6X�:�7/��ޖ��ӶǄ��Fl#	��My���y���H��c�16:�	�|:U,Qd��iD��m���O�5�9@�[�~9"F�B�.��zJTP4-~�&�+v=la��;,�ML��9s���!X)!T_�UG�F�N�!Ot�����DED�]s�amc�~�i�n@��|���B,����6��;RX�2��~Bb��D�+i0J)"�y�$D�0Fa��r���X/�ۀ��5)N��A��
���1�I��jJ�R�ǧ�hڟ���z��*�0������Z�%S�Uǟ(�p�ø�J�)��tߒv�B=�Hmܮc��TcӇa�)��o[�j�T�c6�3WA߉��M'��*�"��v�]9�^w�GJ)��~���fIJWPP��N������љa8�b�ZĲ!<;Qz��r�^M�'��N�AJfu��QZImr/�*sSH^)3Ǒ��*z�� �A�	���R��α`G[x��Aٳi6~O3DV��s��@��Jm�D�������zzy��ٔ:~�'�xO�FY��(�$ �djj-�]ئsN������ߕab5���A�֊,GB��cb��b�#<�q4^/�GU8��Ρ�Sd�q����ƚ�K�qUC�8�8Ş$6��_�~1U\�b���"�dmxw�a���Z�)���ɬ�^(�9h	1���QUczGWC��7��u]�"��2��r���q�!�#a����`�q�q�Ac4�xG���[,�RB���΢:�+�w=��w>��E1=�z�ƍ���꡵����l������l2>sv��KIʑ���f��o�>2:�,�'ژ<Z;��C_eK+�&�p{�*�'YGY�8��'�b�[�{���z2i��6+$�U�9�PǏ��P���>~T5�B̈�t6'扉��$�����GC�Xa��aK=`$;a]h�;�"����8�Qa�����2�x�#C�S+�vJ��;�G�An�D~LGg����Ti��&�Q���s�t�a������or��F�ό������Xl%���K��6q�K�`a��4�!�=,w�Za}�4�Q���m�G���5��sV��[C*xH�QIy=��<d�x&�1������:���|�x1���F�t:)�C�F��kU�S܈����N{-��n� ����B'��X�ѥ�jyb���Dza���eVI[��;�i�k�2B.l4�wqba�]�ϕ��{�7��6���+��j�:kK���h#Ş�H�&B�\7K��+Q b�U�Rн���k�t�u4��wU�$�˪U��U��!�2�f��j�j��h,U����V"�Q��֟R��\����@g�н��Tlt��U��#O?՟�6�#�.��ɧN`�/Kb�Jy��9��%Y��������޿{WPQ���C5V�Ž3���K���Ǔ9r���A�p��Z��K�Xm-	D�XG��K���]�`d�|�≮]�v��ϴ1��1��sf�xg[w�>u�)=cсV��I��`����<�����/^��w��������ץ�mkkG���bdFQN"�A��W%��&b���_�p�;j�F�J�ʰb(���T�-�CFD�57�������e^B˅[:}�4n��W_��:��T�r6��-����m�3����.]��_y��p�w�� o���vS�zR:��tU��4t�)�*'�%iL�E'@༅7oCljk�H��Ƀ�kTi�=x�y��tD�Gߺu��e��yNY����O�8��[o������?�_��o�ăg�T�oߦ�:��Ǣ�V�߿,JQ�D�ۃ�h"+�ϔ[[p��]��i�>�T�ʸ�*�0����@P��0�q'���\�d����n�n�h���]p���Pi�6�R���2]z�����pe��y�m,�x6ƿ�}�~�>ߟk�"�����/_��{��{�՜J���In8�7h�2��>|H4��M� ��XPe�a��t�hy+�:d����r��I��ʁ$�
�{�I���^AiyG����b�^
�W�N<53��,��M	}EbJc����� 47@i��0�2�x�LK����Z�Q�>*�*��5���P�g�7F̮6��$��eg�&��X8`؃�v���z&�*������������N����>W���Q֝y�qnP�N���*����������7k����t���g� �8J�(R�T��ڲ����g�~�]�~ptG�;:��Z.�-�eQ� �#@L�$����g�o�o���"�y�������� ���G2�!n��;���&!O��Y�7�J[YW�o������SD6^ٝ��f���2g���S�0,���RN�F��aH�=,Yi3Zrrq�N/ݏ�@*$��vW�����BQM�'c�|j�>��f�0���>�!m-���0�f��  Z�Zl�`|������قr��Ϟ=��p�o޼	�Ƭ}e'<��v�r�֪I[S�d���;�n��s2ĭ��ͦ{ex*=*%�O_�*���d6��������a,鸴0W�� �y(�N��c�E�ȣ�G^?�ǞԐ3#%к`N53(	�V֡򉭩(d��aZ�+y>�G�M1N�Dm\�o,��hIKZ�Wk+7bјΥ���#�=���Nkk!�Hd�^ǩjS�����������t��'�n����:�!H��f��X7�~?~�Qc�&��5J��]7��oj��p�8e����=
NP�<_�V�WO��Y��!�,Gq�ޑ�"s#� ��k5���h�Q��=���[�g���&�"�{�Ɩ�ˌa�s;��x\6�~"� 黐X��j�Q��ݽ�ee�4c��%��M��ٳ�)���Ç��,/8�L��/ʧ�V>uꔞA$�&�8�.�x��|�҂��<yr��˨!�����YiǏTF���[�V�!�66����xz�J�p]��W��n߾����
����R�˼v�b7����"��#���[d|��ָ2�f�l K��Ea�nuڢ�6��S�Vԁ%63R�fR��Cg0�ܠ��%�}�@�����ϛ���DCe�㮲0қw���4,�D�Wm�5zZy�8iN>Չ�u$�v��A��]A��(k���t6)w ݹÏ�1ۭv�C�d��	)�?�d&G�Pi���1�裢N����򈂾��Cݍ��r���+
y��/�6�epe��_�w�U��fQ�FN}����"n���d�,�麛����Eds�y��V�\��Q<t��*��am��ҧ����n*
c~�5��/���VF��գ�P.6�qa`���Mf�2�������UB"����*���*��<�K|�qxQ��F)��g�WZ!1��� ��MZV�"\y�F��*�����nE�C����-��$sv����������4lof��軃��̸����8�-M��FaHY֠@�M��ֲ�B1�-N���3���	j.>�c�L�R�M5�����.,�ό,_Dj?fL._���k�a�^|��J	><OYδ|v�Il��8 ]C1���6d<��&N�겓���,�T��8���I�eQ1�<�s����Çx(�VWW�_tn�T��(�=�
تw�
�~�"$���h���N�8u���;w6��p1��G���������#���P��?���o����3��
����H���W7���V[t&���:��e���H9���<+�me�-s���9Kˋ�9s���Õ�؄,��Y���t��_�哏>>v���o���07OB��w��uJ�f�1��
��C�icc��_�y�,n���Vڃ�,f2��������ͧ����ѣ���}<�x��)Y���n�����j�5x���Ě �`/��aX
�� ��Y���۰϶�B?(�!�).R]^�<�x��Ҿ��nm}N5��V��<r���܂�>%��̏~��^�Ê0ߌ@���c�[<��'=z��'�L�V)��q"�㰲�����K~I�Z��,|.��&}U�h (��q����2x0�'�.�n,܂xv1�Y{n�� ��*$���VE҈�b ��qD��c'�4�N�i"*|�H.+/�0�d��wE�alH��]�y�VR'ҫ"�=����_��_@og��� �����dm��.�hg0�̩H��a�¸kD�іQ,M���Z��:��xd���!
ko� �]s��x��u�If,Q�;Oҵ���c�ic��C	�'�73T���)%�Q	�Q��� EoA'�9��q�ga���'ƞ��d���ܿ��ebc�:�v� Ŗ��H�В�ƈe�Y�b*�t���M������f�Kk����*��Iw���%�a����|D�'V�ߛ5X&<�w��o����櫸��D��񼿛�{f�Jk�K���lt�z��G�J�:�����Ye�	�\s�w���^�)	h*�.�xT�Q��l%iUd�
��ϲLQ5�0���d$�܎�uB*W��4��e$�s�][�nh%tP�D��2�:o��iU-����yf�q��aI\��ye�O��
�E�pxȇ�)a|O�8�X�_��_N������׾���_|���}���~y�$~��d}��t<b)�$�Χ�z:��mm,:���C~�qs#4��5����nZy��(�����u:ӱH��i
���)*T¾ű7k����`]}��J����e:�����+��0ӹ�����/��šC�朧t�\)�]��[<|� >n��K���u�P��6_[�yuEEZ5��b�j��\�ras,���\V�����<��
_C�]lMܩ�pq�FS�Ԧ}R)QVۊV��V�v\CD���,�{,Ѻ���I�����!aЊ�RFJ�W�j�|����N�׵0���@�����A_� O��dȖM@b���nOP$����Y?=46=te��Wh�hn�(�nJ�2�Mb%:���7V���&�Ip�=���qU�GJ=8r�t	I��"�j�K��.�̓�)�Ȱ��%��]X�4��M����_�"�����sW����=�'��p��^x��ʊR�(�?WN�����<�F�C;|� V�,H��~�B���-⫇;Oewڂh�是��N�����5���kJ���H�a�Π2�j���\3�.3I\&�Ʊ��}!�Sh��p|������%��:���{Rۻ@%[�Q,��+ �	I*�m�j-�gZ9.B�zj�\�J@�Dec�GfP�,t��<��_#�:s9��i������ ���h�<�2"�Ě,�"�M��c�փڠd<f<~��[Y�a��'��
=��tD��wy+DU�Cy������t���=�ᩬR�3�̓���ק�3�����YY/LՠS����'�?h����,uԈ��Qf\�Vc�-�[��=���g2��\���Y�j�@�[V[[������ձ������Ϛ���{�*��i�Y���Σ�����{܋H�Ħ�9f����!�d
�<���\K��ֹரoS�,v�o��h7�|3ݾؠ�'�"a�{>�c{�ʿ��V�w��g�xw��i�C��4PI�Ѱ������hx�҉a������ީ�����e�n�Б
�l�3��@�����:辴�?,--�.��VjC�Y������ec/~�=/�T 3%#>y�̂x��W�)���+�)�����\�E�6<E��'H��^;�;�:���������
�cEc�1"F����vl]�t��v�S��b4H����{.Үm(l���>�a%Sb� ��E�v�ǉ����5�҄U��v-���D&lny&�bss�u���W�K�.�[ُ�]\\d"��Gǔ���Rcz�!��!����řY[}�������ܿ{/ә!�U�f.s�͞�>m�����_���;�s��Y�˗6�k���**(I�@��Qd1Җ�7np��wd^Y��R�1��)�/.,���)��ꀴ��.��/f<��
���u����}j��̖&���_�,�$V��� �%�	����)B�E2s�+lmm�F� �Èm$\$V��w^�n�?��b���;� e"��	��v���SGq��s��~�W�W����ҥ�x��g��9��BK��ӻZ~���w�^�+^.E8=��j���G|�#G��>�{�n��+YZ�!HSY����ĤL����#����}DN��|/%�s߾�:��|�ͷ�~����C����޿�*?h�W�OUan;�b���h�3Ì�#�Z�>��#4��T��NT2������%�i&*+"�fU6�#m�ՍI��a�Qq}H�����ݜXA���	C��$���6�1��#g�}N�Z"��\����cA~4�D��,�����D�u���ȱ��:�s�ζq�5���;�ʺ�{��c���IcR�;c��`�ʰ!�uҤV�L�Ց�LXёh����DYcX�{�����h�ܵ�f�~�:��I�0�	Z<�3�'�5�Wٜ���EZ�#q*lB%F%'iT�cš�����g/C���DU4��` Uu3w�c�{4���.eff�\�F��n�[r8�d �]#�!E���Ӿ���E{�(Ν��:or���u`����&>� ����!��cǨ�`����Zg��o��Ʊ�G^z�%��b���}|��<~8w��zk-+�O�b���E���;6Uo{{���Y��p���12L�k������WY���Rx��2��&DOl���F�5�ޱy��\5典U^([B=炔fa �Xt�a���U�K����`fS�����~˒}�N������&3�q��?Lc�0�Cc�>����^���a��
�玭��ʐ<m`�J��Ė�Ii��K<�K�n�7��r�)��������# .c�l��O�)��0�a��{V�$����\��HK���S��>Oä�0.9Q�����H���죐��~ulMZnp<��N�ׁ�R��7V��CBq�=��[�*�$%��'�m����J&V��Nd?��O�g0��q�Nt[[��n��.��e�'�~/W�"���,~ٙ|ϕ����ĉ3g���`t�ܻ����c��ɓ'��#��J5tdH�$��b��������Uxګ�pj��\G�l �^âr�̐�	�Q�:�[�(���k�E��r�([�A� (v�"���Lf��gA]gF��Rf�Fy�]�v�f���A�h��`{ ]Y�v��T���ce�^8Q#�6�D� �����ҝ�1~b/Wى%��(J�t0�ә����+'<䯉���rπ���������M;K�(��U�גS�&(�ٞ礅;�r���7�B�C�o6bbET7'��s|�o��f��\F�K��&��!wm�7s��s�n�E'|]@֍��IX,@�p��6�]�����X�~�"e�¿p��KTf��Tu;k���8��8�A�[6�/}.�;��C�|n���=n]\ƍ�[h/��6�m�$\e��Z�97�T� �u�DbX?:p���_X��A��,�b\�;y�%m��Fgz��7s0y� �9拶�8��2��z�<,�I�P�05��(�.�<�:!��/�fٵ��YI'�܊�H����Ÿ�cK�֑���+��O
��Mxn��Y�I]�&�3q�˃S(��.ś_ݛ���6j�2=�JXv}�x�{�1�q�Ta�W�����z�1;�Q�y�ؠ��N�1������L{�W�l
��S��&�<3�Nl�,�I�����]X��;����s�-~L��:�,��2�8v�i �X�у�[��T�Fv|"�(�0�ssq�VyUr�Dk�f^�{�a�[�vvf��w^�u��ʾ���z2�����ҥ�$*k���2Z}�dc]�^��.���'2
�-�iW��[7n|;�Ϧ��H�S������ͧO�xT��衚ա�iNR��KP	�0�J�i���<vr�7?�Kf��	╕|�*bww�pc��ݻ����!��N��8�n����X"�_�
Yr�%�(B�w��"�gO�U]�,�_ٿAR7Nn��7_}�v��^�v��d$+�(n����0(_�@�\z��o�?=��y�G�H_����]�����UT��T­L,& ��T3eIF����J�ŎN�0� =�U,v�,�;ۃVH5�ؐ.���Հ*������۷�ӌ�GXz��q��ť\�w��aRG�$�3���q�>d.x:���vP�qT:§O?�t�֭����W�-g�;��'�ܸqCN��B�Ӟ�DP�,ݷ�ĉS�ۋ�`��d��ښs���䘁.�������a����\X�T�v��E~����-؟ٴ�IV0�(pѡ0���#���-����|Ww;a /[������;�N+��h�J�|���_~��R�2_���_ �����Aa������VT���I�r�juiSḇ�2�;�!�e`v�!7jt����V��zm��n��h���ۦ�eP�c~�S��Vro�9�D!����y`�X)�/O��+�Ŝ����MEJ.B�0�XZ�dŚ�)mVF���pd�u�!�w�a��4�e5���2`�эK�H�yAi��/P�8��
�X%�uO���{���-�?��0���o��@Uڵ�T����WX���V��T3�`nB��8Ĺ=Ýݭ���T$�Po��زV��йbP�L�6=��Zl3�[I���X�!�C�Z�D�=8����<����WX�3+";[��.0��;�;m<����*[���5�`wn��$�����5���-lzojt��|U�ͅϻ���}DlL��g�g�ϝ;w��I�k�*�iksQ��/�|_�p��ѣr��"G�o�'�x�D�F戭j�mCl֔k�m����e�cq3˚ģ�(s��ks�>� �3�3Nf0�+��+W���}]��=��ȐJ�i��!�ִTZc��LxN�u�+:	�#zb�����w�քY�b��ʓD..o�[0�(��Y,���9z��Lu;�����k�٤�]((�n&̋���Q���w���G��u�R��
�I,c����<5(VbM��H3���&w���� ��+�`��y&=���ʨN]��b���3�$�u� ���,-$ps��'��<e�O��OQ�\Djp6��0�C�c�͌*�����n�Ʊ��18��-G�=�OX��,�~�[0�Z�?�J�
O���H�e��5q3���Y7�ʉ<�;Q���Ƃ�5F�zc��IY�I`�^ت�����{<�@ш�&�a �"~{��G1�Fؑ���h�Vg��7�B�|ݼs���Y'C��M���G<�Ҹ���
��?<���t���e����'O�\��K���Vo^�\���p8;�I>���]1��"��u����3&�FX���6�u<1H�8�� �B��Ŵ�� 1�eJ��W�`.���(0����mb[ơ��@o�씹�(	Z�����F�2݊��,�$���7F���NQ�&k��ғ��8������F��4�Ub��blB��% $��y�ɳ���p:��v��*����F�+ZU�t�� "˪F�{HT�<��n�	I��7>AO#swR�]�"2�Ym��2���ѬRCn�{W����u�?����v��Qi�+\����Vn�}�okm/&�S�2*��&�U���J���>��s�l�&�	�<NN��g�K)Mo��ZʭC}�������.�D�/�Ͷn�J#��Dmj`�f�`d4=��J��lY�f� ����ebX��J�i5�Z}�Z�eDT���<n,�@�Q��+13�4�Lj�����t��=�ͅ����'O�rMjˬ�G���y�jS֪ar�n�F�{����EI @���[@W�pڻ�
-�R $�e�z���
�_�L�l�'\�6L&��V��+�_ء�W��͸�/~�>�@��Bo��Rܛ���	hR�Nʰ�JZy���n��t��|xp�I^�)���R4�M���T��p�y�9�b��kB�b[t�D��L�}8ڹ|��K�?{�l�mi��E���@_;��o�����}��~�����<h�j
���7!��:�>^Ӭ�6��草l�p4�U˪A��e���R#��B���70n�5nv:��҃�/���hR�/���?�7��Y�;�^Tm�9��ҁ����{�)��M�(��U����\��?��������/����V�p�������o������U�h�/�ɕs�(����رc�Joi{g73B���y�h���G[�rSaat'�7����~��!S̟���G�N�:���O��_�`P�Rw�С۷o/.�_~�e*Ƀ���n#��bAm ��2��w;��������`�֪ţ����vfy��_�4<�~�����
� t�;x��a��X|��;�u������n�,M`"�y�z���{	����JexuD����ob�k�&�3IU���|�G}4��?7A@)�~��g��ZzB�6ަ�����c<!�tlr�W�g,��k��!WY('p���N��ڦ�熀�e�J�J-�nX����r�Ad��I�Z�٢�X��o�{�tL�!��`Ф҇)l�]_�4�lc}��j�EF���Y*���C���hO)*NW�ej��8��3B��ń��Ě9��;�0���*�n�)���b����
���,6��!4���~+����tY���)s뉮�R��4o�2XPd�vw���I�����12����)�W���IM'��l��g���oٷo��:p6I}���7o(9���E�l���j�^'"��[yne�+W?,oۘF��_YD��l#- 7H;�P*#�C�$p�f��܀��p���;�D,e�׼���<�t����[��[I{�aE�`�}�3F�A��K���V�V�Z�}�Y����wrR�&����8�mP���yQ��%,#F�����///jX��Ʊ�����%��A�!�!-�&��ڵk��)����V���ew~�F�M���
0�f<R[OX�h/+llHa@��p))��!j0�ώv:
`@�G�f^��lh��J�=���Jvxg��������W^湃�=~��Zr�2�^bm=F�ǩ�D+5 lјՌ�#K�{9I��.j�.x��yO�2:�����w/f�
Sky�K=3*I��_���:k�`�����"#�q-T7�^�'�5��c��;=��q�;���Jw�;�E�K�N|���f�1��,Hpexl��"[H�핐)�3IG�Fs`k�'������\����d|��>�~/�=��T��f�,Ч�'qc�f.�	Hn�=��-HY���ᙢL�gg���n�j���6o�}�!�tݢ�'� ���w�8f�]���9�Mht�2��}���$�C�	�����ȑ�Њϝ9�-&w����8`H#�v�DK6����2���&��Bd�}Ε��3w�Ds��H� �9�B�gF���l(��P6�#S�Et(0�l�JVK��������d`Vz�U(k�!�ĤvVK�>�4�Y��S�(����7$�]y�$�\[�hG�;KCUyb����b-kdʴ��Ө_ی�ᨻ����)vTp��G��q:M����jׁ�X=��*�g>�7�а�Q+r?g:�Er%:�+�8N�cl8~/���i;��ƽ΂X̋��J�,�N�5Q��M���M�V;I�ņ٧؆�ɩ���j�heCG�Ս�N�Ai�ڱ��i��U9���"�PȎ�̏�:Y��t�bϔ�Hv]�z2z��C|ک�4�Ɠ��Ѭ����#��dWE��+� �`62D�΂93�-���'id����U�g��g�����Jvm�qmSޫ�� �cD�XfD�g�f~%����N]h)��v��R���?s��H�\��:�P&R/]2�e[�"�12��Ě�6�Sl���i�/�7̙ �l��қ��\<7�t($�	YIc$�4V��5�}t�m�o��J����b	.�l�����{���-�v��f��(�/��yn߾������ӟ�������˗Y'LlKi=�^5�`��p'k�K�qijcF2�J��)1:B	't\�{K�ܜ��XՔϢSM`�2��o�
L&�w��*l)~�ƍ�\�x�����[b�����������#��5ۈŁ][[Ӊ�E���V��B<T<�ݻwq{��9ɫFr�O�����6�_$0�^O��+&�o޼���i��^[ۢAǙ��Alq�+�B/R�^����t��L�v��`��vr�e[�G�wz-��igQ��"�Ȱə���/�1{��w{G���֊%Ǫ���ׯ�~���ܹsz("���XR��>FP7��b}�����/�"�~L���G�w���¸l����1��/z��������t$˼�$���<K����oN�<�-�q�� �fm���Ӥ������{VWWqϿ��/_x�W^yeee�9 |�����s���R�ێ;F 8P}�M"ϕ�=��{�x`ϟ�=�E-WG�2�Duǟ}���qy�\����J;�_}�.Z����g�O�iE�}��0����/��ӭ��'k�T����I����i��o��36J�!:����-i�h���[Z�Z����&K�5n+/x��^[�a��k������q��0�����Db��1�5�=�;�d�9�Z�W���}d�h��C׍r����fW)˙�Z^�!r��7m#6���cf� ��;�$� ��l���|J��`���Y�c��Q�8ŉ 9�7�5�x0Y@,��KiD"�Qhq�d��;�,�Ơ�/��61
P�m�om=�L�0����*��������z�m�х�kjK�9:�#yO��"ޱ�E,��g�x43#,Dy�bfd\+O.����/*�ͦK���˩���l��ӧTZB拾�'
�.��vi:��)�^X�� ztD�\��P{�wyy�������]Hߟd��B�ȧ3�Ლ���4LT�,@�+g�����y�������hL�6��n�~����h<������]���&VF�ۘ��ڄ]���tL�?z�������
GCV��p�pW=z������0b禰@.k�s�����Ĺ��������D�!r*�~�El�7^�u���s���А0.�=����?�ҥO?���-�Q�G�Q����~�����'�)�����(6x������c-5ܑ9����#��sʴUT� ��Q��m��l�_�.���O�_����o��uo���k^T��~Hy �5�$�XgFbL��8ڑ�u��6�(�"L�zxX5:c+�0�1��M�m3!�V��!�k�h�!����:Z�$j��z��Ş1,m۔��������s�1E43\Y���m0�'�Pxa�Q
��Y�P/�޲���>yx5U�1��'�.ӯ���af�=��m����v�;�� ��a2�:��1m���F��OVi��Ƞ�n��r���k�ar��/�,�$�S�~$�6P+�k�ʙF�����r���/\��(L&��>����+�C�K/�>}:��-d�b*��V���B �q&�2J[�� �Z� ���uz���Ͻ��N��ܹ�͕�Y�������h���q��.�8�#wc�����.$�"腕p~���*>I��6Z�R*����I����D������D�j�q��K�,�D!��N��$�<��C��Z�x�V�����а�7��m�'�U�Bυ;mL�3�H�
=n`��ŉ�{׳Z�R�WV2�Z)|t����f��=�Cƃ�["������utiC��2k@��B��`I�ey31̔�=VW�L�4�t�lj����[`���M��N���
y~�mʌL͋����΋wj.I����G��D8[e�h�[3@e�tsm�>k/n/#+�F���2�``<��4�U��wl���.�o�]��{(Z���(�޾Z�bӓȍ��O��Y�B��I�(2��`����#0���G�� ~�W�	( ��.Bd�x3Q���Q��n�,Uѧ��t7��EF����:�����X�o�e���8�����ĨexA~�µ�m��L,��paY����R�u��"��PH��%fl)���m�$�3ё4�,R��q�р�e,�(Qw��R�`xp�8�����{���?�1Wl?�`���Jf�U���,~���:������K�c�;�n���c˳�X=1�n
�!���H�_,&B#��k�k�BW�:ڋ�˓��:��b��2饗���Ǐ~����1"��Vp�����`��,>t<�&�_��tCNJ��#4�3K�~H�/�p�������a�$i����t�m�[]��?��9���%�{��*Ұ�-�r��5\N96�>�_�zW,q�'N�`Z�EeM�<�EY�c�u!�~�ǧ���	zx�������F�u�e<���/~���>��E{�#�6�C�7����c,�ݻ���p���X����v �[������B��ə3�(�mir�֣�a��)Ҵq��9�E�,xQ�G�n ��T�p$5��Q4U+��믯_���`߱�{�p�bd�Ù�{��`x���-r�x)\�Yx�a��~��ؗ��7�xŮ6���1�����֭[�<K�M~�aG�<2.�Y��;�G�O햀_vv�spk�)|0ȇ��~?�-.쇇'�D���=,�(��YQ��2��E'v#ݍ%j����L����L�[�]�;rN�D]�,���l8I��e5�3v��ի���}�o�~jÙ��0��#�STAl�eL�O1�RZ�5��A���)a��+������qgjd�Xs�A^��]�������$�u����
E�X��2q����s�.��3>$.�.��K��OD2��Z:�-I����7�	�ƫ@3įHlAd )yt�u�"Q�{h��`b�+7
�ҕ"����
kV%���S��{��~���/��+k�u�#5Z�ʚ�)9�!Fc{���o��y�n���0�Mvs����HQU2Q�{����ef��#�ߖ�,�î�h��V AJsF�����LwYi�0������]�*FT�(LY�PAT��o0#/��'���U��1����k���;�&�_mX"���7u��0&,�rk�f,CG=��
� f�h|�HQr�q��������G����r[�8LH�X|R҅H��������L�Za���{�/p���{痏3��qX��}?D��'�³ ���` 26W~�ϥK�(f���)Z�/w��'�����]��r׈���u�ǎ�x�"����}��b��6�T��3��-+�q�����L��B��C��K�>�|�ro��ՠ(�Z���3������b����;V�9�V���2�8�����}��O�n�E�cv�A7����X�v,5@U�eo�TE��e��l�+�?7U��t`<�ڼ�Vjk^�}���,��H�������(��sK��xmc��xʬ0D�3��d�.t����=�V�<����#�<���0<#������A��O�.c�TKmF7�_�V��S�\�]�dr�bˉ���+�o,���Ҹ!��l��cä1��ۑ00�e7��1rD�d�!������+H�6 
uB��G��P�Ύ��sPwEUtڝ:�ZpP����u9����#���9?N�$~�Tj�<�F���Z�:t���۷oove.G`j�\yD�.��,�$� F���h�CgXm)~*��݂x0E�k�
�6�����_�Bˬ(�(��D��AĂ��[��Ni��T;E������ ��<�?����ݒ
uX�&J�?U�oUd��� �vg\�*Ш,�'���u��J��Fӱ��jr�c�b��Ί2
��!|� � ��"N��nM�C��t2
�P��c�e��Jj�"kx�=I�
ܡ�2�Z�Dœ�R�R���q=�(]��r��S�ţJY�f�,�a�B��5��J�QEI���CEB�.�ʼ�Uز�DS;S�IUʕ��Pn-�����x �ٔ�RX�p��(�UW�~OVU(�'86�TƁ%]E��i��nMx�Q�T1&�r�`t$��n�-+�W�4 /����f�R�?X~;N#H�d���"����(��ܝ��Tmi,�ඳX1�z��x��(�eM%(�a��VA�d<t��w&�*ƭa&� ��
"��u:�x�8�*��ǚM�P���Xq��qpbDLq�|:� ���-r�T6Ӄ��-��k=v<�b�Y˄"���MSi&��RD���X(P�.����=�5O,Ǔ�uc�	^W���Sdi,��Ƭ�
��������m����gy��%��M��#9J��Y�m��x����d~!$��BK�H���v	hK%��m11��AjR���wӂ'���_+���Im�wW�eB�Pu�$Z���Eoww�����7�U\��\� 3j���DC��2�{*�T`�:tę�,�Q�M�WY�+ЂR#�"������pw7���-�=s����瞬�ݼyMl<"Mͭ�G������\�\R���(\~�>�� %�I�!3���(9/ER�a�1fF�4W"�H���+�7XC�|�̉k׮G;Y+�Mƛ���4wT�"��<���ɣ��^?���O��< ���_x��_}=��?����_���=�e���v���.	�v�0WQ7N�6?}��P}�&����ֳ��һM�˸au�&:s����m 9ь����
,�1�Bʮ�����u66���N&��l0��}toZ��W�^�<|x_E�)�*^|���ťv�35���Y�ڃ��ֽ�[;�e���5��	�6
]����n����w�wGi�L��JJ;���O���o��׿���w����/f���^<������O��g�^��۾��eqay�3~��+�*���w5-8���!�K����=M�O� �$��wB�V��
�kK'u4�F�)L��|�����mŰ׹�g�>��le�*T� P�i�͍w�kk�?�������'��dn^�ϱ�ԨB�Y26�:�@��m��������Ga\ط�rh�ɕ5X��y(�nSn���r�c���uȆ ��MG���O������O>~��|������V���>��[?|{e� ������?�c�zq-PS�N�U(�_�/��Ϥ��62򸽘�^���$�>�h6���K��V��D��	|��p������]�C�8���5v��:j�[�N�HL��A�\_��A2Xp)�'�
����,?t��9�(j����92�l-���+��Mh�d��*F��0��[ľ0��u�6��:pKP˼�`|�P'��1���K#���'���g�*�Ȉ���^�x�S嶫�¼��R�2cKґ�5<��3p��H�^�XvC,]�6qE�x�)̤\J�+�ְ�cY�����p��b6�ٛ��t�.]��&�������z�m��qI��;���t|��f�3��ASMgӺP�����P��.�S����p�f�u���c!<y.B��$�(��D�g���<m.�����6U@�D{�rA�t�S�Bjm�X��^���Y�b^���� �:���k�x�}K��-��i5N*�x蹹.u�U(L|)DT0t�c�����d��05�������G�=}���s��ΛW��=���G�m~���t}�/HT!(��dG���t"f���t��81<�'���z ���|*��7�y�G?��+��r���奅�}]�{����۷���;1=�O�:��������T9�q���PԛtGe!���i2M)T\�����t�u,��]���T�W��F�=,et[:�s�Â�ls���f�v��c֚��*K��1N�c)���js����o�FAG�ٳ���<�+XI��p��O�}�gO���·[��J��LG�a���aּ|L�@,H���-�{㉦-@��R��`$�	<��o���*��oai�������T+��v�C/���~e9�g��yv8�e]>~��ɓG��bb�9ݮ2�?EU���C��+8�r����,B5Ť3NM��|�>~x�֭�>�A�G�����8ߕ6�qR�&XD�6',�����(��ȣ�#��`��=��0Ě$���@�BS��k��0$7}9��p�̺���:k4ԷX?ぢk��%��"��j��qRH\C�zV��6�
�HC?~���ښ0`pta$�O�]���o P���q��&͖?l�:n���2�@�(\tI�d��6J�V�D�a�E��dl�ֆڭ0ٙvoh����Hw.)S������XN�p٥��(G�`O�Q�>����k���U���tk7bLןÚ��X/��^m�G�*��,���PEi)��C��C��d}����W����?�Q=ݍŗ�]�bI�k���	�<WRV4�X�n�^�D,��]������{��oڝ���M�%hx~iQ��pBg���z�٬(�y1��D�U�Km9Rg���	�!�)���N�d�h6���J��"3��� �e.���)fIj-#�U�zF��p��q�1d;)���@�W�8���W���g�J-�4͢,N��h��8���ŕE\�����|}cu���;�̋��4�8wu�m�R��0���$Mp�kvO$�_c>� �r ��z��b��̆"ѷ�l��(������Yc|nM���
z��>e�`���k���`�F]��
H�]�>hW,�FV���bz�*J�i��m�l�t��kJ�4��x�� �od��T�m���z}q�E��ti�o�=ǫ��WS�ү�m|'Yx��5�2�D$W�>�)^jI�q��މ#���XAUZ;�i�P'����@���O��[yŕZf-ر5bTG���)� ,���{��"c����`�3Jxg>vd2ډ`����??R, F�g6*5����9)��c1� &ngD��!��
�Xt\ ��l,<�mc|���1��D�@'��������hI-�ihz���u��Bn����=���D輲�M��w���E!�ݲ1��3U�F�Z��f����&�ڟ�0��!qe��L�>|��ԍ�������yj�,�
##5�|�9�p���ўF�@�!e)�񚅍Gt�^[?�������S�N�={�Y�Ke���akH�w����]�xqyy���!-x�?��?�����������/��0[��#ßK�>�v����5����N�%���%(Br�Q&����Ǐ���hg{�䶒�R���ի���ui=Y��N=���i�s��u�#��!���0�+W����w�����{����Nr�z}�-x&z4"� ���OXe��k����ݿ����}�	�~dR���K��-�!*�<?�KŮa5��ё����&3�J�+ֵ������Mޒ��R��hZ��&@\�]��8!j 0�JGC�8;�	����f	��rBW�/c߻:2/�B�>��W_���BT���@��q;���:7�4~�F9����G[@�)�?����������$>x�b$ܶ��z��pd����o"T�֬�x��>M'�h?��O�_�!�ғi���R�0b�:��ƞ,�R�A��<�W1D���l��w�#�2u��V����7/�G�3##kh*Y+��XBg-5�97�Le� {j3f:�މhI.�����	o�;w��1������V���S9�ٓҁ�!(��KP��q�@(�3R�J�%�GԖ�P�P��C��1�*5���:U���E�̮��H�|�'+��e��vЫn�5[8
&�f(�~b<��ѓ!�"��Iޠ���D셼-b?fhY����nט/]m3�0�|_dtH�����šY�����9E�����r�a�KT괰��9�#LƼU5��Ёå!��q-��*f������gb�6ޱ��?�}*@�Z>2�F��ȟ}qq��{���믿N6�֭[���U@��:dQ#C����s��{?������3g΄V���ŋ�ݸqcVJ�8U�TB(�S�bL�8(+yF�Tz� ����5i�A�  ��IDAT�Y�����+ ���[x����'��&���d���\�~���hIc��[K�
��c$���w�S)���I;���7CC�1��r���=}���ݻwq܈��F`I9nxA_P#2N*Sw�N< a9�po`.8��_���8_|��䬳��z$�,�_��]9������R\[@�Z��P�%룔[ʎQo/-.���p�X��7>~��v�B#�$� [=�]��)iC`�e�}�]��'����Q|����'�����tègXx����5I������Ku?[[gRnL߱M2!����E}Q�`7k�]+��}w��R>�?�Ї����)V�cL��^t�{)��=vD���4��޼G���yf͌���l*� �l�dʏP�xi*�F=�n�jz�8��f,V���q�Z)�%�-':�Hu�}<&4k,��qf�ӧ�����[�8�l8�}�����0��ec�;�8cS�{E�Q$+~
����y,�y'Aj�H����y�����C��|���?do֬�{�!mLڤ*��}���b�Kp�l�C�kÖ�:������y�;w���_���_���{g�?##��R�'�wUV� ��a�$��u��;	Uj��@J8�,����DY1U�_q)�<H)�Ab >ϥz��K$X�^����9n#����^�[Q4>��3��;�M7��5������I�)d��N;���NQZ��T�*Y�w�Yd*j3�N^��D�=�{ې�����`���.�$		f���V9ߟ����8�yo��F0�� �(3���$�Ijgg���j��vh�O���H�p�R�F�b��>Y��HR�ւ�E�,� �2~~\�xȗ��5xXf�]�R�+;7��p�1���X%M�U��FF����T�mR'.,�G�[��&v2k6�l��e�bK�z,�ڸw|�'�Gic|�J)m^�u�W꯴�eC?�Ig�ũ�~��WHs�|�]W�Z6�bN׶�[U7����c4dF��xJf�Bjnx�4@=�lUZ�p�Pk:qg�4�3u��n[���|"�U*4�i�B��&��J����g.� �Ii$���[S���J�z47���s�ϒU{h��	��z�k�����f��,TtKK�#��Co����	s��������f�j/�s�ߌo����Y�]z��jVNCNPΪ"�����e$���?Hk�p��v
��b`{�s�:L��Ng�z�����ȑp@g{�>�.�T�x:�3�F+5�A����В]��J�2�����xaq~n���q�P����12KF�Z������ձ��F#�'�z�f�^m41���@�4��vޮ����{�}��7��ϝ=���o�=Z���d ���͟���>`k<���/^�����߭�uX��u�ށ��E�Ōu����F�~4W2y���~j��vG�?����h<I�\�|^43*�Z���uXY٧�?���v�޽��y{�v�:pf�'�n eQ_�{�f�K�����nl<=~���~�3�z��>��0B� ��(:Y�kw��� Ý�N�N�<)�Q�]s��*nd��s���`ﱧ#�ު���$E^��uW	��R�BM����*"�,Ӹ�i)"U&��fh*�{�K�v>�I�]&-�y.J>�|��~j`@x����@�0�jJ�4��#���0�ȫ���Ey �2���ekW�0�j2�Ԉs_��UG�i�%��pK����_}��_��W����G_E��'�	e����1$�R�	�����3&������+W���"�&�S_<��]�
�j}�ՕǫO�x��:��܃�,��R�.5��#I���j��,TVx�۸���[��!�J�Z�R0�뫯!�B.��>��a��>ͧ�We^����!���^��n��R�{'u�Y��H���$�t�Q��k���j����>�[�]����>��L³\�tim�	C��1�#�N��گ�:sK-|bY*�I1>go�+ᖑr0�����{��ia4RNs�\me�-k�cx��ꐀk�Nl-N3l7x�#���f��$�;]��]UA��6��cc�ܚO�X׳'�k�"�R��d �9���G<�c��g�6�0�~�%O�3HN�S��%s��	k������^��G��:��Y��]T��`�i�)��4q;y%7E���Ho��t���/�w�)�I9�W�:����E�����~{��!	���i��&i.��e\���Q8���9�?��8q���~�8���JlQ�Y{������O��=~S�hU������ �����D��Tc_�6�����]`u\�$��-t���|�;���믿�������t@�
�����_���D0�ޅ�2�1���[�O`\�[
�&u����L��U	�X����8>|�����L�����0����q��������H����g�mp���~���Եk�6?����](�p��,e�h�Fb�h��2},��.�f`�jQjx�
J�P���<~�$�g�!mw�O�I�I����U��榣�T�q�K��.N�>�����"s�R��,>�g̔�F&�*�Eq����PL��۷�g�^w�y7
������|v*��1����6k����6rT.u`��&��x O� �n%��ehC^ԅw�2�c+���y.8���|՘DE{9�ڊa����~����[)6�mj<��	���m��<u��=p�K�|��1.��=/��S��L���&�,��f��B�:�G�pqT�F��o�*l�his����~ܰ�
����Ec���T�U�̭���E������X�"�3�t�z���8���fbu_g2��������N�l�'��IYӍ��Sۜ��8.k��k�i�j��Y�;w���;�������?z���E)��w#e�k�(�W=,C^Jkk�nEqV�B,��"���JDT���B�q��̧��Ԧӽ9�p+f=�y	���b�D�G�9:��_��hڱ38~�`MH���]O�X�(��'�S����]�l
��YJ�0ݣam7^<AU!y0�%.J�zh0����?3� q���߿_����%	E�=b{O�j[O)O �[�	e�&r娱,�b_skT ��^�,�=ő�UoN�O!���������K��͡�mg�O|/��&	Ͼs�yn�����H�S5��k�^
F=�#|�x�H�v�=sݜ%�m(�$��K�@i8ޛkL?T�n�7�s��!v~k�S�;�9��.��ƾ��a�=)�|���S�e��1��	2&(i{tO��͒�D��̵Gch��`�T[���Q��,�i��n)lJM#���E{H��J1m�;i��DDq�Ke�׍���[띝A����iG����Jm�����ϩ��@�iY���me�W��HUSi��`�Z]���J�Q�F��Ag��m�`�U�u�L��oe*��ϔ4s�x9ܕ�!�dO��Aex��Z�
ca�"$���S�1bpC����3�d�xwnS����h�7�%s�<ĭ+9��=b_��W_}��>@l,���8�m<Q��!������Y��W[#����.BlIjM��S0���!��$&Z�S��,u��/g�n;S# =\��?2�nhd������h����U��+E�����������<E�[�X�ͭ@/���`�Xt�ر��
���z���"��"A���7�Cナl�.��T�b�R���B��� _�|j��ҫkEGB�_���pK�����/~�������] ����1����駟�p����-k$X
Z��;X|;>r������N�#���(��Wat��1���H�E�Y��������NO@Ѵ�j�^��NW��b�ŐƒM�����,�����B����}Rah5$���#.\�@�cٯ�̀���0Q�=�*�3!QB��=LK���^ �I�H��3
*���'?�Ƀ8t�O>a�L41sd��FtZ,�I��Ho���^X諮���G1�Ҋ8N�{�[�n��ܣBx�SUhB|�%$C2��T�L��!%�hm͐C�$�Tۆ3ߊ�b
���ᩡ1?K�@�ry�%}\hں��[p���Vi�*3&)�����lU��}��i��N���ř�Q�@�/a��4SK��4��a��������K3 �+��`փ��B1��#!Ld�R2f��q��>~Wj��Z��4d��S�n}5�
a�\�s�؛0"|/�j[1�F4���̬��2ʚ� e�Gbd��SEꌍ��m��+�V��A��<Za�ѕ�v�V8d��L��\	�yc`Fc��H���	��Ԩ��di���:�_^ZTC,y��s�3K��H�Th�7v��Aܛ��mAU�F8j����b��jόA�c{:ݕMv�Q����X��sM6���:Ǭ���,tř3gJ嗔���ܪ����
2:x���	y�j���!�3�����ɓ�SW�^ŷ�bqy߽{�,y!Uե%��^�tm�tj\4L1`��B�2:xp��W_{��i�tL_6�-W>��ܽ{����U�c�� �~f�?A�m)�<l�K/���|�!��xd����%��2�ʲ���߰�F��ψ�x9�o���ӛ�W�!�<�aA�~���M�_y���=Z��V���X�N�Q�#��Z#< )"F�0 !0��dp���1����Qt��!�½����C\!�t{�(P+6�'��L���EuܸqCzDb�w��t��0-�̠̉#ǣ
����oǾ����s`�Ӫ����aJ2#^�v2���c-����%WifT�~�<|���~����6�4�ѱ��"�3��c���|bÅ�"0b�V�s�/NMP�\O��B�R�4_�F�6��wPj��L���Pq˳�q ś��A�7>�]�uA��Ķc��Z��2	�u�F���蒧&4��W{$[�=�I\.Ꞥsc�+��q����,--pH��Ȁu����Ine�@/�1�eg���s��FdS�h��D�3^v	�"S�#q����&���� �cV6����b�mj"����gN�.]��o��o�N�.^���%���eԕ)�(��Z�T��tEh�	ਭ�/��������#�SQ�sGK��4��}���g�9��24�1��3UW�5�7�z�e����j��М���c�ݜ,'���,Lڱ!��ե��?�,�2D\��D"e�լ��
im�*1���n��y��m��7��l��V;���h	=V��dġ���d�I�� '�{��Sam��,�&�(�,��eƯ�\GiR1�R�yMF�, W�a:2��Jx�E�H���w"�|�@v�u�HY�pۭ�Ԫ�L�a� ��$�s�ռ��<�_�Jz��Q����ɗ���X�V�έ�@�Œ�g��J>W+?�HU�OF�KU#�����_}LM��pZ�:KY�c�7xp
&C�ii�0�?y�Q����8'��H}w$�kT�m��H$x�I*��:��(�7����s��yY����(�*�
=V����e��d�,W+wB�@x/a\!<�;�K��0��#f)]��[:�@���D74���$��ke�	�CE/"/+&Ҁ��i��{MJFu
���-�7-��-��<4�d6YX\�*��r�4J��y=�IL�GV3-���nN��F�)'_�S⊦��4�$�i�T�LH1��gd�	h��|v5�$��Ww�!�P<��G�E�*�n8i���[����� ��c;��b!A�ͦ5��
���v�C3�Ș�h0���4��ř!Nm���{R�U^��e(Z�r6w(#d
���pŠ�8Z\�+W�`�h~��ۑ�VX���3F��Gڹ5�t�
|G�2����3mA�4�щϔ�H�D��r���t��n�O��W��m���q�2��M?+)A��]*1�ƍo>\=~|ce�9��ŋ��L漠������ @�wy��d���e2��������ˋ�ו�Ż����ԁ�
�|�l���t�:�P����0���X[�D�Q�C
i�v#ƽ���E��G���/Ν;����{�<�Zܵ���[�~�駿��� �����������˿������y9�^+�ؐ8N�4���.�?���:�K�eQ� !?��Of��~��*����������\����a�b\p�F�)�3�@��ދu�&|�n�}�6�r�VK�*�nL�BA�ړ�P��x\t�IHk�;2O��x�ވ�0�)��mD�8�G����מf
�������g�}��>�9�&���.�U�՜��<~���TM=y��eum��+W[���|�T��ԝ��jg���T8�Ա�?�s8��t��/.T����5�:	&�)d;V�e�6�f|��G�v��d��"���`,����T-�$@�;����d]��3���*�籞��l�IC��b�ś�e�������E��YdD!�C+��Q7�,W:m��<�ܲyheK�ضY���XA���^�����U����S����d�>L��6!�Q�T[�/++��3�VZO(��
i���Hzi�8yMO�6���9�ۛIC��pMXK#|���rM��U^m�f%̭ ��=+�!�A#�p����!�����"ܩ̦�0��5���
�
-Q:���ȤO���-,��@�v~~�G_
�n+��>T
�堥ky�H��^�{RS�'��s�{��wd��0�֧O�,՟��PK����<|��ȁ���q}��>�@ϗ|����JP���K�����İ��1�5����
dc���$&a�$��ۇ7߻w�Lme�$�noK�-m�6V���m��k���8�};y���յ~O2_���C�Ҁ���vz�����;s6Ie#�<��W_ݾ}�T�u
����VG�f���L�M���}�����o����/;~D�E�`���7/_�Z����s��q�ةC�M+ss3{�1"�D�F',�1Iocc�͵kנ�WV0���f�!�F6z����}2��ܶQ�&+���r#5ރ�Hr���eT,���:}�����?�;y�Ĺs羹|���5�z�����.���3�	᳏=����t��*�t��8ʳ�d�L[Of[�G�b����ۀ�Nsm����'d��,�?��J����8)���}1���u瞬	�ⵛ7���;G����<���GY]����w"BpZ�M�c�4��B��`���b�3X�_�艭�>��k�x�.��L���M����f��Z�{�"<z�hyi	nN���hh\Pk~�ܕ�U<�婖����(����2vm�����##��mT+�ɡZ������q�/��Rl��8�l�p(tn�� IGuq�;"��Q�iiS���p����l�h<�م���3I�_��s
"�}.��\�����t9j��q�ϲ��H� 7kٜ�$8[�9d�c�%e��7��23�����R���k�uO��2ka���Y�TpO�4�w�sd��n_b#>���(�Ŵ��v�c��	L�����.n����y{������ǃ�����+��z��Q�\a�Ӯ��+3)���iG��I.���-��Hd+g��` W7���YI�eD�����#�\��n'R�$��Z����d�`q��Řj�I�׸ l�Ӣ{���HmF��^�ʻ��L�c��æX[�YqJ�-��^��D]�~gK:�3NJ��]��M�v4�f�p/)[[!��FoA�(ieU�c,.�����+���j�i�}c���PN�~b��	�Z�(jI��{���.�]*ߵ!�#-;���Q�k�z�u��_�pNϭ���Մ
���2YV��f�	�+��o<.Y#����"w��Si�R�:�x0H��Z=ľS���J( sX�Lj�5B�A�[BɌ����:�����+��.s�Vj�Q�L�Iu��dQ��_�!4UO���'b:�1���}FJ���A%!&	\'��Z���"�4�u xn@(�TM���������,{�P,U_��q��Mxiࡸ�c��<�V��LM��~a��R�Q�OR�yCR(z��y�*�1?~�h91.!�*�i('l����S_�<�އ҈5����b�Ҹ�kC�{t�<I��=�j�(�6�Ȑ,^�t�\^�1����8�If� �A=�S��
��qRظ�Ȉ�����\S{�K��(u����� �=�H�-��ΌIǑ�E��K�����m�
�)'��-p�kB�Z�X�)�ӢA�j߷��I�fORh37��u�����50Ntf:����O�**���S��S$;�X����Sn|̎kBN<���2����>|X����_��|��g�83z�nߩ��{�/9�|���`���n޼y�ĉw�y��11\�E~��_��:6p"Aw�����O��($*���,�p��d�E�%�;��*[\hA���i9�R�Qilo�y�X�B{����`�����X�~����\��"rK����`�a{g�����{�
o��&�lx��|��o~��G� �N���z�-��v��u,]l8t&>j�_�.,�c�������\�W�e�u&��7VάΑ��$%��0�,=Ѐ �֫m�@ozԋ ��<� ���h4����H�-�dw�չ���r�u��{�����Z�P���=g��a�o}K7c~t��Y��/��L�oaN��<��Ν}��VV�5�4G�����oll���7��<��]57�
	2�U�nGX�'�=u��t��L�ںp��񄐬�Гg"H���S����!��/-��8��EL��9O�	?����>��v�Q�g��*K�)��\I�M��v) �ښbS������ð�Y�@c���ٳ�q#����JcW�-r���Ү�(��XQᮮnC @���]��!0��`����ϡ��U��8Ϩ�`��F��Sd�DȌ8i��vt��cO��t�p~_z饶0)���?f�+���ţu�}�{Q(Y7~����Zq(<JL�Vk�"�,�gg6 G?��֋���{2Il bc,)��Dd���P��ZX.4fq���8�֯��ʵ�mqY�&Rn�@�'�7) ��!ppL"t�>�C�5�snsF�Od��ޝ�ʦ�w���ġ�F��7q�$���	,���	Y��t���L��ח��p����h�NCoT(]��u^��x%�H}�6�Gj�<өw�3y��Q��k�/]��%�V5;�r`�PU�T.��.}�yq_��@����-�F�=��OHGY5��<Ŕz����V�-��!Z�7��#,+��J��g������*�;�n�a4T�Mc��``�r��h8	��t�9�VK�-��w�{+�V���	"���ps��P��`Q@5�׮\����ZW�:2�{�ӃJ�]#��23�`������	�
�3ۘ�s�ν�⋸��ӧ�>�G�x�y����wVVVނ�q�O|��F`Mi�&b�H�~�)��T(}I�'ׯ_����М��b��p�E���2��0��H����"?8;��;G��tTYY	��N��r<|��o�1x�m��l���
�9"[e31<��oo7um���Sh��.�W��;R�1���)�?��-fY�U�9|X��2WSV����)jѮ&qbҾ��o�NFK�qpY���Ӹmɐ=^�lJ:ib6YW��h�'7-a����(
�/����څ$��u%�&) � 4!������9E�D��O��9��'�!�cC�s2��8��չ�)�9l:AA�?GR�4��.y���	G;���:���xj<)sZ�	�����,�΄���Sg�HBb,�<�~������q/z,���&	Wc��s[)�/4ܷ#��H�j64�ym0Z�����V�:eİ6��/}
�S+f�70Oh�D.��,�UGl����Ts�Ɔ�t�5�$�pa��^C�/v4\d�>�p��Cd��U$WN���j�T���rX�xXpM�����|rj�ԩO�lk��ݷ!��ja�j~���Ss�x�7D���w<Hˡ1J�����j�s�"���Y���O������B�6jB�J�&���*��^>oB� '{<��E�D'�ZѬ�U��g����^��=�
�\�$rAJ���N剦ٛ�����F	�8����;�W�������G�|�s������Ȋ@����uUg����b{n��n�r+�º��$�Q#	:��w���L��RVM����C
��a��J�6���(��H���~��=�4���x���	$Wv$�Ĵ�<��h}8.8���O��EH�J=DU�!����"�Q\POPз�� ���
*}>�=�U�C��,������S������P"x �_A.	n}�޽�8�9�L5E�֖l�����XA���b�1�9EJ�n(�y�a��?UC���`����-z2������b{S��1P!Ih��<lm+���%���]�V���A"SPNQ����H����G#�:AIt�=2�ӈ�\�z���۲^�;qڔ��FF�O	�xv��Q�%��}���&F�늓B31�F:�f���Km��=���Y�ؘ�UX��t2���]v�q����.��ܦR�Ť�$���-��g�a\*�ָ�(K햣q�����8>3�9q�j�tZ\7@k+Ǧ�wL>�tXDlƪ|�մ�}��	$��Q|9Aq$��i�W�ʢ����6p╚�{��Ã�v$DidP^�v�V��`s��n�w^R�%��3@lT�93 �`����k���P,���x��ɓ0��R���~�ml�sg�=��IဇM�0^[����0� v.|p���۰n�>�oy?=� �M1<�tt�J��m����_��U�$����֭;X�3g�U!����7S�_F'���j�?t�Ӥ���$f�w����x����J�E[�
�у[����/����
���aOUA�1�����o��ʕ�X�lR�Qu���w�yG�O>	(dL�.�h�5����$��!����,���^�[���ٳg�7~�_��H�Z�&C�9r�g���^�ɏ�`m�&�Ჯ��
���_x����^�BFE�r9u	%�,}������=�ru��k�1L+v4��c����"݉��:s�̉㧰����y�ݝ�SO=E^y��\�裋����ի���O��t�/L:i\��ˉ�D��jU�qp_�O���b�^�r���,�z������/�~��j��b<?�����ﰊ᭷�:�����e��T��_��[��A��t�[ ���C�5�}{S�qH5�d84��� ��-U����'Sq��r*�d^���7��j�B�l���g0oΝ;s��)V���".�ˁ�}��1L�Z [���&c�ӿt��vMYV�`�
Hm��I6��1�����V��zK��2@�����2�έ�7��(`O�V_d��	��+�E�Di?-�&����^���:.g�RZ���6�T?��L�PP0T�tQ=O�\earfum��L�X2�v����_,̗��@�2��y����D��XuO��Q`�`3�ӊ"��;z)�A&cce��[�,�۸�r%�)J���)��Cô�
�x�(��KEX��DU;r����[׿��o������w�4jwRNx<C=�O���ӓZ�2���6�" ��iU�OBmFq�������%�֏�~�۩��Y!&�����"ǿ��t��J��n��1��.I�(��$��t�z�!Aoi��%8�u�s[+~��$04
wild�8�U� ٹ�a�!+@�1pF�!G~c�E�)��ĺ�`l/�<~�����G���r�S'Nt�����`W`5����t<�L�Q2ꙧ�ZZ�����=�̴��2&��BldG���ϝ;���ϓ���QB�h	��7n^__�8�}m��,�:�>^iL߅Ѻ��2��q�A�5WVV�8RS5q�L���}�ў'���J�1���Ě�N�����@�1�@_8�X}�!�R�.�7n���`5ޔ�Ն�IL<�s�J��F�.�d	%@�ĪNv���Ѱm�4�������V6�	6|_]�ֵ�ư�QV*���q�%Z�����모&t�qkl�V�� ��X���fڦ�q��PNG���;�no+�%���b��ݻ���=�ӳ�\2�����b%Q\]eX�j�ↂ�M�R�sq���4
��<#���0�����hx]�$|�+M�f��"���M
�X7�$��������ׄ@32���t������8�2�*}��%���V���j`�x5F?�S��/��EVZ����N�M�-a��*��2I�����%����f>�J�^���}�Gpʼ���8���J�qnpn ���C�������B+ۚ�����Ui�!��T*�7cww��\k�@�ؐ�� �b�z���eܸ^�WX��y0L���U�Ҋ�f`�l�MȇR1�Ԓ�iUdh��ʓ#kx�i�j���y�Y/�Z#��CԬʗ�wb���h{ uN����'W�܆u}���}��w ��G����}� �A��ӼH�K��8MZL����"�\uA.�"EYG�oN- n1=VMVm��P���<�!0�+�����I��M�	FƯ�Ӭ4���a����hJRmĔJ��N�G��Sޢ�)���Q����4�QωP���S��Ƭ����>���zO=�4<
hw)1k��i��^����.���V���`g �l#�,�nٌ��ƕ)zh��IC���J�-�.3�-0��2�8M��ބn��ʐ��5����U�V�$�7`D��
#�B�0������$s_�iKS�D�T��#�C_��Jt����Se��,H��4�R�(N6��[u��~����T7��?�p-G�0Q��.�3�r��E��$�'�F��ݻ|Y����5S�[�;�p�.�s.�|�M|��;f8mK�B�ڄK�W�Z�X���`ΓP��0b�"s��+q�Jk��y-�cO.1 ���0��F�J��y���R�3}����D��:�׺���(�+��&ܸ7A=�8��xz\����]Z�g��_a|��*�����q�[h@ T���+QH����	�v� ��N��U�Ш��xGQ�:_j<�B���EI��4� ����
<��%6�P<�<׮�H*Y�0���@3{�������L�a5�@՚�b�1Q������y9t�63-�'�|��?&i&��No��
\X�ɏfڬS��3,��sec�ws?�r���̶�y"�)]�~��d�q��[o�ŵ�qÛ��ܼySV�������,�Zv�������H�jXc�Z�N~
~ˋ/}��~ԩS���X)�`�~X���%?�*Fwׁ$a���'���G�s��Y-���1��:_g0�It�:�6�y��lם����^����o���ę�q���W�k� Y>�����
�M��fu�a������w8 p� <��o�O�[��'NH4ms���A�jlŇ0�O=�L���t%z��SO�aTՐ���1'2׃��u�)tQ�Q�	Î�;s���XA��cD��_��;,���e�wX/���ڃu�c��}���ｃ	�t�~��w�^"wӊ݁E�N37
C��"�c�m/��i&QEHoL&D�O���M�"�{���Ԓ�u�`~�~�{��_�u�%1F<�n�λ/���d��,a�~����N�hF�.,/���g?K���v��]��_��c�N����_�%��W�W�D4-<���;��g�9ppjI8�O?��+���R�@�#�П�.��y�����}o}MN�8L�)���/b���߭g��#����ԒWkB'��Y�n�s�u���u�@��5����1.-4Lẹ	�kɛwn�����E���1�t,�;��t�2�[��Z�OL�p��80��_��F�6�q&i�ѢH�j*5�)Fи�*K�2��Xiam\W�񵑒R(��&���3�����Y���c��B�W�"(m���3&���2t	�1��b��G�h�X@��݅7a�A��گ�<������&�Da�ǟ�`��w#l7��3Vc��)����I|���1~�˝�:��2�Dhe.�?qd0���~��q*0�/|LC��#zj����ٳ�8��=��T�7B��#+uwp�H������R��5u��P,�1Y#�S�KK۷4~��y��g�6� R%Ҿ�x"x7r��R��P�	wa�(V�Ab@�a;�K_z��3�����l�FKy0*uՈW�fXA��ӧOA@w@� Uh)����}�E����	�56�e��
�_���8;��Ĺ"4
%����ь��� >���d� �hvF�,d��۴��!����vp��ǐ+��Eo��,��t�ȢŔ�ըDQk���-�I�������"N�<���U;4�3μs�0�����	~��59XZ���#Z�'b6��a�Yk���K�`k�
�����f�50�w�<]�h1`�U��UOfm.T&\nJ3�$��\�B���2˱10�dl{Ƀ�cH
F��n'<8t���D"Y���$L����$�0�l8�0J�O��9Η��Wc���J�x����E���<4��'��Ƭ��oN�s�%[9w�S��w2|fW'�!0�Z�åJ"��>"�"��u\�Ⱥ�i��õ�΢�w�Ǳ��H���_�0������Z��|�uK�Di�{�Sk�,�7���<G�`I�J�S���	�^�;��}NcN��aq=���hX�Sh$*��uj N�!QH�cؒz��T����		�nᅀ:U�|�@�
(�J��xoe�w�P�X�d�h��@��1�rz=�J�����y���!1k+��\1�=���s��.A��0޺2����p�P�Vu�I���-Ũ����+��:A���$�Ҁ$��(�U)�#�	w���`'}G����#G��M�g���z�+������Մ)i� ��?�m{���*?��wvd���8�]o�V7�록������'������;�Qe������kpA�)1�N1���غ�[��1���c��>9�B��l�IfI�/�2g��: ��w!�&��s'�c|0��5}�{��f��,��,U �.D�����*���~����� ��3��q����a�PvZ��!����| "?yM�ǪZ��6�8tk��x��	�n=��!�@@������]i�{l����c��z&U�t�v_K��R��g�<�裏��?������&�7X������7�"�FA����Xq���h}�ھ�:�^��I}(#8��R�Su�%�iW�q*5�;��0R�Ew�֌1���F�qŦ:D���y��ft�r��7��@�9��ʵ��߱��u��$��ؤ�I�	*�Vk�)R�N��EM)\����[����hnK��� ��xX�t���-��ݻ'�]\��t?�(���ge�Ҳ������R0_����ѯ�>��'�(LT�8v���K��$�Ԋj����a7gJ��yV�r�n�����sc?��Sg�TR7� HT����N*hG�Jo^����r��%F*ś�������Y��A2h�a�2����@f՝[��q<���=���V$A�K�2+᭒,�T+I;]��,,Ϋ���XuRچ���3ψxi%��ʜ//�#����|�����+t~���%�1G"KS���̸@�$�j1wÈ�8�ۭ������ۯ���׾���ܰJJ��n��#]�R���<+_y��~��p+�~�m-��̇�zRdg'�O������-77'�i�4�&��`�-�l��'k8�X�ͱ㇪Z��&���'�4�$�*�C܅�$0�J�~Z]�1Wb6h�Ҁ�~�-a����cǱF����u�s'?uzy�����������"^W/�5�p���~�ػR�ٓ�,0�ّ=�ų�#��O�>	����Ꮸ�R^�v����w�ܓ������U22�����4N W�+_�ʋ/����F���'�xw�*!;�;�e����GI��ף�<����l�B����|��'p��x�	��ׯ��������O��!�˗/�9s��Ge>�#wl��x��H��ӟ���d�� l���qq^Z�N$��S�LHW�t�K�c,��4n�6�о�m#���a.AL�u��00~*5���&�&�.����^�ڵ�bЯ��=�5m�̊�D�M�(U-�����֧�_M�?��h�fw�K�׳��Bcsw�/����Qye�o!	�{��0P(wa��
��4�&�b�7Fh���[S��O�=IH�+ږ����܍�A!ܔ��ъ���I%F�-&�j���7�������}���_�s��ʝ�w����	�NI�
7(�0����uwSCh0ѣ\k>)�gmW�R>�g?�i�� ���ҹi6VE��;;[A��X��y�ܮ�>���7nL�bN��v��4Nŗ.]���[<��C�v�c�J�g��
�|�Q�mO׫%}<�͍5f��V6���Ɔ����x�X�xƅŹC�!���U�� �ee=���P� U$�������i�1ì��48}�twn���ρ&�1x|�ĉU)���*ZGҭ~s�g��:�z��*���zG(�����D+f"bXxzec��7#e��>�3��;���n�f,�E��~�ᇡ�q5|F�E9ɖL�&�8��:�D�2�/�}Ǩ��{)�d?��s�=�=�xxG�����'����n����$`�:�d��i�U�;vduu����at����XFU�����H�]��V~JC�m]D�sK_�q�h1�2v���թ��%[�����R���Q��4�uR���)��S�S����)!~}�.4����L�uB��`T�����ѷz�u�x��Kҭ`p�#˅�4�6�R=b���G�Zj��~�a�-.$��8��-{�9�G���r�����f����s��f��$��59"C�Q6�kcp���ݳ�=M\����&$��aY<)����tNe��'4c ���/�3�I릡�U�iH�Sق����2&���I6�oBmNv�Zf-!�h �+�0�ϋ%�̅=��F���H{]Iy޹="Ìs�P>0ZǮ��#���2�N]:�#�0�}l�|�5����{K�*�������|d&o6�;�}ۭxȭ�`���V�9�yǭ���-2E�^�vz,�\�ܓ�����Z;8"���u9�������p4�پs�&�bqI�8#�íByF|��r�r��PM������-�la��۞���8Q�<�i1��nҔ~�4�h$��ti�N�%`��'݁_�;����Ҳ���&��������֯�ux2o�����
jY#�`g��%:��f#���I��$��6-c�R4��yݲN@Н�8�����J��X3h�/K��,�4��Ag��=�A�=�pmE������������r�_�y�Ě[���x_l�Ufo|���Sb��	�v���y�H��L�EZ�e2���9�,��t�c��Wl���L��ǉ�Ǝ�`�3�ک��[���т4s�޸/|�8�D�/xt#m
�4Al);��6	�=
:،�(�P]�LyY>�Y��,���ݘ�����f:;PP[���V˘�\E�F!Q�M^���272�le�~�K�>����������\�Z�w�c�����<N�<�0��8~>��Uhy6�8G:-b���Z*�=�*�K�111^�y(�/'���ϑ���)o��<�ia�Z�-'�Z����#;|ҏv�pz�.dg�d���lP�I�
�@Txd���_�s����¸\�rG���N�&8%�Fy��`<����bqv[��nid4�i���ݖ��|n
h\�)�
��jhd�����iw��1��R��g���3�O�eX2��p���H���[oŎ�m��x7�����h4������^xᅗ_~��1�|G��ҙ��6XK�;���c(�%��`�k���u����̙33o���68�,bĬI�c����Gh:'�֡ ŐVWW�{�o|�����C�#���P�o% �ݱRx}�?�<�x�����y���o�ⰼ���nn^�zuskC�x��r�~���M��2ӿ|�ں�p�l�`v�G[��7~�q�YS�����eI$#ϣ�e���O$��̧x��L}��ߖ.���v��nB�L����M��N�"!�@�:|X�i�c�(]�'����I�����x�ȥ�ɭ[��_$]&#�na5C����%Ú��'����]A�_�B�	Sվ��N�MbAY��GjKFr�j�Q�y��;����o�?��{O�L6U���e�i�2M�/3�*�M�j�f���:!�`����QQdQ/gƤ�� �l��fm*���Iq1R4��&np�����19[�/!�)CoG�J8
�qyVi؀���E��aߕX��2�A��-7>�¬GJ\�Gh��n
��|B;�kG\��e�y��\���TKc�LR���M�DUV�X��Ј�u`��Y�4�(]Yq��2 ��?��?����@��z
�����'��E��yˊ���&�<���a��s;��h�Ԗ��Et�(�a8ъ*qV��N`,Nc"Ӭ` H�m^S<��^��pM&P�g)i��\�]����OD�Xأ���ܥG��F�^y��L����x��u� :n���2�ǒ�O>��������i �KA�cƤMku1T<iGQ�ӼPz�.;)���-�ȵ ��3��둍w�ݘ��n�bT&D%�32�lon	�k6�6���%>�qb�4P��|�G��կr�_�ɏ�f�8 �j��bO=k�?���&/���V�����A�Lu#�`~N�kb�6������s��Y�}�c9Pl�Gdq_�Wn�Yݖf,)Ռ�'�t2���!�ɳa��և�B} �7�-7ј����y�O���Z�\|S�\
�7�B�E#����es�2,S��K��)��%0�]�
|*/��D�SD�⹖��\()�:is�v�P���۷kcJ�-���T�D~�6���>ꦩ5�j3�[����R���zX�����a&�XP�V��N��7<5d��F���;��4��a�y� �F������2�Ԋ<y��~��E�$}+G�Q��i[+�qq���-..��c<.������PY6��4�i�BčIޗ���d�G`�=(�=�������RV����&��w����g�V^��J�>���I�PX�c=äXɗ[�����*ㅌ����8�L�������[��=�{)���؄�?��XgIlr/P������
]�"/��&Y�u�5�xou�MQ��ՠ!�s����4fg�?�Gq��]Y٫�FBc'�ߤ���<����ܖԌ��t���xhWF٘(
�M���/���Fh	�3"'uώƢ���BbZAQ�kUj�������F���9l��'OǰݓÇ.-�[��Y׬2B'4�V�|S�:܋�{0@��0fX��*���eI0����Ը�v�-�~�J��MB���ĵ�4k>L԰E
D>
�����A�{��=F��"W�iU�X�,3�)j6����N��Aj��+Y*�`KlM�ںal��)�ǰ�'^���T)Q��n��1�Vj]1���\�H�`	9U-�y��%�����ju&��[:����IbøJ7�8�ϵӖ�j�U"j9�vIT���gvQ����V�����p[j������WD�#�u�ש=�u�j^�dD�p�Z��cID�xP l�G�-���8��=����m���&I��%J�c��L�WO��ӑ�{;gϜ~�sO<v����ߞ��:k��O�J��+�H��̦�Ɛ�jqh5�v��?�Y�N�"[Ø�O�M�餰�Q#����KWu�@a�Y�O�4�W�>Ci��R�S-Q�x:l�l�H�$�x2�'P|��][X3�ү�ߗ�����lT�kI�4N�*r��b<��r5EFA!�v�|�l�ᝡ�F,�,��NndWE��U�*gx'���WX���5f�h��eE�}�n�$���Pm�zcȩ�N!3�|��'Wv�J(�}J�����!�v���O[�`��W�hT��{ׯ>{��zԉ&��ƻ�߆;��Y�y��;����v��m+{=����`#;>ի_��믿N o�p$��g%��wށ�z��YxD�Ta�HI�����N�-P���V�s����-TzNs��9:F�.
|�LǍ��g6���?�n2�P��.�xy�:V;�mmmfq+��o���FM#�V)3_�I8ם�'��T�mEw���]�*;v������0Dݺr�aݴ�|Z�-�]� t~iy�����6p�}��k��h�.��ƚ�(C5�xܴ��f�*���"YK`��A~V�b�aܶ�Tv����4"��5υ���co���������q_»��0|p�ҥ�荫7�㞻;2�T�[��e�Ŵ�I�h�meE6�cճ�R܂Eф"���e�cbK��nm�^���'�x�O���l�5�4�p8��d���� ae&��9N�;��0���r��Y#2�����Ɩ�8)ү�����I*;��N����4@I���O��[�b�Vh ��!r���6�jޭdv����_�<������W�H�
���2~�i�MIú puj,X.���GZ� �����+��(��6E=w��&=��[��r����O�D
a��� �T���'�8��Cl�R�1��l�&�J�����2N�zt�Ө �	̫W_�pJ4)ޠpg�BM����Ѹm0�tt�Ƀ��ȱn��`��)�O�At�d�ؗI��r���%�ac: ̭8,;[�����������s�<�0߇yes��H���$��Ě��I6�JB��v�|�&�=���ߌ��i6]R=W�ykgG��d,E���@�:�����O.�����;�$�c٠����تeQG��F���847�ml�Zb�$�<N�}���M�D�˔�Kp�������cǨ;�-ˈ�	�$?1�	.��Aj�66�ڽ��?��N\�hq����;ݺq�o�4d�ɏߘ�/�����N}��SO?����19v4vo�� E�M�<�᳹�������&�-��&�>l�z:�l��D%��>�����_!�Lby�c#�H�R�W���4���0�*K�,P�}�`Xn�J�-��]^���a�?!�:���a�Yw���w$���X���gf��psf2�)��o�W���X��v�J�����u��c~K
�'ʩZ1M2妥	!�2��ٻy�f�����۷���a8�;p�ǟ�/��,���ʭ�U��Xٍ3��,�����WB8>1�ׯ_�<��lК���t�+�@s64�1l�4S��ڔl����v��̎3�CLt�����E�$*��6�7��oonQF�/.0��S�.c-��ȷwTԋ	鴈�DYј=T��
��Ԅֹ�����L��b��ae�:)�u.�+��TV�S(�"�k��]�3�H:ij�F9V[s�ԩW^zI-�������K�#�S�]�J.��c� ~�s08" g���3g`�҉�;8�L���k3��Қ�T����O2�����F���qd���:1R11�6�ц���հ�A��{��Bw(�S����/�Gf�<�憢���sW1��Ude��P���c��~��Yii�Ђ������P�DH�R�I�+W�̓�b�DnVR�(mN�r�k�(K���Xߩ�����-���R�!�VB7�YM�6��ZNtю��ȯ�z͌o��+Qdx�J�	���O �nƆ~�Ӱ�+,@��Ѧ
���
b��I��b�2���^<#�j�1�s��<����商|�b�	]fqDQ�;�!��t/�����n'Uz�YR�=$�d˪uԑQ�EjaWf<���k�z!Z�'h�*�[��	��O�ava�
o�Z=�1d�-#[��mp�`����ke4ygM���P�\�ò��V��[9:@m�������,g����ʺ�	^Π�]Ԓ�F��(��F�q\	��Xnl�\�q���iyPњ�u�2�(�/Vh�����R%��<��ه����5��&-	��G˱�����΍`��Ϲ/Me��_��m��L�:���(+��ݓy��G_y�˗���TC��!�ͪ�~����~�)c�B�u<D�d�f75�t�K�h�O������le訇Ę <{3;�܇�}*��`q��<_��Rk+L�9��=cG�RX����&���uR�.W�ޠ�_��ۏҐ���� dV�ĉ=�.~��=�z��%��v���ʺY1�J������6��С���7n��XK+թ]1��|�Mv��{i�K���c�&���F3Q�1e<���T��FQ�o���\��3��GFP��i�5�^���,�)^}���~���u*�^����NG��ҥKǏ�wI6����s+rB#�S���ŝ�4R}�a�F�����?��n$W���Ç���T�hRP�p�=x���eI�\��5О\�0�v�^��>��W�����9�3��|pS�B s3P�x�x�6h���jj8�=Z�_�h�l|�����/~�W���3Pj�d��?z�h]7hbB�eG��3
���}��]�,�9C^�D��d�bM^C����ì�9���u#�t�\��^���`W�lU�����~�᷾�-Ŭ5�j[��Uٜ�J�)E;�4���ż�b��f>++�ǃ]nl"%b�3�%}��X`K�J�����Q�	��F��Up/��Sk�h̪�L�.7�p��;���|�n��,K#�)g��&�4u�@ق�M%E�JI Μ^�Pk�dkMr�]b�Q�E.��J���� ����M�>EC6DT�G�u:�8��u���#7� L�u	S'�@�[M$������O�W�y���2^�2���Q�e�:3�Kr/����shdR1�f^W��G�U�@��K1K\����qY=<A���q.�OS������v���}����9En1�`\�%$�-�[��ZI�W�A��ϋU�9ݿ���������W���6�KK|��,�XACO�ȧ�
��L>߯��l�:iϜ��l�V~��<�$l<��^?���H�ﾋ�A�r�Y!E>�VK��1����JawG�B�Oy�6���8��ٱ���M1�P��5E��#mNn�@���9ΦT�SO=��5��-�Xy��U
��<�|��9u�ԓO>��BW�^��YH�dU���؄��f����uj5�b��f��\�K�,V���nĳ,/�b��C�iBFJ����<�6����-��;w2!l<)��4Ep�u-#Z��un��a����[�T,w�*�rQx5)(D&��H�i���^�~C4Z*!��E��ͫ���)�"�\�@�	l�%v<�ţ9�$��;|�yia+K�w<m�㜟��z�������]k$������|$Sh�	&u��D��A;*D@���TT���#\&` l��<�'B|�ᎏP�P��V'��q3GV�&��s Z��t�(�YQ{���saY2���������u��募��]�xqe���d�)vQ��Q��Tr�FG_C�G��?�����ȚgZ5Oq��E
m�/C�q+k�D�HkgC_���V;�&�S�p���#��/vv�sK$ҥa��,/���nx,f��ݻ��_��_�uJM��Wi��A�����U>�gm��Ҙ���gr��32�?99n�xD"7[ZV��V֌�im%�Y4��a@�}V�ֺ=�bd~���"4���rq9��U���J˨`h�{�!����Ǹ��=�B���M㨶�	����̯��bq�
k�"g@��>k宀E�O�N���
�6�.Y��2� Zi�ѡ6�f��}�+؉U=&�#�`��+��<��p��c�71���	t1V �QN2�ͣ�cQ���!��ܣ��.�+�I�<��bk��ܖ	�Lt�h��j��0R_B1���l��Z޷���%]�����������4Lc���Bl�UP�>4*��(�J0���m��ꄁ
#j��2�	�g�*9�_�4N�f�f�A{�k����/�R�R�Q����6���>�Jv)��ǂs�CU����v�_�v3�J��B�� �1��TI��Q�,/n���T�Oi��*ĆnȔ#S��X�򘇇���W�ȷ��i�B�鱗3%s
�d6-([�D�6�\!�
�,�}ui�[�-J�Ï�y T�2���i�,����J���,�T��=Q�pM�h6�,4T�`h�*��Xi>by������eʥ��a y��\�]�	G�i���ex0Q�+U.]C���`�R[���p�K�@W��
��4��
G�%���[C�?����%��G[�K�ti� �1�����DH�;�P��rF�H���ie4H\d<�94��3���'x�Ј����х���M�zL���j�~�N8E��ψ���2Q-�-ţ��8�������B�pH{]!I��$�G�q��z�pm
=NV�\�!b��
�5�k��;���tzsS�L�=�: "����?�0� ܕ�p��ɚ��SMP	�����B_׵�YQge]���u�JW� x�G}�����	o���͛7a�<��P�,,������A5-j�Zr��k�¸V`tTK��f�Sw�֢+�X�T��i��$[��ѦbM{��HHi	�%������G�Mag�I�������4�^}�շ�>O�PѦe `7�(��r�*\��'O2���s����'�����+XZ^TCt�RIg.��b���d�෇ʘh{wlY<����"gMm�=x�X�JT�ď�敫�>�?�rW9��,ZHq����O��׿q��E�o��*�'�Ʃ�./S@���ő����3ܨ��o��F����d�� U���@����z��k�^~�3x�}��<�Aj�(xIK���*�C��!�8=��
C���'���
p"���Q^"��ݞ&9�5���Wx(��:b޵��S���Lz���ﮬ���?i��L�$XX�#��������RZL''Х��x�8��A�z<�ЯrI��B�	�!!��o��?�T� ����?O�']H)����&��z��]t�cāYX�ʨ6��S�Jiv����ڮ,$8�6�eLg#`$+j�v�Y�B����Y�C���Nֺ�Ҍ j�!c���u�ɲq�vD�L#����C���BmGK�@������M�7$�]�F�H��T�.R8WF��K
�ܡ��ik��jU��7$��3݋��FQ�껉ȫ�i5u�g���z��^�㚹���崻O�aY��ĺ&3�v�x�Y�LU�0Z�3i���j3�P/C�I���^��-��m�4k�J���/2n˵�-cJ�_�bC���PÙ�u�WȂ�B�LqRq�+��P���f� �.�/��0�m����o{�Ϟ=�ۿ�������w�|��k�n`����U�A��m)ءQ�y^��0T.s��4�VV��X���j(>��!Y�s���]\�{��%�B`�Í-�],Z���X��]ZPh���fvS��,E��G���q�Sr�f3h��|Z�g_bζ
:1���2�RWJ�da�!}�X^�/�p�,^�t��]ǉ��w��W_=w�p�����P�5:�0&�+铝v��˿���莚���wwο�.wo~��k6�̭��/��xT�_�9�VW.�=�T[������G�B¶YY��f�q{PO��+W^�uZhO>�$n*!K�TB���zl%�f�Ԯh'������^�ۉ`]t���y�J2���\Oe���-=�rZ���}������D��I���oY�Y>	�Y����Y�9"^���@��;C�V`3rg�Pc�C$�4U���\(����*�<=����L\Ye�h:S
?;w���6���W`�:x��n?,��KK�|D]6�r4U5[���3�et����EdD/�vvr1B�W2c:^o8??ǔ�{F��q�)	VZ�N��� �6Tj*�%|��{��ʍ0m�v���+�C�f��U��[�7ٓX��^��|U���xE+�m���K�F�=�q��LH��M��"�>p����{KY��J׆��޾}[�z���_7���/�������K�DZ�N�{����V[�6��i�I���w�7r�~/���f����oq	Vʾ���<s���>�����~=yXm�;�.�]��|)���	�<����]4�#�Q4�(L�a���kCK�2u�*��v���>
��m��35L�e{�)!\h��/�f�|'x$�/�Cq�V�[��ɥ���~�g�F2�V{8�v(vGC��j��ޓ�m��:����9�V���y	��#GO�E��wo��2X�C��0�IF�Ņ%?��NfOkbc�j ��p9��Fm�\�����W��c�<^YM�{n�:Ҧ���ى����Qܴ��6�QL+��7�<��Eԫ�O��ZƤ��P���� �A*��)�U}�
��|:��k�yX&!��;� <���Ȭ�pa���ZY���س�U�gx�\󂞛���ׅQ��`��y��(�e`;�
�j��	�K6�u×�P
SD�3+�Cȡ��)��(���r��{�Ĳ�i�'������X8�#VYgw0J�[1��k/�+����\�t��u�-DE]����L�T�\��e����m�W�=���2�����Xp�􅮭f����eJ�DV�7*fx�D�FM�T��瓷jKM�&Õ)7sK�w(z���s_V�6�eɱYiS�C�/�o!�A�[W�����Ew�eL�t�*�Lf/#��z�}l��@U�w�L��B+7��H�reuk݇��~���G���T��j� ~�_�.����.�-D�_�*|F���&2$�Ěi$Ɯ�6k"5��O}�S�ϔ��i���{�_��_�N�ǡN�CIg)�o$��FM��%5���B��p�����Dxħ�`���TV�<{�E����/׈x�	:�ʱ�n���b���݃�6\S�-��0)?����t��ߧYI�%\i�>|1��eI��K(��>9���I��v���u���t�h �k���#pW0�FE$���s�>���Tj�c<<�Ç��W�q��ΖPY]��l��1�)rU�*�&�R)�����Y���\�vM�w6Ck7DWM{�4l&ܐ����ss}f������G������������~����Cg�'y���؁�w�4��߿Cb(�����>�Q�k:r�D�te�����r���G���&��Xv]��h��| w��_��� .�������Uߋ�ވ�>�a��� (5g)��r����D4�X?;?�@G	='���@^-/�nJ���#��jwRϔ6��HC����D܈��a*%��Q+�z\ +B!L�I�5]�/���I�h���?�#6B�pY8�Xi�$,���2�S\��WM�&J`M�y���V<�����t`�x��a.���ؖ5��һ*�Y�=�Ȋ<B���#֍$��U����DF�)y�n�������Fa]M(�e�灥�۲f�DX#n������<$fw�q��7��V%lB��>	sL��GS�lֽ-0��ޣ*��g��:i�U��������r����Yqw�-,7�	���R����E��+��\������_���c�~��~��_�*<G�CB�p�p����F)X��j�ed�T(!�;��jf}�#����J�����d}U+kW�i{��&9��U&H~[py�K���$a�]Y�&(�)���1G��=%d9�/�*Y>C:�W)�{d=�q����²b뤓td���5k� ����ߟLEb	��Ar]<��=x���[^�LZrx��W�U;�%L��N ��C�ip�3��4Z��"���3�;:��m���۷oC��;�e~A[1��+)�w�`�o]"�.]��,5�J��L|h�A�����Q-�;�\����ݻw1Ed��׌��r�
$q���K�^"V���[UКZ��{����� �ռWQ)jY0b"�M+�cmw�Ȑ��|�d�D������Ʃ'X{���w�yO\��m�}�V;źȤ��I�[T�|�{<Qw���#����'N��;wW���+++���Xa-�)��|�K�RK@d�`k�fT�f9��+Do�Dr@�#�x|,���ӂ��Wp/���0������)��U��puF���7�}*���p�Š�N���2��yq��_���3��=@�Z�'G����DO5��ر��_���qbu�p�2D�X1�ZX� ���Ӎ�� ����]�x��~;�F,��\�\��2z΅h">�^��0�	�	�uH�����<�1��RU*��<��s7�jC��-�-I�F����� �m\j51j�������La��)�r#��h��+�ZZa_e )n�"����M=6BC#�(�iFò��������ș��"$�����[c���Z��t ��r0�P�xF���(�>�0By�2���ffM$�~<0kT�������H���SPm�x�G�ڿW>5�`��'b�R5�8H|n�2��� 4�H�^�9�Q,�0�r�TZ��{R�ߟ����'�:
����S�����"�|����"��^u�q<�+���S�������6�$�٫��ZZ�li�l���J΍��w*���ۜG7vK����y\�c�����Qۚ�Id�^�~�H+�BcIk�v����(�)G�$�߃_e��~�Ռ���Ky�~����\��#�[�8h�^�B߫r+��fڶw��?Z3�5b���2RXY�h/�P���?��?�=np��������l�����5u�U
S�zB�n���I�x<�<�'����rT�:����P�a����`��R0=�"�1��{��}-k#I4A���*(�(3=l��",1�a�o���Y��c�C�1�j2L�U'�&��ILr�l�+��P���g�+C�CB���긎�}�����bd���VD���E)�55P-cJ����$�.x/�b��w���#*�,Ҷ���!���a+	=��r% �3�H���h�`Ρ�C��v��q؋BU��p�	;�?X��1�aŃ�]��-����S�*r�>��CH��H�/�_�F�P�����G�t�*��� J�[ORɗ���ZA��442��eY��<�E�(Jn�Z����B���h/RP� *�(�6�8fA����ð���/⼭��D��؃�@uLGӝr+(���?�/���/�(�H�޼u�:tHH����^f�ԩSgϞ��>/ۛ7n���������^Uғ����c��|�I�6~�����/�]a�OS\�;w�/�~��[[�޿w7
�[��|��\[�j)G�0�lR$�h0���@] �+��rJee��n�Dڭ�>��hR.�SZ�)�#����Ք��^���D������+\���h��w�Ŵܸq��.+
iOz��GX��|���NB2l8��$k�Y�6�{��6��ح�m�_��Z3%%�op(���0��.0d%����"��?��1�U |:�uq(;m�,i;�1���V�V�Q��C���^���Э+h+؝����Q���pw')�����U��������ei������:�.��[7._���~��[%o��6��s�=�gQ �l���z�=u�.��:������e�G ��u�x�ȡ�҇�`XwL,f��k�9�颾�M�ڋ.��'�j�S[�tY[$m���P��%L���V-
F�����&��3���v�pXH%�5����ʔ�
'Q��A;���N��ʘ��'�Z���?!~������	�,yVm�;r��xyZ$}r@X���Gl�8��G�7i����#k�Wq�-�B*� ^�C��"�&��Bݥ���Gͬ�����:Qh8��Am���DO_dy�@CZ���>š�T����t�m�����8���z��������;����\��������~���o^���`���>�GВlLTY����5b#T��gv�Y6��1�����]���B�l�`�(�`������H
�j�kB�+���Ӆ3�k���n�UVV�^�>\#%�bFWF��g<�(!ԺȋinM���`p[���ʝ��U@D�1!p�S�<����G�^����^8uZ2�ұ0� ���̓�+Q݇�nno�?(MNa0�����&iYs��B�l�����u3��0o޺~��UؖB������cBwܹs�Ǜ�5��X�7Lއ`�hS]\ߒ��xH;0�Oi��<�K��������;u����7o߾;?�(>�Jt0�Ng��J�F��t�Ĥa�,��w��]�2��!����<���Q��*��``��0�,o��\�;SJN��0�}�+���ο�}LEi�}.�F��Ȟ)ʾ0���������w�����~F���f�>�~us]z@>rPrd�2x��N��ӡ�vE! ���su���`�g81RoF
h���-��H!���pD�a�����?L�Y���[6�*�H6�H�U�SC���1RB�K�>c�!�Z�߉��������PE�FfUkUDi`���&|���< �Yrv�wS�@ڼ��P�0)a�Y�ㆎ�ւu���V�xO�k�=�Z��ؼu�����}|f��+�i\)U��A�
s67��޺u[T��{]2��F=A�SL�sa{n��i3�A��ֹg(������bn2ix0*�%�T��X��A~�u(wNh5"mk	�V�8�&g��;���,����nĆ@t��kR�1?L��l�M�GZ
�x�Fg��T����V��X^�#b}4��CS����TG�.,,a�E�p�;�@�e:-�N��bN2�H���u�$�*j�р�� ��0��E�e�7�����g0����X@�F����u�G�3�;�f�K�d�"Lb�3������
g݃�ϊrok1�)g#oV3��Y�P�up��j��c@{�ʔ��ȥ��`���[��	�6N��JYi��t�J=�E2�6��q㵶rN��A��~�
�C����7&.<���x���FkB3J��s�N��[ϑ�:8��\6�T~�0q�3FYI:s���*�(Zț�}hh��|�����g��A�����3��\^^&4�`(�uT���ױ�!1YD@s���SǏI/-���F<>F
�[�
�@]�EՅ7a���}����6��*KƘ�r�_ܝ,*�W��溱��c���Z���|�2�����C��)��yN�M�1��4�~��+a��Ӫ-�!���"�XN�����ne�f8��pB�2T���fC�,�f8g�A�����n!H-(aC�V�u�����)�J	4@�'�ҵ�4M�ԭ~x#Y������%���b��d��8	��U�T4�8�I>]��a�MBB����iZ߻�J�$�=���b*_�{g�n䮣�6|�ϣ}�v�$sWK,}�=�/L�;��`~�-���[T�&��O�G�������]�p�6�>���O�1�s<.ԙ&5�N����������*�r�����M��(c#��_i2� M��f��=��a��_/�uj��z��  ��/E=���I\X�41-P�,�5�`b�I��?��<鲔���j��&�,�G	 �ɲ�nO �w��[[� ����k�N���<�o���8lbX�Sl�fL3��7n�3�]�Z/��v�8��U�큞2	���P��0#�qj�v�P}g9�zYˉ!����Ov����E��燍�������=#ݕ�b.A�I��Dz��!�7�7������#���ϟ�����0�.�/�n�!��[�z���\5���@�.G��b]�rE;0
&�y��'�|�`1�����3g�Ԙ�z!��q��%N�x≃cؗ.]W����K������	4-!n��~p/�����4�x��X���"�Y
xSht���E]e�J>i$�van��%���6p!� Z_�z��>�t��p<��o��F�E�������þ�#�%0´����-�K�~Q-��St����|�3xjms`��Ξ=��+/�
�ǘ���}�g���#���ZBJw�2|F�B�#.(v���Z�_V��P����h����&x����j�TB�ZՅN�,$�c���!$i5ٓ�\D�N����0-29�Iw�ya�:�JN�ݡ0�;d�R+6�k�]������0��J��x_J*�`�@�Yn5�%{�G��*���r���0�=+��ڌ�p
�F��K���GK�2����������g��h6�뇾%o�?�.M��(қT����'��HmN�$�hd��r`o+mH���>�T�}Q��W�[��,J��׾v�ʥ?��?x��'q�}������w�wS�q9�����q��*U��C��K��m�8󬡦�G눻Q3�"BFe��6����"�_l܁��Q��z��¥��k��,�(f��PW+%���Ff~�1HXv�U[<#(��嶗��P:��L����)����!p�P��`&|�'(��!����j E��k��������e���b�Y��j �·!�DI�s�iy�ǖ���d$��k�C�CD����%�aC�C`r��C��gr�1��Ycn|"4M�=76�=y�	{�AMؽnЋ��rRk��0�j���l��\�ZaZ�|���XYYGR���,�8������~@��M�{�c�*m=��w�[�j���u�KK4a<i@M��q�|����˥2'�b}oݺUknLc�L�41h�����Jב���KEGV�W?T~q��Ov%��9��v��d(�n>N�=�7�<�0�]lX�Ě�Fk�=���ty���4β�1�/������!Ҁ��+�>�T���i;��{�!H��oI.���Z�|s��(���z�����0Sd�¡��
f@�$����<�>*�,a�S�B�%�	]0L>9X���jN)��m=X)�4W=���'��������.�px�*kAI4%�s�ᧀ��a�Տ���2uQϗh1~=�փ���L��<���95bSW^$�a7�YW4��S�4�5q��oe���}"V�r�#B�p1d���!g�u����<�G���m�J+��5=�65c��;�@.��P''x�>�__D6ܻ�"i7 6!f������R2�Z}ަ	'�4JE8�����!5��*D�ρ�<�YAu�;Ա�Hfx-<�&$ס䥬,c��g�Vahn���Je�S�˔Z��柷튌��6�T�n���X;�$
5��X	ʢ&�p%�qHK�����ڽ���m�}�߀���sϱ_r߾t��P��L�r�i
�`cp,Xc��S7�I�B��K�K��eqӕ� Kr`Z��bC8�Z2<���.\T��U~[I�i�;z��ѨD9n��krl�b��9e4,GP������t��x�~�<ym jf��R���Ի����ᬫ`2��پKP^��^�~9&[y���Kq~~me��)<�Qb(�8T��v��Әp:�D_cp��׷����yLD��!�Įì�#�^��2��kb��<�n�m}��7q�5a*����r9{� P���)r�����%i�8o����.)V�2��_��X[�l`�|pX���K}�ڲ�n`�p��'O����e�ߥ�CYH�J���aT0�q�L_��>x�r��K/��O?�Z{0���ZI�e���#*6p-vRx��J�ևFg�Ý +�	�˸,��I�:l�x��8~rWi�y��C��Js����^�T���iW�Ac�/ZM�:.�:H�z}{���QCĎG8�A�/.��r���,��P�a+N�NS�+�6A'mO�X̰��3�;��vO'6�ja׌¸�D�NP����Յ�ւ'�����ɓx�z�ҁO?{F��[��N{�����cؑFI��J�u�t��Xz��� m%�v���u
��%"����`��p�5�y��v�Q��� ���������'Q�0�Y^�f7����,� F�#����w`aQ�ܓ� ����/��(MBH�Ӓ�Y�aS�vW�^�{k,3W�4�����V������a��� 3�%������d�ߝÞ��p�*	��QrП���ӎ�b\�M�1gj5��:�e^먘H��9Mߌ���z0�nb�oߒ��x((��L	@��xU��{�X�_Rj��F�V	S­oݿ̈́��/�Z�$�q�H�"���'w8*;�cr!d��6L��7��{�����v.���X���g�]��gNBTi'e>�V9���0��Z���o���"Xr.Q�R Y�6�V��ݐ�v�p��Z�\L�`�-ߒ2���U��;i<�Q� ;����|s�ZM�`{c�Jc�<��ȋl<��V�C_M��|��H�NY��|��b�QY�>Y��
��DUa�0[j|���g�}K�������E�-/O�������K_��t�A6�����"�o�z����7o\���,5L�}'e��S1J�?���W6��^�%�Ӫ.����^k4��2�R�w���έm�o�n���_��+���'�'��T�A�׷�U/���:K�(��*�٭���rQ]@��y"���vKHv�pa���j��,�gǢ@�����'V�֝��Db������o|p�m�\�)��xz��k�@��������G}��������]P~
���'��2�5��w�����k�p�>e�KO�%֨��F�G	91��$yĜ4
(�)��T}*+�� �t���`�˰Em�z	+�ՠ�B:�a��1<7y4�8"�d7�{]9D�x5�^�����f1�^׹�?�y�SsuU�#�[E��k�ҕl'�A�������!�߃{� q� �����l]ɔ5X��FR�(��M�硺�3�sַ��>�)ˍbթ�{�5~�[=���6�c����.Ϛ��$�^7*�ᡸ���hZ�죁��X��8Er09����]~Vl���d��@�z�z�������G6�cE������(Y��gUQ	��E�Oݢ�]3�X�.�o���r)�$l�Ig�~K�!����X]L%�q���j��P��w8Bg&`,�d�Æ�y�B�*���D�4����9&���Z^.}��'2����^"_*דP��&��K�q��F�p�WVĔ +7�X�]Y\b�p�@�$`�,��ao��������/���O�
_�7�w���w߻6�����T+� �i���	�m�k�.��3g�S�[�ĥ���l��Dg��Z+BV��ma���s�C3�K��d*f�� O�� �2=��9�s�Fox��x��+^5J��h�M�6�JT���;(D�J�TLǮS��ED�Ԡs�?��*���w�t48�T�����?q��ZX9~lM��>�c�Ee��(���ޜ���	�m����=���X��$;/G�� ����-.,������w޽�޻r���"���C��(����D�D�}4<g&�!�4����As�W>��3{z����vSy$� J������z���4n���6���Q�������P��!I�f{;�����\B�<�����1ٚ(Ks���]r<�Vd�EO���Թ<i��W$?U �8N��'#���1�$JE���#v9|)��0��D9�Hʭ�Q�����V��JAc�F��d�;�o߼����Rr���k�BV�V!�6W\B{�7/Vb�8������&b1�y��:؜D�#�ٽ��sL\�ի��z���+&�1�CT�3�9x�&+|p4��6��>)4�w���h�;/�@��( Z��6�Q��+�[�5�M�ۊ2�!���9��kc�"p&� �K0�JXi��j���փ�\��mv�;�
����S-��JXk�[
ɰ�~@ҏ�6���F�M'ј�V1H��q��0�a�E��	UI��q�;�jul�H;6<���k2+$������o�U|�K'����Z�[LR$�f��,��K�N1�p����}��`�XO���(;�"�.��u�p�YoJ|���S4DC�)R�q9�8E�j��3�DF�f�����D2���a��с��*�	�ݯ�
�oz���\�@2���*m�٦�m�.���ȢQ�Ȳ��<ma��"�˄��<}�"!T
_�a
�0���D���E2��^�&C&��r\U`��Ԋ6�[�H+�*�X��+5�Յi�dZ|��9�z��(s��{y&�a�Ã���P���A�M�V�b�rIl�ׅ�y��@h�<J��H&c����;|I�$�S�i��"�f7�z���fv�I��[{Q4���@l�ͪSHdy)xt�X���|�N�<�h���`�]�]B��Q��c�&���;�PI��y �a-Eȧ�(�4��j{��!O��`��1�O��3�L�*z[�xjZi/x���M���V����)!�2�d��`�]�^�^f��  yOy1X8�&��sV6�N^�����ϙ�m@%�p(~'�q���r�����[tX9�Q>I��J��2vQQ"�$�z��Z"��r̂
�6���\3_�bB���d�A�[4"�ɣ+�%�e
U��cs U..kN,��2++��\��"�xZvv�mǨ��l���~��E�2��|/��ge�^~(���J��zz��+A3�N�����YyN�W�C�^���Ӊ�VPѕOʽ�*��ceg�s̫��9��� 5��Je"��N�P>@P$��`�'N�Ր�m�t]+,�޻w��\yq	&e���L����Ҭ�
�у#��7n�����H�`Uu�+՜����j�l�#�4���U41�&���t��%_¡���z�.]z�/^�HI�;���?����R4�E���vx%��r�$�}�z��E��a��f�`��&�,3Xb�*��5�2�<���d�%)�-� ^m���q�m�Kn�"���86IqZ��#����"=d;v�𠿰О("L�{��5"�u�ԮoF
��=��y��h��}to+��9u
	q��Ç	���PM��"]��W�y�/��╫��k~�)�F���@��&A�뗿z��_��(���^�QW�"�g������#o=7�� ����h���>�8"^��)f��,�M/�x%륯�JI���c���K���������c�1���7on���$`�v�&�/_�t��6;���./�ݿ����r�!�*��V�*�V�7�"V+N�"C'�Q��h���ӧO#��$�������������Je�H��£�,c;tc����{>�E��É8`���S�LM����}lq����wd��?���/��x>���[���u��V�0� ��{寮i�&�s���G.N�d\�C���w��=�3U�O�4��&���46�F�RErX���*�>�8�I��C�g1lG��ٹz�|����u�Aɳ��z������{J˟�'1�R7+1�����p��Ѡ�����A�*;��~�.�EK�h�O~�U����7E����_�����pQuL��bo,��4Bm�ɠF.��$�O"yf��2����� 4�J������[��+ܺsw{{g2���8�K����y޿vx��(G���ܸ�|UQ�7[Ї��f�L�������_�*%��x<��P?5I���J����J��ф��.wou��s����LQin(�wB<i�W___g �xU��s��Z�Р��ć��Ɓ���3�d�f��BJy# va�'!#���aj��O%���n ��š*l�a�\��˩���tu�_.*���Z�O¡��O�O�xh�y[��!�g��X�ggFl��!$�aO͌>���m5b��Z� 0-P.o��8;v�e�:��6p2�g��d�lۗ�d�M�*^�FȲھEV%��ry-������,�`�	���Y^��F������4����ދɴ�������8�����a�=���3�գ��믫lLj��R�yL����j����1���&����h�u�4g�J3!��]엦M�`�����d"9}Šl4+�_F�����rq㈠�����՛�c��T�4'f�W�O$�1��V��`�7��i���c�t���AaG���D�~�$�<�ڳ"J���2#P�b�_��F����#Џ�\P{pxD<?�|�6~����s?�)����"J<�܎�6�-�ZL��{Z�B}0qfægQK��%ў�A�g��54|��zs�*z��W� |�8��T\��0rҋ �X�ϓ��C��G{�|�G��ߦ�.�"O���I��<x�����^*��eT��4��\_#��&����\�W4���(�J8��h��Wi/�#�#S��cn��gX�,��k��q��i�t�O��٫�jl����BO�Fl��6��I�J{-�E�pVj���WB����k�r��!E�l�H��k�V�"������YZ*�FL�����#��ojs^��vR�X�]C���N�2=��i0׈���K/u�+� 666D*�:S�P�paM�@!��1ìB3{'3�w�7,L�1~i�+7����̳/H��emf�k�f�Xj�<Y�[왖�	m�.0�z.ij(-�-���^	��M�]4wf�tf��V�:x�셡Y+�Yn:������ SH����ҳx���h�R��<\g�Q��f����)<�9M�<��b��桳7��mǀ�v�H-B�|���r�mR�)�@���y �_9)����DE$G��pߵ����
���}J���'����r��''���Y��T�������13�a8�'����sR9��'t�w�#��4��4���n9�;�u4���KJOi�ܽ{_�F�������>��g�ĕ��.f�Ms�aQ=D�[K@%5Mxknv����`�J`*qp��r!��b���zf:�o�Sl�NInR��OMJ����f�t�3��x����?�*������0�L�8��y��$�d�C:C�F�e��3_�0�ϯ߸F�`}_�F���z�8a��b!�.twv���E��S�E�w�x#)�Z[�ă��(a�_�'�
U��\v��JJ �,۴��̈́�� �L����������!���jܽ{�-��.)�],�Ν���>EJ4(/��_�V�u����*��.o����^��8��F�����8������'Ϝ������*l�䄢PP�?Q�c��ȇzNѨy�ss�N�"���S��vU�c	T�ȉ2�ƃv���3��O]<��o�;�����88�Dzde(��Ib�3��
`�@��S���ŶN�Ġ8q�"��� ;�V�
Q1��:�I�Lk�j�իiv�{�D��0�ɧVĩ����Ӭ���w��Z��e�!Z̲T�)i���^����}�����B �lmuQ��?B�t���u��;�&�酓[�����a�}{{w��/&�A�'J��ĩ�E����;�t8|x�v�D�����*Gv��'QK)d�0�:j:��ڛ�)p="�It�
�֚��J��G������x�J#�����'����V4>�&�ypp(������;���e4(*V�ri�'����@M��K���8�i� p�'��Ț9�j~�����.`�3gҁ �{#�[ G��T���Ź��W��>~��c:��D�����/����7��.>u"W��Fd*^m��>�"R̄�8C�!�F�5f�'Pc�H���9�X�uy~�4�c:��8˝(�n�����N�:~��Y���wn��w�핕%`�w��#�)�%���:�᱉ɛ_����Q]XXT6U��F�����
��p�x�����J�}��>%�)�@��jܻ�H���`
��_��_ݻ{��j� 	�fn�)��{�n�¹�(�8&��K'Hc�M�@!��=q�D�WĮ�eO��A.�1��B��|��g�i%6���-{��S��,-,�����8��Ւw�57ǉ"4����i�r���<-NE9����Q�e��f^P��l����y<�3��$�&�!R���W?��]�|�����lu�lJ�!*w�����	��q�J��%Hs�+����K�ϟ9y�����޷eŒ��4���l�I^��,�,���˿��#�y��}�nm߾}��<S�}Xk4�_�uL7��f�@:XTW�"�;^[��5�>t9yI.gA|�"���Cz5m��
nJRq$� ��p�X�}�D�/˾��r��������*4��^�!ˎ~j��R@��O�ZA�KC ��F�:�b��,�oW}V=A%|.�Fs�d��U��P���;���%9d�t,B.�X�Y������_\YY�-`���o|�Yo\�r��)k� ݸqC����]��.����]�F걑��V�WZj�zi
}�%+IzJ����'0=�t�������`U55�|�CB���^1�6�f8
�g��|.�p�FAl1qM�m�m��G��V�}3��n�Ifla�Ƒ֏- á�\	�����BP:r���d05���<�C�����k��C�)6b`N�V��_��z��������Cs�s���ϊ�����5p����kq�+�_�6��dI�9ZX��������%�/E ��8��!Lt�#
6O��L���J�Ft9��r0-��d��2�J9��ʘ�B=3��qq��N>w����x5����	;ODW�h�����g�W��O�|z�&q&�s��� ����+e D�����7on޿�hiY4�PwST��_���<������*�>Rv��`��Đ
�_�	����V�H���t�(@�Z��,�_�����"���J>C����ronI�õsb�s�� �!�����v�ˁ��D�ۜ��uH�}gFId�M��5;v�rz��l~�(��C;��0�x!g� Lef��,cGd`�rJ�Q���h�*��k+����`���1ʣ��f`�sm�0s��m����2��3��Z�#�(v�ʜ�K:f�2
�N�Qgs��e��P I�ņe�ϩ6��y)���|f<�kh��$f~�5����a#�yhZV��.{�\]^YI��/74�=�{0A@�g������>���YkB��Όpt̨�p��96�s�|�h��T����̸ÒJH���Z�����j���8˚�2R�-w����D�|�h���I�Q\�0��Qklt䃮�i�=�V6��i�ב+�`�]��図yO&�l��VG
���ഘi���k�����L�����wנ�l�=0C�l�.�a��KF���܆�6�a���~f��r�f���cH<b3ш�],�-	������(�8�?��#��uh���J�2�s��qD�BUh%��$h���P-�X �1�#�f�8�OM�('C�$Ba���VU)?l7�#dK5x�\���d�L����pH��i��Q&ʭ�=+�^A3+_�����3��t̴vb޶���.���Xh*f����Wp&l�.�^Q��!+@�Q��p��=b�XJe���P�uX�-L���̌��pP�F�$��Y@�gf��$:�r�����̴��f�ҫ;|l�BY�`��$ň 7��6��lP�G���MV�g;3�*ufjѶ�ƬXC2B�� 4�V�]d�KG_�3�'Ԓ|l�������k��Z��
�w�2�x�B�@?�Z�ūS�a�ry�%��X�����2�ʌgX��Y�o_s|%o1�J���ڳ�ș��,=W*e�[�n9
��3F #;�Xn%��M��C���K���Ғ!�Y�1q8�
�:.t�,�@�҃���Pg���UJW���~ѳ��v�T=V��H���]�$�7��e0��Fn���t�*��S�%/��3ψgC�$?Dʦ(���/|�����v�xU��O�((�Q��T+��XLU�Ztɓ���+i�J-l+Ne$�	t�dz���4�L��3���K���jF�u�`�;�KȬ���T�u�ˍzK�y�p�E�}Y�EOt8e?��aO�X��'����m�nMj�:�U5�Ѫ�P��Vy@R����f������ cd�\�]��{��i�?<�܂H���^6���r�����ꩧD���������x��o�Z��?0�a�e�Q-�9sf}m]L�D z!����l|�zs���M����)�yj�N� �S�@7z
ju��{��)��s�α��Q&��&4���������/�u�Lq˾	�$Ky\�[]��:��ш��
�W���-��+W-ݛ_��˴X�S'onn�&ß���{�����n��h5�My�����Ct���@�j|�L�
��c�k:9��O2��ؐ�J��e8-�BT�f�$S����Q[VI�A�����?���:]`�ϝ;����é����,�0W�W����Y����A��k_62���]|��nܸ1E���L����M�Fm|�?����~&2���dw��ϟ?//%v� ���@n}����p���D���;nllȽ<��R�� �#Ԧ����23dF�aY�6Uf�����ǅ�L�}h�#�)w�w@����T!�4�H�V��?�!>y�,�W�.]�$k��~L-lt<�>�ƓM�����[���3��O����T����ַDr��Z�y���e�R�όH<7Q����>�h)K$GN��!r#�J�$撋eO���N�"/:*�$�_��e���K/���q���r�ʿ�Y�^�mZ�W 5��k��hTk�?��"�\XXB���W��A���(�5�bDe|���3E�.r��.�"�9u�|s��,N�<.�/�3v��q�WP����ľ���'���|���ݝ#��׿�uyY��ã�!��e��#�օ��k�HIaCS��oF��u��t�#���$*�����x0[���{�Q�QT4a4��-�I?CSB�m�F�����j�쉍~mH��F�L��cä������&=���&Fr�sKj����=�E�I����'��~���_���������V�7����[����ޏ~���O_yᥗH���W_�'�M���o�����;�L.Ȏ�B� ֐b�Ә��-cҧ0X	z#\����/1P�˝A�I߰.��nA"��ņ�m�:U��,�DW�U�gW>2C�<'3�*φ@����O:�7ZL���}�CL+�<Oo~MAU9P��ǒ�J��o���bf�Z�"+���!�W	�N�vl���
�+��&Y9�rZ���Z��`�?����'G�>8+)r�b��F��8ڸ3�"����T��a+�0"Ȩcv�Z9��U�S�TPɄ=f��x���o3�����s�H�M�"f�7�7�l���T����*� +[�JrF��HI�3O20�Y%��A����x���20!&C;ZP	� ��Q5@�����	�d�K���lS�@M��i�$N�j>�&�E��1��hI�o=��JABl[�Vډb�k���˸ME�$*�>���_����JY�D1�.W�=�֥��Z��-#�(ImE�����6癎��N��M��1pג�df(Da�:���9pLR,��j�R�M!�@��=#Z-N�`CӲ��U�(��QM�qt�h��|�C�]���?b���|���$%�?S�KV���'bUiζ�v�z����E�u+t�=S[��-���.6L��9F��e���Q�XI��������T>�.�+�s��6��@�O�����7�"����b��'�+�6�F�0�)��WbHˌ�c��P�,qH��*�xdfW�h��(��*BO�5�O��M�l��@�ǄN`�wvx�D����´f�&1Q ><��#!�Mz�A�Y?9��i�K�ə�)r,��p=X�P�rhb��-����+��1��}3{+���~mz�%�6��ɿ��Bq�d26�%��I�MO'�[�RK�I���C�5?�����Mu�?w�5��
�M�8��ׇÂ��+割h�!^�o�+���M3�)L'Ju7o&<�*��VK�ߔc�����\k
��L)?CC$ow�(�������,�}:"4��2m�+���)w������˂.�;4�i���́R��,��F[�t��}i]�s�R����R�3o��+�Ǣ����z�<`L��9��Z�|#w��W慗�Wm�1@�ZN�KuR�>�8X�,S�1+����أ��J|��Hs�'���_2�(h=��f��/א��ip����C
�WVT���` ;-n�[�)9_��-�V`�C�ı���O������G�cڬ�\mnޝN�i4��J�j�jV8�����]/�U
r���-��͇�}7__[����V�><JY���(���띖X8���ҵ��4F��q9��L�3#�d��{��ی6u�<$,S�gN%�����r��z�*��p�`���
4���N�E��3���ѣ<?�t<gk�V�]c)��9�2���y��hms��{��@����������:��©cW/����VA]����ي_��S�O����Μܨ`�ڑJ�Yy�Z��c}az�}�����Ǉ���s�+��8'�$
�i��z��K�=�,�4��w��������f����so��C��G�?HA"M�$�6�Ff�VG���G��<:{r.;��6�62��[�'���Hh�J����a�8F`w���^G�A~ *�z��mq���Y��O���xd�t���w�����{��n��0jA!�þ� J�������p��{:�3�&|$���B��X�X\;)����|��������G�����ZRJy��4���=�-PN�9w����~G��N��u��v���_?>��GA��?�՛�Y��Ǐ/<z4Y�5�d�:E>H�Q��88zTozG��څ3m�q^~���`��{שּׂ��m=t����iv�W��q����b��b��~��Z���QO�Vm�ה�={��Dn[[[�I�Q8�sT�.2:��ƛ�t:�p�x~�Tà���,�~��:���w�T]'�ݸ�@�-J�f����#8փ��)e6ILK���ਿ����,L����m9����X��6����PӞ��9��Ϸ�v�h���-��'ϝ�GO]<?#����˓��k7 x'Oc������7�֪��$r�q��|���	���3E��Txp$��I$�Nl޿��(r�}p�	j5v���ӿ�_|N�j�-.�&�C�&�>j6�N�..c@�%��kN�9�68�sM��`�L5Ic�Q�~qi�4�H�Wʺ5Ŝ�x�,�X%��{{���3��$�f���G����i\n�r�Q�$#�+�wEZ$���jwn��?��EN:
]҈�}X]]���:ޗ�x��H"���J�w��}�����5�Ϭ�&1lW����dk<������/�Δ�����ۓ�O~��'?O)J��Dѽj�r��
ĦM��$Fm���ވ�[�7iSx���q�u�]$d��ʁ�*��tW8I�І �&��A�4�6��5�v7I;^W%B�J�,c�s= v,4=��G����|k�\�·�]�5#��)���H 4Mp|A���hH���]��U*CUy�5š?�����ի�|R�r��O_�ؗ��'NN�u ����0#�ȹ��Y��a��n^����0�;u�Z�C�/?'�3�����ey9a\B�H�f�a��c>RNM��-z]P��+���];�����O2�*2&���l�Ϝ���W���&��b���P
��m����L~�	A�Rr�VC{kr'A�E��:�9�@C�����gh��Xf��(3��aX���J(>b�F���F��Vuy%qlD���w�֭�x��D�9�) �
����]9�W6�j�^��f �~������k++"'�<��k���O���;w��.��lz��!����p������nei"�P�ɕ�'�6s��`��
�p���"���&��B�pd�ܹ�����e=�,衣"o���=�W�;X���%�q��q>NV�32��2����U���_.#O��V]��GR��HJfy�2���wz�9�PTa�m�LaB1{2�a�屼^����������󸞨ʸ��J"��j�tjs��
�2Z���fl"%�@��1�
�P���7L�0�j�hT�&�T�gy�����LI�D�(F�L�l�$�Ŧ�����cvR�p�ץBU����%	읙<�tjh�e�k�v�_V�^�����Tm���&
��3,�[�Ddh�F�h	S�����C�|�_c���R��;���7Sb%�?	*��M�mw���Y���<�B���[��!'+���}��)������[��X#��#����j��&��x����R�.W��&fԤY��×�_(���=bz+7c=J�[���[wLv�"�S��X(��i����I��<gn����VN��QH�ϐ���C�Tλ�*�)�.a�y\	���c��W(�Xb�2��`�;�C��$Q	�6c�M��ש�]���s���'8q��.���)���˿���:�2�RZ��
3�I$Q&3z�h��$=�*O�Oު2����[��w9�+)^�<ϬM���'��b�����J{�����[�� �{'��掘�-	-fj��㔉T��CN���x>8j�K3��!<h��VlJ���7�+-H/�:�3����z2�3+���3�{����B�3�V&���t̘$Z�����B�l`n��0'��^��d}k�a[xqLJ40�6��MQ�U��f�x1?g8q��S���W�9�3���r�>�8.i�&��/��43�ٚ����#6�yQv3�:�'#�� Zq}�����ь��3g���䕑�I��=G��c�����0y͔(�;K��d��|���*V0���V�2�$�d�p��\˰���>�"�u�]�7$�d�d���%�&���w� !#���J<l�qST�H�s��I�5�T@��3.RN_�-�+++�6f"$>�7{�mYZ������C���0�1s�)6���=��)X�C��I3���&}��P-�N��lh�����-yٳΞ8q��i��2J�&��t���) w��D=Q����{�c¢��*`D���cp�y�	���h-E)#�����6P�5�]s�o�Sಲ:��<`Y1��ʥ׮]؀���sx���ut�;��ܽ���UJ�<���/��b�y����� [���4����1(���$Ur2{#���k�A N���ƴRB����w=[��)]X���*����@`����P;L$'���e6�O�9#Z��菾���~�+_�N��#��Ա�V���$+�:T�t���^�I��[��}�%!A�A�8��C��i�g��hS����˫��Ά�$�и`��j!�`Vd{�yD6�ד��?����)j�����{�O������4��W;;X	�ĺK�����g='��O�
N�ټ�~�R%��������@yz�ũ����ِ̬�y�+W�@Y�������W�q��\�����<�nK�,�D��S>/�S��c��կ~Eĺ�/���ҭ��ن���4����?�D"����.\(]�
�WVs�Ghd>��YLʭl�K/���2#\3�*ҐN[�h%x@����ǚ�:�]�t��w�?��'3��rb�&�zr͍�:��S��h��V�6��z�C^�?��?��O~"g�����죧q��V$^���J���ssrHE��:БaU�xG lm�t����G����[��f�wF1�@����h'"�5Q�0+�ξ<<�*R���^:��.�/w�'1��#� A5#v�{E%F�v�Żx�����E9����m�DvP�d�y�O-�āXy�)k�h\���y9�R
q�@OW*"��e5�x�m�����U�O؎�ԠJ�=��M0]�ܐk��Ɨ�����B����Lۑu[]�$ŋ�'���la����m�}��s��\>!�+�] ��d����S|�@��HR��g 3�C����9�9G�q���0�����kO���@��O|�zR��7��37(E�5���А���7�.����'�1���W_ŖU���w�j��P�ڪ3}o��l8��]��h�}��؈Ԉ�R�8O��Bß�LS��C��)6�,�����|ޗ��;+!��e���al�@�����p�3�ɐ���d��.׌K^��i��專�8}���;7y;��.t�ȶ��z���� Cf�#4�`�-�;�/Uđ��G3���@h2d#�=��'u�j��^ē�c�k,OY����
�YT4Cf?)�rF+�TkM3�[��vJ(.�gQ�K4F`���u�D���%����hH��b����B+q:���a�����L�=A�ܩ(	��1��Ju����;,���$k�Q��8~���20׏?��f�mg{u�'C�26��j7��I\\^pM�:S���OuF-������$I�BܥM��DE��F���Cŵ�Uxޓa���z����z엫����ia�Ҡ�LD�ㆾ�=`�>�쪢3J쉖��M�f��^�h�"4ݎ���1��Ip8i9$��]��t@[)�;R�f��_e�ʠp��)/e�;6��7�r�ڿ��D~����9eC�H���; 2�Z�����'�]���U�����|뗬�0��)�����^fQ-���	�F�!��U%��KƖ�\3��0�c.rj�9h(M!���{��5�M&:�}���a8��W>��>ώcJA�ז��|'�Gd0�Q蘖J��ւ�^��d43T��Wǥ&t̴�</�<����B�tS���%2�ӑ(w�o�b|A> /e�d�T�
��"�k�fM:���\��M��x�[��>�m�=���8��"O�P�������M!@}��.,&��s��.��Y��Vd,�������)r3�HG�Ď'ɍ7�y��A�x�xs���/V�&�0�D��� O�����A.�^nPl�w^��P����P$��)���#�8�shIn���@�de��j=�@{F�:+�V�Pt��E�Q�wa�����N��q��zrM����O�y��i�tU�jIᶱ=\� \"�T�����
f0��e�.8k����"F �a��,h��Z1�x��RKt�5��v4�xr{ps)V�;P��W���b�c�'�H-�/O�[9߫~F�V\'�C��\�\9k ��~�ǻT�z0�GE�!��j��t��x��RK�V�M�����.�n��:@F<���Ѡ(��LY�(�XpGY�
w�D1��1�ʤU�PRg�Q�m���G��G��e�"wP��T����f}����U�V90-�s-ǡ�
�}�`��`}m5�ܽ�ha)���tr��p$��Ր��������݁X5j�:u�� K9)ߔO����2�V��:M%�H�Z�.Ή�77��iϯ���{�}�1�����%v�r��O�XX�5C��hg���u��n����8rq!�	�� iY	�Q���mll,,.�_��'��8yc�x����oh��� ��l봾8�aQ���d$���`�DnO�������!���^I��@O�?}���R�C1��
wΫ6[���Et����)
��p�ם��?����?�������[[���j���hS\�8�Zs���8����Ш�>|��o~_Nqo�|2G���g�1�-� ��&4rN��"A�ߨ��G����N1Z�v����NS��M�M��}x���\q���������7�O�|$� ���w��bg��eog��V]�9j��KY4Lڹ����9���?��`�ߛ=�s�D��ˡfj���k|9�?VV��)�N|��k���nqO�"��\q���>p�O-�<��λ�E��`�����'^x���N�=���i���߿�#�{T�1_�hy��?�y��+�ǖ�$�I:�w�\�|��I!�P�[���Ȟp*���ʾ���X%Ҭ���	QEPD�o��כ��1�:I�w���P�&#���ΞZ��
�3�-�=�\d�$/mFCT�6h+�6�4�B U�l`��^��t�ls�$m��+/�B�.g�nokT��j��m˪b>���U��EӱطW^~�QA�31��7u��H���_�˫@����iOu���T���x��4W� ��y���9�/�]�)o��l?�4����U´�DA��ݻ�{���P���p����kT��Ş+��zu)\�a�+e	w���ͅ�ydj(�4e#�j(�dfZ�C��#�mmn!�6�˝`/���W��wo�C�y�_�zU\��7���c>�]���������'�&r{���S��5�M���������#������T;�.v��O3�`x�!B]�|b��hS"n��7���VG����p{���ޖ�A�'EJ�hvX��Nˤ�;��`��pv:aQ�o�3�Gt�	�g�ʟ�ֹff�2����1���0��1�/�̐Jy3�t'�l��1A�����jd���X�
��ڱO�����;*J�)����*꩙V�|b=����
��;��_^Z����}.l�>�Oʩ�+����"�)�y���Jo \VvT�g>�q��_�?���w~�wN�:!{��k��e=��7��=<C�.�3�U��һ)<��`�wv�r�B��@���jܒ�)D3sC~-�8������%.�������iA���e΃�L�dnК��2�1��UB�C���6�ƾB�!|��I@W�r�8�vƓ���S⟬���-��w!9�ڱ���?| ��Ro.�8J�*��G��Y0g���K�.˛��ƚ���)�V��ؑG�>y�~u=��D��`OYt��G�B��Cȕwvv���DI���zM��D����yn��N�h���'+��@�[��@3I��@^/a�{��������v��0�э�g�<��ؔ3g���lmn�r�h6������B�s���}y���Ge�)�p�x�󼌁K�_���i��*���,�d#8͠4�Lb��3BW��"�聞"k��/���R������FaA"z�B�@����P�4�CǸ��F=
 *�4�c��$fZNI�'`��,	C�ҳ*����q(OM`ƭPI�ʁ��%=\�82��ө�&�vp�����In�]���*Y�%�#.+F�������!�&�8�[�V��&�
�
�����όff����}ߠU,���M㓞��
��)͇^ZbS���#:KD�:u��WDBr�)�H:Q>�I�Ժsmq���Êg�IҴϬ�s�h.1�.����ܹ3{{����WB���J	n��	�:�yU�w��ӊ!�|�$`Ű�RQ���Ү���
� 0w`����8��+%Ϣ��&Zq�ɥ�bنK���'7���0���T����d���5B�A�/So_�3^9w��[h	����A(/�ME1Q�j���p<�ث@%��6 �i���`���9�C�Jj:��ؓÁ瑹Z !���q�na^v	QT5N�=q�5�2+2fb�~!/��8��+Mu�	\�~(aœ��"˕���k�~�`ފO�(��ф%��0;�&��PeXT���u��T�5ͽ�G
�gq�����rK�����޼y�RSQ����~���O��D�L��U�o\�������T��͜i�`M�z��s@��c��/�H>�Iz`�!Y`���h_��C(�*\�zߜ�F�����j虊+�C���j�}��4|��`2�
�f�uƢǴ�}<��3LV�Q�.�ZQ����B1�d���̰?fXf	�-Ϊ��<�B��*� �Y��[�b����؟��a�Il�Qp�^�h���Ez��B�&]P����<ˠ)�2�c�(���qm��d3�J8� ܑ2���ܯJ9��Z#�� 6��"b�!���!�,�Ȫ�p��9q��7B �Q�crx5b�V�`X$GC��B�xEW��WR[�PB�G����R��
I��[�;�xp�:?�a#y'K�{�DqI�,O���(�\P���-ݺu+����B���������w�*ɺkL��,Y��Z?ğt;\[�+�a$�;w��SWN�͜(�|��G��jf����#��bnú���.��:�j�1���\���--4��c�F���`&I�Ȼ��,?���EtEy���˿�{oS#Eh:+���c��D�x��VvX�gT�$����r��h�O������ٳO_~
�w�APN��T�n~����VO]��rq&��I�,���ɓ'��`Zi4�?+���흇���=~���3�O_� ��'>���es�R4�&�c��nhn)������Ivj�P8L�Q�O�g})���������e)\����3�����V��z�7~��f"�<Z��Ϝ>}�FU\��ǅ9e��)�5j��Ν;I��ۙ�����VW�!��ů~���+�"i�r8���a!�ԥy�I���T���{Z�ϵߨ��#k +"�e��	�˱c`�?ܓ�z��W�3Ͽ�yh�������:�)KD��Xv|~gv��i=�$g�����y����w�Ɛ��E	u�In|x�����o߾-w����8:�٬�H����|AO늕j0b�	����B�::���b��Cw-����_���B�[�\�+ly?�� �)�^�>á�r"p^q�����x'~t]^�ʕ���?�ɛ?��it���C��;f��중R?a���w��
̀��f|�H��~�/6D�-.��:ܾ��H�K���n�<,v��:��)�7�?�����cǾ��/_ߐg~t�<O� Ѳ����ַ����SO]�tI�����~���֮���l����ܐ��#�0d� �,���M�n��D�ɧ���TlG��ًOi~����"�KАK�s�=����	�ί�}O���o���S�/����#ru�uVW����Vnoo?�| +O@і�
o�����f��TO�e�G)�$́뇟�ꀐ��U��*to��>(~��bC�ߥ�����e;q2uf�<�O�ż0��gt%қ�M����"F����y�˶`k�-�0}L��h�C,S�a��	�jQ�4�g��EM��X�F�v�/[�}6��q�O�^u��|3X�	s����L�h�k׮��_����W_}U>��/@��k�k\g�z4ᛪO5[o�1���/ɳ}�_F�HM����k!�&�?��Os'ӹdS}�2�Be��?�ge��r�f�N�I92�e7�0f ˟�?4�B:�/ǔk5�À&qa�|y�Z�i����y3=.�!�`a���ZpO�F\ܷ��pZ�
H�V��g���'^�����y����;R��ݲ��8���w�ʮ1+7M˦x�C(@��D���):l̍�p˟����W�����E7��W3u��ݛ����{����G���[o6�o�
����f�	k2*R�сO̪Σ��-�,]l
����k���<�}�����ŵ�?�|��]q�䇴���ԭ�xI"�Zi�z`�d@&�[~);myBy�� ��q��D�y�c��ϖ��rk�8����J��W����aL�1$Y{&l��QYlFn����Pl�������l�Fe�%SE�}F���aR���<��s3������*��횃(��6�ē��#;�.d��"T�N�" ����빡�+�ִk��C��=��A~��c�k~�"���̀"�zN5�H�6~�f��[��%���T%̊_J�ςh�쨾5��Ef��	�L�s:3��PެU�MF�3,��f�^����ξ��l�;�����w¬+i+bC�H�bvIm�߰i�&m3Ӌ͕�H05$���-�f����0n/�q���'SCf�
"r�Y��m�{�]�+�����&�h\�9L�1�OI5�ݮ<�v^Y�(���V-�0�#�-�����q�%�ɵ�L3�����K�ETr�Ĥ�@����,Ń3�Q�1S7,_�����lH%�Y]��ZH얹^�������z��6��$d&+#�oS�mAw��L��YE��R��8��z~5��L��t�X#�4�>z��������֦�Q2�6	1�(��	KQ#<<��+�S�<��Y�YU�'4G�<�,KP�,��fJ��#CO���%k=�8YV�$�l�8�m����X>��s=?��r����؈u�?qƓ�'H�b0�9����b5��\� �fKeف\sbU�r�
C
RG*�*i�������xr9D�O5���������Xv���G��nV�mM��/X�,C>)�����s��"%�<?�GG#�����*"�ʼ�c���i�LeF�Q���r�!2D)���|��;Z��bbB<�|��������^#�r4��S�8;guy~<JB�`[1��9I������(Z-�άE�1ތ�Ȉd��N�S�1''�@�W�\lX����ώc�,́��������&�<s Gi�h���Q��.��&QJ�S��J������z��Dw���\;��Qd�.���	;�Ė�a�V��5��b���b��J�r�N�p�J���>y�����n�1׮�Ae�����A�p2N���cQ�uL�����lc\$��Lkj��e�I%�?T��$�X��-�:�� D�&����39^X]��T���j�w>�u��Ɖ��NG��2�@R��$�N�P���Q}��&�$t<5��H��J��t$E�Z9�����ɹ����%G������8 �1�8N���jgY3�\�Z���@w۵,��5X��t,��\�/�ؓ�2��D�<Ʃ���o/���Ғ��T�s)�-j�ԓ�!Gѭ�R�E1�����?r|���s'�_x�ٛ�js��Ɖ�S�N5��H����c���[+��~?-tPxೋ�:�U̿��x�tr�e��'�٬�^PZ��,W��VMlB��s�VÁ���C���έ�KKk�-'/�z�@�9_�ڨng�X���<���	}YCq�GӉ�?OC޴�mw{�������"�&;}�T�^}�x��-W�J�ת6�h=@/�7q^�Sd�'QFU 俢�ÀI�Z��*ϊ�R�����?�����V5�?{�n޼y�����^{n�QA��h���Y�L�Q\D���as���9N1�U�s�{�����ﾻ��@"�J�_8j����'N��������N�i�s`��I�� Wy9���6�ut�;�?��<���R��_��'_�S^o��y��ӫ��5�G[V/�::��4����px�������0ss��Y��у��\�Gq�����N�t�<�o|��ãݟ��m�j>Ť��**W	�|O�c���=N����k�,�1Eگ$�
*{�Fx��㫯��Z���;������W�^u�کgQ�L�G�; �K�||r�֖�$����������(X�d�ְ�D\'�;�qr~a��_�x�x��N���7����ǭ��4�@J?���O�!i�t>��oQ����=v��#�k�3�=����5�5���s˧���������ܽ{�����+�&�㷷�1E'�^Z�k�������׮];}����s����-e<9<^��6݅L��ǖWz�0�6�)�;���/'�=c�&^/4S8��8x�8oni�;����\����h�vXC~$�'O����1K1�����@t��nO�Ӻ8GK��	�$��ų����a�kg� ��Aל�mf�^����Y��6"�м��y1F>,	��(Ǭ���(�i�,6�5�[�a�fr
e'���:��L֢o�,?=�eϴi3�B�\����5Z�m���&һ����-�����TO?��Ǔx�j���?���dte�_��$�@����@,����7����<K�qO��XL�n��ʫ������ʟ~��o��n(��Y����z=��<�šӹN�@V��Itj������c+�^}��k��o��v��.1eX� �ʎ�DYh�<kc~I]��o%�r8Un��6gD�2|�gۃh;jU2��2�\ytؿu����0Y�l��a��v��C7����f����BHVY^;��o��}���ڱj�.;6��+L�z<zȚ��}kg�5<B"J��뭼Z�(3��iBt�|�Is�����0O�z�f���#���z=h�����hʪ� :���+s���� O��������y4�:tx��?�ʌy��a���H��teiE�����`�@n��q���#�/--h��,7o}t��s�α��և7>�Ԙ�ʃ��C�Q���yQ4�~u�m*�g��8�S�.���_DNAIYm����Q?�J��K�Ж"�Loll�
L�D�4i�=�b���77��pW�fi�#����T��dʣ	@^�p5���,�Ͷ�����h�� ^�ȕ>dy4>��Fc��1CM"G��_LiR�L�p9|`ϰ^�U&F3�5#�Fe��[����ɿ�S����f��)�b���n�c��rȉ�+����� �)�'O(�i�;�a5�2��������X��.�	MW��"�H�.�=���=7PY� )\��dME}�@���e$���f�hQ���u�JTŌ���\GUA����4�z��OKZ���Hm��͡x����ڕ���º�r(4�&M�z��U5����QCZ�]n:)���O\�����
�\eY����x�i U��a�r}?B=�ө�	2B&��,Ԫ��V��6��%
�oe�$4��+��Q�Q����FQݫ;��f�	=�(�;Lǌ��<��iZO(DQA�f���*?��,���'e�Q�c�'w<ӎ��H�w�3�+{�g���Lo2�<�B~���m�]Y�4q6Θۍӈ�aI�l-S��:��#�-�]"ӓ���ǔ�5�u�3��ȕr����p��T=)5��=�d��l�*q��2#d��r+am2ގ�ڇ�(~b`OE\ބ��<x�@�rh����3I��GU&�Y�rPFk0�S4�ęO	��0d��-+�Ƈ�cF#1[D�M�2�lQ�*�N[l��3=�Ci���H�~��d��vW֫0 2&ȶ&f,��rjOa�8��y�|���|o�tcI0��<��2����0XJ(�%͍DN2���z354��,�.�S�@���maf0�n �
P+D6�}�+p����'E�Q����o����k�]�:	l���</�x�x�;T�����x��*�	��f��3R��`[�bLB�A���q�T��_�)�ZSyDy^͉��DC��,�h��Ӯk ��o��g�O<kݮ�yd�$6CΚE�u�M��)���v�%r�0>a�(�t �!�j��{��Ե�8�Q:!aMh:Vh�m�t6)��df�5���6.i^�����_ݾ}{4��c��G� djZE��߸q�?D\O�fy�o����p=�X��(�~�ux���{��z�v�����à�3^o��QѺ��j-%_�Q	��y�*E�BA����0�u�*~��ʗ�$�x����ĄjN�,N�{ｷ|��Ri֑�v�Z �X�������Ԟ��ާ:}��$��*ԁ���z���o���f�کŜ�T�����W��O e�}0�	
�V���@*�f�Q���/��R�[u�Rsh�\��U8c��Sz>��(�����H/,�(3Pqk��E�����*=�w�Ӳ�f� ����J|����^�Cr!Q!����18%X__��t��Y��톢=Ā�����2��"R��zL6eg���͛P�ʞqx�����$��moo߿~qAec��ju�^����
��Tg��7��\�JKGO�\TUB���c����/���<S�x,�3T����wE£ZҸؙH��C�� ?��ܼ{��s4ړ8ym�TuZOA�ur�[�u����TaN��&j�Zf�d��S��)�l�!��Y��Z�o���]����R����k�����}I''�("{��(d�b30N�hi~^ls{����^]Z=q����M�Ǐ�ڤ�.�&Ѡ���ϭ�:@oh�4m#�<v,�U�SVR3� �D\rϩ�Oc�[�fQI��H�%Q��>���"Q�������D����I�N�4 �~{��K1it�Re�� RX��ı�ϟ9sZ�彛��y�f��W^~�ʕ+�πW�E�)�~㦈�h8U���[��B964�4�	�rS��m�\
G�w�^��a��9y��n���Z
�L�E^r�R�0�� �[C+I8C>z�@�j`�@��I���x"2���r�>��Ef�OK�>�E�^��f����JΝ`}�Y'-��I���x����y�>��C��7�H���qN=��0�0�U�a����G�����������O}RT2��i�g�gD����ڬ
R�/!ۻ��x�אS�W�Wr�W����Oˊ�>��˾t��|��pu�{kk���
��56^ZX�|���	�GS219@������U�r�֔5|����=�"B"/�;7��6�g"��t��(T(�����H���1qL̅%sd��0��dI���������O~2��={���Ңz����lB6`}>��e�j%I*g0Sz������D�����������`���9*?b�A6e��S�eTiv��熿���1�q�b�VVV.\�p��G���0���xq�0��t�#O��aʙH�}Ċ�W���$�N���k��������v~��l���ǭ�MLJ.r��-� <���K�mb�tc�E��"�`_�R�r�jqQT"ݒ�v��ߨ�8ԵtPm��`%��k�	���u-�J����\�Ξ[s1�V#�<�"�y@c�7�'������M0�d2��������c�1�P׈�#�BnM|nh1��&+��\��2w�r�LZ�F��*�ί�� ���*�(H���۴���"Am�`_�ᕅE0�$%s:$��J�W�)����#ݬ���g�lD�3�����p���L��4G3a�{�b�d���W���R����L��g��3M<������~��%;��$�����[XX�FC6rل�����6�0�yL6��>�K�P;i�	�%PX��
����t��T�+;���N�����i+&�&�"���5֝����D`�=���E�O��v`���Fʹ�b���
��6gJ3��=lhQ��#��!)g&�%Ħ���g�V1S[�aDI~y����03X]�kwxL�PHR3��1��8�鄒��A�F�@�e_ܟa�#���o�z�PY�������g$��1c0�3n��i��\r������/Q��Y��B�^i�P��W�TZ��]D��F����	�l���
��!���Y �\d��m݇�>hKT]�掋*��]+^� �� ~���0��m�J�z;C2�>��(T�*��xq$�3u�Z�Qd��9bt�'C�����!?�21����i�F��~�����J%F��)Xgl��.A�
�5����e
`=!��M3��ʴ]��k����z����5�R*"[��AH���@Z?ՙ��T$�L�y�I�g#�gԛ6���$abB���"G�>D��`Ji���8xj������1��X}Yc�a��3|	��VӬ�D�T%>7�/ѫ�x� �X��_�Y�%:�X�,��۝�LG�(9f(^;�&A=4�@��eVT�d�!���
k��6��q�>0����,��j�Ӌ����mTA�M�<t%<	��I�(cBJ�#�&�t4�^��t:�s��`p���W�z(g]��٨L���h|x�ך[p�H�	R6>�����w�-&R15LI[D� �.����+�cr���x4����A�?���#Bw�O��NO|�2�\S!�u���<y)7��i���Ey�����&y6ן����/��}�E�zl��E��ވ��Л_Xp\�"�k0V�^@W�߅��LDM��������j�������nUݪ�q/,aC�`8$5���	�&Z�33OR�A!F�C+=�[�hA� !�#�����;>���/��CM".˜:�����~�[{��rK����@ԑ���-9��NS�|�r�fi���䠚s���y�k�S�Ko�jTT.��ו?��
v1��c�aa�T�Y��V�:��Q�����<�t[��������ז�Ή��R�4}֔u���x����4K�(�J@ e���c�2���g��śY>�����Ņ��]��f�+�V�ĝ(�EߋD�;Y�XCQղ2�� '��E�<�|�rB����HYV��ь#O����\�h<:>:ln=h���_zʡ�	������7�������b����+~C�q�2��]�,��x���ݝ��������{������6V����pt(�h\[��$GaV�N���{n�d(�M�/2���i;a��=���k�@����J2Y�@Ձy;�t�?�s�fᤛ����qX�xx���&F��T���5�8YF��G �괺��'�]J�t���;7�#T�K4k��7�����;���L�%9���]F���ǁ޹�v��Z׌|�"AlP��JӘ��h,KK���j�Y]���� �^��l�O<yY�������^{��v�ь-�o�(�I�β#�%`Ǉ y<�ە�_��|���=��t�������I<ˀ�^?{y{�!�lA�EN3+�J6H"O�7
��Ѣ4�w����D��]i��R���a�_:kF�������K�Yr�����^suo��|�?�������^���⢣�z1/_�g�<�����s"?7o�tK���[7�v��Y~�������0�lll�Oܿ�䵍�).Ĭ̧S���d���.�/������sc�:E���ɜO؈�V�%7|��&vE�|�ʂW�X��d��x�_]],�平�����?�!���m��N'GVi8쓮b�l|��D��cN���K�Y_[��������S��I��믷⑈G$�1���V�XN6߉5�g���Y��W�A�� Y�����-��q�>~�|�d�3W�_������b��,�� N��,B���9b���w2ף�xI��q�|���.l�=�,jƆp��<�+�m/���E>��LZW���"�[kd��y��,�"=�y����UY6$S34�}��[{{��0���
H�X ]B�d��W���~&w�&�7�x��n���K�P�?��?���BH�J;',}qZt64~��s�����Mȓ���_v¸��_����'��H�8冲��tb�n�0��ol�_�rIDGu����H鮴'=������E �m�]���(U�f���3�5�	R�Z�H� :�4帤��ZQlfs��l7�˺Ğ2�J'#j���G?�q���*X����uS��k��I�)ނ��.\�,ݼs[n��O����������ﯜYs�x�ۧ^J�!BlU��x�J�Iva�q��019�<��G�N���Q�t&6DĪ�hvZ�;�]��o����������O>Do��EMS���<�yN<��I_���M�!�/~�O�SKK+��r~vm�#��P&��\f�̙�����'��p<F6��ڃ"�$-t���Ϝ9ã$_.!�k��h�Q�G6������C�s��HP�I�����{��URάФ��4�-Sp��(M��W�f��R��:A&$�c�����ZTŢ�]7A[Oa���yg-A7JI�t6���<M�L���ɺ��\U�	����`���_"�Wi2�H�f�k���8 W�}]�ҷ��z��,ea�2|y�X'n6[J�*���P*�0uZf�vH����*�
����"uZ��ۜeI��䈐�%F���è#N���$�ƃ���Ud5ӽ�vƹj64_���?����0�e�P�i�栝�!���jo���1����D�MRQ��i���_�Ġ6���b#\��S��D�,ͩ��)P�6F�'@�XcI���L��ɶ,����r��G:�[\��P��Q�Fb�U��a�W�`nZt3]�ɬP���� pb�U�����ͯa����@����F�4Q�9H[톪�R<��tdK�Jχ����P��9��h<H�Y�8^l�G<~�E�&�t{ߩ{�8A��r�	�-�3=���EV�qX �:�
lN��͍ڣ "����2�"T�G�W�N������9vN���[������qŉH ĤLeRex|Te3�sP9�qY)~3��v�S(��wڷ5�
��3�U�}��'W��j�\��#��d�v�qb0K{�๚���fB4�_���6���lӉU(��=�Y^n�S*e�lr��
(ub����^��>(�>���̼]�G�3L�wJb��ul��c�S|��Q�ah3w�J雖O�@@3]N�`FWF��gˬ���S�2���J�	�6[��[X��k���Ю��ؾ��ז���PL�_��=C��G���nu:3��6��l�:�kU�U��D���x�{|�SSg�͠��`x���v�609��4�����`n��7�<9J�j7�n�u�3��&'ҙ�r,��@�27D��u]��ފ��v �"[�:�u�*Eܰ�o�yCc�Hβ�ċ�wCd�k��071�����յ5R7f�ʗ����Vw�k���j<9��,)���c���������

h~U޺uK>so{�V��Z
lUR�
C�XU��u�ЌO�	ϗ~<c����������h
�E���r1j�����=W�\��O\?��C�D\O�5�ȷ�%q��q�!#�ڊ�z��M��Z���e��@D�d]�T�u���s�E�U��`�(�Y���J��i�s^f���I�9n�=ܹs{�3�v�0&YYYy�p��ޛ�\�V�^"�N;�S"D$v��pq��E�..����n���~��rX���YY��T�H�!w ���u(�8��2=�U�\o^҃Gѩ�<��Ğt�G�B��=�'Tn�^��o>x�w.l�oll,-�#Z[^Q�xL6HO��+���$3���-ڔ\h��[Jc�ח<8J���0�~�T�Y��n��fz'�Xjq�x����#+2v����_��c�sm��M<8�FK�!qS�F՝*���L�@J����G8��]�i���\n-R���u�Z'�f���-+�v7�3�9�Re��UN��zђ�)E���
���HWŐ���˗%&L�T���ZK�ˎ&��
��������F�9t(O���F�t���8�4'3����s�=��Q�JF6FK��{�4O��Q�F���J�A�q�^2��M�9B'�~����/K�C����! �/��;�����F�-JӑȰ�V�8E..���_�EA��%n�*�L4�ֽ���\K�!���D~r��U׋�
j���(5�Y��M��4�W��ȘqXe#�4��@S������y��(j������<��O?���Q�[]��7��$�~���g)��]�rY��~�3Lo޼9D?P��h�IΝ;'{q����F,�����Q[qp�N�l1�.���^!�H�5������4���6bؑ�²��������QL�\�{��֘�*�]6G�ϳL~�uC}3E�)6�;冲ǎ�!P5���^�EI0O�6a�4�Z�h��*��� �չ���~j��)����|��<����E�t�0�-�2�_�\"zh8�e��gdW�Et,-��~�W�W�/���j�����~�[���O�HQt�-U�G���E	�YY��������/7{�-���ٳgE؞y�_��W���l�g��!�K���n��a�m��l��<GC���L��ض����U�Z��:+g�Uf��o�좶�o)jV�z����BKG����uΉ�ʲڲ��{���Y���C�V6��Y��A�㉁�Y�7��%i"��ل��tp��r��R�iZ��&��S2
'o��C�A�>Mh����CF5��7ƾ�U��g����f�t�r
~�q�%�WwH�Rag[�����6�d ����p�a�uW[|bl�Dl=z�)?7Sۍ�jN;���h�WWW�k&��&�((�[��:5����i�j{�
�Ѡ����a�e�1t6�>3��<3s�#a\�)KGX=%�w"G9ᩔ���Y37�CgF�T�:�ѰyE�Ga�� �D�t��7�,]�:O��#M95�as�L�k�?j�/u�J�Ҷu�*:W�!���07��E=l��H�15�F�(Q�8-��.����˩2��*U~��{��Z�ʮ���I��\����=1�z/�U���*Lh��Y�J�&�Z����`�%Own�1��fW���s�fZB`ZG�|V�XZ�����	!�#"���^��NW�Jgn�߰���'I��,���G���g9yBe���x�p��ݻt��f8:e(�$����f<vsM˦ *�"'7f���)���)���|_i6C�Y����k6�YW�� �f�E�+=�$ %Etf�
����߀CC�g-,7��hn(�S�z^��5q�2�t���k�?�̴�]�G�I5�`(����J���a4�'`�PSJ���x�	�@4:��5lN�Wzץ��&_����s2�*[]h��+N֡��qaO�1���[���}��2�'!�|����a���M} ��0A� ��u!���k  ��IDAT�B�mN�$�u��t\�U���7�����t</����PbD�6L��3��;�O��r�n�h�~Q�Ge,�7 H�s�2�\�S)D<��h�A�Ftz� I)��
=ֈf
�?���Ņ3��C�C�隸:�R���-*�&���Q%��w�:��4g���/��X�K��(�@�XiP4��@~�(����>k{�VI:�u�S�+m��B�����U�C�4�(l��YR/�S�����_q�U*K?-n(�	�x������L�V�2q�q���tc	���G�j���a��L�|�ᩦ��,�c5�j4��!��e�#N
	Ϙ� |d�b� �h�8�������pqj4v��tiOc!k���@rfE�3u��ܕ$U6=��T!*��@�#K�N�&I����x�^\pPN	e�"7���d{�����'�ȗa���6�(�x�2�d�-�@�vHf�)�P�=8�#���,�@R�rHEɈ��,*���+.��`� ��{
��t�zi�"e����p�T5�f��<�s�fB�i��������4qd/b�uE�[��mn<z�5�d�?����PU0�4k������ ;��۷=�'>���	K4�y��*��"Zn����d��lI��D,���H+.]��$���F-5ZU:������k+�;��g�!¼skyyY�j��G���͍+�`�[����W>��$M��bci�x�>�d:�*�ݨ1Q\7��*�"pI�d�������,�;�N'��w�%���Wy8��p�:��bX��(t�Y:U��=\�I����켲k򌲰Y6T��f��Y6��i��դN�'�?�77ϊ��k������[�?���xr��s��q���ȟU�,.���K=P,{E��l:N�Q�H'�l�%�Y�\@�mO��
�Y�۾�ˤPn�XY����A;�f@��Ή���O�&��+mDYʬ��ǀ<�tw�`�N�[7x1����|K+�d�E�v�GG'+++ˋK��"]�����$<>8�{�1v�An�#m�It��l8�+͓q���4��d���nO����ٌ�p�� ���揧
���u�Y�ސGCѳ�=c�y]p��Ǉ�b�d��o��k���rm}��{����㏮]����"6U�:��s���!���zr9^ �B�����_LF8�������-/@�T#n�!x�E�w�@��[�?�,��!mQ�`x��v�GW��ɰ�<����� ���[�0��'���H>Y<�I�����V�׮��}�J^|��ǇG�+W��{Kb9�Ay��Y����F�����n?�!�)���ŵ��huu����&��[����'GC�$������A�o����3g��A��޹r5�X�]��8���9&X�4J����pum�捏�y�Eg|�����ytg���F(m��g�m5�0fa��g��:���8p<@*�,���������$�{�o�	b��t_�(����L��{�qpTn=���˯�eTg-�U��k6�W#�v�E�m�Tg�辺�$M�Y"O7�3����ʖ�=�����QN��a�I���(�h�¦����fr+#�C�e�@9<3�@b� ��|�c�6�y@[���k�x��p\��gtL#���B�?;#��k)��Y���&�{4��P�kBo3�����i�C��.�]���#O�P���●?����_n6������$͚��[o�����:���+7l��@���Ã���O>��eD�g����8E�t�-񋎏Q�9:�VVVs��d[��ۣ�w�!���8�#����ž'�6P��&8��	A�ul ����}g���$��F��@U�`J���o�Gɝ�g��^�^�>j�����U�i� ���� Znaa	������DB��f<��y��W�p��q�@�1�S	��qL����d2�iտa]\�����N���Ώ>��҅Kd�~��k����'�ZQvz���{?�����ob�PN����:��@�YNЂ�ڟWT���m$[�P�i��p�H�;��g��x��v��v�aU`�����|��3Wg�1�"����o%��?@G�,�X���D�ȿ�J]�tI��|�H
;J8�m.����@��N���[Oe�=�uw!�{h.ݹ3��S>�� 2I�'}�79_�����oo�P��[��:�2�JE����uS s�Cҫ� �,D� 9ۏĤ��=�M	�]C,W���p�5�`��7=������:�c����\ג>s��ui:�Zy�D��n�j��������ѣ����,��J	�<`:F.�/t\���+��F�d)����:'��ϗ�VdC��}�؂z��c��s���s����ΰ�ք%����|p�(����*<;6���Z]@?@��Y+4
|'z��,��h���T$ym��ά,*V�/�++pu����`a��6�ѐ�e%�}N&�J���F�7e[��(���9"I���Di1�y+j3X*~Ţ�歡;�0k�\E��d�ͪJ�;��im�#�taZ�<S`�#��j̤�`���"2��s�J���d"W�e��xf�^i�����b�2��W��DUV���D6
��H���L�=�V�S�W�S���;.��j�0I�D��t�0J��>Y"C�k5 ?G߃��N͕�3]�ϪY��%0lC�h�&�qU#�P��Qt)#�/A�s���yճ^Jfx��RS~j�w>8�+A葎I���^Q�!��X_4X�{�DY�E�c3�u�4����u1�Y�Xc�9[u浪����� ��ñ[��hy[L�R@�6����6+Db��+�0O'՝+��͹R��;��+�t�i*)M�3�b�u�o�'6��6�Ќx�a�F�?6�h��Vv{]���ƒC��m>�<h�ޒ�f��<���1�l�D�aapL��&��i�a�ab+0S�,8������V��*�b�M��s-6s��Q����F��$���+O� ��k����ǵ��t2�u��+K�@���*jl�CBS�D��`� 3yϼ�-SP>��y�U�"23+�i�`n�Q�c�'��N!�O�T�,'�ZXX�.B��_�x�s�bBzK�?���'�X\^�� ��}�*%ra'�3�竽u��X#�j
�|�����ݝmԸ|�aN�q�a z�vg��,��I��s�Z[��o�I�W}�*�����Pִ��!HJ>|�~��xZ��%�b��U�!����-@�Xbx�vyR��!ߞ����-��ۏ�'E�Q�\nL��\n�B����B�1zyD��?�ȶ U�A4گ�Lw|�!Tá�|��Se\���B�'YOy�k�F�jˡ�"Sā�t�<�q����x�=0�Ofy��yc��4Edr�����{�(ў������D����.\X[{���˯�'���l����D7�-Emgԥ�Pc�P;� �ZǱ�J�>[�<�fܖ��p��q�1�?��U�eY:F���V���O��[T��ݻw�=�{���C1�����lչxY�f�m4N�.�ݶ�qLa���	�����dw�h
�������}7aM�C����{Tn�Z�޵v[,H�F�<��hU�2�w�ݒ�U�����.T`^J8��2�ű�2�\M�^����Z��ߟ��&��B��$�k>�Mn��P�)�m��A�8z ��hz�Qg�Ȋ�=|�&~�ﯯ�߼uK�h���s��%9��t��(�������,��˞x����A�rVЇ�K��p�5yhi(AqG�5f0Im�]{mm���gd�g�nJq�����Q`h2��B��rjvwϬ�uz��W�r���ŋ"�{ǃ_�򗗯>!�x��HI�A�.�&Q3�y���.�݈��Jt�?^�J�ݖ =�-���2��7�A0����iI*�����i�ԥ�(P>ɜE�7�
'�~C�.�S\�����t�c����e�	c��T�Pݿ_V�`��������i� �d@�/_V�#m���)�)�mooϩ�6F�4������]�����d����4{یCZF-�8h۬�ln���~Nm,??�m{��4��CQ�gϞ%�L�Fe�h���f�$��4�َfi%����ڟ#ު걧5@�&C<T�a �~l���:`c)��[��1]&��k0��S0���~��4g�����o�36��m�3�B��s4V�� �������ś���w�����,/��������6���-�Z�;;ʓP���O(-���/��t���D�xϲ����:K*w�<�4LN����l)zԭ�<���ۤ5E�H��ڵ�i��8ʐ��l�g�J-�i�יA�k����[��A �Hy]��>��w��o��l�8K�FK;��ؤ�E��T��zH�8zLݝ����H�k� ��U�O�=I�Q�l6�����9d��v��S)*��?���tf��vW�1 ��T�\im�޹ݖ]�u��>K2�N�,�ߥc�R��r&�G����և�G? Z��nE�<�����eEw�F3��WV�н28ּ,���;i�!͔JߞM:iW������#���@_�r�����4�4M���]�켍��^��e$F���m�('�-g�� ��)V�P\u�O�Xi�<�e�	�ȥ��T�B�1�
�(5�����dE�`44o��N �F�� �����u���
- /��7 ��`�=��9uM��=t�fYJQ�n�ܔ:�8M��JFH^�Y�j:x��t�c�f/��[9�-.�(�� ����C���X�d�t��S�K����&�J3K��?կ�:��Df=F����s���������4�`�K�rw�r����p
O�5r����v+V�,]������5o��b;0�K�����w�}W%��bW_5v��la(�\C:13���hѯxF�i�ɄQ���]j�����ތ�����XH�gz�mD�.�tC濋ǬL�ۚikR��VZcZ>D������rl>A��ʄ���UhZH'���5�
;#k
6/s:B�����jk�	���1�Hg�ī�#XY�pM��=��<�WuL�|���:�#�6Ы��\r*yf�F�W� �?��A�a��=�'4-��WQc-��(T� �T���-+ fQI��� �0����A��SOO���r�ഁa:�(��sj�e�s(IT� �QH��(v��t6��B|%�#��xV�P���<q�z �JW��B��������]��e�[Ҧ�ʹ�����15j�R���g��:��馴�o��3El+R�\�u�*�I��X�|���7c(�.m�kfY��Zg40$3�wf+��x"m*��m��i4]��<E��r�8ܢ�����W��rO�۔����wdz��?�LFLy�+�-�Bo����=o�\y��Q�� ��|��Z���/I;	�g�4��߲:�4�%'*�7�m��rre�eõ�۹\�T�I蔰fZ-�Z?��TG>�tU�#;�̈����H�����ƭ��_���݊kx����z��-!�BC��1������c����G�}-;`����B�^���~���(���#`����*?��D���d�Nő��T������e��b/����UW<�&��r��������x8�e}ƋZ��#�$�ө���kk�>�wxr$޳<f��L@-e�A��h����{�7�i"���Y��N�)�6�z7X�ՃQ��q����F=?�iAz��3@4��>���l�?4�tB����16��,v;���չ;KKr��'�g{���$�r��G�te%lb_�앳H"��ɱ�(�	��r���>�OG1�=z���i��O����Z��8ʳD/�� �'��F��|��@-�#>]2��M��J�[]%׫B7.�j0�z�Q�[�,�ݿ{oia���,�%�rw�[��������v7�D�p��� �˓�y'�'��q����S���i��RTi;[��k�K���Ң�ma]�Wy<���x���7��z���b��jS��=0�}6�p�Bߨ��:��)5�I���F�ݘL�daBk+��iFX ��\6�E2��ŧp���BWΣ,�ח�9<���bq����;<9%+����9����ܐ��r��p�CWLF��%i/��(�w�,i�T	��0uo�ɝ�����(��0�e��ݻ-:a�у��E?��^�s�ƍ;��}���H���c��)������Ç"_h�B	)FJ/��8�fs�L*�͓�� ,� �i4<��&q�(%ٗ�>:U'�t:=�5�n���Y��� v�X��t��+�	�4��KП��M�dኈh�ώ��ܽ�n��V�⹳�>�ĝ;w��d���������O?mnv:=���G�d�S�~�s$O$�O��v7��q����z�����.�n��	'�&�D�x0��:t�\ѧz���3�!n	�4C� �NXߑ��-�vڭ��2��'ͳn�)j5����f�����=���j}�/W%PrǇ۞3��c95QwE]�J����ʢˣ<z�-
\Dt08�w�f�$��#����s�k=���׳���H������ѥ�+r�FcŹ�:�é��H�{�?!���5A�	�U(���XpG�������[�<�$ʆ��:�A�B�E[縚K��O� ;�UL��H��`��+�oڑ���V�`����fk�6��w^L��O�;Ǘ�J����5� ef���S4]��3�ה��5�?�~���4_i8��n/�;�D���}�{������|���敫�}��'y	�{�Ֆuπ�Dշ���Lq�67.����oݺ-;��/=��E�Ϟ}�&��������]$�~�"�6cs}�6p͏�t2��|iyuu5K���=����y�@�2XUs��a��熟�+�≽��}*�b�L���S�I���7�̏����f�*�v-Ph��:�Q��B�*�A��uS刊'#� nC]����3q��
��f��4���ź�����"=�V~8f:����~�'ov[]� +o���P~�l`QV�i"�--�FP�(�(���S)r'��e�d��މ֑�:��(�b|rr��Gt:�W^y�翴�~���"r�z���0�Ӹ������Vy.�1�rt�+_�_ �S�V}̿��M'�5+4���*��Z�73�r8�^�V0f��73�XX���&>���eB��ɰ��Q�x����t��=Y@�;�W�[�#�7�F%�(eG��y���~�g_>l�U�1��S���{��cW���O��a�aA��z��;����UMQ�+-����^�!L�jܜ�㐞��c�}���<,j &�ȭ�Ծ��`4��_�+��h4�q_:	���嵫��?^P,��0�ܩG!S�W3���F�A�&�����
���Wh� l�]��Xn�P3o$�c[M���D�Vh��ɏAt��q+���h�D>��{�v� }��ߗy��g!-���S�L��x�(lw���1����d��{�|rn[�� ޞ�������4�f�¤�h���/��$<L���̧�a��iR~!�ۊ��	2Y؊���L�9%��]:s�5�2���3mF���JP�ؙ���V�A�a�uw���0T�IE"qA�[ʣNĶh�G�buy�����cQ�鎆#u�1������:E(^��гV�gim��!�ĥ��J�d��,�l:�N��  藽���E��k��B���4��\�	��geQ8��K�-q��k�#�'�f@D�X��@�%��!i2E4a1���V&�<#6E��%�7��
l�����	̶�嶟Y�H�L������R
]�:w�����aц��umX׊�J�G�Xo��$�0����@d����g� \S���V�͌�܌*��|M�f��U��&֙���5gǴ�[w����4�[��f�m��1� �y�|z0�a����� i����	C�@�8�j�,+M�۪oI=����`0��?��|�;�]��/�?�������;���q�9��Rz�$V�� E�����_��7���L-G��@��Q���`q�Óȓ���O���Tdrq�ӂ�E"X	���)	�D�K�J
�H��\�*���h!W ��y��β\��/��5
B�Ԏ"��Kloo�m�ma�
xyD�����1������ݻw�_�pJ���{�9_$w���F7��#�5Ia԰n1̶z�dMff�0S2Ř����T��H�F�-��JӣZ�#|5�+��`M����{�4w�x�յuG��C�E��O��m�X�H�moi�ds��dLu����i"��(٣G�-�խ���L����c�	�"f8��<eh+}��y�ȃ������1��-�h��Z�X*1��F:����[ F�T����EKѽG�8�%0��c��nC��Q"��P�� �?�1�)�D���g̜:s�`ejz��W�Sԍr��=�l�bl�!��Q��!"u+˘� �d�M��-���;;;�8޸qC�^[[[��0����;�=Z�9!����β��@���E<���=�#�"$��� /Gg︕򈥉�BΨ�`�K~�&��� ��\��h&e����w��x㍋�]�&0��^�Le6�$���t1a��dHU 2s���Q@����v�J^k��\��.�cNk R$�g��$o�:�*-A���7�_�ϞM5�A#U�t����{S�J�'Kw���K�.-m��'���)�w��ʋFG4ш��Yأ$�O+��F�WΈܼ|1Q��B��U�1 [�bT� [#?�� _�$%X��5<f��nkԃ5�IQo۩��`\i#4_T�Tघ��݅�8^{�5�n��O?��������o��v�q6�$�D�r|�|�����է�~:k��Sф����V��I�}�	,8�=Y�}���"U��
E0�b����D%�?MSR�9sF6E'��܉�����fD]�GG@]5|9&a��<�.PE���ï �*��4�����<q���lN�My
$u:���!x�>-�f����jm%��XC�rR8��.,��H�$Y���m9�ZdB���o�^܄��(�c��*��Çr�)<,�Hf�x�����0���(�����.��i��1$���t�-HkKM���Z��1��4v��"�J63t�|���,V���EO��nd}���~z>��Χ���JtT`^�9I�_Ս t�<�������'���o~sA��_��W~���M����dv��������W�7?��G���Ϳ�7����\�����o�+Ǒ���o�}�n�p^��Ű�'�����!������Vf���Ye�ԁ�F�C���l��^�y�u���g�Уӥ�єV����]��W�d�y��a���_v�����J��+<89L�H���(F�I_�f�����m����"�E�5�G���ĬV,�$S\C�q�dR����9����߇/w����I�u�����?�������]݀��,�]f�V�P�Q�j���{�A�e�9�X�v��M����f�Pco�����W_~��g�]���=-��O����,^%���/"	俖�YYY��<+��>W�p�~��˶bI��e�v�u��+�J,��g���DV6��Gu�@SejJ}�M�J����M��џ�韾��o���ܧ�[qf<4 ��e�9���ş��
Jp��&fi�FQ�;�\����xw��?C	�!�{��/�%KqU���J��OO�yf*S��Wq�A��	�Ր�u���l�|�w}6"�ҫO-`�K�8)��Rd5�IC	tJ��>9��R�;��\�t��*��q2��~�`�p���3��k���E�-0h8�0����%���T}emc\��C=��ԂlL	�D�'�_}C�M�!��ń��Ӣ���Q>
�FmJx��L��b�(>��۷�g��G�nw�{(�@Ĭ�ZQ�s8n>���6mDi�b���R��ϗ�(]'�ca�|ݥ��Ҹ�dߦV�����fQ3bئ/i\<��o�g�K��6�b�m�&����ϱUI0�1��e�����[�$��F�
k��N��YJ��ȱ2�fej�M�8�\���Cqe��I���4�2l��m`���>���q�lj�\�T���:����uV�����T�(o�{h�ZT� MIل�(�8R�lV�9²̘&v���UVK����#���?q*J�����˼ԙ1��ShI��N����_���>��Pt�$���Fl4��F<*����n?�+�N>-9Zq�h(��銧ʨ�ի$��|Ǐ��1x�F�h�������*C�S42� s��G�s��
m���e6�괲�-st�5"WV0�N(pq�G��T:q�G���4���$H(�<C��ļ��c_��� -��|6k��FY��t��\(JHr�s��?*v���7�!s
'(댤x�x���#�
��[���TpX%Ov��i��8;���t6n��i �v���l�D�j�@�8��u X�3�N,��Vސ#��>#bd��:W��T���6i����e��/#dK U���h�X.xꩧ�������HJL���d��M�u�c�u��0����v,�W�|O��ĪV����l7���񶆖]���u��pb�}y�a%\�t����RKq��)JJ2�]Ps�7��\]��M$GĦ�Z��c��4��ڱҏ-���b/?3�e�7���w�V���d=OƓ*�:M?�� ���G��^U�N��F��i�:�r��T���v��j8Z��v;v�����1�dg�v��$���W"���#��5�~�'��Ř�V鴻kj��|r����g����K/���^�z���p �ð��xPep�J��^^���jZ�ߝ%�4qә�����2��
�
c����h�N	?o����(�8����^�j�����S�aC;2:�VwaQ�}��jN�j���~�]�~􀨈Qy���zq!:lV�p�����3�o��F�Υ+�O���F�uk����>h�A1�S_� K�����pW�Z���pђ|�Y�5}���L&r�bٝ�3K����Rs��m�+��jVQ�m% ɘq�B�N�}4�9�����?���u�T�l7ě.�8XZT>o����]�~�/���K_}9�:�ά���˯�?:��X�[|�0*;8-t���,ȑ�D'�,�Gi�V<_ihX���N�˫gN���^�ŕV�&8��R�`^(�����j5����Aϯ?���S�4D��dr��n�	��#	��RV`��WW��VS#��<��?��ߘ�n���3W/I�(����� ��������s�΍4eViNw�,�Lh���{�F��� -�CѬY�\҉��g7ּ*��2K2uvSD�;��^�{��[��%�
��$�Ts����������q�~����h�,.6��=8:<�~��70G8jo�����O~�d�'rV�%��}��i
r�Q X���	��\C��jm��
�;ͶB'4;�`��x�?9�+��%��+�	6�"K�1:���x>�g��� �Lˇ'��f�؇a2@�V�%���Y���;�,v���+�y�]���R���0������ߺ���_��j�ם$�o$�K��V�����n
*̪�;u�܆�$���';����=�䋽N��ǝ�=��$����p'���2eZ�� :^�����1Y��O@By��KXųQ:�[�5Q(��4�l6�~�~�;��x�g�tu�ჅNcg� �c̽���B�x:	N�	G���ѣ��}p5�>F�g��ˋ�]�����DN9+Rq��,v;=��vv���CoVL��V�}�p�	�+VcȭH������l=�l9�BM���1d)�u�[��S#���Zh�Z.�������Z��*��W�F=' Ҵ��f0�z{"U�ƥ��t��n	�Lߐ:9���l1�1�}��Z�PH2˂�|!�Β͞�`"�1���P�%�x3�\o7�#I'<��JLq��!��g� �VK_�Tc3Č���������<��U�rי�H���e�N�*���b�WE6G�r������������ǮM�l{����IŅUq��,l�G�$��J���3�Dʏ�pk{i�̷~��G�>�i�������͕�e��Y� ��(�^���w��i7��ݝB�?��:ԎH�3/�zAࢊ�s�B"�T�a�ČȺ���1�)J��96ȯt���jҥ�W��r��ʡ�Y�W:l	D��鈎��@������`{�F���8)�_���㛮Gb����8pYa�
���]V�^I�%�(�J�A�'�I��Q�A��1%�a�\ʓ:?�4CO��w~�����w����O����:&_]z�JwqA��T��1����ç_x^�BΩ����RQ�l���"SS[����8
PQ�M������zj��W.���sŗ�}�V���4��0f��&�w��l��V��k�����#8��nߕ������߹�q�����b�5�Z�5�+���̶D�~�J���f�[���9Y�'�x�����׾���ʿ?�6.�����{�۷o��)�[rC���l�=�U�w��4�F�ee���(��g�1Lqt�(��D��P�
Y�N�+++beahKm���]�?%}��������X�TL��A���a!�=	i�V�Т�D}�FSg� ��=ͦ���R��6EQ3��Eyg�f�k8��"�� a�Sܿ����	��UA�l�YV	k�8�CQ�2��b�o[��ۘ���13!�5�j�����a��iS��9�pʜP#�D+.�)�����*	��j�0t�t<7����>^\Y|��'Z�W���7��~V��ä�I��i����� ���(LFME|X̜�7�Q�nYă����n�S���X�&���e� ��vdsp�A����J�V��b��|3�YcY�t��sR1ٝ���c)ȬdA �� �-�������w%�AFF�����t� });.��X{�}7��t^��Q�!
�,��ݗ$ �I2̏+C&� k*��*�ԃ�w�契8hS��F�9͇�+K=�������:Q�8G.\X]]�{��rjZ�>�i�E4�`����[���Y�K���%^�J��ba<��&��>=���y��t�iJN�,��fpا������=�rz�v܌U*JJ��pΝ]_���C��D�`0�t�q�Z3��R����Sʊd�)|�Wwih[�R������;^iz�N�r0\,-��%t���ԩw����z��]1r*��ͧu4��>�:���Z]�%��f�=$sަ����8���9�� �60�iE[�!�����i�IU�9B?V䷺:r!v}��"퉮������F��O@b���0� �18OM!n=�CV�Mdb�܅���k%撺�K��cL <��jҊL&�)��k~1Ӫ��a��~sa@�����0��3�#���"0�˻��0_����a_�E~�#�n1�J��S���s�='�V�%�RZ$�b���Y��2Ϭ��<ۗ��6A��G}q��������XSd��%q����^���o����?m)۔h"� E+i��C���~�&��L��bv�UX�h|"���*~��������5̝�<�t���#=�P$�[��C��1��Md�"�e�V�ߜ�u���v�8���/�!��Xv�0W�!\��ԩ��
��R�`š�b`�t�Q���ׯ˧}��_�u���?>�V����V���,��/7��D\l��c
�+\1��=:Ӎ�JM�@l�d̈��)���Hmk]Ÿ��J���yhEY�͊B�L��y��.����O^|�UY֧�{��훿��o�t{�������3P����v�j)g�(	���f�{�m�5��V(��*���$�T�	�z���Cߑ�~y�����<��bC��`�^�~+��E��؟������[��V�h�;��K/mnn���M����#[�ְ��c:N�4_XXX]]���Xu/]��.,1��WuH�]'0��B~���!���9��&�"l�h8!�J&���H�AU�tx�nz���ÿ����׾������Rݽ{WG��[[[�W'��������Eo>����YqE-v���j(��L��H��U�h�k=3*A�H�g�p��J,u�yW��;3l�t��b }�S��s�]��ln��s�4ee/]���k�]�qG�9V���Bgy!=����̬��l�)���1��D�����M4�uI��%E��ia��1� Q�����tC��1Q��
r�Q݄�9�^���VD(_ZX9s���}����k��<>ځ2W��Ё������k�K��f�ҭ�˫j�N�\!괨�X����V�z�"�anb�[���+%�סBQHU1Xm�j�@����?�s��u7/_�>��c��\����N��'b�]����9Q�r��gϊ�9H�
�<��Vń(}�����3z��S(L�u�EJ3�j�����D\4E��j®��S~Me+۴7լC��v|��_����w�3rc9
�<�K�/�����,N��tR���ѷ]&L� 1b����T�������~��gH�r3V�F�:�p�V��|3N���"n��b&*�Ec蘬��:C���1����@-z@d T��J1H��,L7	a�n�7m:�KԖ��o�V����>��c���7�}���A�$P���;��xA���e7_|�EY�����Z�f�}�PO\�)��E˥1�6Mc��\?�*����w1����<�[��FA1�\���t	���BRr�h����O�_��Z��!��N0&�L�s�E��M� 8"j�9�s����r��k�ةjfѯ��fX虹ϔ:�]��g)����2���F�M�N�9��2�1���EL����p���ۡ#K-f�w�QY-�]��nBT:!l�2�=�7 ����?�v�q��"?r�yu��"륇qݚ�Nh`�r=q�hoG!�"�O<����s4�L�S#l}3Ǡ}��yg�Mp�8��i0)��fb����oܸ!_cL���-_�c��<,�*w���P�]��*�C��5&��񫏉`{q�ʫ�b�X�'k+�e{�S����P�4��zu�QĤ�#�"�933A�^���#�8u�UG"0��y�lq	g_Bzŉ�W'��5�@��Ԍ���s��f�Z�J��������'/��J�	4๑||��!^�SY��e�-a"���*�Ir��ͻ�F�a�YY&V�JO�� ��E��Z��o����L���̤���Q��䮙�嘮d��1Bi�,�i�*գ�N)eH8ծL'�i&v�����<���ō�]߀���l�8�<�2�Yݹ��Q2Á��-�^���т�)���Π��ֈ��V���%+�`�W����\�t7��H�ۃL񐳩Q>�;��޻��L�R����H��)�֖}�<Dc�)1�Xj���f�1�w�6WE=*�[�sO�����p��u�i��#�<�m:�����B1���j��&m�g�/){V��_�jA�v������傧��y^u5��q�(�9��u�۶m���af��qt��4a��H���p�B��m
�N¬��|��-%��9�� ����ҥK�}�D�R�����Z�h�6�$
�؋�
*3����z��J����oz����DQ;0�Y=c.e��&��$⫑̕�Z���u�[ӥ3����$�z�z�+xTA��K{�n^��q*��8l��G�W�/�_�~��� s7Eh0S������To
f�O�>c�٩S`�ΫB>CX܊��˯��N��R1�y]���[��˞���d!��<�7)
b�,��xa�.�����;�V���<W>Ӎ�$�q7j7��h�
�w��x�T�W:M�S�K�lΐ- �kP�j�,��]̴� ���$V	+���rú�u����N5�(Rg9:!����KR�Z�VϮ.�,�ٖH|�$y�.�ﳔ\N�������O-�<�B9ۄ%<�=���.`��-�Bm����i.�KW�]��\�:I��z�m٩^=ԍv�a:�jr�B""��݁�1��RW٤4�؎�KY�_,����d�'E�ۙu����P�b=֮3����D�n�����SLA�`i=w�)-ڴ�X89n��Ӯ�::����ĕ��}�δ�:
�����a6+#f����)"$k��ޑ���ޖ���V��Sy4��|
��j_*^��J^Qb
�b�L���>�<(�	7�^�A���I݂��D�r�ŵ�K3e�rH��z�l�:���q�p��H����q����i����ۘp��,�؆+W���%���:b{��`�	y�1�4�B�0�i_��V'�y��p'�~e 3%�+��$��y:�]�>��.Q�Y��g4�[��"K�������׊� /MR*��A�`gg��g��g���K�d�nmi@9�T�JT��<Ӏ�*_�䑫n-`A���ɍ���	�8���ΐ�*�HNJ@(+�ֱ/H�Ô43�S��Z��*j�
�Q,mU���^��?�K2I�׮]�r����3K�]9��/�W'�"�tE	n���Oj����+��R@�#r�A�b�+��t,����&9�2�Zq�j�I� �0-��䈀Eo�m�F��=m,Ĳ����*���ǣcLr��O~"�p���N?�����Y=����U�]{�)q�'��"O1P:�Y�vfqm}9n@���Յ�ь�|'#��k�W��3�Y���L?2P��� Ǩ��W:+��4�r���'h�lJT�&֧�'�H���o�~K�1n_|���O��?���x��^��s�J�F�]���i)�r#^\Qz�(����5���VWB � 5Ӿ>����ʏ���&��k@[3��M\$����xu���V�,�?A�Y��ST��p8N���}�?���~�W^� ���>�~��d<���T����8��S)��d�ޞ��6�\������3 5ch�&�WK"�0�E��u�h��Z1��Q>�&�:���h�J=�j�u#�����9�[m	�B/���y���t6�8�&�Ο�w����M����z��Yn��L`��yU�;����L���WQ�	L�'ssT�6�Aǰ/y�˜h/�0R�;�����T�L���8�|Zy��&���A��r���9���8f�7s���@��'�%f.,�Ǆ��Pw�DL��6�����?��?��?�����/��3�n�B놎
U���V� �+r�y���?|���E���7�p�}	&���ɷ~��g���d(:��˕Q\>����ѻ�{��tɕu�U���j�&qsJ+i3b�}��@�F��,D1��l$l�Ųh䃫o�?�l��eZp��[dSY__��N�u���JЦpp�:MR��i� X�E"�9JH9)��k2�,
�`���-KC%��a]��g��x+���kL2�S>�ť3D�(@�N�:H�2��9���+�1WjU�����
��DL$vE6�(	��E���٣�����f4Blǿ*��l���҅�{����T�����J���	�V͚�6vE�⣖M�rUǺ�� 5u�q#��?��[o����?�|��ߖwn�oVyurt<O�7�+e$s(~=�1g8�J*Qxq�J�����

�=*4G;�a���* �ˍF��Wbdu���,t���h�����oH�-��,6Za����(�Şz�g���(�D�Ӑk�7~���!�W�dʚ	#��6�"� �����׮]k�zLB&+���ׅ�>�[���fmF�\�Ҡ7�����j�J��V�=n1W�ﴸ�[d��v۬0_ �򢹙� ��ƚ�Fm��D��4���WXə���_��)���B���Ea84�ˁ��l��gSc1�s|v �c�k3P�5�xKT}��|jV�8���)��Y�ݟ}Zv�g�M)<�h����B��W/d"I~����R(�tKUv$����Q�	<Y �Sa��_�����1������"`�&HX+����k!��pEr�����9��9J�	��E`q�=�v�NN��,\т��4�UI��h����k��b��b�G��NM-���Y��':+�4S��T,���K���&��7t}�~ވ�Y��cq���,1_�ѣG�v,�q17iww��s�{1a������XN7'�!����b\N���l�M>�:�%�O��e�$�� �>����Ԍ¹���C���w�Ⱥ�+ܑ16<�6�OQ���D���R/�K�]&QX��%���X��wB�o�!�W�O��h�M֊{�g���!�Lۈ�It���8J�a+Z�aT����'�Z�Ǎ��V�O�RJ�����{��⥉�������	�?�w����V���)�mmf��O�Ѯ4�Ap*E�፞�o�u��TU.\`+��A�*+N��Mk@A��-pM�vu�c=����=�9N5�'����ŷ�sװ0,AG�*�Y��������8B��u��5�nM��Ƞ�3���.CJ�@�S���	8\귝��@�[��V���_��փ�u̖>/C�&��Ug�Vb�ͭ6q����,�2y�<HPSy���)�#��MR#I�%SH`[iC���!D�R��ƍ�p�e�54:�pypX���zs���ymN��m��,kh�D�n>�
�t��.:��9�f��TU��E��g��²�nh�]�+ع�u���?���o+�xq�+b�X�:a4��7B�p���28@a�ː*v�3�8^=[.^(q��m�4�Q^�s�pTѾ��zƵ�`��1�;�v�!kTr���b�hYN���I�{��}��g�<󌣙�kמz饗���K�	N�޽�T�Vt�9�۔���&�edE�(*�����D�x1J�������#|,�3��QVm��b�0�Fu ͺhu����,���ܿ����p,�	#̖�I6kwwWE�b�"%�kg�UO].����A#&;oS������f�2Ix-����h,ZhY��)����L;��ŋ�"ߊ�l�*MH�J�Y��!@�č��G+����k�.\�m_�����w>�@h�G"Wa"Lܣ�E ��o�zT�v|Բ��|AԠ6��U�5�bu3߰��s���Wm"[����W��З�A,n6���}��g�i���}��ꦘ��������?�}�6� ����{�zY�!�lhۿ|��.t�4�"�@�"������5�&tfyZ�45Ȇzx���-��O� k�K'�N	�4�
�\�A��Z����믷6���־��ړO>�/��N�d*_wo�"
 �����Uy��v�u�x�N�����&bgM�衲�^}$:�<�4X�a������X�<a�^^����N���nG��9�"���@-ŗ�I�]�;�zF̫d���~����mf)R�6_`waX�CC�o]�S3�O����VS2<����L	�@�ʰ�Z��1u�´�ڲr`p�tP�QS�̱w[����b�R������cՄ�EU���#�f��\w��%����ǖ����=����{�����\ʭ>zpOv�E�zɧ}�駽Ņ^xakk���^YYχ=�<s�,����f��Ts�t�����3M�E�˛��j}�����d�4
��d� p
3Z�F�`~ʳ��I�a��o���9X�5&�"3��S&&nA"\UB�����`w�c:Q��,q�%�"��d��rG��vR�#�H��*�(房K�Qd��� ��'?GD�
��_�� V��?������G��W'��[�Hղ[=�C^&�:�������#h�|�^�#j�<3��5s?m&���]e�ay�:8���S3ꑊI�z������_����&Ez�ĸ6АC@!Q߀SeO�y��|��Ey�Y��7�|S�����ig��B�n�U^͠��1�&M�eW��>�����Ȉ���T*_�a4%f�+++�����P��f�`�f�*�x �I&�23�><����k}��k������ry�_?����^�Ś���*����G'�ĵ��v����䋝�@WSB2$q�y
x�tV�s���(:#�d��.�Qt)y��B�P��"���߇_z�N���ț��]�!��(
��h�G��0�Pa��$áH�g�}&����{y�l���<�ܺ \�� ���e;�QU����Y�'�#R�z���2e�d�1t(�(\sS��JΆ�rG�<<�8�@B�5H	�'[���cF�� [9 �6�=@T���Tk&���-֩Q"FV��S���rWc9;ÐR�-�_%ĸ�u�1R�E$j{%@�p=����E�`�Q�IE��_�=� �i�P_\��Lۑ�������������ͬBwG܉��A����%Z_�I�/H	���NdIS�����5&J��ra�k�;0<Q�zh"���`� �2�9��O6�zu6����*�����՗8>�뱆��*@��5�c�-=D�CZH�,*n+�w&���H�b�26�"R.t�9"(Q�R}��}���q��.�p��mL����C~u�3טH{}͉աC����u8'��Q����f]�ғmڎ���nm�S�k<���@#>�gi�3���Ɛi�0?���E↶~���pT����>.����<�ɢ�uY�)�(�ނ��m�'��'���fFpG����~/����mDW�(����H��xcI��TmI���ͬ��ڿ�&H�Q�E!�#ݴL |_$�$+;4��xn�e�g�c��j���^��#K��
U�1DYsU�i�"1�د`��;���$�OP��s�D�Y)�ӡ3T�lKK������'O�����sm��cs1�ZSű~��=�
7:�x
ͮvQ�I�Y��n�������Q��9�t�<9�~�U��7Es�q���Q��W^1��?�`P Wp*<�7��/y�r��x�P=�9��;��ſB���.�O*��E�_YW/��/{ۅ�����G�p|�6����̈/����Ϯ%�Dt��X@	�Wș��ֲ�^�c�7�$[	�]`{l���Qܗϊ����99�������Rc���^S����mbjD�hlZ]K{�E 6��l��P�/J�RU���:))��W_qI��N��F�}��.`kj/�k7�oN�W~#���n+6����r�\�R���,E�!�'Ǟ�攁3���(�Z�g�e���V ���eY��h���߾}�X�ʺ����4c[ �����r��.�p*�$rx��v��	F��0{ң���P���svk� ��ʕ(�Q�T�j���f(�'@m3���P�kpy��ce;D��A?8L�+Y���i���O>A�����3�(�yW��l�O6Iᦸ�U��*��@����"kE,o�i���i/ê5d�b����*(���x5�N3���B���&.�e0]]��\�F�?:=~����F�U$���N��U}	�'O��e!o��2�N{�׊�(s���-�R�T�N�u�q�	|�J�y0��Ȁ~�󍊵?�z�����������t�m
����l��$'��>����VK9w�xT��w���dG~r��d��v�ܺ���syR��^,\W��e�bW*+��F�ZOW�
��H�������A\=���`U��kͼ0#C$��=g�9D+h� ǹ?�f��d��[,Wg �m��b�~Q՘G>[qS��Ö�x^O>~����Ͽ"��G����_�������ϟ?g_ƭÃ��U�9T������ Y�n2�M�� 3R+Q��YZ���%"P���Q�a�&&�����hY�o�`)Om�t5�\�r 	�jQ�x�����~�D���-V����]>:����+�ϟ=}����b6�ܜ��|$�Aw�{qT.g�|7�[��h�'ǫ8v[��bn����7]����H[YT�1�碮׫�m:���->�-�^��a&�8I0A�ɶl��w� ��}��Q+*�%- �Ze�n۫�����}���)f�J\�z�Td}���`;��C҇�OP��T�t���\y7�&��oQ.��&N0_��E���9�̦v��s�aL�1��1k��\��sa'�L��^��B96dEՂ����#�P���u(���G?������ַD�$��O~�O��O3�O[\"y�D��~�ZT���}��/_Jԡ�[L0q�����a/n+sC�H��@�]�ҕ&��b�S�=g�1�}�E���X�vG:EQ�L3��巘~�Zi�) ����9J}�������j�Bg�u. 1�U.�!u:�����t���czD�Ads�!1�Z�E���`�)�M��\?7��Y+e���SH�D�`rV�u��-7����������0k�گ0�Ea�̸Γ$,����N��BH��qZ���$R�������jq8��ϵ��+=�)�`-������j��#�{i����X����_J�!����'?�я��g�|d�~F������|�����t#:�)F�ٳw�������}��ܹ�m}�����3]j�N&L�p<���`��,�p���{�E]��F���/8��,F�!�p�΋	A�q<��̼�"?*�Sk���M���$���3�TS<f|4�Yka�V�����S�t�!!��g�Ʀ�C*V���:c�������˝�$�ɺ��%}��7�SQ��L�1qȀ0�Z�Ѡ��
"�ҵ� M�:����t��		ez�&�ˍ ��L�D��p��i1�u�Z�D��CS<��M;���0p������"v���E_��������޽{j)z<�s�e���ￋ���Cֶך{"�E���Ɩ]����<e, �ע��I��G3�-?�����,ڸ����;OӚ�--�����<�N�e�r+6y��q���#�;9���'���ä3�&}y訶��a<1�i�b%���۷hA �)j���jt� ܗ�c���������s�Ew:�[3u�^��SwU�.Ћ�uU�<RX�H���J����`j���Ptt8�����(���H3�U<��9�v����(���Yq���UX�1M��~�\�%�գ�a>����M&j�1wao�Ե�DϤ���]�K%��?|����唶V2N��i�x;���Ob��:�4
�"���*)tA�����Q�]eX(�r$(��j@�5��T��B1���5�*o��C_�*�Ą�!)3(vb��|�1466�9��~��P�`J��!�S���"*5RM�7E���J�5�L6)J�O����˛`�DRY��b뱪��_�"=�wgEŐ�	�L���g:j���K�85il=2�� `tF R����6� .���z�5�F����l�l�Zs�K��P��7�J/G=��W�F��	9:uθ����l�j�>F��%L����z�d��������RL!
��O?}��k��L�i�0�Ωb	z�d�����DY1���A�hȐ�^߭�R��Lm�
�_�z:��a�z��n\�\.z���~���hm�<��f���\�+qddH���L�1ɔLz2�0�5ދ6�~�6\��� �b)Y;��R�YL��ˇ��aSi���-uv
�Z���NVZ�3�|��Vo��#S�J1%�����/fs
xW�O�{��Z��tm�a(YG�� |�O�K�QT�VGClSU�(���u����^o���ص6aV1۝����8���ܾ}[���x��_>|򐵸MX.���I�8ڻ�0�9���VJ��%��q���m"����ŋT�b��Œo��h6*����_.W���ѩ�
~nC{m���9��V$�z��9�@����
[/�8�� z#N�^7�'�@ڬS}QO��Gpy9�啟�]\L��$Q,���_+?A��}R�`��A��R���zh�ot`b|䈐U�y�e�޼ysy�`l2�B[D����5�ǟ���� �2`N���(ޟ�?"��?9�r�D�c.���Vi�4�p��@�!���j�5�i֣����;�a<,��MW �ї.���j���N�X*�	���v��x�u� ��߿��>{��G��7n���($�z�r�����b|�Hl��v�.�UT�Ϟ&���+5���-�֠u�!J�(�&:��{�e��eEx������~p��'���7��� �D�\�@MK�Qqv��莠�r���NM�iKQ �ܺuK�S~~1%��C��0S��P�%�S*TJ��@�X�Gm�uP;�X^�z��_ʝG�Ht�������)����=�լߌz� ���tB����V6��qZ����ȐV�ll-�A{��D61�*�~s�f%LR�A��uY�ow�5�K�=
O����4����rv3َت#�M'@S�H����g�H7��g�#���*m�|�\�o��o����~��?�e������j�q�"!���//Dc��ٕJ��t�l�.�!����3��cc#��~iW^1y�~���Z��yC��q��h�:���c�Q�����v3�E�B���4�,������BI��-
\�v8�Q���ϟ�>8�1�V�h�h`��Mg�N��1�}1�л����g�y���~H4h}}a���y2,Ca�@iJW�c��1w:���]�8;GYH���e<�4�L=����d�'�K!Q`p�W��������n���)ԑr��RBn[
��V6?9k�l�N���7b���H�+���������b��L��<���HY8Rm	Ҷ��n�Ț��r��aX��d�~��tqZD�{qc؂M�m�1�<_X:��BML��&��Kq����������ы�O�G�����1���ȼwg�e*1:�u��B�e�={6鮨*��3�էOVY*E15.�Ǐ˶�y��������-,��	[(�� �Df�|� Zw	w���7!�����n����Ip�O��3/xőqD��ʴ94��S��O���]������a@���2u���a��{c���� W��m�~Z����%��{�����_�e�t�b�@O*�S��.8�A�c����ȇ޹sG�#�)�j�~�)��[Y7�����=�*�a�^�e��2�p�n�?����x2���@��H�9�r�♨Ea�+�=��oE����>},�1�?�yf����}lw!������ؓ��2$�6�tb�|���8�եB`�-�
uٙ�mU�gw���)���B3�{�s����,���F�r�De�����ڢ�L��赳�KzY�_t��2dF���)��%�v�XQ�k3f=�e[��	%� �!�6r���`<�+e�EAu.b��v���4V��A�K��M�&:�9���E�"�[7���8`{�@��T8~P�جf�R����e/u��)x��X�N�q�:��ba�v�Q�i� �kq� {l*�u��\��v�`E:����3�\@�v�L"��.�@;2�J��c�S�^�W�P�f�z����u��E]u����AV�-Wl	!�`���]��(�e��&'*|�6�Uj���ޝ�"58/ۢ�a��U��3��~wp+y�D��5pSz"�mQb�^о1����aZ��X6�J{���5!o-�R�S&���bO-�qu#[���)d�2���刄�>,����h#�jBV{앣��"h�V٩X�J��h�v��!��/+4%:5R�I�����}|��gł]q�i˿:���o�O!�G�3�U򱘭R�őf�ţef\���G�Ң���A9����(�C�q��!���in�cP�$�ó{3cKW�?u9N�In�dá�ipe���-1=!S�"I�$����:�k2�Zv��/�k��H�7�b�{��Y��oC̀�59��c$�>;ǃ'�OY�)��	���x; S�	�����z�����6�A�J��=�ܝ�
��"�T�Hy4C����K��5Q�
�J������g��Ѹ��g���_}���:8>zYh�X�.��r��� wt�<k�f�y������7D_��o~�b6=99c�ωs���}cl�/ꨨ+;#��-�c�yR���LǸ�{lx���:@Fh�+�n�&��.�Z�����ĺ/Y�R�Y{c�\D�ĄN�pY_ב���l�3�f�I=gT��?���1��i��^�V���$E����۱�Ag|���T�}�M|��l2ي�nowB�}\m���')�MD�)*�u�����tB�Bq��Ώ\H�?�Q.�%	\�E�ו�g��p<��;;~V��4��[���d����<4��"� ο@bb4��ҍ����S�M5�C��k�k� 1'K5ƈs��ŲE���cpCAP7˺�}���R5�T@�᜼E"��9f��AD�V!�Z��r��R�Ԗ�j�^�+K�\J{��q_�z%�&�77���,��8mE3�.O�����+]�ĦU�)�T5li�O�CV����&�nh��m�����$�7N]�f1j���+��bq
����}��\��b
􄲋�S��4��̊����'�UIH��ͫ/������ф�q���Qt~��>�<m�Ս�]�܋U������["b$
��<��* s���ߓ�����@0��N�m��������ut%��-���ţG�>z&��A����i�	<�DU]`���7o�8f*�:2�^k���U�|Q}b��������B��.~��C*9���8�"�e�
Xc^�g7��b+�כ<6���ʨ�R��S����1�H���<Bm��C0����I��V^L��ϟ?.��ݻ��m4�bn�dҚ����|��[["�jN_Ҍ?K����w����ǣ�w>�@m��ry=1\q�g1e�(�1o� 7��*��if�&��J�l���]�{���b��ʕ�y��܀�|>��"tD�"��qw�
�1�2�+n�d�oj,mZ>�e�*6
���sC%2O|���"�C�-0I���v��l�ԛ�^j�+r`�j|�%��u)])�ab�bO!Fd�L#�AB�Po ��{m��xZ�Gܼ��������Ϟ=c3~��$��4�'!|�9R�D�a��&����]�8I�JE*M�
�%��2�#Yj[�����zww��X�؜"�	EL��-�W��Si����ܼ��9;��<���������������{�f3��dŒ�����hS�V�eM�U�SHS��G��	2��1���櫭� ���r6��Ջ������],;:����8o�qL2>��`��-�)O}1]�i\�����_�.H�#u���rc��L7�M�r!�����g!8��|g`��p��~ѽׯ�Ru`�O�+,�7�X������*8�~C����s�,������<ͽ��b�fF�j�����O�B���?�mJmv��DP��Q�D��Jۇ��<8��ó2�"O�Y�2k�SgQ���8�7oߒ��	�5T�p��N,�ݻw��Z��̢�"r1�$á�:2��[����������oZQ���2�B�Zό��7� Ǥ�Ⱦu9��)�ш��'�$�n\<�0���-7�<f[�a� �E/x��!K�s��jUer33�H�O��*m$Ѻ� �.j+�*�b�ޝ_ 8����ki0���!��j��G\$ŏ+�F[�� `"�l `��R¥Hو����T\I�OԔ��ʍ��'+��556�z�F��T}�	xe����m��H�r������S���JX�k*U$���&���4V"���Г�����6u����x��^V�Z���b�^�l�p�.++9�ْ��ͻ�˙D�r�ww��LX	�l�Fv����G]\�̱��ӓ��60�z/��	�;�Z�W�"e9�z��7/��U�F�+^�X̿,�&�Rv|{��{�����9gt���H�4���*<�M�_R������բbk� �����N�V�F�,R��mg��B
��9� js�
�KP�+m�s���(�鯯^'���C@^@��(�Qf*�j��E����4 �Ja����~l��x:Ku;>�1��Jir;�O�_,
0���Df{4$kRm�xaӾ������6�D����8���E�j�ָ"�|��o>(B �+uj�5�gg>����ׯ_���?������RA9�F��8��ɉN����0�m�>q.��{(���.G�m�'�lGY��k� ��m���v����lEҥ�Дt-�N�rG �	٬�2b%(�eY�k;��B�WA��Nh�&ul��D�_�c�{�1ώ�n�t����m�Jm^ �	�B��D�@��h���*��2,Q�F���S�9\����+�
�R��~||ً������S�]@�@�|��D�a"Pǆ��Ao�
u2O��j0� ��=�b���֌����& c�앾9��`�k�ʧF!:nk�.4�Pô���^���
�\v�] �-֥B6vQ�� �����¶��ߑNB���J�$6�{k�t�����$���k��ڊSD}�C�=D�afA��������U����uD%[,�P`^&��m�J�����Z���R�7��FUn�4�<� ���Z�䢄\�,G�0�D����Z"k�I,�K� �?������c%�{��U�r˶	�.�$�hg�l���A����M��3���aiQ�p*�������ʣAp�|���;`]��<*��]̤s�
D�����[c�����kӡZ��R!0�M�|�x����En�苵�Pw]��p�L��^x�<��R�0�ԡ�j]1��Q0�|0�G�a�����?���9{�՝P�T=�̆�*��율�f���JuG�:C,��b��:SJ�u{�c){��B�g[����{Q�]Y��Aqf~F��bj�F��8 R�Bϣ�9�.�:�O�Jl٭[�0R|�'��rvrr�P�����)�U���/�D��,,WJ��B��Ű�v���v��V�k���On���i��khZ6�uhK���/�ӗu�&Y��h��d���DK�r�dw�����a���D��#�o�	r^N{�i��\�ay��d�Ǌ�����C���,1�>kf̗5��A{��kc����?gO����
�FJic#�b�{p(�y���Jl��>x�@�/����ٳg|y,� �#|p�����m��l�l8�A�x�C�Y��o��oE��)�x��Uj�k�RB>]���@�r&�	`|��=�V�KB�����"�6��zZm$<=����3���r�Ğb��S�!s��'H�S�V]2ƃ�_�f�7Z
	�V��]��ݭ�X�İ�k=q��<�DR�;2/BEA�Qg�	�*�l��\e��\�2�yR`,Zװ#^�#���m�_���V��mdYb3de�i����?����ٺx����7o�Q�y�\�e�?���� ���T�M%����Z'��R@����v3U���d��,�����CƱ�ܓ��/rW<k�8�^��R�5��ĳ�y�V>T�������/����>��.eX~���X�ơ4�����b�J�����m�T��>o��'[��,���Js��OR©����4+��t�h����Cl`�~�k82�|�F���6>�y��P��t|���f�F��;g:,�<>�X��$g����ƌ,�r��Ր�� G�~[c�_���F�)�hV�ͻ��Ydx���(��?$
(m�x8�!�I�٠B��v��Ȅ>� ����j�j�������*F���>���Xх���ޑ�p���8?���ͭ�$�E�<�|Tf���~�|/�W�.`4kMyIV����+�c�� �rA���^RK�]�j!U^]Ցn���oe�W�5�!�4.��n��o��v�4df���7�=<f�g��ߨ���وu"���Oċ�Pԫ:�Ӂ��Sg秺Υ���.���uX9�����.�쉤GD��|c5J?tQ�:���8�Z��ӒY+�д!p�a�@��x�W�^ 0��+~ TJ�0�N]�U��A5�g�Xݰh���o5UD�l��{@͇1�*QcM	p����Ή�%p�	�ej�~a�\��m��xa|nʠ��(�֚�3q��P]�7�������u�����ngk;O��ˋ�p�����n�]���w�"��Jg U�P1/C����=j ��d���: J�Vk�+�(��*R1�?���>m��@�vdP%��(W`B��ln��D<��0�\Cw:ה�j�"x�)[aM�N*�+o'	�6;����q���B��llp���F��_�[5�q��q,��v�����|^��3�%���@�q�?٬LjQ�X��.m��m���q9v~Vq@��/bWÄ�q���4�.�e�LV_c�7R������3�C2C�a1���G�����U�ou�"W���:"x̍rT6�VB��&(є&�nܼ�V6>C�xU�9�G������18zT�ʹ�#w��;��~��-W&�cO�5�G1����تP�ѳ�R��2���r�ՊI��i�jS�4��JX}S�`*��]\��j>�sc-��
6��C��+V(�u�${���`4����Z#�`g륲�����g*N���f�����P�Pz�,JG�i��4=�ç��h,���~~~:pɗ[�O���p5��y$�ޑ�Mp�nܺ%B%����S%���:�=6v*9�l;���ZM�a-����\�ζK�3�%��i9e��8e���S�Б�N���xq!N����8���@]�{���RM�+�k-B��8� V�^]L�8�E	��3Ȩh9�:��xRَ�Mo� �<�	5��Y"����m�g��_#�a���gl��G��Ťb����j:?����-�f��[�6yX�G\[-<� �����136E�6SصȖVr
q@��(#ŦU�؛y&���{��H�sq��.JY;�Qw��iu�x�]����,V��^�-�0~x%,��aV�/��UU��X+/q�ߛh:�/�[i"����X�%��!j (��cxrvv1z.t[(�.�s�A���s�����x�3��Ҥ��k_C�f�!eD��Z�(&.�'�v%�1'�.f�*7+rg�r1���k���$��7���Xl�C�<[w0��VQ��`��|(�Sh������ַ����D�v{N�\?N���v������7/ϓ4�l� 2�W��q�LS�?J���^t�H�";u�`������]1O�t���)[ ���޾?>=�0�IղB3����-���1TА�3bD&k�|��0��\o���Ĉ��j{M�/�b�.�iWE�:�&Զ뢘&H��55㙳���A�/'�!Ub�L:�d�_+Yy��,�y�]TXjL]�zS'�Ǳ��Nj�D���Aaf�iz;c`�vw�����0s����NK�!� �jU,�}�s+Lb�}N
-!���qt�|n���X_X�f�2V�NfE�\鼸ĠatިX"�O<1qU�Y��k
�z5�G���N����)����ވ�`f�#��G燆���s���~�w~G�Q���ླ$��-5��|���vG��$�3��I1zg�=��:����œg�~���	�w%��&�R�h^�L���,!0=DjKy@Qq�4lm�ҍg���_pd�t��!�[SxF	WV[�����r�[��]��@�)�5�C�����m}����fk��j?���T�L�pט^*T�N
��b.�Ȋ�$L5��K��fz U�\�T�{.��a�/�!�soe���H�O-+�ₒBT;\�&ߙe��KTTl�t��ߐ	J��������ރ엜q*y��GstWd���������e����ζb�"�/���3�P�/�8�g[��Y��CN0WZ���0/^�x��!��o߾-����Y��즗s�8y��g/E���l�L�=}��G�)��z	g��E{�m�����׾�u+��P#Q�K9L��E��s����O֫U����P��j�ȓ�Fc��-��1&l�Nsq�Kf�h��Y�u��~&�R띩��dq6e?%���A���$i�g�q��DVp_�4�������9�Г�j��C�4�S�=0_L���\+6S(T/�:ǌn^g��iU���9�̎�ٜM��l?���g�"a���3��T�.�8�Xq���i�<��
���=����5���ꇉ�ޠ��Y�3s���[��+)����D����:���%��1�N�������>�ZL���~1�=���W�V)7KG���<����HeK�7�@+���C�E�3�.�	n#�:kgf3�f����;˅"`B���{��E��X�BfY<��z���:��脐�PVF�E�"'���nv��2u4 1�%�bP�̙0|��TFQ������/�����ҹG�r�:T�b儙��1�׋u?�c_����S�O9o���X��t}��
I�]I�]�I�8�՚fd���F��V�L"a�To�jN.��!�#���dvq�A+��bwtvt�l-�C�z��Mt���(�|$F;(�Ν;�LO��:a�B�.�n���s�*�e�����}���0hv额�λ�ǲQ�)e�54"�p�d�8lܪ��S[gt6���/�0���F��E�`j�[C-��쬱�������ƈ�#�ߩ.�{��>}xK�"��˙����Ě>�y)��*�)jb��Z�F	z*�Kq\B�+�Jofs�B���R��{���Q���b/)R��
ա�he:c��:P��i�{�?'���`0�*�5�������g(�1��+7��lHw�9��w�Z��g��Ԫ��IDFt6�(1Tmj�8�ph���k��RA�/��h�~p��S��:�����Zgә�}�d�ۭf��i�3�W��4��˰/_�|��;�ZL�SD��<�3�Bg(t�.j�}$N����s�µ].����U����b�=1j�&'��b�CmA�s���s�:��	G?��L5crL!@]��@�jڇ�����8U��\�O󃍁�αFY�Ov���/_�i/@	L�� ���N�ƴ)��{Xz��Um�㇊;��u+T��H�"O.�٬7��욄Ecd�ӌ�6B����K�x1 �Dӹ| ��-�]#���������Y�n>He�'/��1��߿������=�7ӚR`rpxd�rل�S>�t���$�A/i��$6�oz�lA�-iv ��D���]ʇb�o׽?z+��/0�o��w��5�8Oґ��ٸ��;`��W�`�~��(�l~C���X<�PI#R�&�{h����.N�&N���u̍�{�!I���u���@�3�s_�^��Jk���!�D>��9c.Oc�%%uQ�y2�xU��IEt֞
=xi8�蘍ԡ��ˑIa��@Yg�ժ�Mnj���1D��J���6	�B����Nj�'ةZ��[ۑ��t]��+=��QY/�^mlj�����<�z:��Y2	jB�����V��# ��C�@�l��^�v�����D޹�5�&�|ߡ���DK��z���J�<����� �8�BWm��B��S�*�F�S��sc��~��[t�(]�'�Og<nnc`��5ј�f(N
"o|m��XG��~��#y��Uew�W�ӟ�4x�lPp� E��kz�":c��_�/�f{�������ʃƒH�������FH�Ċ�n��o1׶S��i�]�������3�m~V����<��)�qL�1xK@�g�z�:�:g�I|��Nۣ��,VK���nݺu�������W��kP���[�&n�ڐ��%���Ǩ�����?���O�YX#1�3^
7�rE�(�+����q�_(ݘ��C�4�O�����������ed8~PȻ�n�}�V�W{f�F�_�q�%ʹA�&��f�ꫯ���~6Y]k�(j�q=ù���@m37�Ð=�6���@N���?����D&!�f�8�}6>&�\��3�/yj9�U=���'5dm��̈��SJg��gU+Ѯh�Ȉk�o���~o���g)��Ǉ���m6w�⬥:I�܉nc� ��<���"��������"�B΀�l)K�ҲH�蔿Z�1F c�c*+l����µ�� 8�*2DsX��͌6�	���0����<�N�7� ��>�qw���JD�]��/���~�ܠ�v��7�8=~�P>�k_�ګW�����7<x �+)a �T�Jn��ӧ�?�ŵk��o����?�9S'�����x�ƍ����w��D��'��a.����"C]�t?���1 �Lu�.Pg��`:�� 4��Xb�5����[�M����Ln�§-ν�c��h�.��$�b�[�l̟qaV��B�G-��b��g�:D| *Lz	g�i ��iuX��5��!K�4�2�q�c�횞'���s���?:��L��B>4�G-��6D�1S3Vm㬼�mL�eH�w�k�&q��%J�OF~
!�iF��ڠ	� ���GG>�͐�i���:c�%�E�U���ԭ�Nmj!6Fd�SH����%��և|k����Pn5:���L�����eq�,��]���`��B���cU���t@����7�;�	�k�D�E�����C�[�:��ED�7����\��[Y�Z�,R��n�qg*�p�z�ۘf��~�U�hk<o��1��ڤc=3��X��S:�+�����|��eE��_�d��
��"-���uJ�dr��_?�_^\���wX�>˄)�	ԝ�|D��K����l�)��|u��m��#;G��� ��3(���N��(	������w��,���k�j��$��䓏>�}���c�T�HRU��4���u(C�N�k�"��U�Z͢�G蒲��nv�3��V�X�%[��ɏ���J��\x]�Hd^�u�t�^REM�%��"Y$F��\�O_��M4�3��C4� ��l�Q1%ɀ�2��Pư[�ILD�i��(�.{n�XcW<�,��jg��Y�'�+�X����kj�6/4����Br�L���(��A
��^�o��'wv�l��X4�|Z�3V$��M�~%�+���1��gIb�B��D���i]���\Z]�j�����X�q%�5 �����x�������"/�K]��Q���p���(r�d���y�D��N40Bk����rfI��2ڙ�Ӛ�o��]�}m��;[.�F��r��8�K��v[U�`<�6�Ч&1d�X-��S�~��(H��3/oS�j<�j*Lä��TI��:�m��4d㡧R���A/����D)��2�g��]���b����7�:��V�\!y!��u���_�M������r]��^��Ȱ�aiJ�TŦ�ٶ��h� ��J�@�ڢ3�$Ü����g�Y[���^��C�!$V^J��ɓ'Ϟ=�J��v������k�&�[�����rr����C��\*x?P/���l +��=0$�i�:G�NA���䎨��7��h+t'�SF��8�������g���?����m]ɖ���2��S�\�}�j
���h(�l� �<:>֎Qj��u���{�n�;9	�uݶR�=V>�x��$a�|tt��U�W���T�RK�j�Ćp&��+�G_}����h�KYIE����pW���b�/P+?�7<$E�A��e'�?��1_Lk��Fv#�o�qȝy�i�}���Z]�\ē�`��$Y:01c�I�k��t�V���&����[e�z��o~S�1q� c]���p����J,��b]9�*[�l�i&�I��B,fcE-Ai}����.��P�v��@��{��	�:ğ��PNP���W˪h���8_����k{�$_�~	���ݣ�ɇ~x �����EN�,VJJM;��;�D�Π��q,�|R��Ѽ���,�,����)�A�i������g� ?���X�;�3�G֥� ��P]�m�9��򡇊dbӉU��*���G��W���䭕s#[�,L�"~� �������>������[����uC����q��*I8\�F}�2�B�#��|cwr�d�@��O�怱0�e�6R�r!�-�S!A'��� =H͌�}9Y{[��*!U �y�!b�V�zVc﬋����Z��bE��Q�[>� �xӁp9���k�h0#�	�ez��}(
j�Z�n�zwP��Y/�!�FX�3�**�x� A�͛7�H��������Y���pK�:���ulߍ7B��Yg\�~ql���ձh5~)�J�ݢ32� �n��W5�Z�#� !VR^2��J�dg����e�OR�%W-%����禤��ͰΉ�3n�x̞�t=L��N#>��X�
�,}N����6��N�Al�[y�_��_Er-Ϟ�x�7j�ؐ$���Ǆ��X�[�����_�v1��������[�v�**9;����[<ˬʄ�MA��S��F穦��K6�c��6��<V�`bݾ�t��W�u�G��
 p�(�f��bU,�1�����2Z:ߠ-���z�f��S2H���8Q/L�B��f>q�,
�&�V>g#E�ޘȬ�\��
��*o�@����)�������b���Hv_�<ӑ\g����f����-�K0��F�����eŰ&��c�G���P~�������?�q2�h�˿����ʿ�.w!�C*1\�����_��t%�����
|p�zr~���S� (&���uiӊi��AY�`]�.����9�mL�JN�u�o�yf�	��#=wK+ ���5���A������q�]�Q�ڔ����7!���������D\3�$��`QVV;��{��u��F�OH=[.W&��<��A6��eh�W�PRTx�"ce����g'�UQ���q�l��<�.�-���R�CA߭x�b��k�jlpt�EdS7Y��ҧ�ۍ���C����_����$W����������j��$����C���/�/�>~"Q��r��7Ať�j��0ϡ����LJp�yصF7��_�b6礀pZ����[�W�c�ڧGCY�5���ӏ&�$�����Pd�ɟ����\(�j]ˉ������Ti�h���}���b�#,��X���b�f!"�<
���<�sT+��Ko^��˾}�n��?��51I#�lr��r�:F26�m��yk<���[�ob���#}�x�9���2זz�'4QFO-v�8��
o׊Xuk�xl7����3H#�A�.4`&���NJ�a���z&"?���i�(g]�P���N3],l�dbb�E����?�"�:�z줝�z�H�=d��ވ�a-߿�j�j�vw��9�r�d�NV�U?��0@n^�oa�Mig#-�ҥQ���y�m�Q\&�'�7�VG�"d�U:�) N����>|��.����۲jհ�oGÞ2����g��wkR�1@ͫ�&"���o�SH����[����`NBb=��U�]䫑���L��l��56Έ67��j6#���!Z� ���nd|�!����{�m�m��±�V��׆��3�'6����HB��&S֙$��WNd\��߆���5�{�m��7��.�D��T��r�G�B�u���S��ܗ+E���e�=-I�Jןu�FG���y�=�d�K����_@ѦD\�Z
2�d�c2�{��-�G�|�m��H���i�F�Ɯ�hJ���";����(|�x���I}j���o��}	��Vq������Bp��k����~�ս�=�D�i>Mn�,7o���+"D�����J{]���ʪ�4d`0r�ummJ��%���Fj�	��F��-��
fl$���7�[����KQd�,RB.q&d�Y2�!��P$���Pd@<Q��X'S�(Z��ӣ@"���_*�Ä���.^?2�E��&Oc�Z��m=�6��r�Bǹ�y[n0�1/2Ҁ��4�a�LF�=:>z'N�����O>v�ķ���܂������Z?G�A@8��c��o:�ᮚ�'�Uj��ÈLzN=��J%_-��,�aDLnH�y�nT�K��J�N��Q%N��~���>}*���x�
�ܢ;ѻ2=�r�^z�t�4�׀;��Xצ*C.�U��:���b�Y�֣��PR����G2�h�Iˍ��F-�� 9e��q��{�dw>�sGOb����"��~��Ӿ�	T���1�󩷡 @�x�;�pg���\�38�d�޾�eUj��<?���"H��0��9�׼O��]� �G��r%Rtp����|*Ě����ݻw|t����%��d}4�cu��pfb�S�v���zO�j��@�&*�k���p��K�akkVRM5$��}���$B�H��m��u��:~�^�L�6�ۘ)<_@f*HM[/�K5y�j�.Hś*�Q�Ib��V��q�.���:�{���e|5gl-;���M�q[/��Fs�̔V="x�G�\~,.�Ge�ʗ��%Ҩ�X2n�RM���rND�2�u��߇�O>�̰���o�	aR�h���w꿾zw�������Z��!k��N�-C+�����r�A�ܻ�7��!�H����nf�m����bJ.$�ZkԢ_DD[�1�!2�=�"Q{!��l1}�_��� �W �LPű�:+�D��#���au�BVQ��_��o�A�*CC"A�R�iN�������&��m��0��xM}䆧�2�����-��+A���Z�8t�ӧ�e�8c$��B>%eEN_�o�e�������L�m#FQ�}�+�\�z`/���G��p�3d���jHx�'/7[v$3���6�E(�4�û�v����L���5̬o�w�X+㑀j� �_"66��:ՇN?���8��Tt)�����h�:�L$���Jg yy"������}����.<lQ:��kY0�L�%�奈E���Pɍ�c>>��~}�;�����|��i�a�u��t1�K�*R�G�w�R2%M�$��̅V蘋Ɯ��ʖ�������Lq<Pe���M�+.�p�#K�;�>�Ġ+b�'��V}�.�_b��/:]�N�����ǌ�Ƴ�:˒+�#'�ua��#K��܅�&�બ�:WF�� �d�}�3�h�((.�H������L;R%:�.�r 6����s��%� �E 6���"�O�0��Ȇ�D�?
�(�/���ɩ޹�6�>�)7F$�/�m"e�2����@���~�bO�<M��9l֝�7%<ܿ��� DH�!��s6�Da#�j�7O}��䣷⟼}wL�?Z(��j� �ź5��ب�ɻ�Z�H��k��ă@�GuATu�S�u�ל�eq�� 2f�	�T�������Hɖ���G�AW�yo��x4j�fm��./E��=�ѳ�OQ�l�TEb]-�om�0�%�p;�z����T��޼q(�bzv*�sq1.D�I9T6Z���N�Z�V2�n,��4h��J�N9C�7�
+f�m<��J]�^�BF���(	<�dj���z�Qq?V�z�a�G ����y��rem�]�\hc���� %��W$֙$%�Q~��'�gPJ�"!��W�F�Ҁ���O� O`�.�c�KY�v�l��K���_����骚^�$&?;9}���b�x[��d�ǩB�[Wn�x~yr����R�g#׍�~�"h�����M��p�B���3�#3*�	�%��d�;�{bkYrx�T�����F��a걾���l�@��o�p���q4Q4���b0�p�S
F�mL����ek���m�u��~n�Z�[���Z)���i��8�6�/Jw�v��(HX���v§fd��1G�$Z�R���$�SH\�tFg`��y���w`�Eb���x�U���Zov!A�b��J�Y�-�$ײ�n)����K����U�,�5XT�����f��v�żZ-����q���rv)�'��&�em]T��񲼤㨝8��9D�M��m_���]"g���}x탬sb��Uї3�U�^�钺JW�AT�a�5� � �\Li��I|3K�&{�[�3����,[j�;A�G^��3��,���ʱJ|{L[(�*��E_%:K�諯�z|
,���7g�u��l��,��3�I�0=�+��m�v)�M��6PrWv-��V%J���J�D͏�Q���Q����r�@G�L�$qm�)ﻻ�Y����/H^NǼv6�6�[��g,�����\�ƨ�����G�G�0��ؘt�dkѮb|���iO4�V���1���3�F��ױ�RN32q���h�$Q޶�������_�拣�c1��Ȱ�C|]� ��SLש�i�*���/��b�9BI9�V�7 �C<5z��,[�=��bł��M�C����q.6��=QHoՕ��r֡�>�گ��_����O~���÷o�"0�*#8
��2zQ$;��mPΝj��E�Y��¸��bg��������}lY�E�":�
��`G����"K�� ~�d�-uzzNm��`�(φ�/� J'$h�#�w�C����31��������ݻw1 e�ӥ��4�=ͯz���[����u%��$>�潍#�C�лN���yU�sh&&�&�p�z��H_�ӱ���gy5��ڍ�O�	�C������.��v
'�����m��k�:h�p�(1�U��NW��3%
gJ�	%L��+_�b��2R�Q%Ӡ{����eA�X*���Ƙ���ԏ</��$_�΃��c�}���?����O�>;9=����6�Q*g����e])�����[��D�؛5�Ej7e��X�S������؟r>�]d�Zu��'�����6#'���2cf�S^�R�m���ZU���[2[�!��G���qv>�/� F�᭛䔀��;"��#�Z�������R·Kl����L�E��C��̴�s��;m�|����bV+9H��R"�s6�ݼy4ݾ�^���?������TP�>�U��[ ܋��R,)-�l�p��}���Љ�YD���56`���
�a"�<���Aq�X�4~��z�h�scp���g	H�V5���b�<3|�V�����l�Ve��1�٢��	��E;:o�O�o�פM3��Ԛm�/:���J���P~�k�$*�PD���?::�e���C95L钷k�XM&u�5t�Cޭg�4O,���ڵ��ptܝ�1�V:����I5"�]݈/���+uޘ}q57�R�I�mP�+f��C��3V���T��Z��{�w�����b���g/�E�o��Doww@|V@%w�[�����Wo���P[
�׭�m� �[7�z%�6s]1�1�	�;�i����Ipx3"���G=� _|ȹ��QN(�x��{��CB����Yk'i8A�*�sqj�o���=b_3�t�E;���@�r���%�����:�� ����R�\S)�m</�*-� �2[,օbvx�=(�ot�CܑXc#ߓY۬���ֆ'8�C��
��y��aN�w�"Ht��0�N/ȡ�����O*0�B.��&�����vm 57�P�L�v�S��ɑ7rj!e�� �PQ�̆���g�E��l��0�!>�d>pε;2��j#%@�����P��k׶0r�D�
!�R�<Y�d�,���<#^c��;����&nK�L866$��_��8U�}?���3��[j-ge��hjaĕ� ����)���?���D�_>߹w�ާ_p��-�}��rEJ7�s��Pu�9���h�+&n	hO.�i��9_Gij ߵ�9hZ�P3�C��;#��@N�	ź��b�6��r�D!�,�H��Щ�Su����.B�������n��#�bO�A{ty���,�dk,K'�ٚ�~��/HE���<��_��O>����0�� ������ى��H4���^f����wvIJEWjK��U��P�6)�i�x�F�E���0F����	zn.. �M��IW�lƪZ!���Y��xc4�ĭT�r'��@b]�N�[����-[ �����&�6V��������Q �\I�A4�<�x����k�������qo����[�h��d}E��if��l�=3�20�߇�EJ���h��"�b��=-�m�`P��R��@�Z�}F�ʲ���UdyKev#{�'aS�r��@M K�5�Mx��|5W�]靐RL7�Ϝ���X4ʋ6�ɹ<��S3��Ҡ�u_�gz����S�	`A��
�![bk���A]T�a�^l}�\�ĆSM�ā���լ�ۜ�v�C�����|R��2�ژ�'�P>�+��[�^f/�����~����?}?�D�a�Cx�"���ҷ�c)꣋=�+x��m:�>� �smgg2�qn��F�D�C<�"~��qJ������n�)G���M��e�v����b��w���$��2���)��β�u哪�������H�j�{�<�SK�'�:��+��-.5y!���a�1bd��h�v���r/$~�Wʧ�������$�+�E뫦<��M�L�t��kE�Γ��Xߖ�ڋ�@S�[��*r3��]ޕ�sm�4�fd���^�Rl�_���+ �uI"dٗ8��������zL�Q
6��EQQA���T��
�i�G':�2(m��z�N5�s�u����b�� �+���쇸�\�~m|k�r ��ؕ��F����W�T�H���ڰ�/ȧ�o޼����kM,�/N���y�㖦Wԙ�sd z0���
���	:^G}�%o� ���\��Y�Nk�:��ݲ��lsƚ�h�Q�._dJ�$~���������+�d�q�����CQ��{
���);�����|A�)�YPH(rr��Z hq����'20`�m�����Ov�Q��Ҟ����ߐ)��7�l�����ap�����?�*ɚH����JY��0G4�>Me���`��ٙ��K������#��a�s�C�^�#3�]��j�Z���:�g}.{�mQh�g��ߓp�勧"]�.�������Y�f=�-82L;g�S���Hmh��s�r�&J����Cg./�"���������:f������Z*��l?XB~tQ~)�q��燇x^�@�c�0�֘ac?�a��Bհ芶��zdl�w��oTȩ(գ�y��"ΞSgU���CE����A�,}��0&�qZ�� b�8g�B������*�N���x�Јa���@w����G|�)/'cZ�T3�&6P�|/�n2�;��/�1���''�lr�R���`�^ �����to0g��݇�����G}�����������������+��k5��BB�;{��@��ׁ�˯�8��{J�k���l@*���K�L�V��2��A�͑�sU�<�2��
�ɽ�o������n�y��Po5�)��Ƹ��7-����:�1sI(�D��*zq��\\Ȟ�NP-���Ŷ�'���:kK�*r8�DU���H׵�n'�F֟+R���t�y��"hH`N��U�k�N��M'o=qFZ�RG�M�y��`z|��B}.~��jq��{�Io߾M&; �+�8o[񹽀�bN�p�>��{W�j�/����.�ǁ�E��=}�TU�����`��l���0�'G��?��dn�Y]k��6���@�M��~��i��C|[������E��c(RDg�K1�T,Њ޸3�7�^��{p�J�{���?�.�Y��r�wM�ndCL¦�.���,:#��l�##Vj Q����C2��*#�ś�Vn����yJp�L F�k���G�(�܏���9�ɢ��D�5�̠2�R�Y�J�ly��(�ʈ��C�*��g����o�T�r9��y�.!�f&�p�;ň1��k�N�����ϟ�˂��6�,n���p�,3<��O��*�w�������$$�	Cs7u,]����X��G>cjta��(�\�PI��5�l~����:�K��C��ڵ=9�+�`kN�w'����8y��j��Ōs?v�J�����q��L��
���' ������ᙊ�@&�3xx��?�L*�ɢ�p�*G�&�\�Iww<��!��2?�.�R��F�cg	��O��:=���������ַ~㷾��YDT,�
��U����_6�r�V/��cYgq%���/�L����"�8�:�j�5��c�G��x~e)�O��kW ��� �ԩIVrj�Q���1�'q�5`)��& �:q(y��7Y==8B<�M�o��h4����g?�B��9�\	R�5|0���� ������q�]߹s�ѳ@tsg\�Y{�(*P�EW���� <�h�j�)�,l�Ũ����E{�l��^/.I�����@�^T媁d�'�x���?�'�~_�X,�,;Fb�'�2����t<�4��i��h�q��rL���@	�Ɖ�Gq�^M�(6�y�gO��W��|o��y�n��$�s���<=���$v	�����͠����ۆ���8��]�(r�9˰ȏk�u�����F?��m�������5
=�P�/tbg��ԏA�:�_��@��I��1�/�ayvo8`2�C	9P2�Y��5��G?�^T���JfEN������%:=�8��V6"�YZF�r���^�5��߸�����8c���Z����X��ILH��͛����_��{������舗��n��r�駟>��������������O�{m�tx|�����X�>�s,�&XS�	��IhcPҙתR	ZWQ�y�dv?�vH�,��ᅜ���}�vz9'ꊡB��S�穅�1�|/������{2��tA�#x?��OK��u��q�gg=S��Gn-�at�$���mDgU��`nHu�H~��
���r�%��O�l���{C>���I�"DL��Y6�\r�����3[hxز���^f��TҰ���:	h��6:&��T���=�3z��l)�rE�`�䮆������8�h\-��}��p4�e)�b���}/�LI��Q|�����]���7�������S&����7o��IiH5��A���� �z��Md3:���rH�������=��=*�y�B���_�O����^�CX���P<~����h���N�J> �)�M$A���Dϊlz��f��8�JL^����g1��<J��U�UQ�\�uk�3E��S���c-�&��E��G���?:���PA�"����e10eQom�u�e7��ť�@�>��7���:y*�ݠ?J��A�q7� �,8:��1��qh#ˣ�������`�"�y�|m	_�@3Őj�Ko߼B��m������D`��@�wi��a�.�G�L��u�pMv�s��ͻ$N{Yo4˩,֗ ��"����Ԝ��{�㫦��Zu�RUC& �Rd��T"�I�c�B�Q\>0!2$�N\���(��c%@�,6p:��12���*��h{N��>�/���իgϞ�qE`LOz;�g�A�6ӑ�Z��@w7JT�Z1��O:H(+�� 
�/��*�i��HP�j���kre�I�&g�h�,Fis2��z���r�2�4�� �9�I"��Fѥ������|Z՘���G7�hUÕ�q=��\��*=Y��jQ�Q��0;p�<�7�~<Idp^vv3�У�0J��^Ӌ��k���8�l�Q�\w�d0�e���PRe��K�m�e�Z�7�Iْ�
�>'���߿��=��o~�����\b��	�a�� vV!n�]�1<E�N�ߜBg|�M9��X�{�\��5��w��!��<8}��̙B�;J�����vZ�\�`3s��{͞�����>���sE{�b7�]ʇ'��R�
]�?�3O�$*7#�|�S���S	dT#���3EO�`p||��:;N��r9R"*VM����]�fld�Jغ�er5���l}�ZuI���U]Jx�5t��c"&��T��-��dMl ���ΚOeH���dl8P.�Y����t(]w��B�Is�5��!s�����e�S���W/0Q�)�Q~��o��O�~tt$�F,�_~��.tH��eܘya�#,Bu¢��咳J�{`1���I�p���A��O�X="D�LŊ�	ܞk8�N쑏����X������E�˦X��sp����Kɹ�㣡��e�[n_�>OQ�3����1_.f�y/�>	k�ϕAld�t�lJ�����05��X�xZÊ1���R��M�e׵ع>}��j��w7f0 0C�#?I
��O��>��?0�*A���!0 @��io���|��^k�uΩ<��W1�S��y��s��k��� �I�e�u+���/!L�xa�Z�4�˟�1����c��斵�`��Z�&T;�l�ڙ��YN�$�)�k��\��^�x\%˱�~��%�����6���8)��\R��+yg)C��i6�/)_��+��0c��;���յ���HJV˴|@h�qo�cqB�'Ǭ_:�[��@��O�J�̽�=���k�.^�H�w��?��?�Z&�����p���P���0�0�q:e�y��6������ښ�C��ZvųБ�%�;��d��]{\��8-;��b��an��,���x6#ý��8����\����,ϪY���i5-j^q㫶jö��	4�S�e\��V�tl��Wk���&�I��_�����T�� c���A��n�@h�g�g_��o_�yz(p.����-z�B�/+N�#.�I�FH~�tp����!02F����*E�o���V��Su��%��~�h�tᰬ&���w�
��I��md9�V���ma�n�h��6Q��f���!RL��1v��^&h&��ʙ3of���*\��?�x����H�Q��RI��G��;dbI�%5�R�g�o�+}_ވ\eWH`�1T�S�]O�i�����?���VlLk�`����R��-���@]p�+�ph�@t��x]�\��p>��<U*v �
#�38�k��: "�Q}����7:p��AE�&u�DDzә`���UnFx�X�[���y�<w9���bS{��������q�<�Ox��%:���W��j��d�w���e_*�/���A:R7��f�+��"��e������kt���`��tA�o�_i&n���{��~h⬪l&�9&���MZ�K�[��9��6x/0r�5����԰�/_���+�̂6�V��qK���"PXV���������%x׶ݸp���_��>� '��O׼Ѻ������(=E�W�#��Q%���dZ%+M��\��i%_2����Ƚ8��e�C�2����9W�úe�C#��R7��9w�����K�[�a�����!M���O��ֱ�h#����2��`�������3�9-�^�p/2�Ԕ#G�<ǂ�h 3�$>�Y��V�ɎGTB�&	��Ŏ�2�nu���-������cqV�{`�/�5J���ϭ�7�I]�$��&K-�pm����8r�b����{������������_H�\|���2V/PtOeQ��EZ��@��-m�.�La�t N��*��
%�C�T�Xk*|d��"��Tdޕ �v�ӌ�c�{�#(��ٔg���L)Ұ��H�SJL�����˱GGF���L�3�B� p�kdl�0��̑�s�*�o4��Im�S��3>�ڔ�2P���F��W6巣?�*ٗ�:�M���b�1T���\����7���^{뭷�!b{��#;�)��5X82b.���|�)hZ�����-�=Xl��bIڲ��V�f�f?iD�uez��AW�R$܌�Q.��2�7��[l�V4��BQ��{��O��ܕ�uk���ڀ�U�zX�m�wN��e]ξ�9�B��4�Ӑ��0K���� �P�Qʈ\	����9�{����v(n1�;#^���Tbro�Y_������6��EK�϶h+��P��Ա4yҺ�muZ��e@��:+�:AK3l�)Jmr�c<��i%�Ν;"/�[��?�$Ҫ����e�窔&ĕ� GNH����֤~�����L�L���'T�� �qX9�,�N�XH�"q��"�p��CXთ��|�ͳ��0�����j��{{�{������F�j�z}n�`������W��F1gC�K�hϞ=c�����'�P��B���GX9jl�0Q���<#����֭[�ԧ�~*�ŝ��X��V+G��;wT�G�v| ���h��%nJ�/s����E��g+����ʉ2~B�\�~n���B��y.�L���ʜG�Ԏ,,X��5*9VVu&�HJb׮-�q,EVUQl�������Y�M��cA��m�����OxHdL�8C��ȣH�1��=��pا�ȇez��-EJ�#t<9�X���K�K�o�y��Xg
���Ǐ{CA�A|���ؑ�������>,�m�`$�B�WΡNsZ�5uӌ�Q�&�)�����v�3ο���[�2�![=x���<W�q�?:Ѳ���bH�ry���X*���V���殆�8�s����ʵ"���-����I2bGj��$84tHvu`F�"8b� �D:1�+=����h�0�X-��K�4/�ӄ>��*"v� >������J/�5r�w�kEӎ�>�0K�}#;�˖:�#�\���>��:���	�e�� �&.�g�?��ˣH'<N��=bnZ��/��}���a�?ts���:,���b�˂��L���;_}���Rh��>� �_�x�Z��Nh��>a&.�'�kI�J��t���>��d"M9��,�#�#��L�a!q4��1��}*�R�и��>����v��hK�B<9��_��|r�:�����9j�`��r�t�����{7o��:�H�f��|���W.�д17�(x��ݝȌܧ�9��ȧ��n2��DQ�b�訅e��hu;�׫z�B)�^㖁�-��Tt2��q����wĝ����:s�����5|^D��E�> �$��
qPFi����0G��9��,ΚH�"�����I���]��B	`#���t�Щ0��+RU�6C'�5�p�ќb�rڤ��i�&�R�0BCc8ۇ�A\k��3իM,R!@UF�i��&=�IB���p?A
����R��Z٪9��C�B���҅^�Q�:�BIC�U8�o��EKy'���K�$�K���	�L^�(���L�Ox"��h,���x��~�iK��쿡[�/�!&�G�ˍ7���vem,�l��y�7||2;n�RD��$�
C�#Z�IB��Y��TE��t���<�Y^y�]��yi��hY^�����yu�>�m��ZՉ݄r�F�����y*�\1�x�3p�\�@�?�Wsα����.Q;��ne�A��3����5ك�� ���~�Y���f��u�z�Л��صر&�
Rm�ʓ�N���$>K�T��]��H�]u`�
z�U����͞�i�e�j�#���d4<M��H����O��?B>#!�Yx�=(�*6�]��1���g��'���nuQC���s�J�k#Ĺ��e�2l��a��xM��8l��}�:xE�%�o|�<����{Ch����v����yd���zse�Wx�zF �m�~J�l~㛿��_���/.��VX�&�fU�EI�f3����m�����DƱUu;�Mj��Z��I�5C�Y^ADeZ^�e2Ȃ0��CӨ?i��Z���M��&*:.h4�nt�U�z�Q�z#N�|6;T�r����^ÍNN���Gx��l���Q���"O�6B����O�4�*Ms#��yH�h��x*.>��[��M���+N%�ku�t�dP�ŬZ�҄�H0t�L�E�U;��S%��W��į�
�۵S�ԡI����ޓ���cl��3gV�֏�����`euu����U��VUkݴ덶��J���
��[?ض���TaY�REvK5H��\޶
�wgӅ�æ֑��T҆e�&��t84=h���p×��3�xg,<�VeІu�ŋ���'��M=o"�����ӄr!��h������ɚ���\��YGA?�2G� ks}}:o"8��T������*L&�y�i��%��d��T����d�sl�kW���<[�����h:_�l���/��&�uG0��|�rD�wek���U^Md�����]��?8:$�Jp��yD�R�0�`�2�A�&	����Լ,�I��p�3q8;ɢ	��O�HD�}�w���Q{����r�l1�vJ��m�cu+��E�e���R��pW��L��<|�������UPT��P&��%,T��Oa$���͵�鱴B������n�,�R�y��jOЅǓ�����٢�J�x{�a���VM;�����6i$#�q<�$���nBH�bksC$ntS��-Ƞ�h��.�8�F��24Mf���C�b�&Ľ��"Dfg�y�a��m����"�U��b!�*��z��g6���y��w� e�W������޹wwR�O�*>»��D���m!�Lx2C0'��t�wZi��:R�^�;�h:'���(V��E�ĳ餟u���vҶ*O��'�~���6�G�vwG�;eʳHno 8/(?�5��=�no<j�i��˸�Ǐ���A "q�5[c`�a�M�D�m��,�ZI�ko����LGT�=�O%�o�_�$,������1u^.���Tiwg&��d�����Ɖ�o�moz\�� "N{�EUa��爤J�5�:Mf��p 	�������:{��O;Yϵ�}h�τZA���㰋�M�l6X���
ȶnj��La��'�P��q�m1�V�Y~����#��8cЫ�3���dc��5��[d�����:+�1����$�Haŭ�5�������Ç?�����۷o[�D��d=��";=0�瑒�Yڌu�h�&�֮Sۗ�Y�-={�_G:��%���O�Iue	��U�p�����&�G@^�Z8"���h؅���N�!R(���:�sqjp���H�VW�<h��!
����t��I����)��f���F���E����#鎄�R21s�b+`�at]ǲ�;�$24����9��h����E�/`zi6�b�;��=(tz$vԸ��1��,�:I�!NL�	��.r���Z�4"���k'�Ӥ+5'�v�WvVu�lH�m��Ҵ�%�>�n�3c��\(��������!�Q0\}��Gy>�q��>	��l��1Z"��2u��ىɠ��S��<XƧ�q����`�_����C�����gϞ�A�^�����c�|�ρ�p�ۖ�g��"Cr5�+*��Q�H�D	|9�T�J�������g�JN�t�
rt;P�У*Ҩ͒dW�I��Bi�AӉ���pܼy��իX"��/���]'q	�N'v���_@JRE��)%O:-������g�YUs
A�$9��6��i�o�2�a�-q�+�P���NC~�kZ"b++W�\B(ux|����ņ�u��*� D��.j0*Q8I\���XhN؈b�~� ,�l�p2m>�F1���F}���q�'��t��(��`��E���R���!���be�H��6+���!\]Sk�\�gu�Q[J$���:U!*�x6�N���ZQ��������x�������o�I�����R�g�P�
�!Ĺ�����A��Be]��-��\����>��G��j�]�A~1�r��������1l����4R�D�'f"P��h��<�G��o�qq�L��ޒYn��M������{7o�8sf���T�.$���I�Y��G�-�:����2��.�X�J�@���huMPB����bq�������d`�'P����!����S�ӄ�"i����E^�B�m	o���NR&M8*+�P�v&ki� �4�A�19A����U����%�`qi�ٴ���/t���M�	�>6뛛d��Va���
-�Z7��������:u����7���pg�,�^��܃~��;�7n�@	�����QkhjBjt`���
��S)-�S٪_�0*#�J	փ7�)
�e�-�6�'�\��i?Q�ը�-�wmIB,5�(�2a�m��KDc� j�xcl"R/�PBl8N�'4R
=W��믿Q����+��K���b�Ǽ�s\�/���]��޾r�,4�gw��W�����L�j5k|�ʵ4�!���0!��"�����F�-��7�D!¿/'-���UH"m㇫a�pa�,v��@3N�<�a37�|�F�Ǘy���?�.熜&��g�i���*2�A)vt���T}���|Q�v��c�S:n��Q34+n�C���YT���⌯�z3�����I�e�{���>�Y[��fN�R�L�������c(݈=����uU��N��q�:˦&�Q�ÆXB^Yd/�<\�hǻw�~��G�d������!
�r��&��ed�x���c\W��v]��"D��a{�N�Y�R\���:]΢�+�����|r���8�.\�����.]��D� G�Sgq-M`ω�1˵GC�K1�pz����D��tj���D�Ƅo������=�9UWC�5HI8d�4�[�t�S_y��0}��g;/^����PO����=�	\dI������d����G��#m@6
)����^�V{��S��4���4��k�t]p�u��G�4+.?w��[o��W>��|#��΋]��	�3�j{{r���,�{- �b��۫t�<`H��l���I|ɚ%�L�G��4W�c	��J=|�ǵ\_���$�{]�Z��+�(�8���X�l �2�+�3�	�a*�.\����=��H�D\:�حV(���FF��Hl$aR�t�OF���R�I���ph���Q!!ͣG��z��Q���T��]�G��1ɎM$] ���Fƹ��ʭ?��?��������!Ϻ8�����x݋��i��О�b�+!D<R���`j��ľ.1��GOh���$�Jx^*9T�k:��AMXgn2��*�6JͶ���Gh	�q��'�Ů���/��]�u�Q��*�{c��+��M��u�S���M�2��j����R�i�)�1��G��ֳ�]y^�ir�<wVՖ������dh����&��hѢ�P��d�D`�ڍ�b����
Ob>���H��	4�n�O�%�1"����[N,�l_Uj�� Cm�o<sf��7擣�a|B#����g�Pb�D��QHz-�ñL��Ίu����H�Y#���Cr>\���Ї�X�	eѫm��*�q��gY�M�3�[֚�&�wμ�T��V�26�ɹ#E�@�0E�_�����ՕMY�* ��zڻۗg��*VL`���Ԃ =s���A(�qӫb�yG�ZN�4u�[�pe�m��F�Ǯ�Nv�;�ǖ�����,�������h(��'',>qwxk��G�7��"��)�e(�DO��"���/��/����b7���5<��P��͎ǚ0K�u�YE�x��ؔ_���ϟ�5qN$U��t<)^�{���FbrD��� ��X+�.<n+q3@[�y$V4
[�����c�2�_��
�Б��r��t�8�������d����M�10~t�lUfv��mR��[eH�2v�{�`5���W�׏���a�:��:�9S�,	sf���b�,KUp)�꺑$�B��S�\�F�ڵ���<���)����v�3���p�G7F2�5\9N�إÉ�P�!N�7�+:ΝgsU�Q9�Q$��_��_�}��_'*
���7�����Om\'S�z�x�T&ˈ>ߝ�Z|��#�W�����W�������}�}Q����{���$q��%��D$5�����Jx�/ل�|�١u�A��L�����Ó��KeX��I�`����:s�㝫���8e�B�<7���դ���_,����9h����"�3	���Z��\Y�b��R�>�20�i�r��r(��%2+PLwВ�Qn��s�X��v~#7�ǧ��S���n�,زc��؍��ˊ�j�P��p �o)U�����=W�M�+�6j��=��a��%��rۅx�G2���M��r�Р��B�J���k�w�["��7+>�j�1����菠�(G�������0���P3�n WңdXH���_���]�r���&��6��	�tȡr;�.svU
��#j�,�������]��|2�	cc)�� �S�Ů���ALb�L��o][4��)���a$nt����`>>8"1b��O��2Y� #j��7w�'�*8���ڇ�o��\�4ؔn���]��!���9�r���B�f���֍�5�3�E���o���h�e�����r�OV��<����x�t��X�&��������u�En'G���ƈ�w��xٚ8nm�n��	������u��-s;��b� �'�D�++F��N��qEU�A�s��w{R�	��_���k~�ag��w��1q��\2҉�Y�)@m�eu���w�����/j\�\�˗/�|��nQ�\�����ƴe�s�����88���?�V],����)��¸��/�K���[>����K_���PR�Z��Q,��2�QC��
\D�8ܟ5�/�۪<Ͳ�G�U$%�"��L�܆�aԖʢ���$׍�%��*]f�R�\���CIG�2��bz��=�B���m��FO�d�����MIPa�`d"���\0ޠ'eJ�����b��K�oZ{�ؠe6W���V��N�ӤG`kY���@ț�9�M-�;¤.בhѸx�
�_]]˲"Ua2��gh[�S�b�kx�ζ��}	��l�5��k�b&�����1�T��z����;�#�ɲ�� e���`i�6Hn�qy�>��GeeI��*\����)M��'�$���������QNwq��\ٯ��ץ�G��^��0Q�~�~ ^����KW���|/�<y�1�D��q���T���%�n�`����D�,������$}F4�t�DtO��^S`�*������ɮ�j$AI��B�>��͵�/"*�����#��u��·�5X�~�*�T�Ҳ��=��A�D��ߠ����f�u?|��-6I�M)���Y���o,&la�/Z��K� ���C����p�kŨ�h�7I����e=�bQܿ� �%��Ek�艕��ݽ��	�����jşi-S�`]�Ӥ�SV#����걽�V��|A�g!>?�<x��P�f�o��
����G���43(������d�<�b�uv���6:����Gt��v���n>|��2��XDG� ����ܘu��]�����e��(M	����uS�"GQ,t�v�[*6����G#�wk8����+%�j��~�p^��A��9a�O;�ݻw��_<z�agg�ٳg�����hδI����>�o�׌�c7��7jl�AN��Q�W����W�\_���i�Z1��:q2���v���B�g�~��Ϟ=׊�P|�C.��Ry��݆Gn����z3)�INM��m;ҡ?�yNCi�lܾ}[A(����C����b�6\��ZG#-0m�ϱ�`Ëkk6�U�	ё�t�ي�7��m��S'p4꼸q��ښL�{��n#%ܓ����M4bxq�{"dd��x#e�W��ԃ7�z)8��')Ց��f.@uB�->O5N��ɞ �:��!�T'S{��cd�>r������gE�|�ý�=3q�(;8�L��:��A�:�̫B³4�����ݳ[p�w�v�=���^s2�����;w���9?؛�����/�� �b�(��,U/Du�Ev4��W	ݯ_?�f�#A�����a1a% �;�-��V+`[1�=����3uBY;"�P��Ϝ9�@nww�,�b�X2ٹ�/b¥u�~*H�~"ǳLu���0\���QL?��I»����~��/��/��6]��O�@�ٮƵ��n,�O��t3���b�c�2��7�x��4ū� ��a����o��HB��6�mg�4'��v�4�����^���2�י�cZ��ص��:?֟n��կ~uu4�z�2\Ry��7��dJ�V!�q�L�:��n8^G|9�2۱�!����21,g�C.���hqe���i�Ҹ�}����\�!G��X��}x)�1vr�3Of�Y���zA�?� �`<8n�R��U�%�д��)�z��^���w����_����{��ޭ[�����>��?9·�>��jev�=]��+X%N��6*=�,�s 	I�Ű�}��TprRx,���D�q�`����2/N���1۴����v6�g�&"�ż�O?����^�?y��ŋm�����RQ��v�1Wٙ�*�2iZ�;?S��J���s|�FC��z�S���q|�5\�O��\G�xT;v��3v�O|�(I">���o�z}��ĵU`i���\~i�5�m�U��$L�k\}�i�P .�k�l��;�|�O*�y$���{�2�5$fEG�
�K.�Z��:���<yp��tm�Z ���0�Nd\i����~q�v��D�=�~���o7����|:�
��>���˗^p�;��*Uw��i2"7�����/��@{��_A� &�[�ظ�*�����,��
��N��gb"���t���]@noos<;�b�$�h1�-�o�8fq"4�$�+��B���n��b�W�Eև��L��EM�Y9f0��CB2n@h[Iq���_
��x�����������?��(�ݑ��H�zd�x���=���t�!�L�ʰ�3!��:�l�S�@�s�m��~�����cx��^J}���>���|����I�8�GB*C=���H���Z
|���:�NG&�@��i
I�%�Wy�Q� M�'h��l�u��2bB��Ӌ�HE�U��&��Ъp�犦��Z��"ܺ��|2U�)Kk��z��X]_7u	9t@NCALh�'�L[��Ri�,!��dW��.t�k��Ci]-��pt�CG���u|���N(��Z.;3di@zPoY>]�}B�
����	���KH����8-���\ǩ���ΜH��}�������'�[W���E�h	?i�8A)o�R��,���Ǝ(�u���]vY�|��Y�A���_��tHs������
��8��.��	��g���˟���	u&��f~I�)� ���26nF�~�t��H���+Gu\6e�X6��O=�#':ߓ��4��^o�.!"�wѻ�|gr}�0�)TUdI�4ʷ�W�>�}��(�|���ʌ%�Щ�[�Y��Ξ=F�"~s�,��:�2��Zr�����nH1O�w5���T|��@������m���nq�[ZbF2|@�拓��2=YG���FDo1��jO�t)W]���������o}*Μ��="L	<4N�I.�/Y�#$N�H�G��i�;V��4uպ9�&��>@µK�.�q:q$Q�˦1��삀�$�Aؿv��UR�ܿ���{|?�%�g�Б�W�5R�-�N��'��3�2g.�������JFֻ�T�ݛ�����l+�k2�s���ZBJ.����I�e��{{�9�֮���<ҡ�0ֶ���^'%˃�^U�9c�yVX����<�P;�������{[�O�5K�4�$eE���7�<�~6��A��Oݓ�A���|�Ei��F�ԥ!bs3Є���$��7�s��O>�a��WiGP���!���RV�T�*u:R��"��YT�Ri�a���Lm�")b!۝(9}v4�aa&�䶰�q'�ڞ�� mx����X��,�������۟��񾌸�#A�a���o����_��׾�������|�����:��)�v#��b�K��v���0z�g���Cn9}��ѕ?����]ؗ���?��!��y��������gd��Ou&r����N@s��D���%�����X"�b.�y=z��C�$�d.���yE��J���i�#Q�4�J\U!���Ջ�]M��]�al��hd��ݸq�O��O�4���=�{\7F��pkk�ɓ'�O�I�M0��g3A"pD��Z
X6�N��L��q8;8\'vS��B΀j����ɣ�L|o vr��1M�T���&��{���v' "m��;!n.Q�(�z���i�'Ǉp�+�T�ח�{�Fx�fH��(y_*�X�oZT�^�ڀٺj���p|"Y:>�ɋ����/r�R��6"��c�gA	���R_d���)̕c�����T��<�<udS��}���%S�ay�P�C"yz����A\��N�#�kn0%�J���iħ�A��8�E��bN��dƍ�U��8�[7��g�g��C�$Y<�7��Y�T��d�_��)t�h5B�����q���D�bI7�i}�j��YlO{\�[p�$�ʎϲ)�q���e��l��?�1t�+�ؘ�(���-�@E���ب���5���SF�J�G��]��A���eC�'�8��:*�Ѝ���]���A%�ZE*�����F���۔f�A�$h���ŕ��i�Gac<���]����>0;�Pcm&�.ŀ۷�����>�_��?{���2x�G?���ܚ��P�P�<T�	\�d�['��`��[��w3���ן4��h?9����ьr�q�����,@E ���C��f�����������|Eٲ1��jW=�S�Ѣm
v5��|E�j���&�GL�,��J��$��ߙ����G}��8���QR�h�5�.E�?��b��b�ß儠�!*j0M���ŭΏ"nCRB2�A5@����#e�Ჶ�0סp3O���1��_�f��"Y�����M|���|*�����w��^6+ձ-e-Q�'�}�FfTq�ɂ
�A|7����9�#�r��t�c7��{��M�Ʒ|��߇F�@��?���*v�@I�BG}��e�\�Y�`��@�Ox6|	i��+��B�@���O���lR �h����Hf<�W�a��Zд�!(Pk,��9�R��-�V�9<�*��Hx0D�f\�-Y^�����O�Iǔ���v���6��ŋjd9�S
��p �w�����F2���F"_X[�iI���U�ˋ��
�4[����"��V.n%ƅ��;�+�L:;�?Z;&��L���z:�;0wC�|YH����=7�Gfum@�\�X��q3�kE6q��G��T{Y�'5��p,����X'n��Onȝۜ����U��b"�X!���qc��tV�>jrP�)���dS��b]�i�����d{����AL-�6�)]�~���SO���5���̩��bכ�x��w$�L�N]k8��:r�vL�J��a�-7�q�8r��Ò�7�Û�^�629�c�?�spuC�I&
�f��t��qE�kA���Op�<�
殣>Tb�H���4�</{6>Y|�Y�
�j���R�ڲ�7�Mdl&Q��R*py���j�~��(ס��^��NoİqOl˶�0��m��D9{�����jhY�Z�D"6��>%�պ�q�A�iҤV5�Y������i(�q�6�����XT-b�,�"i�H;�`4����Doi����::<����FĻ�����q����h�6�a��%��d���I�/#�C|T�J�^j����kiJD�����,ȝ(��r���Z�a���2N���ur�t�u��OA4�a�r�Θ��F�R���,�=؟-���Zhjx�L�y�Ν;++kb�������W�M2����{�ڌ�>�BW�X�؍�7�蚑v`(8�޵���Hg���P�DGI*��H�����wA�T֑�M����*�ܻ�|w�	��٭Ps���P�VJċ����E�^Xt���X�~g3x�v�n�{��[���-�A�I_hU#L�/��eurx���C���?�S/ğm��IN~(�x<�L���9#�m<��i���b6���+"��/�@�$���4F�H��1�F�E ���@���!�A]�z�=V���D�L�c��N��'9�L�I(!���yZ�𰱏�Y�Xg 	:w�>�|$���~��`0�{���)Q�'�L�е�)�p��Ν{��������h��P�x,�]�5*(Ņ�ہZY�x5^���ɂ1�^��-r�4)�O�����V��I�%�מ9�K��Hv�x��s�_�~tr��������|>�3�>{�|2C�]�~���*&�q=�kO�����E/��4��6�4V�kU3�^8G�6nH�ln��KJ�dss��`cqa�9��ǳ�,�^�vO�w�W��~��w 5�or*q7�ʹMYe=H���e-��9n�͊z}z���4�c4����9���o&o
��ee+�6�8���B�N�ʰQ(�r�̙��3�\��䚕n!q7��j�v� ��؟��t�d�}�r�΀�7E�J=r.>�K
�߂���N�m�bI�L��٩(eU���I��)�֢j�<���������֖�]~��H�¦2�����>B���uh��T�Q��gy'�tV�?�w!`(2�5W/����ߕ)I�@\\*%�a��l�|���&��/����M���'��Z��⎆�xX�NUk�C��v�vݴ��r���ϞE, 4`֡�f}��Ã#U��n6ɹ[�q��#zG�#���-+֧T�L:�25�X=���t ���sݼTZ[fi���2�2M��B���?� �c��w�Y����5��gG�vx��X|{u�P��ҴGZ�H1>|F<|K_�G3���#)KG��S�3)E�[*t=׌r˥ye|"�dI�Au�:Zm�V��չ!�xF8�Վ�/�tݾ}[�7�����41���8��k����8�I�t��EvV{�s�òN�� 
�����q!թ��Dn�癞�w����Q��2X�����ْ����Гg��;|�|8�?��q��_�7�a@�8��te�����}�qP�����v�� U��>
�vgڍ�:H� �`���SD&�7����7�À�����J8��Ա���TW,� �F����{&��l��'�&�V|d>�P��`ׂ�I�kb�g�Y䣷��j�܂���G����`t��w~pp�o��9�"��vp ��8E��.�S=���L]I��e��Z�C�D�5i)K����ع�Fk�/UW�1��BG:��C�<vC&���f	������m
 �[hA�P�LOiN+�*
����Ul��Ǻ�Ҥnd��$�$�B�n~��C�@=5/H'�2��ȩ����ï�%H(�S�5��v��>:>�?8Lt�N�v��0�NU���6 �}�f[�Iɰ��ϊ�|���zgϞ�ƣ\Y,���m�<[�������wE�Ê�'�c�p�ej\�:�M�^����_��͛7�ӡV��B�E�\U<H<ޱ�Z���Q�5�i�$��A�/f��vvv�t��aZ�'U!���}u��������y���+X�ΝGP�2�e�˝���I�H�
h�\�P7��'�W�&@� �X{"PV��	����Y���S�d�g��w^�Ca��٩�J�Q�P�܅ �@�M����C���J!�]�瘟�/�N)p�)/�2-:����DʲLs!��f	�!�\��>�O+[�v98�����}�X8��K�0�h�EՖMDh���7��=�cx��&�.�{�քM����ђv��bӗ��񵟆h� ���
��h* ��v	[8���Y*����A���Ze��u!�S9�����>����"0>��3-V��-��.\�%!@��$��N }wo�	u�ް���‣t|纓Dq�����ѡ��D#ᡤ�NQ����m�s��EH�$�QYU�\��Ml&�:�S7�W#
��A;���	��M�0KM�ܕ��=p9~2�%�s3,Ϡ/_G+g\���#��}6ե7@˴\�y���@ڨ�3��BG�K=�������]N���G����#��he�����d�D2��C�!r}�eu����R;�%�ԃi}}2�mO�J�M�REv��e������w���tV�
:s�'�-���\U�~��`P�&��޿s�M#�lQ�Q��������d:?H|_NIK;i���FR(aߨ4�K%���e�#dtcd�X�l�|j	NXt
mG�q)��u�Bj�F>�-��؉�3k�ԯ�I�%c� 3�x��~�8�R����������6�w��8�U�4�ʊ���/�o��¦�.*=s͹���s��X��fm0	�W�Tvr���0��k[�B�D'����ё�.^����h0���|����>��R����!��m�� �9t	+��@���t�f�`�Og�-{���t�����F��2D�τ���dUqK8�����o���:EWs��֭[�H+V�*�5�gb]�l8�J
۸F���$n+���<zt�J�1�Kf������8&G_��4��7�O�q�q��`��5�����XB"\)�Iy?��p���3x�i�ڄ��Ϟ={fu�ɓ'=��"�"�|DP:~qƘ��ի{�2����)��6�U>����N+jkN���Pf͔���Td�Q*�(�&Bl��+W��T�6H1���j˂�@{����n����>|�ȼ ��ģ�x��ϟon��!H� ��:��T�%�[��r�H}�c(�}M�"oA��D������5,��aQgeE�b<�#n�N��Ɂ R_�u,2������m;Z+�L����A�]b'�b�-��W
�59m��ńE���6ޛ���S�����ق��싁�lT�A4ro)I�l�ٵ��Ү^���o�Ҏ���O~���#�2�z��y�V,Iz���J7�Wuo�v� (LV�.u|�.e�D:t��*�{���d*qq�҅w�y�����w�������?4푦3l���w@�VCb%U��+'/޾}~#N#�=�Wx��彽�Ǐp`��jǒ�m��G�1Đ�������/�_���C��j�߲&�U�����ăD�����H �M䠦��@Q�aѐ@M�CeS�2=IRҶ�KkXW���p�}����Gt��94�ܲ�7���a��>%�q��<S[��t�ߨ��Lg�m�X�k׮�8a��-78�+3�����=��G�c"�S���4�<�����s� ���2��c��?&V8�7�{�����(6�^V���J�+��S�L*���2M~?���d�N�����˗�VF�!�ˬ�[[�o�L�Ruz*N��5]�˨��(܅�c� �U��;N�#ղ�B.Sf�k��$]}}.y|���gU�P!Q<{4Fab���QyrYb7�������Ij�j�l�2�ӂ��(����޷�z��a��O�S6Nz�d�h����*K�8��/sR���g����@A��N�D�νK��O&�nm��#��BS��V#�x��â���۽�@5�H�@ۺ]��k�qz���̍#R�ݓ�"N����S�������;�HI�L��8p�ǵ�Xz�ĵ��0S�Pd<�M6�>��{C��W����B'D�8��*聁�E�,���L�5וk8UV�H�����YJ6y@%foΨ-�1�;-kf_���9V��&������+�FV泏?�w���3]��\��H  G�3�����"Z��H]X�m��{�ڏp`r�q�cא�����+_|��`�H����x���Lb�0@��gs���^k��UX�z�b[ �al���"V���JV������N��j��t��H�k2�4�t�}�k�k�l�M��E��pb+�S��B%N&�T�z{�������NQڮuN�M�@�!��
H�c�(�TX�6V�lҒE�x��񞣣LmwK_Ko���yI*�P69�d]ʡ=�����@��ҫ�l.�j�rl�?�{D2ryC��iZ@� �,/�AQt�Y���yo��c��:8Ec{�5�"��� �ˊ��:�M����Ox�7Z��t��n�j�~�Z�JbȚ$d��XȽ����ū�O>�2x��� ���ǉ*k���.��F�;�+֞�V���S��d�ZS�x�E�R�E�����|<Ӽ�0��(p?8��҄l���+4�S����v��=�+��`�>�]l8�@�5�.K��o���1H\�Zk�e#������`i��?FGer�9����͗��+��.���ҹ2���Оܫ`[i"����u|4�v��ї)Ɖ��ӘhI,�7�r��(��T�����KLJW�ڜ[���3'	�ah���
۬��S��x��N �ݔ;��S�c����pum0����ĜLŮ�|Q̭��Dui�_���^A4���Am���ΛA��,��'�Ǉ��4���^��HF8�
�U�E��G�J�aդzx��(�M�ꈀ/�s��щ���~���@s�N����C@�N�+�����A)*��	|�OTUU�ʘ���R�n�뻥h�gG��ɪtA���oDѧ�|��������߹s�wx���:]��Yܫ�j�;Ԥ��y�����E�\�����]kG��o��&q���w�l��Hi�ʋ���3
��9'��0K:��1�+���+��p�?�6#<��kc>����!�|u׷��k^�~�Y��tr�#I��#��}�O=��8�q���;bE��h��1`;����UP58{E>g����m�v�r��ͷ���7��`<�F��G>>9Ԟ�$S�:��E�P�k��P�B����?�	��S@�w:��Z���.��+��|9�ɲ�]��  ��IDAT�/��Jr��DE����{��rM���-�[��������+�.��[�w���GQ�����wvWV6����돊�`��L:�	�ي�D{�ȱ%�R�OV���1��t��ĸ�]��Td3N:a�� =k�A��]�f�p�4��p�N��z������܅������{��ͯ@Y���)B=�BIe�ŉLX���d)+2yvJ�hqU�;��2XH�*C�R��j+9�^,j�gڱ�y4����FVru�� ��j Xv;�����pgơ�M��aɒ�g�_�xY=���ֹ�����<��B�dI��5x�l�]	����	��qK#��Y;��S*�P��4�.`j�ѓ�$�)R��yQJn�6�(R�c� Gc����w�.!�J;uc��D���q��k��Y:��~��=}yp��ݕ$J�/�I�|{�@]g��@)�ڂ���m</C��8��9Fs�rڻ#F�"�F��Օx8Q{��X�8ͪkS���vhD*o޼���~;lͥK�._>_�ʍX/�k�s{q��� kdsCax@c��A�;�}�	����{��?�]�vM�m������O�n��F�G΋"��@6���?���E8����z�^}��s��pt�X�3�D�m�~�o�&�����5`<*� FI�f�HQN�6����w��C��g�+I��M��H�tJ��d�E���d��}j��^N��0@aS�x�ckf����2%Go�)���\ U1������d��8�|B��ո����?�91#LG��Kh��Yk4���:V�w�7�G���@�䆡�07�ݕ'�>)���L�u�Lޕn�����5]�[�(G���P��V��z�IR�G�ƭ��!\YʐƢ˅/u��Q6��1$��!wV� {Q��^--Ү�UB&ii����L�����w�P2Dz2IG���I��:Z;�Ď3+mʸH�1#v�����(3��(߱B�VA+M���m�8��=�Ԩ_����pp�y_u�,j��W�Q���=?}��������կ~����/��_���'O|���Ԓ�rJ��!B����n�Ư\�t��Yf҅�ke����x�j�Τ:`1��� R�0;&�e=���E
����N|���ƍ7[ě��[i�{��O���n���]��xX��2k=�Cی����C��p`��{�h�#[�#=�i>o���ݜh/����m�?
�n֡���gRcO(WR��#T�f<��g�ʶ)CJ���������z7�|t$f揝��$9{��!Vv�LU־��?��t���v��v �Ȍ�X����ӏ��,���Օ���5Iռ�燁X�p��>X[q�,>���L��ܾ���/nCٚ���/�����#���1Y�k���%
����ͫ$T�r�L�T\���5���~d^��?�����=�N\��=�t�ݻw������_R/b�E}���ڏNe����xb��ۍ�`71ܤnO5B��*�KB���V�V�o�o�(nj#o��3Ir�S����'W|I�l-�,=K���ɱ裣�=���A��G�V,�.��L�Ѡ�\[��$��O&u#�<iO����K���*>���d8�x?v>�6�Պ��ºs�濔>����EQz��I���R���8�
IhfQF�-�2T�lNC���5� p�Xg�f�":�o�E���2��
k=-m�})���Bl*��!��2���wV��4�*;yl�Zp�&�/%ݻ���i*(�v��$���n)�m�)����g<8	��tf��9�o�80�lig�>9��D�aI����΋m	N��������?_'��.�u�{K�}3�ƚ��jSk���t�� -lr���ӿ��lY�"���h���@r�0&��_F�!�C��V\�A�Q�L�3���Kw`�'��Y�S�$$���u�-4��M5nf.Ř�J��8e��o�H�v��)q�����mx_D4]h|}�ul��w���W�x�w��=�K�b>5��̿������4����\%���
��ᕸ�>9�4�9��E4�b,eZK�����n؛*�����c�����^E��{��u���e*Y��DE��[]�x&�{Z�X�8�xt+����6(���f	��S�0 �����ҍ����j�!������x%�
$D��=��V\����9z�v��-_@`H�C�E���`�����N���J΄Wg��P�i��z���2ݻw��Y(�Q!:�Vl�?	�M|N�}Ҏj�J6���L��:�����|�M�Q�6��TZ`�Q���Lv��y�h�i�.�@�䫯��1�x<S�C(��W^���(�ǦĢ:��Ē9"��a�Bm.�v἞6�x�i\���$�K�F�X&A��4,��6cYؼ���;��\���h��t�W�d���/\� _
��X�G�~����'¬4U�<��hFtyP�~�V��o��(|@6
	+b,!JX-G�����'�d�fY20 ΅��I���?hs:svdՅ�cMno�A��ج����)x��F�I@.��i\NH��&M���B� *
�w��m�C�q���B zZ�l�0�ݯ$u"H�W���aa�hI?lW��g6�;���ZV�$�7�p��ի�n����7n��裏���I��N�5Ux�/FCf.�D�QE@ҜL��gQ'UѶ�*��<�<��B�"ĘB�J3��zDku��Bh����Ǐ	�a+�9t�n�/_�t�;�>�胧O���ˌ�8� X|����AQ����&[���*Ϗ�(�)�V�KIEK��i}���j��5�K*S��Lj	�-��A��jx*��+��更;�έ[���Tkw!Yh�.]z��aOÉ���N�Ok+2b��Kxw-�q�8DE����L��X[Zg��L �g�-f��% ��X$ o�����}������S$]~���^�2�t��o��v�Dh6hM����~������>�	;>��h(��c%��������>������?؇%��/DUJ��.8ϑ����E�㗕�z޴h�������>�W��Np��y��?����*P�T��25�/��M;aC��3U!��5�B�N�D���%�>2�B��5�(��]i�<�F� DW��d5�}ėr
!/K�H@����gc�w1�M,�rɍ�[{hR]Ggț���5n^j�PC��Ds\�Y+�+�3��3h��8�KȠ��4�ϻ�na�t�X�m�[ԓ/�f ����ѿ�j����b�)���O����W���[uc:}Qq��p<��}�VAg��B��M��Ae��gǒ/�&� ���}��eNA 0��I���v��q�kBG��|��q�X��%r��<	�r�w�w�>�Z�ʕ+D�����=L�--�?�|���ir#҈/Z__�-�|�]N���^]SAхV����Y�\t���K�{w�%ٖql(Sؒ��,c)�Y/%}��?�����N,�>��7$q��8i����^{O�i]������T��j��U0_�KR.(�\�7�]�!+���;�L�qH7<��Ŕb"C����[�>$��\�s����x��G�?����Sz՟�Z0��+��+C�;��h�����勥�ֶ�D�T�,Bp�p������}g2�/��Gq��&^�9Þ� c��O~�Jk�gΜ�5����Z��:��8�h���p��+(rq|���Z��<	8�?�я�E�f�S�U_�9$������4�Q�`^�l7<�ˠ���В�D[�̔� �tI9����8bYz8�����p4���B<R����1C�]x�4�a�\��.���ꅓ�5�,�݅2�Q6)
~5U-	A&`xZh#�I�Dv��V�q6�/�~Գ0&d��$����`�l1�&Q ����|4کұ�R~��b�7�/I��(�����DK8'��Q��4�R7=�9
o,l�Ä>_d\��l��[�#&���o�qw���^�v�H�f��˗`({*Ґaj��*�爖�B�H�⪵��w���W����?���z�+�w�d)A�'�]��y9�f��t�w�U\�'NqLBB�,�,{��w[�"���Ԝ�)Z ��l]�vP6��|>aϣ#��fXW��du�0v_L��r�Oِ�1���N�H�k4�,T���O�g��M�9s��y�+MY!���f�S��%�B�CV�j�dj7��أ���8��_l��'�䳵.�|�>e�k�H�]�	
�lZ��Ϸ��a����q1�_E��@�u����oQX�x詏��ZmZ4n���$�@��I�F������t�l֑x�i%5��������d*I�7a����3㩌sCsa)u؆�kZi^n���WO�*Ϻ��M*Ci�ʰ�h[mj�,!�m�],sl�4���*W�R3}��pv�X��D��7VRz�EM�O��_"Z�G<�`��g�x�B���'����̥-;*��(V5��n?OK�،WU���C������I7���(����Z1���1\ �J���`q2Q2� >���W�С��6�8�� d�%eR[���2�v���ho��'1�T%�jA�hjZ�2׵��z~���l�b�\�5;a�u%mA�ٕ��ų��n]�p�2��MQe�D �Yosc��-8���B��&�͜}�k��x�X���J�b����B֋|��NR؊3A�����R�2D���t�Z%�2���H0۝t�?�LϞ=[4'���<S��߭ͳ+#�[h�6�7��
�� +��qC�1�;�~G{C�JB��D&<9��O(N���3��TF�1�ƴm�c�Zn�a��
} �O�ҡ�l��_�v���DZ�jk(,�x��6�zq�7��eӦ[g/��������~�O�n���[�	�@W�:&XLgp��4����yjJE��9m�X(#�LVs/��*I!"%!Ǣ��(���Sc���.;�체��i�J���%������ņ6�o�����ׯ?�u]Z��tI>[YېYm��'�v91TfK5SN���"+�=���X����k�5p��!j�߼ߦV,+�	L ����P��po�3�ťH�Rg?
� ~SG2���W^{�7}��G����]�`G�:�OaRM%'Zn���N��h5�a�l�^��fs,���E�ȋ?��t�{�y������O��d�3���3ꪮB=$iqᢐ��i�/-у�3&M��~�;�=������3��� |��l��fw:=a��F�ٍȂI���mq:�Rda_g��,W�&�c��m�#<���32Hg_�a�g��dr����bg������[� �SƦ>����	��ż�M�˗/�Wd�_xe4�*��b�>��~}0���~�ua���Ǐ=Һ}�8�����P�/�8�WuW�)���h����xz|2����������O$ȇ���X��g�U���l>��!��i}��s$�(����ܽ+-���\��Y/99�j�>��R'�I�j,�|LА��8�z��[�,��5����7���;N8f���ݣ�ۍ��B�J�ʧ�+�tv���D�W��;r�l�#d���+�nvS�H�|O�M��c����ʂ����Ô3�SC����߸aw���᪶�O��/1��	��"e�M�#~�
� T��G��Ͼ�������������h*�srr�|���<~gO� �Cvݍ�3�&��9TL���|i���r�Eކ��jU�p�m��o���9�w�u���х��X�5(�����K��Ai�@q�ŷ�Gh�p]�|8�+���� ��j�a%�q���>�NWo,F� �$2��h3ra��lƭdM�����y���g?������?��?��_��װ������w�q�O~�$H���ӇO���[W�\y�R8�����_}>�i�/!KJ���9+�lΉv�*�!���Ǆ�(s=���[�u~kms�p$<�+k7��8t�`��d�밲���6�Wϝ���=�~���~��_���?��7��Z�MT��t1�1 [��A?�Y��ՀO4�,j��"܅��-��g6� "Fv>��-/[[*[�>:8��%��ϒ8\̪8��/S����������#��1�����gx�}Ƨ�̂qI�N��R�s˸׺q�\�&�lNd" �M/�f:˯�V/_{A��l�lu��PD�~oT�w�=x��bJolnJ�C�5����jc�.�ˑs�=��M�e��������R�/5�q��J�$��*�P������w��ꫯRi�=���OX���4�ws��^7�@+1�D��4<H����p�)�L�6�K[���Gn"p���'}x����Wߕ~���|A�̶:LR�Ę�@$-���ncyNH�s|<�߅�!���ci_:�p<�~�Ɔph��l�誟)��t>Ͻ�QC�EX$�q�ѐ����	�ٔ�u�U�y��(�l�-�G"�Z�I��^$��_��di���'�EZ7��H�&��*m5�'St�FmA�E��m�����Ы�6�d�l8���P��VBY��A��c��{7�uOfp'D�L,�(�6ȰHzF�m�:aX�m�Zj��-ޗK"���Ӻ�zB��e���H��r�jن���F�j|G�r啲͐���B�8�&�X9K��r�߽s��rw�ŋ�����n�x���흝xv��7�Io!nm���z�xΪV�F��������:%N-Έ�_"<e�;���d[Y�ʑ:E�����
|٨�#���Y��Q�j�m<ڍ��ƃ��R١r�rk��̸v��/t�{|��︱������s�|���$�ܰ�`	��3�~���������tȉ��`i�V�4#�]B�����q���Yf4/��>	�����0eNe�Ik&���YBe�N�-DZ�L��#ݽ�u�аG3J��ڟ�ȡ�D?�K�;�
� 1V��t$1gz�"[2Ue:��01��C�M�⿙�Ù����z��q����^M�]י����������@�P4���G=����#:�w��w�"�!ƴ�Ҍ�C�� ��@<
�}UVڛ�?�Z��;���0��y��������2Q>|&����u�fZ���Y��	B���T5g��,B,�T���cq�C�x�+�=|
>Q�E�͆�+�j��\��l:s�ȳ���(�T�T,���g�b	�g��k�'�cJ��*Ān
S��+���V�+s�3�2
��z�j��`�R�IR���~ ҕ�ī��Jo[&˂s���wI�#��M�(4�ތ�q�	4S�%��&P4���I!���Iq�)9�ipM
������1�
ӛ�hĂ#Cv�Gx�7�=���qC�^qv�:�6S�a7���!�ޮ�fR۟��tAHv	H�35�S���?S�s��4!`F�=����.#=j'W!���s"�Kq�͌ �����3ޤ��#��?y�qE#W����XW�`�΅� ?αcrF�����L���AP�ҙ�s4J!�����*7]C��6����|A�5��z��Ꟁn��5�r������~%s�4?��"H�$ӱ��!�*1��
f��u�R�	���P8����!M��RJI!��Bm��k��2T����),��Jk��_e��:B�4j�֯7�"9��*�����	�������-��ޖO,����ޕ�`�S\��s�&S�p�b�&ua�yZR��p�6�A0�
4�EqP�n��o3lR��n���$pea�������ΩS�
�/Eu��M"�J����bŊv$4������j��w����dj��Zn{"�\h��et��f�S�"%Yj-�]�/��BO�[�����"�/�x���V[�w��|�ҥ�?�q��j$L� r�u�]�&�`H�vQ� �&a�pðG��0iL�g��+I�����Rz��.4Z���?�>��3�(W�^��H����XY�m7�B㸆�/ȸ�1�'�T$Y�q�ț�[x
r3��&�U`\g+ʕ�*�����/�N&cf</y	78�_���{��)ߋ� ��尩7�k�&��4�����6�����n'}rQ1E��4��Y��00K���L��L�(?����aZ�19�Rq�s����n�6�N�HO�vj��*��a���n=�ͼ������՞?K�5���^������#m�r�fXjSvr���!��av;�A�kx����L��E�&�5�Ja��kwn6�EN�ڏB����!�H;
��~q��щ�"�5l�"�T�I���nGO�d�Ȁ��[�H�ٟ�n�{��މ�'�����{���������tMN�
�1SF�ʹٌΝ;��������+�|�ѿ����3KZ�0����3Œ�r�m4�y^�
�d�r�>8�#��E�9敘�H�̼_g�c˶��!�w�,PW��D� *Ks�Ҁ���d��4�<��ݯ'���(��6|���8���G�f�lafZZ��ֽ����$����DL���?�Vf'��a�Xs�k"Å�A}���΋��H��Va�K�L�X,+��s}���A���C�Vd�F�� ^�����C���c4��n��ãa���Ei�su�ԤU6�e!?�㈰�lh��s�:#�,N���˷�w�G?�^p��e��"�@�5M�y�`jEm�����,�F���9[m��`muW��;�
D����a���嗗WV	�aE��r8֣Edom�4̏s�Ȯ�GR\)���l��|=|�Pf�eҤl�ĥR,��wPr�֢��<e����,vm�	f�U�5�`*��g�U�^�77ՀG��]h[8���D�����SЗ����/6V��&�t���6��b���uu����^��=��+J8^T�tuz{Qߒ<uU���0?:s��^U�b	K[�D(�O�It�Pq�QV��]��f�}�G�@���я�����[�ˬ=��xϵ�/dtH^~��-29&��M����\�8u�%P\Z���{�QDP����4��x?�3]�К4�(�'.�.`5ǻ�9l�����(� 2~����n����9�e�0��bj��$���K�b$Lx~�l
8*U�G����a��%Y,@*üJ[�$��s�*\_���w�3/i�\b�o���A�7��j��:@�i)�_�u��\�)؇�Ң��K���bGX�����=���*��C��k�J�dɟ?l�y2�M�w�=x�&N�|,��Bql��_,d��/�lZ�I�`�`ӳ�p&��N�Y(��t�?�{��Y�׉�&3�3\S]C�E�~<�"����'O0�"�	<�wp�zED�(�1��,��]����z�@����Z�ǵ]/O��A��/IF������:uj����jo0v��j
�r2�s�[7>!�t�����ݐ��G}�E1����Kа��(�ƤRN�"��ԅ�%h�.�ޱ��0��y:����.^�2�#�����ؤE>�NX�s�ߑ��%3(���S�5��rM1�G���DZ��@�n}^H�c�+���6ih'o��tg%��a^"~�*�$ִX�s)&�d���?}�^�� *nN���]��t@�8VJ�B�*�f�"߹�O�C��A����_c�k����}]ɺ�jX"�s���Sq����Y^t�W7Ui�T؄�u���13�LN�I����s|eJJ��J�%�=?KRȩƂ��bg:�2��4Zm榧)�{�s�E`x&D�{�����p\2*��T�u0�[�N��J��b��L�qe\�߷/��z�g31$:��&���R3���*T������=r�R��g��������޾�8y̎�����-M�cHuM&�0�Yc���T42�W��2�ױ�h=�j���K<~��W���\!�*ʺ�$�͖±(nS+�)���,�±�T�J���<mv�'N���}G�AԈ{K�N/�ɝe��&o"$,Sh*��ҀT��p[J/Aw�ә�Me�LU.��\~y=CS��Ld{ggO�W����c�7��Q"�lvw�����-x�D�3e��Uf�񕶏YzVAL��G+�OR̂X��x��26+�̰�����V�0�DBC�f�/�����۰$V�bv͸Nl����2q	�w�=[[[sa�GG���:����F� ;_?r���B�Rj![���_��_�{?p2�_� 2U<
�����p���3�;�w#�6;���Q�uLbZ��JOTD�gt�����1���P�+2����h���z��u�m���9��$��;(��gOݻ�L���M�Z|��q��t�6���j�@��W^_][�����:B���ɳ����#W�G[z��U�'juZ2c[Æ�H^�
7O9�Q��h2�LSE���2Z�6��+�@�(��q�L�u��� ���v��\poo���]��+�瘭��NN��m?�G��;ծ���}�i���n��~`��霠O���+�:�
�EU��p��U��n�1�t���Bm�,�jT�le����ר6]�z�%�:��0�S�0�+K�T�C�Fd�#�f�l�¾-��oȡ�ҳ��h�^٦6lM�u2��.�'�#;7STL����m��1-��ɘ.�d�5z���O6�P�s���+W�p\,"�~�����ǜ�3��-���xf�y�.�?��Ò�M3��g&yM�{fn��l6!U�f�bnLQh>W�)P�U�G7��vU�T��#YP�L�L�DnJ���6�m��s��ԕ���WW�������i�����w�%+�$F`"X���{�G�E�����k׮}��_�3��K/��z���u!
dpV������k����ϟ?��_�|Q;
]]���c���lҝ��陹.�f���9��A�Θ�2i�\���<tt��C��x#y�$)��m �f�]�:�΍%)E��x\��nA=�/c�Go�	9�����j��R�~���3�
��q.�T%g]���lL^͑{z��m=Y�:RW/�kbw6���n��W6�|���'Z}�	?{��K��*�9��T� ��1b���i��qwt_�=�%AdQ�� 3M|��M�@��z�nR��_'�`��B	���lDS��p������lt���t�Oue"���?h>�YJ"-�ݕ�#���++�z1�?����nI�Ј�n��l�������//llk7�^��7�T镙�k��!L�������@��*C[D������s�Xb��n�;�x�{�K`����{���c�i�0��Ϳ�ס7NBvR�ϧԙG�p��M\g���h D�o������aga��E��m��(=֐
3��f����Q%t7dX�l|ݾu�ĊJ\)#�I���p��I�D�ْ,�������V��9��-��I�Zm�h��(�=�e.�3%�������#D5+��N<�y��� ���v!d��vZ�D�j�N(!����̬�}���f:�u��\�F͕)�/��4��+�!hU�T�3>��CH$��̓�n�D��pP)}'N��)Os&Z��OOaSJIK��*��$��hZ_�8�zt���$[���f��	vK��S�0G}�RI�z�!ֽؕ\!u��_j9v�sjQ����9��7_�?5}��n5�f�;�������1o��7����=�c���ZmeND`S��a��8I�d^�'O�w$��l:d�A������4?��V��ά"�/u)�/� -����������;�aQ�͔���8sêW�Me �ѤW�U���F�Tw���R�5(�L�������FVs�=g�ſڵ*Թ4(�bei�vALP��Gf+-�֝��������j��e.oe��#���/�J���@�����"��\-���8������S���"����}��d���C�?~\�4;]h@\�������߿��W��w���� ���q:�B��;y(�6����O�~�嗿��/�;&ZU:}���q��I���/?�%�
�Y��(Nr����V��<�2�)6\3d�SQ����������^<��A��a��R�+��<$⮹���x��ʹcjz�YafL��.P3���s���I�H�Ce
5�C��Xɱ��1�t渊:���8i�l5a�`T�7�'��ݻw/^��ztC�WMS(�-��e}�$rlV["�uU�F��f2�UzD./���.zM<l��Ҡeɨ���M.]��+߫����	��#V�!X[�\�2aV�����!Dӂ����J,E�A,3h�7�uN����$��O���gi�y̢�|�]�e��L��� R�Vs�8��M�z�]):5f�E�#-sey����;ju�7U�]�,�~ �R3��W��kJ5��T�0D�9���묓�5��e/�9�SJ)�)�n��t/-IĒ�q�4��� �����r��MrܥdB�#�&�	!�b��	�D%c�.\�<?aY�pd5r/Mm\����+iQ*ϧW0�8U�kj��z�dʍ%JR���F�3�U�C���R����=�b��$t<N�V��9�����Y	HD������vVP�h���:LmL�3c�����v��ш�������Ո%i2gR*����O)���m�bq�%��i�/�r��hw�֭[�!��u�]P���P^�9n%]����\���Ll��h�@������W���M�'���h�fl1�'�N�S�@�'��w��~�������*�AR�]�,N�"\�������7p��>��LclG�lM!Ur?��֯@�<䎑��|�EP72
���2���X��&UTJWrQi���!E�;��ʙ0O�j��)ET��7m���<�-��~?]OQ$��p̜t�������M=O��",�������B�v-LC1��D�L����/2v��%.����9lFۊtexf�.�y�����d�0�3�)�A8���7���/M��^�rb��id��_ �����Mc`��f�i���3�G�9��^]�9?4�1LnI0~�-�WUXp("?x��ƍ[p�f�$^m��r��`��ƶ:�~���Y�����M���k�a�
���ژ��9V�쒖�)'W��0n�&�F��ZzM�a[�8%m�xp8��)���t.�d
�ڒ��n����T���|���w3��o����t������Y�,�2������W�b�!�0��N+�B���>��\cfuDC��8��!biP�I'BV_�Md`����S#���IO�#�=�$�UAr�� ��.c�����+++o��~�s�	>��:�sRYQ�.����MY��?H�r`��o�>R�����:��1y}>���鼚��_U�K���&j@h Q���p0�r���������#ň��P�����t|�uRJ�����h�p�1�_�@�
R3�ѐ䅻+C<6�D�E�;��g�������k2�*�A�o�a�Ɠ�|�k�[�U��s��t�`�j< o� [G����=���$]S���2�����w��+Ϟ=�&� �5�-���¹u�4�lV]Ȼv�6��ʥ��j�㹋�\*_)mg�wA�ّ#Gx��o�LQ)\��,2�N�Au��_�v-Ҝc��[�5j$'D�Lwa�ĘZet�H�9ֱ���7n0����9�%ym|�����L�Ϛȃ
��^�$���VL#�hB�O���B#�yF3�S[������!/
kn�Y�t��Z�I��7h�ڵ����2�ӚS���,�%"k t����S)`�5�As���66�W�ï�x����>�V��Z{Tsx�������4NQ��#�,�:�Vn�rm
�\���n&J��k��L�YM��'y��]�I,���u��� �����J�u��a�F��@��j ���L���,Gd�x^&������tR����q��T��4�cB���Iֹ��f��N�Z��'�O-�*%klRv�oA\�d�F�,�%*�:�#�m>���$���zQ��T9���B`�ӺzA$�ʢ��7�����&�S�r�Z�ګs*����4Ri=��ޕÍ1�B�,5Qnh�2�A�)K�C�B�ɩ3)���o��b*�TY��n�8<�*�@�t!Cq�Y
	.(���s��&�(��Mk�?K��wX`��mX�d�_�2�jp0*J1�r���_�*��SɅ5"�Q[8��P�a���kw���*XC�rZ�w�+�-D�k+�R�	�$=y� �Iڥ[��t�$M��	�&NBS�s���tgg{8��n��]��Ka���_���>����M�x�zf�!�Q���,��g������wBZW)��U�M�v����k(���+���CѢP�Ֆ�@�/�,+�h1�*�M��2V\'69�8�%2mC?�.��擧��8�*4�ܴ{k_�5�6�M����Ҭ#E���^NO�B��a���8��t�I���5��ٕ�^�f:y���o��]��|1`!K���s��*�te�����,r�D�a�	'�b<C&-��\6Щ˒��U\.��i���QHٖ���.�h<L]���ե�oa��4�u:�n�u�1=zK\a��#� %�@J0��
��roa�;5[���m43C���b?�L���		�c;���Z����l?�O�a����I�&��\0�{��(ĕ���N5�]l�0�	�l�6;�;˫�!d�W+�R�+�K��݅n�I�E������9�ܕ$�D�5�N���y�݁�~�|��R��S2�?/sS�)�����OW��f�	}G�q��P�^�ܹSǏ�'�s�T�:A����$���#G�7���{Q0�M�v��ٳ�\2(nwW�̱V�?6W�p��bY}��N�����ܱ%��PaX/.7Q}��������Apr�h���9~���cx:��V��hkznW�"���/1�5�V��Y�,T�#g>+�{2$�"�\a�{��a��S�\�T��]�L���v1�>gd�m�?��:g9Ԭ̂��υ�ʌSj�ջz��?��8?~�ꫯ¿���Y<�:�;��e�xB�2�Z�������V��2��"��`�H�$S�Ɖ�H�{M��� ʰ��©����)�X��hЊ~B�ٜ��v<�?� )`j$=�GF���z�9�I@������K����+�|�4[G�,u˯=�ګ��|���LV�*�%X�N��KՄ�3.�Y����⇭N�tک2�Gi���.a��Q%7�����]vJX��O��6MVV�M�2I�Q�N�������-��Pq�}*q{����YV��1,���A4�+�j
�}65cQ�����s�B&�5����o`5|ef�Ȑ1���!c��[��oݺu��%BH����J�Ɩ�5�MgR��t�0���1<+�����I.a�T���Q��3@�rM��n'�Q{t��1���E_?4,c�8������i񹆬�2ˏ_�S:ca��c��B{_�z��ŋ�f;�.���{;{��P#\�R�BE��p,�	ɞ*�2�(T�=���̂H�gЖ�)�����5	V�y5]Z���H��<HW�rI�0XL7�V�P�� �ǆ��R&�'�d�M����ҞB�qel����z ]h("���#�F���0'�Ny�Gl"������>�ٳg������G���?�[2��̤)���^}��NG��X�����'�߿���A�n^���.�{+++6�$}�����vvc3��NR�<��kA�
G�<~�"�q"��f�.�n�<>]V��;w��鳐�B[|%ߊ�(9NHK���^GR���n���:-��a�#ϸc��A���cfPd�HTNn����b;666�z,��<�Mbyyl�]]�]�#6�/�mf�)�̜ �åi��f�*�g-���ʄr�SCFj�v$٢U�͛i�HR{S��F��NQw�77�֖Ebg�p+C���H��8	��x4��������vT:����l�!=ll�l
DF!�X�3g����Q���K8̵`���&�챭�x`�b/ ELI(Vݪq֘}�>_�/��RP\��w�yG���.�C!��x�	˞\�'xA���).�m?q|CJ�R\D��.]�T&H�W/x���� 41�GHt���1�{��8��ׯ_z�E���pJ�D㾘���*���Ԇ�T�B	C����!ut��jx,>�I�#��_��PG20�w��V����$���}x�,�3�j���gQ&$�px�i�&rw�Y��R�nZ�M�L~�y�XQ��B�W�s�ޤ�ǡ�C�F�L�/3Q��X���^�^���jX��쬦)�zC6N��Ja�ө�� �1u����xy�.���PH���T��'lh�)�����T��dQe�x�Q��76���
���
ԝ#9�L�~�
]�mA�Ⱦ9�W��)l�*��A�/�(�(�Oxz��L�������3��;U�����ׁ4���i����$U#����j˂��n`�*�Y��ii~�x�g?��H���)��`q��!G��x6\��t>�n.K�u#�U|}i��0C߅�?j-Y/�0<���ξ��v	�`��:��Vt2(�r�����6�og8��#�c�������,i����\X=��5�]�g>���@(��qxоW��y�@��T�R���L/���u&_?%���.���4�W� |˧�\�{2�r@�
��:az��#�xA]޺���R�߶f%��\����̙3�{�
����J{�\l5��̻1Yx�<3� 
Y�$���4t�^�j-��ٙ����XЅ����1�8u�lҮ'y���Yz��{�ʕ������eR�1MCu����GDG��1�	�$;�nV*����:��ԙ�g��~���ռ	�"��Ν;k#��8v��(��)�Z��)��h����D/Q^�i("�x	�D�O�pM�4CoKCS�Q	V�uB�:�c�Y�o6��P��f���_��_y��S���9ٓ-k,���H�����,��NjMz��M��x�{�Ec�-�NmN|�t_[8�S�����@"m�u��Bf�If�&�"a��N�#?�N�^���˻;}�Q����������
@��3�^x�5c~.9rC�8��q�M�\A�]��pkVƑ4������z�|���4A����	PʨUJYV��ս��%J�����z!h|���O��g
័/
k�4d\2N�Nv�M[��X|�ʠ�
m`�uˬaf@´lV�Oth2����`�.�gZ����R���f�+͚��M�S�C]�>&<����7����6�X�IX�!4!����� �z%5Ձ�,AT��v,����-��Uk�7�8�h��2��Y5�`U���dD���<�J%�l�>�>sXXF�������߆���{����]��w��Е2ʏ��O���ž��Xj�� �M�с�)�g��h��F���{q1��y��b1�]U���3�ŋ�J���w��d4��{�٢����Fz����W�
W�t�2&���W9�����R����$0'N�8�k(C����(��U�@����i��5ѪC��a��s�Z�Ԫ(���t�)��&LӤN��#�<y"s����kV)�$�^��y�h�5I`e��&�^7�)WF�?y�2ii���vu���0#z��h
����j����,��ꝋZV���������bzt�
"$t��3T�L�^�t�` ��lgGT��%rAvY���eأ��U|"��{�?�)�������p_\3''7Ϳ�����!�K��աP����*�$6t�ih�֌���Í�x�;Zm<8�g�}��k��~��=B�K3�#��i��>����W08o6{t�9�M�I���¥�C�ܐc�r3[������m��E/.]��|3�7T�^ΐ�h��>�^/�c�Ts.��]��̒�;yK��u�JG���`�56_v���6' ��ǅ���iHCPwT�FM>��F2˥�y�~�j�S�,�`XF�4��s���[(Q<�P�$X��3�c��Q�X%���Q�xd�����!�ZZZ:}����w���H��wi�]�y�����_�n���`j����}����>��䡼�7^{�����χa�wݻwG_��ţ�o޼����v�,�!�F
T���r�<�
,�AY1�'9m�!��>؁(d�jЉ����'�M������d��$��-!�rB�D��T����XF�ǇK�;���5~�2�ۄri�<M�ឣ_D�v,��Ac�Xg���V���è�Ml��a�=ƒ2m�t���S��3fY�0�ߛ�i��q�3|�d�'ګ'��Чb�&K��"X�xe>�1p9~g��5L�Ťؔ�-���	�-�w戥E�*$����˻�~"�|�"��Ռؕ�F��Ǐu���	����sNBf]�KSc���fP{i ����
q��'���'����~��ۼ0w�2�oTŔ����'�&�J�"�}3���DR?��KK���ތ�g�&59���A���.e��w:i��ՙcY��X�Ҵ�Ո�Jb�����=FϞ=�I�4���Y`ZeO�<f�XP��O(\��Z�RZ�w���-��L:���χ��M��oMfc´933��2���ֹ�й���e���u���J��WZ��-��9]�x�Γq�9@�w��y��z�J٥��2-��@Y��f4�!e&�g�{�+��v�ݻwqR�o㛿�E�e����e����Φ��]�N�u�[���|!��Ǆ�BY��^��"B�LzR� �t���2*g�ݺq�F�;vloO�ZFÔ+8����ƑOt��aS?K���cO����\}9*���gO��_>��g!��6�JC���Li��v���Q](W/�L�>�k.0QI�NX2�y����3C���_�3�5�S���w����Ye��r���4��B'�fXS��95����a�OaMtM�Tn=Bh	�y���7�Xژ���R�Ճ�K/�f3�����<���t��!߄=H�^&�[��6͡�VO� o��NV�TB����1�3�w�kB'�D���x�H.`������:�|���Q�5,���¥9PWR����յ�u?qy=�Ep��tEQ���pfc]�lt�#�#5��FY,.u.�gEUu�lV೾'��I����$�d�	4��u"�G��a4HS��G%��w��svq
�{��'�|�h��Bw������q��*e��`ﭨ;5@q�NdkYY��.�l���c�8�����?��?E� +x�܅��]\
��T�Jt1�c����o���m!m�:¥0<�6&��N�6�����Zu,,�&�<�x2G�f��3Aҕ0�w��c���y� ja	·��v�ʥ���]<���v�����&��h�XIRdBq���n�M'�N����Pm���L4��+#,_U�D��ѻ�ő77�J@��>W�˚��iM�r��<��w��ݎ,p�LS�/\���p��O�����n}�!�{as�����~�M����'�b��f�)��Ë��f���t���tbxv{��+�\3��H��2������&��,H�[
�K�+'�=������|��G[���L�6kgw�������8!��̃2�����;����6v�yp�CxHK���p�t�K��x
[�9<�v�8�^�1�RЃ	,�0P�2��d0`��k�a+�Ԉ�8�Ϸ��;�xa��W_ݕP�u0:�v,;�`�bY��Y	�,��S'�ܻ{[:��$���C�ӷ?��$��c���!(��5fA�V�t���ZH�VPw�*s�_w��2�JN&�E�K�M��j�������36�3��8��3�(�gu�=J~�J����խ��z��YU�BG�d�C�
�b���J)��'EM�#%8�DTk����~�n���T(P4 �.d�q��QV��0ǝ���K/]}����>�����vdye}g�ѣ{�oy��Iaؙe�솿�vJkN��<5�*q��ҭ�|%�����Bm��}2�L�3��*���g=.Ib �1A�>z�(�J����8vjYP6�tǻ�����?�������`�eb7/\Y���i��pЗ�����s�jyqiks�;n2��Q8
�0�M E��V�Sgϰ�Ǒ�Umi��l��#$�i�[��[C4��S��J�rٔv;�|�LqtN�`0z�t���ڂ:�Xh��_������_�zt��}8}��G��;݆:�20�1�Re�ɘeu���vB[!�_�׊�c<8�6*��.� �
��&|�L5�3�6�-�(Lfv�������e�X���"!�_٘�	�G�`x�|��Y6�3�see�ԩS'O�_?��3�{��Ԇ{:��k�)��D:t�4:ڜ��#����9�Fl���)͊oh����r C?.?~��i�����ye����SM�ގY��8��u�}�%i#G^���v�
�i������=2X�s��B���J+tH�����0g�M��홙 ��K/��f�+%�=��P!U�Ԃ_��K8�,[��
,u;,�#�0�T'��y���Q�7�����/�N�>)�l���ou8�:�OA47e	7�����������_��B6���=}��端���o���˗Ϟ9�U�۷?���<����Φ�S�!r��:P��-�)���'�g����޳M(��.>��p��a��WpWwo�a���Z���V�$$t
؇�\�0�<p�!�C�ƆG���@۟:uF��]ɒ���a+%T��+W�?��4,)fŴ�ne���nn�P`��TyyN)<8�\k3D�)C��t�l���P�j������n�(��7�13�X�v��Q�^��R��_s�����K�.I�T<�~��2ۇ*��$,�b�
"��-��Y]�����6Y���e��8M�t'XM�pQ�"��IYi2>Lᦍ�:l�֖�^7��	�h3d���|��vX�2�����+md��~��湨H�4�I�Ґ���ϊ�pH#�UM���BE�߬C`�ǩ�?��c�rf�y�����2���@��_�jә��G��(�V�׭�������G���C�K��y�lł��&E�~�sͨ_�.j!���_|�O$��uB��&�^5&��SD9��7�����.[�N�ȒBS��2^_�d���jn6[3����]ث��2fDR:��6�T.�d��X�������P�U����-��a ��<	q ;Z��
� ���d���!a�N�l����DFL��Oi~.�`�!4dY���]&���I��1(���J� R�qpc?\>���g�wo{gkkk�?H2�~�ϰ�/��� ��*���{]5�Hz�*�bJ5p� 6�J!s��Z'�~��|V�|���97,+�SX&9fϑ�p��͎L�a�7i`1<���-�x2�2�vw���9���R�ӂ8	�^� 닸z29E���-/�G��O�A�TL�cyY�|����<[�P<ZZ>"r�N�`5�O�aB�b�����c]7������,�,�h�R���O��:�P�$��Js�iE��L����TUط�1m,pQ����6]2������L�*�)��L՗�
�5�A�3
3������I�~�u�m.��7Ԟ��i�m�Q�:�u����^�����u�S3v�E�B�θ��=�8y2�}��C5M�l����4ᄸ&�5𛽽�k���K1͠�yW��������u$"��m>��o2>�*��ͤ��f#�u�������k�i��Ӿ��F!}߮vX{2��;�'"x���S�3IW$9C�ÉD��Xb�8�Z}�)�U/4F�I�*��qX����S���@�N�IB{}�������{��*
��h��S����]9nUV��ѣ�ED�LO�����y��N�:����Dk���,��0d�tD\�tL��.f�+p�]3ьƒcX�����^{�\wA�E���{�w��fԖi�� ӊ(��܄"Z�-�D�����Ƹ�|��W�|r}���_O�;�OA
5���9ՒQ�-G}���L�k�S�C^�9>��F����8´��z��W����Q㘴o�Ν;x�S�O 2<ql���~�Ti�+;�"���-9�G��/E�!�d6��+�{x{4Im��g��Sehh37ʟ�̿JR�+G+��^e�hD�B�;��._�V��������)����MT���PW@�ੇ2���KR��z��j�deڗ;e�=�:�\Y�DG<�p�!�L��k!��k��Xf
'�*�2LX<_��HWt���^xA�#z���zw��R�Rm��%OY#�@"��hK��G�M5;T�Gu����g�W�h��T7N]�2��a�
O���!��7sJ7�	�l��d���͗�ϔݩۊa�5�]��\�6$[�&�鄣�p�|DPee��'�"*Ô�����A=�}������;�� ������U�LSU��6��쬜Y2��������f:�n=}tK�}�޽WVW׎��?��������Ǘ/	A�Q4�B�@q|���`�'�p����LD�c�lm�`޴�IHD䔱GN�*�.bgb�tC`�`G�1P�[=LY�e5���63~Oz`�L2�����:3�t�?��o}�O��O�Sp_�Y;~����zҔ���}Vns3�9���T
�]:lF�����~���סmG��D_��vI�K[���HH��G�>H��w�tp�%A|0L
# ��~���P5�(Vy����d�e�iK'#c��^�E�.�g��D�N�%~�q��,�3G�8�1JKD6��L��b	I�؝�{x��q�۷o�f�#���D;s}�={��Ei�U�U�֜�����}��G�֭[�����y'�Qba�f���Ur�����/!!TJx/����g�h��z��N?T���b�~�~�W^�e����o��.�����R����G$-�3��j/F���f��_�){�嗣@��L�weu'�����`����>zR̨�8f��MBz��Gi(q+3Q�2C�0,F��g\<3!�! 卵� ��jyy��$��E���1�e�ŤoI�93c:Ś��)�j"�����yj�n��h����[fm����ݻP�.\�̙3�#/�õ�7�|��ŋ�JP�z�+�>��ݞ;wN��4���
P�Ăh,�[R��e���!3,�h������x�����,����x`��}�����?0蠐0�'�k<qx��A�ܝ;��--��
�n҈31>u�O4v����q'UY&��6>r)�-c�h˽T2���R�e�[�=�|d��v�8a�r��R�9$hu*��I�O�/y(/�e��*te�0KK\����?Hoi )}b33�$�5� 7{�	�'Я�+��b�ĕ��O5�vFǕ>��$p�EʡPIV��b�N9��LB$c�T�*�[�o�>���֦��04}�
��i�d��E�¢��┆��U��PV�(fxL�2�>�,,��:�qe�m�����p3S��R�w��_�?@�-B��IЌ��3h�'����͋/]��Ҍ�P�iDM�T�)`D�b�h�#�!R�9֖4��	K������޺qS&��5�ܫ/II(��ׯcYN�>���<����X�:ҙ��-�����[b�	���,��fI��εD�h��$�`Ztu�V�e��J�]�l�����+/^-Te3�d@sA��Ë;K�By��QL(�<ap��(J���Y��c�+�f��J�a?o9&�	�S�(�L4m3���V���T˞)��_�_���8~��8��������"����?��������#�Ѵ͵��L��<�2��=p�h�_n� ~pX���X����G�LTn&���g�UF�v�l�a&�ڵk�(����'B��m0�ϫ]��5�i���1�T	grj�JuiHDZh�DR�P��TE�9�[eN�z��]��4:�B����L'hŷ9~l�[+Zu4QI����,-�t�I�V7��Q�B'�t,��d��f��㝽�����,;��M]S2FI���9s݄��g�fs�uQ��>y2�S�N��jsg��q�ֹm�q=�ӛ���0P,kz�j:�n���l�D>E��`��S�`��O'�!h,�4"��9��%�0�yl0�>�7�cK!>B��X��
��s�3�����D�ኾ������8.���1Sfx��0��� ��-u{8-�%�C�O���Ғ��M��A�{��:l�!��e��&� �B�¦�a1=wVL�Q]!�`����� �p���KĂ[�`���>+�ԧ��4���d�,UkK˽���//�bww���/?�/@�<�:���%	�ҋ�V܆�qO�$��aS������9V(_Gf+��*u��<�t���:M��F�rW���pƦ�N�O�>���p*�oui]��N�F-�m�)��V���tz�N�g�p0�Yɸ��VOvZ]�n��zK=	���*�+*g2	��`�����Nwm�*4���3g�����7z6kz���=�A��=��u[�=�e�6u�./
G���$����\B1��B�w����pk6u�m9���$�7Rdi[�
�+o!�3"y� GFR��#�P�OG�n��x��ZnK!'�R�;{��,}��z*�����{��ݹq��l2�l��+O�Rt�DVL�ӐC��5�&IЇ�3���VV�$��úG�p��&C^�(9��q�o�xg�+D���j�I�WU��`����2���/�	+�ZU��Y�c��~���lw{���˛7�z�XQ��Gz׾�ͽ����|)�<a��!|���ǣ��o6苳�Jl����]IR8l�H��?T�a�ɨ6��������l��~Cy[��h�xۑ��YfR��Oh�X ��Vi:��6֎
;������\�d2�˙�A�����a�������n��[c��FӽM_��������7��^����ASs��$�:����>��G�
��{��ʉ��v'�d�����k��QU@ =� 苮���׉�MI���+R+��� /�fY�	�����}���ً-/���O�/�����������L�����{���,I���)s:���,�����9)�z�Vw��i7��@b��������d��P!�4g9����ǃa���t4n�6!�ڲ᲋B��E�kI�鬄J//��]��o���X]Z��ޝ[����ʕ+'^���?���?O�z,��?�|����'O�Ԓ������}�Q� ��JQ��P��l��&_�
Ck,�����¨�fN�r�dogO*.+-���L���Sc�gZ���Ŋ±�,������`2=vl�,<��p;�"����S�v���[mG��`����;������nX!nԒ����n��A��h{�`�ͧ�N���!����B���`5-�����_,ua�׏�P۱�7���;�V�L����a�i7�
�l8���Ih/.��[) -�0 /f^(,�~{� &�2LFEZ��I3lM3'��x��o���ˏ>�|e}-,��'O�?y���~�U �]�t�7�rZ�����X�Ѹ��1�!C~&l��G��x���������t�<}�	���̄M���W�SW�EC(\�E�,Bx��B���i�=��Y]Y�X	�>�2�����6[�#�W�o�n6���^�@(Xer ����X������y:��Q��3��h�I����ĝMS*1��l��uPV��1�����l6Wf�M6s���L�Ope��ZMI��I��]<v���_~��[V�&��~a���璲��`�]0Adh�H��t�e�N���:�	��������l�Pr��T�-WR��R��+����[%�xu��T�1��վ�Xϔ�F�7ncA._�l-##UBV�|��(� ��h�ZJ�����A����w��8���t���;c��5�����,
��W>�!�W���/?��VƓM���v
�>�Q��T0�����#�^XͲ1b�$O���S���DG���rCzC��js|�BQVaC�MQF~�C�!�W��6����E�N$��/w!8x҃]��F#F�;Mq�F��I�Աߗ�Nw!&E�@]���??y�,�۞*�v�� X� d�2}�� �ƱT�����=���������'�Y[a��ŋϝ;�k���~2=�#'
�<�]�t	˵���95w�$�ƂC�����O��1��Z�������^W®��!����_@���e���p5~Z�5�� l)��Z�ok�J��A���ħh�I��h |>B��m	�k���>{���ç�p.��!�=	��bm}����ϟ?��W^���*��,�c&!!<]/���Y֙��R���	�ӄ!4��h(_��
�mű��+|FހJ1�6��(�H�s�UgyF��\�L8볆��:����p��(�*�rP���1�@Bg�DF)v��hvqn���n'�C��h�z�������y<3���"����:��3P�Z�B�U��c���	˘�����4z�p��.ͦ���<����&S&醃]xYR:��Qs=�����7t��o�`og28H�#ı����MCD_֌U<�߽̌{2,׆�p-bf��z���(��t�l�������"�^lߑ���gN���0�",��TP!�w�Yi�	��7�����:>E�q>VC>7�f�a�!��U��G�.//4Z�F��$1l�tB�g^��xG:���oJ��VHZV,{�a������o�A���+�Y"K%�)�⨅Xc����8���+�K��sp�`��2�����p��|�8z�T�z�[2�p7Z���$W�w��+a�[��3�Cq�⸋Z�9:��WXB9�/���q�WN8x��H�2�	�	���v��BZ� d�_��Ñ�� �ffF�o�J�	oW��P�@]A�č��2]���hqNĻ���7/�����4h�3�J�d0���>}
��Bh5�<�ݑ^W<���)�S���8�I�n�-Ij�ga�)\X��f6z��|����W��.��T�gڽ�\
�N��˙�t<�"Y�ȍ�/ޭ!h���	B�d���6�A1��bH�L>J��Y98���&���4���.�
k2g��/��]���K�v'l����ӭ/�FX�m���,yn��Hq_��-Q��!�f����:m/ᴡnqu~6T��@�f������z,��G �>�=�UM�g+n@^���K��J:a"uuV�f�I+�PEJ��n�p���ikK�N.P�I���9�+Kxn�ѫG[��j_Xa��l*��d�Z�y�J��uT\�ci��,IUf����	hY�`U����&�/o���>z�H1����H����z��%�F6�V��ö�P[��2��l4�(�����x����2��7F�_���X�ٮ���R���Eˤ�6LkPnzc-�47�[�/0���	.�3�Ē>y� g�G���Zk�~[���$�-��&���~���*��UlRS�,��-�\�v���y��>����Ba}�S#h}��F8�=q%�y�;.�%��yv}���	���?-*�9���Ň��o�f����_��_����B�������x}.V(%yi:�GS�X!�v�{�����1[kg�!�2:���u(`�^gsL�\Y�L�}�&�����(�^��_|Q�|��O��'�3�o޼���ä�(�7�ׇ
�ȕ��0�����0XÛϕ*QI�`� Ǝ�F֠��N\��,���"� �8QDw6�+/�}'���~����:���*4�����V"-��&��P��ln�~���,��$�:�ז��;��>&��d*��Q�><=����U�*��<���'T��}%����֢k��*=5�>.�ưS���m���+�����K޴vK���P�E�!>Z�}�\p��ή"C��n���r���y�۬�f,������:d����Fb�"
����ls��Ji�#��r˯=Q�j������S�BQ;}G����ϡa�"O���d���6��0IY�ab��E'�r����8��!�&%����P/Y�25�)�vj�����w$י��6����cǎ�9#�n���ׯ_��qO\���-.����-"�R��<y��駟.�m�#�GyT4м���YKh)[P�$HgO�DDVNu�7�jz�����H�|U��L�:)�k8�<�=\Wt9�H#�nP��G3��~�7>��h�._�#S���PQ,�Bfm��C,�#"I$�7b��,uI�fqF\����������8$��)�Srm�ү`���x�`(�x�X�>�"G ��.J��+g>�m�e���m={v��	/n�_�忬����O~��Z��������h�ླྀ=vz�j07!�f8�q�a�;���[&��T[t�Vc�u;$�$��6�hH/�m}Vv�E�5��DB�
���OW�|�W ME����[�b®��^1�
�'�4��$�y,�A�EJ�g��4cG^i�eġ��ѷ4���1�hD�Π��=0H�2}���:�4�t�,��[�Pbmhq�'��1G7n���~�5h��O@�t�i�����yǎ�_�
"�+�6\A�e�������G��?�������zI724T\��������,Z?\Plǚ��.��g����3@9�R�湚�B�)UΒ�ud��>����y�Y�i+�;�架�I*�s���jn*� �y]���S�3� ����`.E`8(\�X�q�æN|3�%4l?x�g���+J =�䵋��䄖��"�����~��_�	~�����s,~��,��,��,�jFPGb���?�)��w~�w��o\|�<��I�˹"9�,ẅK~��^�"�6a�&looן)5yM�"��u ��2��E�t�r��tDz5�z~� ���!�,f�֣�9jG�V��2�:�����w��]h潽�����?����&$D�D���Z!p��G�o�Pr������Pr�,>��lW����ۤY��[���'�iq�>2��m��:��n�ȑg;E8s�Z��������!��P^P�p�1#�sEZ���pT�!,%-�k?9ó�λ��V�E�׎�%��A�C=����rt�o�:��R50awK��1!0�z�Ӕ,:5��*.�ɗ���_JB��ř��1f�S�M>7�[�5�Q"����H��}�����lz�$@8��s�A�_x��$��c�y��+C �)�Ec�s�߿%�� ����O�A��3f�ٿ}�����4�ip��˝�P8Sg��JW��.�8�D��O��˝�'4�x��Q���g�;,��K��VE��K���5�Ӯ��+0�˔V�v��G"��]a	"���#|�NGz(�ww%����ZY�>�I�4�x2I���5�K����8�MAV���#æ��>���,�������賨���S�^m�������ӻ���	���_�#�uUp���R�mQz.t2�%����B�T����<J���]F�hl����Dpw�ݻ�海��v��4m|��<�֓�-�s������u@m��=��i����Nb�Oj�0,$�(e`�;�&�0Ҕ�h\8���ړĝ���P|T�(���))��j�L���#��>(�*1s'�a�Ũ��I���e�BjR�,	8�Fjا�b�
e�[�0��,�j4���%.�:'��H�9c�2~3|�f���Tp���t ���&�'�{�f��f8+=�L
��f襍i��y�V媍=AG�N#�+c���r�I��}H�@���ǬѨ��ܙ��$-:�"��,W N:ּ�z�ʌ)�A0�y�)K�~��l��l�l*���e����g�'�����"ie�jbyɼ&�z4MZ��0t{o_�t#�&�U'��JS~��z:��<R�-K::F�;*���T��P{�`��Vi�0J�5%I�hIG4��@�t69��Q��u݆'NO[�,d�/a$�.#Bv6�ZOQdݑzu)������*x��݈�S��B�?y�����v�?l��t&l,w�?<�2 ��p:K����ԛ���'�oL��������lD[ۻ������+/K���	���k�KO\!(��v�����f<ӆ�̲k�����8h��8?�<l�k'ĜL6����5�I���ȋf$<��T�����N[�j;j�ZI2T=$s��lg�֭-��t7�Ig������v�&�N�9,I`9>U���"f�f��%�g�	KK�H���+H�B&qD�8�8:�V��p/3X�чPY<\L�� ����ؑ��/���S��sP�2e2.3c�!�G�o?~����o��o �)��s���'�!B���F��֑V3��N�9����U�+�%g��$u�"r�-!DY���^7�/�9pO椉��%���={��_����.��(�\U=1���W��+�a��./tԁ_�>�@�������	&�]�|���W�zso���_\Og�q�?~XԐ"��1�����-�����DO)��P��r���):��ufyF��jq�8��M�y2Ϯ�#��2��`~��\\�D���?�x��}U�s!��!�Μ�����Ï��4W֜����󧏟�z�9��B��j��n�A��ѹbC������d�)�R�B�	���XX����e�s�.�+SP��0S�+h��llՑ����U�)z`2�B!���7ߩ�m����T�wK�
�t8�?�zz��'��������/~�3������5z�
,Ž���qָqƽ����8�f��m-.I���`�8qΠ�4��=6Qr� ���Ҍ�P�]��z=)/�p����mq*���0��+���ݻ���gΟwZ�Α�k_y"�������v�M����r�#/�DL�������F8Y�D�V��k��ˎ�D��K˔�Z� s�He��s��ɴf�9�P���|A�FA]���7 RY��פ��#Δ+#���*���'����������_��Kh��v�UP����ЩN���4i�I��d2�j�I��d���Zl�;q��tDW�
�*Eظ�.,t堹N����c%���t������ *M��W0���*�z��F����6B|t���0��FTT%�R��) 䐲2�*��q)12fCGk�;'x�����5�����(O���Gc��85�T5W�)6k��c	�"mk`�dl1����/ZO�q�k[����jP�O�~Ϸ7ۇ��M[!�є�S��M�c�D�n�C:���}�ᇁ��M<x`9"�9JV��ec�!���_�z�Hh����_����ַ�}�ݟ��>|D�z~��p���y5{�R�B�j'�B���S'"�ª��>8DH���u��p���Lӫ_��^-�����c�n.;*�J?SAIv�5�|ҙ�-��Љsf�V���p���"�I&e�M��l4��_��� ���K�T��
�2k	^�%�9�����2$�7�Q������/������<y�4�A,e��,^��� �E�]]^�Ͷ}�l�W��tڋo��+/�t�6���'?��������́�r0Og	,���2�s��4IF..�@�����-0�ص�������;�\\[[�7�1��<y[�����	U��ǟ7Z�O?�L��r�f!�HFL�W���}M
�Q+���#I�*�r�Mͩr����%��Z��Mb��},,!m�]^X��S*�Օ�%-�(d�	���O�m�wq��P��QK}��R�3�Ei�c?��ā'�6�^U�����y����_����4ܒ��n��G�y���13Ӝ�����b�_z(j�'�Ҝ���ꨋ��jo+6�?U�yz��Sp��Zǅl��Wϻg����O�:�/b_�Wd�Q�/����o��-�$7�݇,Lff^0����y��=�	l���ݏ Tl��-�k^�� �J�M�3�9���R�|�#�^�v��^��JQؠ3��T�?~�T�ÇT �(?{UN�
���ҿ�.�	E�����A,�M���R�:#���e)\E��E���y�yS���x����7m�캮���ce�(�0� �Iq�(Q"۴mwtGG�C��MG����O-�#Z!;d�-��)g��@����ʬ�x�^k�sN��p����w�=g�=��6n7�R��Ib����@U7�.-oJ���?���#lKN&���>���ݻ8,,�F��vO�cX�I�WZ�N�|g?㻪�2���=�b�瞽�w�߿��l������/_���>'[9��3���3'��k��*6U��+�a��Ҡ�S?m��F�V�H��W���;�{�a�[�j��f_JDӸa(��/�-$�+e.��~dķ�wPr2�-�DQe���K,~B�X�����`BEJɀ�*"93�5���}��$O�'�x�l��v���#1]Sx	�<7x����w.^:��r�
��$���[@H����X%�22��&�n~�;OsɃ�Xe�YVW��l"vL�&?	����`�<�_`IbaCO�{��T`i��l���ze2�RB:���M���U6�l�f�:�aA��-�ɠ�n�������9�O�r�d��cǝ �O��ٔ�����#e�ႆR��G�Y��yW�x�t�n��D��U"� �i�$(���G�jA���N�3O�l>4Gv[���\{��u3a5(֘�'Web��"V(�S ��	{��W�+K��M[��j0��(�Ȼ�Rc�Yu	�i����I�Y��e�xÅsa��9�:�0�qRe�zݹ�-Vfb���-?I���3�����v<�c��yP"!�.>V746�� �]+�s96�f6�U�?�����<"�F��r��u�1}�q�KG�FM���V��,�>f�
V�J�9�'b�Pw��{��������ϖh�8'��/����n�������W�:k��׮��lA���/�$�
١e!"~���fڼ�����Ri����DJ�����R�baeեM�ؘ�,��0��G?����ԑ�n{�a`8:���FmP�򬧙-L�&�Q;W�+�T�l(��,5����}CChpJ$�a��I�U�;���ҧ�C �E|-�������/��m0��ކ���'w`w���2^��6v�(��<-��k�V�Ku�t�@�6���L��e>��c�$�/_��W�����nݪ-����gԃ�j1�4̷� �P��R
�*,6�<��+Ý�?��?��Ɯ�l��%b0j@�~���%���6EQ+�-=���v�ɓʺ�=ٓ�	Ϙy�0���</�b��q�\-�@�S��r�<`9����5"~���}��_����=h��/������J�ƗW�)��w��˩��dO6��Bԕy��e�g�pc�w������IB"& s?�U�RX�IT�x��"��&lm���\~�N@�/V�������??w�Z�^A����/�MYι8X��ĊJߥQ�)�V)�'o��\�-�D[p�iw\��w�J��M���4�v��T>n��RKՇ#���Yz��[�|����O~�3��+�����~��_��}��ß�����+����v�*tv*\Ij�/���D�
C�oF7H-< �
���(3��h���0v:D����JRhF����N�&�2t�_k&��NH1K.2��\�s�^Ž?��?�l���?$����/T�2Jʔ�
�P���D���0,|��ԪJ?@�U��9�N'R੟�(�.R��	i6��ww�d8���lH䊷!�{*��:��=�)$����n��p�'��<�np��l��4��J���ǲ�PC��;�e���d 1p�6~榞(�F�>�0�P�o�P\x� ��))m?�E�$e��Ë�J�`%��z�	����/�A�J��v�S���v��:G*'��?Vѥ=� xQ��,`�fo���������!Q�3x÷���_����Xb$6��ʆ'*�3�S��S]���8�^��%�x�v���i�I0�u�,m��	L�u�p�*��$(����?�,��gw�gP��r�$Z�������g�Q�z�����O���W��*Rx�j'�3�;�y�'O8����lf�f��!���Mv΅���W���a�Y	؃������O��?�lnb�t���)m��R~x���6�n3��"r���Maf�ATN�������?��&������/�D2����đ�Y����"2��Ck���h�nl���o���k��K ]	[��}��ױz8���ׯ_�_�W��QK��Y�pM6�:�\���[7?��駷-jh%�O�������w�D�R'�Dod/rr��_�|7v�ƍ�>�L�,#�$R��y��v�x0��M����M]j~�J'�1s�^cѮ=̀��r"���]aL� #����ﵡ%9���UF:������m�<�`p��*��;�C�-�ꞅ$�N�'�$�S~��Ù�}���w� `����O��H��"��7�.��1������y�J��-�=�ʢ��X����7�8�f=�e9���_���:>3_^�� ��g�W�z�-�]8>YR|����w->�c@z��;w�@h����ad�Do�ա�ep��]#74��rr����x.�J�z��J��s䘍���o��B·�-A�(��%�+e�,��h=Y׹x�^ꈖpc^sB۰����[��Yr�cq�.V�}�6E�T`
�X��%��HAgoo���K/�Z?��Ք#2�ltq��?�D��k�E�P��V��<��;?o7�D;�ŋ��厶&�:H�xB���@N�Џl있 �|�ec��Y�P)���ژZ_Ã�M��{��c��|1�����5황�,2X���%��YB���e-�{p���g�\���[�w8���{;������#�~>~���2az^<��3l�tlEQ%�B�Z[�~��֤]ͅ��-)��A"g�dX��W�3!���������(:���4q��Z�?�� ���`�:]-۪d���Z�8J��Eɚ��8���ǹ&4A(�M�"�/KB���Ɉ�����0���P8���"��v���i��Ԝ	�l��k��b��:ҩ��/l*s���� ,A�.e�W�U}fjJ�b?G!U�M?�V����	k�3��[^\���Y�� �i:��`<n\�L���\�6i�Fp&}'��*-ll�/p7��w���*��`�"R���65���E�����i�CR��:�q��lk&��w��iR{�V5˴f��v��q<wn`Ve�(w�7q {���T�@��-U��B>=1]�񅣡䢟�n"w&��ER�����)�������_��N=:fSչ��+/<��_<�x���պ<:>)����Ǹs�3� p�������%�χ�/ǐ��m����Ʈ�~w�ӄ<x0ǋ�����������O�lm0��
~�������w:ˢ�oVDPjlf3���]lp��|�۴�8�B�s ����ҝ]������u��qA&�V�N\l�{�������J_�v|��~�;w?��7q0�F.��tchS�mݬ�b�=���ͩ���t� ��*���tVK���A�nnM��p���Ѵ�4������omLU�S2K����!�B�V��zl���a���"�A-B �]O����֯<~�W�{�����W.]�}'Mڸ�9�߸��*����l���D%�Y��%��t�Q�<���Fxcʹޤ�dCd�
�-����������_��gw�(�U;�����_�z5O��M�8�S���nR�6F�������K��>��?��oiw��xN��������lh��己1͢n5�A�Vd��4��f���6-�N�m_�]��Ԕ��
V`:a����Z�(<E��`ϒ�tr�ო�ѥKWp`qϷo}�u�'ބG��k_�I����~��~񋿇Ζ+u���{C��0J�!�Z0 �0�j���)����S�ஒH`(�kT
T� 	���J�\q�o.Qx8;���및�31�^/2�]�X�� gd6_%Y������_���ѥg��r���~����}<��"K�'��5m�^-���DO�����]�y��t����-��2�:���t2�B?lln2��dmW����o��"����A�4j�r��A�T���N��R�v���@$~�w?L���׾u�p0��������	wG�/N����=z�(�|��onN��l���0�C�BĖ���]��4:���Ш�f9� ���d����(�4$V�"dgw�O���E���Q�9��W��w�Z��lN.^���_�O�����?��ӏ?�p|���� �Ys�ବ�M�KÎ�U�̕�8�M�bAz��;��(�#I��NQx><�+��%��ll�	I�+0N�	w;������F�I�mD1BE��`UF�u�q#�W�l^�Z
%ұR4�t�k��0��-3�M�;���dg�?9��?�R�D5�[�x� +��S<H�g+�"m��!n�@t�*�*}�߂�W�s�PC�6��Ða�[��e�&WU�P)���(���P�ZeB���Y&ި��
�a��Bw	W�y!��4�\��,}��͟��gl�r�)Sz.�+�v�& �O���8>9ʌ�Բq�ven<�NLn�p��+Br$��>�>SU8�-Ѹ�XeB;�����nP6g>��aa��s>3(g�%� !9�2����]砝�� �T�/H�k)`�NqN 磑+�[tۭ!��z��k(I�e3K��P85�l���އ��@B�8����s���~�_@�~�K_
��u֒��j�r`�ϕyd��F��8j}���r<�ܽ�o���6{���)�g�}����'�'�G�P<�a���՜+uw^�e�'��pbՋXpr;)l_�go~���˗�^-�?����>;�M���ݻw����ѝ;��RPS���^�N>��Q�}�*����:ջ�*@bg?5i�l�)�f�r��9{��9fV��^׸7D�P��`���_`b����^��0��O��Ώ����/�������x��<�]��Ok n�=�@!�N�9:�.��ӝ�� ٖ/m~PW�!�
���u��#��D�v]
�����Yڃ�d&D�mm�,�H��;ws�|�o�#�]��L�<�.�3��� ��^o�\9uc�C&H�8�%���]�EV���W6ua6�l�8�bjε�2�/_��nnnb�O�����b�MQ�#�<�D���[��UqN�N�?��'�|�X��e��*�<9=91�`=?x�$�Be�P ��<��ׄ�P�7#4"B��sܠ�"��e(|P	#/�c#j�@Ǘ�m����\�� {�o �ӏoiA?~�?~��J��i?=>"W�������� ���C�$���������,��f�JlϚ�u/KG��<3h~������n.]:�Ȩe��2�$yA2�+��
�Y E�Y8$���*���Mȉ�(9|R�,��b��>��^���&c����.,T�|��>v)S��Ei#2�3B����t��qګ��rU�Z�gb���\M�
��t�;�Y^@f�o�����ɟ�E���^��U(��Qo�fq��.cf����q%ڴ��2�	��blJH*R�P$��to`7akI治=���U�y�ӓ�����t���_-���5bRR5",�OyF�uMψ[�4�M��Y����Iߺ�J�V~������Eۖ�I�:�!���VeU��!%V;�liuz�0�=r���)���Ʋ<����Q;����4�����OOk�/eJ\�o��c6�hF�y�Pp��hj;����ۄ��\���S�yIt��0;|gmc�vV�eء�Y�j��՛6��p��f�*
g���'ՔB'���=-H���8B�R�᯼骔�2^�~����L7#%.�p2$s�v6�7~�I����qh�Ԉ��MƊ���ܼ�%e�󳛵�(^�����~5n `�y�"��m5�2��_�s�ƶw2+a�Y��e�'7���{�>�(��2"�b�bx[�q�@sV�*=㜶1�7n}g�C��f��Y�*��7����_|1K�Ȧ�yT�dc��0>S���֦���T2(h[���)�D��ߗ�k�YcobGR�B��>;��K:"�BqX�t&1 ԨZH��sr�v��ga�g�J�*h�z�n`#A��=l׹���@8���Ejg�1!�����]}��Gx]^�)�It+Y�Lݵ�RhM�N��0+ʕ�g�W8p^a����?{��W����tneJ�#�!U�f�]�����ɞR������*��"�J,lv�^y�����_Wǋ���w��{~�!)�pZ#.�G���_ǃ�H��j>q���jt���pD�}���{+p�ƍ٣���D	$͚%�nfd_���GTJJ����DDY�7M��IM�|��Ԅ��g����t�whl�x�Q?�b�y�91���u<ѝ���f���?���.���/�?v���� �:�G!#�P03�$�&�	���v�#[��R&D66(?u��h\Y��8�CW�QHp��@t}Iz�a����O���$����,�_�EH��ѓ�^=*W��g����_�p����qSĞ�����f1�կ��f|	䤎s���zem��f�k~�񩫺Gc˨�SsHfu���ZG���b�*�)r��d��.;��^x!.�ۗ/���/�{ｷ�z��?��Gvu��� r�V�(�A�0���a(X�,��Z�Uj�x4NI_9��z%�ޘL��-k������J]�H��L����T%H�����~��_߹p�X���_��Ao���}���O�S`sϸ�~Pph4���sX���x��C\b����H%�2����4����x>֐�)W��C|-,�FdUw�t��}
X9��G'KH��[ӎ9�E����}�7����C{�X=�N4.���u�O����ƃ�~d�Z!��"�U`��]Q�"4�iNbv�\�E�1����?��������q���L��;A�+�(Z��!q����Qt���v����"��/����Ţ��]ƚ�"�9*9<�(r�LboSAO�8��{��z�;�^��o|C��%鷦Ap_�;�m��\�ʘ��惃S�5�=��
B��ݔ��'%n"?����QK�VGggD���PT�U�(�E���m|[��ZjG�<26	��j�q#���h5p��En���ez�17UB�R΍�$X�M��+����s�\��7&̅ _����7���|�_�h5Y��F 34�SV��j	�����6m����8�GH2Dh{{�[���׾�����P;��_��G���U'Ϊ��)���p�6a�>s�������}��+�����K`�%�X:��V�����;[es������RI���·H��R�G+J�J��8w�-rάemo��[�77�
8����k�࿩�^3�+�/��omg��#�8d�%s�p���2��ƃQ⌸	�vQ�	g��H�#r4�gPD�����5�3�y�Qhh�t]�l$�ަu���m�\�Ď���#���h(�[��ɩ�-f�К��6d��ث������YO�ux�׿�|*���(���g�=	��Sn�t3�@$gx:��� �(.�u�������h�lgr���R�
����c���?����<|�/�i�k�_Q��)"�Nx~C$�
�bn����S~[%��v횾Y9�G߹sG�>E�#�bҶ�ZY�ظn�sG؂ϊl����>'W�f+M$�x�;��G�<�u�c"E�ɢ���ˬ7�CTp���u���j�"c쭎O�{dǞUDt��T�N%�WS*��������z�iSQ?��!���l�0I�"��L���-e��1|�>��d�۰Arb�"�<J���1�;Y.y&�_Zc�6��Z�����"GQ���cg(0Xy�>��B�"j�*di�K�P5Q�}��i�O�z�O׺4��/�b������?��7���6��"����^Xc�"�e���_���v6u0y��֎��9?v�,u�_�K.$��B�ˋ2=�����Ocoe�B�B7���u��:��)��FI���Z��da�|���Z�U�$�ں��(��`�����U�d,W)���H���b�p�.��� #L!�1ǿƜvfU&,��-w��䋸�R��1G�Q�G�~���
P�3j���Qg͸,��i�6�5|�}��YK|��-;nY�QZ0
ZU3|0�ݤd����S���C�n��6ծ3F���d*�ѭ�����0�]�\v��f���Z�1vJ\�b��p+,��%�+K+��g8"eW���ä���H��Ud_)'�S����d�+V����5Eǰ<�-�6_��U۸��;er"����/g��W�{q�(�!uJ�'��B� �`�m�zt���?��??}��w����I��������۹x�瞃 ��������O��\�.۸C��6���[h�;בa1<#o��F���>�6��Z�k<�{�3�b��&#w����* �1bo������+$���� �����N���ɘVp�0U
'���i��o�E)EB&%D�ϔ�W͞�^e6:��ٜ+<�1�Y��U�*פ}Ax���Ʉ�<�=)G���-�+�R&�D6����½؞�*�R�dH��>��cG��ҍFp���u	�\����pq.h�Zߣڜ!a$b�����Q+��+�������aɺ&/�-NʓÇ���O=~�`ss���p7⿑9��YS�W(K3Wa�(��y*=�AH#D�!�5����L�5\AϴU` P*<!x��_���oon�l&ma�`(����ֵ+��Nkd�(�lL�J�1X'C���d���ݷ��9(mYZ�8����ȪaǓab9�l�Om1M�Vq�X�Q�~|_�`�V�i�Lg]yqH�pS4���<Q�8��8�s%UռI�z>ys��>�p����8�yooL������tQd���w?���o`�Ν�p��.�
Dn���_>���Xc1�J���1�,�#���:F������|q��͛�?\(Q}�N"<��\ n�_0װ�L�,6�2�-6l�y��*�o�bKh�2#�Q_�i�U�ry����y��?��u6���|���Y?��?�������NP�R����:�����8#�JY�a2��h�Q%$p��d�^on�ay�D�6�s�>�ڄ�Pi�t�Q(�N%K��NN��XnoB�G���D�"?��I��[�~��w���Do{:}��p�Ο��������c�����%]��"=�G	�QP��͍|0̊���i_۠!z���dEu�-v�WDУq�L��4�!ؐ����e�*Hc�����ژ=sl���Q����6�GG�������㗾�u؎(�����ۿ��|v�a�M�^�C���hNǽ��H���z��k��pķ/�?�f�(1Z�%Ԕ��]�Ucy�H�=hZ��ȥ���Ky�B�\d�n�ײ|��4���|A���V����.a7����{�=�պ�Z�[qb,T�R9G|ɍ7������㏃RuX�F��O���unʖ���~�G�ǩ"���]�CqfH�)�T�@i�܍�bE9ͿG%�B5g��������F��
���"s������y[_c.�E��c��\;�+��~�[�b�5�W«Z�գ����?�я��'���FF�ְ� ��R�b����a������}x�rEl�"����?�����ΫT2���ĵ�q��f�X	(A+|����K��S�A�ha�v뛂��T`�'>����4 ��p� | �P,�/�1�Xƾ�F{��\�a�(LA����*�ʤH�K�J\k²��n$Ex���rHq���!�c!���n���[o���!�8-�+Sq�Xj�$S�
�B���� ���IB�G�3x\�͛7���\��X.nN:=U�K���2��kk}�!�|�*��I�2���~��d:5��n6��T=�=}ײַ�x+�����V%�rp /^�<��Lې��>>�����F�J$�"G����|���K_��g�}���C���U�Ш���^W�e�k�
Vu{E��0Tb�b��m=�"�Ve�2��O�x�^�*}��_�Z�a��p�+��,�t8�i>�Å�Iu���<�h����b7X��EN�x��[����@2���,'�<+S�����J�(�k^t��!ː�8Z��P��[�0�A�"D{���g#zGY����Y&����%LtS.��zagA%쉆&I1���jvrbh��B3	yȳ{hN�.g3��'�⼻��Z4�O��3��t����T�8���=��O
��IbC�j��x�7��loo�o99�I�l(t`7�1�s�8!���m��w���ņ�̿�z̫��΢)�Q"X|͸����_��~��7��Ns�:�UOҞn�)>�a>b��bjy�^�
�%�W+&\|{kS<��ΒW^ye8���C9�MY��r�0�!yc]��Ew��h��	"�*��I�K�G��=fj8��_�x�b��i&[�����^���v�B�����E$�ag#O@o��Q8�!&�h�xIas�՛�7?S�sY������U�I$�C}�ҥ�\��8��{ ��㏆c�"�]!v�4�F�e�����DS��'�ǃaϦ ��A��~����|�+_ٝz���'���E{�A:+�V(MC���x�_��)��8vܙ��K/� �z�~���戔�GF<~|�����ѣ��>��#p2;f�~��*4|�f�M������e��H3��ͮ�'�g�]T�q�f6e~B��D�����_�/B۬L'-��p����9�V����q/����3<-�C!�!���q�宅L�>��*�(����$[�/��J�~<.�t�$��aE�׿q3qXʲFd� 1ܰ졍=��1������_+g_�L��F����n��t	X���heg�@��I��X�@�����-ۂC�a D�&BF؁�c`��%2X��7-] ?
��~�E�±g�Q���E*��PN�&��Z��7ƬN�r�Л�Z�|��ڣ^w}�.*��p&�l�pk�E]*mE�wI��w�y��������=�=ՔOQk�*���ګ��~�ʕހ�Lq��R����+xө��v�[+��,&��z3�8�u��7�O���Wb��{�	������	}��Ob-nз���3�Z��1:��v_�^U��3��=��u��'�����~�ǰ����ީ2+	%XW�����&�vx�{�ϓo�P~]H5�zd9UWfg�̱����L�`�;���4_�ODO@���\y��B��Q%Rh�:{=��4�VC���ssO�L��+Ϝ��̏4=����I.��S#�!�������Wk7�E��+RvO8����q��u��@ZDJ�����������۷�Ԉs���祊hJQ�@z�$�G2?9��ړ���&�:G*�P�qP��:�y�w�Νސ���ѻ��@���ʱ,�~*tH%�cE��7Z1<�T�Op|��;c���5��X�u�D@��<v�@���Y�o�Nf�m�l.y�b��Tui�͞*~x"-p��y�=T�����^��L|��U��pw��(ťkW��潏�b���<2�jnK�D��be̫�RG[>.1��u@d�2�l�E�f^$��[��������˜5�W������ǎ��Q^�=>b�7�w޿�@'��`[�_bua�y��\�=�	��'d|��-L�AH��nI�q�:L�F���
�����7��Em�F_�җ�)ēPSm���BYH8z��j�L;�_r#N�:���ځ�ֶ2�F�d�������ciT�.R��ƫ�R���Z,-5���p]�����8�~��w�}��/����.��o{��Hn�\+�gji7\�J��!�U�g��.G�VWS�����8Y�'�?�Y�PY�H�B���q�H�^]إ]l�������o�9>�+><<�y���ڪ�]�s�mR��ߺu+��GQ6�.x�%*��.dv���ծ����kˌf��l�Iܪk,D�R8R 6}��1�l�'����|'Md�1���E��B�3�ܻ"E�@�/����Ϧ�t�ҟ�IR'�;�g���bl��ؓd�;�>��ت�La!��w¾'���mM'����?��zzJ���
�z�7��l�N]R3�5�����r��)�̓����bG��V����O�\0	����Ƭ�A��vZ� ��<�m�b�~X��>ڤ������`J��Zh�n�q"2��Hx�{	ƚ���8��8�*m��C!q�x��_��(��S�J�`�G���K{{{7n�x��W�OxRq�?y���ei>҄��i(�Z�����O��8�0
_���7X)�XԹs��k*���$د�����D��_n�n�}���M���a������)����NM���<����I��%����S��!C�ƀ:�����bG�@��R�ݙN)yª@K��z���}&=&�+���ؠ��,t�xB�t:��/�&��X�;��sȈy��Ԣ�UGb+���F��$����w�E���N�I_��N�>���-��dm!��0�{!�� ��yN��m�|q*��u�ȑ�["R����}S�440�ŕ��$���NxS���_~����[��"��cZ��c7�>V�{�o0�z,$���v6�:�-{r⛬3yr>s�:�߽{�ڵk8�罽���q:,o8��%[w���j��g�}�ҕ������g>��n\˗�@ѓ�޷s��Z��(�������؁T\�Uw����в���Y� �O�*8w������:^x�7
,gAess��A�����?�\]��I��1��M����n
eE�%��[Ʃ:��b���g���7}P�x-Ȫ��F.�{WWC�-������lr qc�],#���
����I�g5S�/stw�4z���)����B9�Ǵh�}e���(U%����\S�����ĸi>�N��">Td1��!���4�  ˏ��H#Wg��5Oc�n�đD�"/G">\����(X�e��	�����K/@�_]�A+�!�5�+�j}�/_66���uK�۴�Y7L~;�%�g!��}�UY္f����}u���,�P��o��,���nb}� Aq8KuՖk�?��N[�)�qI\��|��*�Z�0,*�Y�R�||o�|:��*���W��#���g���v+��QhP��ݰI�K��iD-�U�Ơ�q��=5MB��-�n~nHS4Cv)c�m�4��"�h�M����-]\����@�&nk7&b��KfT��겟;�eE���))R�b,=[����@��9��豥cr��w�i��{�$�r���h»�))�4fG}���3�L��°�=�A�]C~,��T�o�{ɸ9{�+	�S�XJc*?B�1��۝����Х{8�}�jN��$�.C[�V/����\G9\`֋�ժ]��"1Z�A֫ڪ�!�p���z}xxr��Kx���㝝sM�����K�~�/��2�>���%��g������np��:*R��dqo�)"'<�!]G�e�vD�Jh�M`��b(�����U�z;�%��~T;��o�1B���a�TEW���mU�k�%�x:������.�U�ڨ\W���Z�xk�Kk�4�ى�5�kŖ&�,��N�`��W��N@I?��YڳBr���1:�T�]n{�<��r�HI�=�o��)��,-J���I��H
˒mll�&�����q������W,��|]2κ~�#�7!!'���+�q��ƒ�8�8�j�հo��� ĭ�O7��G��?�����
��1�i$q����I[���K��h�Ǉ�rS�,�a�*��9�\��Nz�09�B�r�p�׺l�k�����ip��+w>Z�l*Avr�������V�A����7�،8�u%uCX1�F�ڈU��)�:a��]����`g&�Fߑ���p8 Q�;̉���˝r.R��bw�9�z��^����ற�h��.�u�bl�q�QC�e�OgO��:���6��ñ���L�V+�`>��T)���ã�ì�,6k�L��� q�p(J�����T�ب�d9�g���瞽~:#����T��`�W��[)���G����֯���j��)�֏��^�쒕Ob�c1!������=���NS���'G��H�d�7LP�6S�!C��MS'׮=������!�ޠ���Z�Y����`4L|w�&{�k�.�o��)��_���ʓ=q ��_O�l:φn�L����r2������Ǥ��G�%<�y��w<F�إ��Yr�;�<��j.C����p���dcgg���{�y���Pl���ʰ��[q~|b%&��l6gS�f8�d�"��H�Ѳ�?͸�l�_/!��Z��dI7Ma1����������t��綶7wv��$�cGnݺ�駟�W[���_t'��C>��.O��,EjUX��[u��zv��YɨOO�ds���ȳ�,w/��2�C�#��M��b㽆|����r~r�_����wf��6��h�^f��5����	4��Pu��L��B|I�~���(�Sy���˃��p3�
� ���[�sKGv��T�R�G����+?���m5����<�d���ĦFū#�&M�7�Y�~ҔRrtr2�'��������U�Q�����F��^G�m��׿�7�w숨�����A
D�Z�H�̕M-,t�H=nܵ��"?�5�ll(��ޠ�9�ǧP�-A3���	��r=�'��?9Z�$�R]��I@?b8
n�e���/�������QZ��bɡ[���G�ޕ9PJQn'� |3ص�NP}����2JN��9�G�Hih�αZ;B+e|��T������x��"�t5bq���m�^�#t�94�I;'��1�D�	�4�gȤ+S���FR�p2���/\���L- }�ݻw#:!�K�p��.�M�!{$G+����b.5�������~q��W�U	�����]�Zo��6���xҵ]�,���:����g��v�n���ܾ{��_��<�ع9�llmn=9�|��ÇM��rM�皌\4�rA�ֺ�N�۷�0庵��K7��`tv 7X������5�Q�&�G�j�8��S��#L�-&#���x��t����6�6�;���o(h�i(Q�oK�N}���� ��*�T	s ��2Y�!Q�?R���+��h�~�1��P*}��L�o��u����<1t�K]�PeRLl�e���@��N2�#�d�8�����dM�mzz�����QV1�k�����l�p1&ǈ�l�c�hHz!����g?�ٓ��g�}�D�3�	|����Zm�`��}R�c�8*�ܱ�~._�,L�>��
����:>*�F�$�!�&i6��t	e�����/���_}���>L�_���'��<�$/���;/ݸ�t�ܖ�~�#�D��P���%�s��$�!	P$
??��cܡr�:��o��|�~3[���h���-�R��u4?,�L	�p��g�s���;�3�
B����X��?�������O༓��s;>�*{E:3~�����@�'�[�_$1e���~p�櫯0ۻZSI��L77�T#6��8¥q+i;�����ّ�V��y�Jz��)X���:DDly~��t@�<������ރjh�f���|sc.�|1����6�\��l�b9/��ؤ+K��N@�5a�k�ȃW���\a��œ�}H ���j����+�]�N*��~DO�Q
�⬺�8d �+�q�4]�C�ƍ�Q�1����G�[[���#ד���{1�>mC����ݲ �6�\優a�|����C�.��qr#�Ď2R�8�SWT�FI7m<�j�s=u���:�r���Wd����T�t�V�ө�#������V��d�Y7���3�k�-@�4����L]����Ȧ ;���#��KE�-Ⱦ]/�:�Xh&��6e�<I|�� �j��<_^�M�����yl��#�����^�}^	~�|2�A��_���y�NZ?sjY��3s�R��<�\1�V�n����[@�&���4�K�������z͢��S�cjs*`�uYC͂�#�eL�$�(���G�΃SB���l��eӒh�Nu�6<V���N��܃+u�!_�8z���K/��;���U���D��
���_�4�#r���29��7�n�>MǛ<>~b^�;#�g����P���gY	�=d�",g��ɃR���i=�FrfD��_���s1�OX&e03��]�Ҡ��ke�����E��4�LI���R��i���I�i�������ė�]�����k#��bOS��y��Z�hz=#哤O��X���˭�_��3������T�~@#�w���ǣ0<�*�Ҽ��>i�Z�8wp�����bi�hj��kbuWjҡ5>�$bI�X�����$�c�����Fk�v"�I��A�Ɠm<�G�/d�h&�\�/�~M&S|�tc=WNי�������8�Gz�<q��$�;3�d�˹#^����L���0
���S�SGYo��;J�I_I��qC��'��^
��q~��K��N_[{���`�S�і��VF~����ѻ���C�?G��c6c�0)R�9�|;A��u��^k�h0�ɐ3��֪hmjDL�x����]�f�P�3�k���8y2�!|����T�|���Ti��UO�UǙ0��]	=x���W�P��3��a1R��Pu�����me�kE�3��ݮBB�Ƃ��k���1φ�G����>�I\�+�,�*/c�yJ6j_�0�e]ʜ�8G��i��n��q_�=M�*Z,g�dcWb�@��>u,��}�<�W�M�1Ԓɞq�C���F|�,���"���&����A���e<]	�+X��DdD|�^��ʸ)� ��z��i�f>'6�9<B0��?��H@��r2��\�ц����'�B�h_�vJs0ppy�[F���$�>�$rr�R.[.��=+:��"8ϧ#�Y��O~���~�qpm��H��f����5Vka�Uc��<�Z�K 9E�g�k}�<�?�'��%t{�!"+��|�I�t�Z���YOEPI��D�)�p�"�a�a�Q�F!�ּ>C`��T�&&�iY�.��C�LJ�J,c��(�����F�GR7��_x?�l����w���;��&�k
����*�4�R�Vn򻄼��=���ffJ�-uҲ/^$j��C���{������`��{��A>�"�YH2��4g��w���Q��-k5,GJŲ^�[x�O��������k�[Z2��WZ�kb31=f&�e}V�Q��D$$2k�V �&AЦ�5:^
�(�1��|AV�k�T��/�!���Ӂc��ٝ�Ō=�J����$�fّ�����;�ϣG�>��c��.�-��4cJ�昋Ὃ����ȟ���o���W��?=z�������� ��ݝ�7��!���-q?ʃ��3.��޻w��ի��D5���(��ۣ�:7ɝy!�J��nϮR����t�ckc��n�Z�pO1%I��$�2XjJ����6�� 1�ӵ�	
d�1rn=�ť3�<nl�Rˎ����E~���'G]��g���_,VP�x�$��Pz��r�ڮV�*��U�V���	����b,/$��I+&�S�&C3�[��^��{��{4�]�1'Jc_��j
ı��`9u�m�NA������[��q��N��Q~�XM��C��(�Z�pЖK�����"q�u�>2�=��ʬ�����$����m-T���"�w�k}��x�~oȮR[O	���QM��s8ѯ��*Ǆ\�B,U�@-!3&�4�͝��j�X�$V���O?���pϬ�ڌ��&ND���\3x@ʇ��ċª�:��{�u3fo/_<�ꫯ"&�J7����?�'�DPh���t.��Z��#�Fy{.�-� )<.���|��d��B��g�|��]�j"��~�M����;Ԡ��:�C����R��5$�l�-�{�nZ�@�^���+��<�u�?Lq���(����H����bK�w�3��t[�M��t�Fd�2�vr{�lCȊ��b8�9�3d��`M�*��o1i�J��j����av_��x"�ũ
��U �J+WƸ*����{����*��B�lR�9W���;��.Ǧ�	�x�<w��ZD�F�S�TS��6�{fӲ�u��4�skYΗ��R���x�F0iq�#P����׶��۸��M�N;�S5*��6�J��;<�2|�.�D��5'XYZw�$�Ո-��dá�UXP
M��EV'i��!��	v6�8�9�1�C���eBy�6��t~|���Z�6�,�F�h�K�E�j�Κ��Cg��2��]/WJ[��]%f�9Q�Zj�P�+��i{�K���r�)
+k$1���i��9´��>����*�y��D���<~�2Tܧ�)������I%�f�5n��o4Ԕ[����j9���p�9��$�!��8˱�4��g�žI3{����ըc���6B�X�iْY�X�lm�4�P����9�g3����i��w~���I<�`��d>{��g�.��s+/r�R�p��Vu������6��
;�b���h<G1�ą1��Hd�-;�VX�u;:MҦ��<��O;�.]�Gqc���B!��O��	ϊUh˚ D3��h���K���M��_8�΁��6w�|�w��$M�ޤW�+��>�q����ks��r��#91��^�W�Bo�pX�{���Ë5򨄮�E�;��7�;Y�gvMOZ�α)�jm���ؘ�|�?w����w���_H;-eͳ\�BJ��Ù^�V�׳��xc:�ٽ��u�ÆeV��3.2��Ur,�x�	�K�J��.�K7�r?�+�s˒\xL7]�7ml�L6��;Y�R���, �
�>gk��:}f�Y ��a��͠๨�'���S��s�l�����x������(+F�����aW�K��詹���rQ�ah��\.��?(�g�%����W�9Cq��v6��Ѥ��A#��Yq���:�[L�L��Z.N��D�E�D���d��/˪�/V;;6��6���],�90��榎�,E޷����ue[i<m�ʂ�3nOڬ�4�D��|R��83�G����8ȸ��"�Ө���ѿ��ﯱN�;<^K\���2�!�����ެ��*��Ѭ̭�Qgywgώ�
��^�W��˳�`$tR��412�si�p�[�0p�h<m�t�j?~X7-sX�0N���W%�� �}���2�Щn���~�ɩ~UGFE���,��M3O�$[g���8���9T6��&x�vEa��< �����*�s\YH�tm�=j�js<�aVD=��b��9����"����X���`�5.�������sr��E3&�I
��o�$R,�i�@T/�+�<��5vp���&匶����OGUD�Rn���^���z��$d��l,���p{��ź�K�j/�g�''�3v�Z$���{q�1ʋq���EɄc
�����R[D-�{x�f���������u������T)��L�asN��ul3.
���m�of�QW��M9��v��iT0r��&�Y�t���=UiS��w&�V���{��6$1>\%R,�oY
Ț�O����kR
O�(ݐW�9;A��g#�|ǫle�i�#qI{T����A27��<���c�*ƱP�x������on!ĥ��fGgx�t'J0��a�<���/%*5����NNu۵��3�|1	M�-����6��Ͼ�o}kww�o��o�?��?���bTё����!���|?��W�GM�gńlk7ٷ�_�avV�o�&����>:Җ�� s�(iK�˲�X4�q���-e�t~a:�Jd�֨�<8Hp�ig�K��.������0��A���N!���R�n�����JgI'�������b�K�c�Ο�gL�8�q�'
��/���?v:�޻����3�2݉1/Q�8���2�I!�����>��D6�˗/]�:Ol�1���""�����a��1��C��,k��+?~���1�����>O�O�6̫Q�!�#�	�>D�= *�.rj��gڠp5��X�Ap'8bׯ_WV�>�|)blV)L���C�4����v��j��t[|&��xG��aAu�:0�	O��'DO��q�t�4^�Hx���";ý��v��-�)<�իW��O�to�9/����͛7�����1?B16kϿ�^��*;���7�$L�Jֺ�O��F7�v�3=�A��v��m����H������x4==�oo��eR��g[5{�@��h��U@Bi3_]~:�,�� �?��O�ݸq����IU���ml���[p���.L&p�z�ϠIK:�j��ҥ���1�6��邇�Ν�>�,���fd�-	"���~^�6W�B�Pt��T�	��B��=8��\�4��������7���C���6�Y7$Z��Ժ��������"���T�W);rVGӭ	nZ��b��OO �X\}g{�����������ImʚK��dh5"|��ie�Ow���x������#�i�j7�*���U�P�1��e��D�DQXHd��.�m�2ǰ|�O�Q5!�7F���34n�G��u��Ρ�rM�"�ȱ�ƾ8�y��~N�����'�G�O��T� �
Z5�W���SZ�J���p^����jU%1>!���(�ȋ~/[��O��4�2<^�
M&B��r# �@���jZ�5����A���:~�����hP��M
�]7L8����[nV�<�y"��-r�e�2O�t�$�:�G��2�J"4~���܇`&r�κ��o�o�m��,g�n�1��ͭGoϯ�LI��z�J�n:u��:|a����LF���PH�7�;<䘃w���z���'��y*]b{N5�V�j�*��L�����<��wt!����K��c�(�����B�Ҹ3	���nL��s�B��� jdP�,x^����iCH��0������cZ�j�(��w~|�S����ݻ�~��Sl�uJj�k����''j�$��u@�3C���H�L5ƥB�s\]i�pe@
�e�p�����$�~�xB����=�=xS�.0�R��6�LF:��䦬�N9��`����^����WgDf����#�o�gG�ʓ���^�!��ј�$�-y���m:d_�Pn�a�"�k[�NB6P~4�j�ܩz-���:a�7wvf�����4V�$������k�����}��3W�X,�������?~���a+O
�Q���0�yE��%";Vr�f�MfXN'�&;IU��;7_���B(��uIgg5|��M'fc�;�+f�K��?VLK�hޗ�/w��ӝD�p��D�#.�s�����-c��l�0���M� I��4��.��T\ڔ@pC��g:q�ԏ�2_7�.]�4�«[����1y�u�tgB�߉������7�ĘZߤ�#�P�)�b�P��!��c�f����|��7��Oc���LyH��n"?5+�B=�_M����%LqY�OW�'��XYQW-Y�I���{������t�#�4�/`*���Ո����O|'d�����6Yb3Q -�hՂ�?m��'�SjU��!��+�6�y&ZU���w��������V��[�tm媩��ysm�~e�4TI�rl?þE>mO�Ji>z<����.����-��C��c�$3��J����H�e�'�n���Ȕv�����l�N�`$z5����5��iC��8��r�`@�y�����?:x`e8=�_}���{�\�H���e�Y^.�Q�w3�i����k;�­���s��z�y}L,�bm����d�J,BZ[e�EKC~��m�{�r�ʇރ$��h3�"ކ��
s���S�YM�k.z�@э��lo��V� �QΌ��%M����O	Џp���"G0�OQa�r��?�i29 ������(�i�V�@��/qy��;�w%�GI��P�I�4
���=<L�x�_�а\L��z���iO5,xKlu��7^�7����MFʑɠ�B�7grd�XzO;�I�{�C5
���_�
~����?�a_I?��NO�8>Y�9n꿟t��Ɠ�Ӏ$�����յ݆�q˙E��{I��[�&-�2k��&��� ��.^�G����l�\��8�rZdgeǕ|�Ս<K 7���ۺm���]�q1�����J�*��YP��r֩���W6��n�{?z�:��F�|WXX\��Çfr��<��ߚ�^K�HsL����p�v�ܓNe�7� ,��qX�ܡ�:��^`� VH�����l���^1U�ym�oc�%�eu3��q6Ǝ��\Sݍ7Pqĺ$�\]�>Slڭ[�zոp� t,ތ7����t���ݻw��z����&ޫ�o�_�âJV�tBN�N�q���/8i&��d��΋Ah���%JL��l���~Y�J�R����~FG��¶�Eo�O��O�{	:�a?~�DT��Ǐ�� �'@�>�/_E�$l���N��gU��Ӥ'CW^z���N�FZ��W0�����=tY��~�Alԓة���ʉ�f�H:�*EXI=����^U�G��/�����_�����W�nlLtޭ��鬕!����nC�Y�q�"�2�Ճp9��{H�,�(I&�H�#8<x��	$��Ν����3��Qc�CfF# -�0�����������/�r|���o���ic�>}B�	���Eљ��S�/��;w����'���[�ō�X*�T�E$3:�	a�B������'�M��889u:Ը�4~Ҧqa%oЗ�:w�\�Z}_i�ՎEW����W�@�K{�Z�RR�eMBw0ݏ�����!�k�x�E.�o�[g�h�s���|r);�c,�Y�r�ZF1Js�7�\����/�ԑ�u:;>��IɜM67¥��WU�!��*g��k����|Jؤ��}���K;�CWS�y�|;[L
qۉ�ݜf�}��i���p�������uQYՆH�\���S�v����AC�Z�j�7pܪ^uF|���UD��$j*G�Q�f�,�ɪ�1��$��\;���K�0��F�EU0K��1�r\���5��������+��͉id���Y��<��B���H��XX�iэ�;��U�3�A��@�]m����M�G��+㖓���KZNje860%Y��oi�e�J���SGSN�r-Ky8�����>�`m�l���yG=�8�`}�eB� V'�j�H,s�5䤊�]�B����R*C���ޥ�����9��)�D9ۮk�O�CTПOH�e*B�e9&뿮�/��u���4�����{���o�O:G,��b����0���.��G��8��2�R
�k��w�w������Z���f�t��;��kzT�	�U��T��������f5�i�/������MȌ�4���z]b�L��6��Y�k����_��Ylc��|<~rr��S�䀭"7hl0�ʃ�.��+�9����R��l1_���Of��*�����|��ps�1^�`j|C��;`=M������o��M���F�*g.��Q��)Gi.�8E8�]��	�0�]u�Σ&ʱ�޺5_.�[���V-�F�"��A�Ɠ��]:�/_������uu����d�`��,m��3$��&�8���'�U�.���(����VA(b�q�QˎE�<�cC>r�4q��'�G����k�"���=��1��غ�IV�v6/������|g:݂ȟ�׃>{pV�rD� ��<@�.c����"U�!�\FY���l���mo�{�"������'�sW.�Q��p��������{�VQ'U���0%!S���9F1�G��q���`�{E�7��e�>�i��s��%�O�F�%*9��κ����)^g����l!�Kc�T���A�Yp"�V��X��X�XxH����QOͪ��l8R?7UL�\��� �F	Z���w:[��삥��ր�Ʀ-�<˃���J,#�p�}�Ȇ8�р����DT]������;��~���<١+O"�����_|։�∪�����8�|��˵ꁋ�c.�����"�z�H+?H��_���,r������e�M8֣�&�Iډ,`�֛��I�\�Dp��i��)Y�Ù���g���:8�3��R����T�M���F��y���[v���V.��SQ�ۚ��|��2D�(4�-xTgK�x��.�,�����VYuN�a-�x�z��?<��0x��#����ݐý�.Ϧ5�Q&(3��;�b,g��7j�n�9���xG�Cj�d<��m�ҍ�=�*�y�~R������3��@����	e�����.
L�bYC������Iϥ�|]��r�w�M��*1r�c?WA	tnM�IYu�M66����1��ְW���@����F���7զ��aI�r����W��?�b�Ї�H(q��:?S>$�2_�1�r5�!.��-}6���7�a��N�Mї3���ﺒ�z�z�v!!�Z;�S��$����Y�e�v�[��^T�O.�2\�]S?[Y�l#�Ӆ��� ށ�_NN��Z)ӧfOmqϓ���Δ'���k(��T
;C�՘nk��{�7._�l)����g���%��>����RG/�G?��<�����xc2��ƫ�M ]����d1��h��Et�\�yڜ��T��y�����A��K!��Q*~��_���j��"ܺuK�i(=<�r��Jø%�L W���]y�V����V�R��<�i4�#~ܶ��*���o���έzG̝��:�S'� �oNbr�s�;;��(;)P!����^�A�L���1�����vO�g[���b����<?!+��r����Y(��/-�=��7���?j�Ƨ.\���e�����!�^�8௝��5�YIǧ'p �-+5�
J�@e&T�`κs]�̘��d=�|q�	J�mO+P��:2hZ�vL�;�^�gL!�����ի�ȯ~�+|��7��b~���60^E��"�м�ORv��\�[N×���

r�[���T��ձ�'O�w��,RIH�6ƺ�?Rb�T��꓎U�d�a9��:��g���XŠ�$i}?27����@ Yq�����C����["F`�pl�9��*Dr��sv��nkk���������%-=��ҙzϚ3�*��T���	Za�U�@]���N.���f9� ���~*�W�@0ٱ�(1�a�J�z��\@n���/;��%��]M[����Z��2�T�FܸP�z�tncn�������h=)�6~nUV��m�f�#7M[	M)(�K�M�~P*-����)�[j�^���",T�������>� O
]�F�-H�'�p��w�W�MBP�֘���'ܬϳ��^����r��C0U�>������N��'Ǚ	[C��Hh���B��޴ɲ���s��	�Ba( 	�lH-�I��n����u��_�p��h���Kl}�'�r4#��ЀHb.����9�tg���9'��b2���=g�=����l�&GHR?y�k��2*�0���KU��#"7�"����a؎�Y>Ӹ����ԃe��HyI�QBI�c�0|Nΰ�c6[V�m��� �|�r9�T��	q�� !D?��~�l�,��8KI8и��K{�Ǒ��;d���kp}�G\s&�fpc�QC�_��ܝL6.�i���R�	*r׸04-4,�Ǩ��.���,{e~����(�#f8997%e6F��� �2,��ȕ2�}s����tWFӭxe�摱�bױ�;���
4��B�F�S6��@��ܿB$���Ⱥ�,���.��I_����h?eW�2� ��֝$���\ꫥ����n&��{�/c�HO�����!k;�G�?l[�8�W��f�F_��q1A�Ã�	�T��B�-=r��%���~�^G^�
�>�"��yi�{bO�*	4�f9B�[&�W5�Upܟ��:�����d������X���Į:UO-�
����ʧ1�!5'���	rdO
h���I �AS�\W�H� T�lr�����j:�۳m���kSᄈ�
#��ɘ�7�Qg��+q�3�(iD���,}0{��Ϥ����ە��������M�e���7�$�����Ƶk�NO	2����./�W\�&{N�Z��� QU�H<�nL�~r2��Jn�6B�#������6d$'�mB���ϟݿ��@�.��
xfl-ɫM����4�t>;��\����o���9Nm�&�8�m�'�Y<<�/���["�)]u��=�44xN����cY:͠�p�����Zq�W{�Z�|3���n�^��OGghqn�� �w�,�䥧+�fS��� yf(��M�ҳk�"7i���k��_��tk��6t�f6�73\F���\���P;��/c;�
<b��.�E�O�9�,B1w~BN�*-Z���N� � ���b[���K���3ȶ5�F�!)2ǧ����g�at���IY�H���C�����;w��ܾ�2�/�K8�7���<�{Ù�!P�T�N���<#벷�*�ƆV2^��������p�YM��o��[��� |��'�U�JN���!e��>���$QW{�r�����:W&�#Y[.��ʍ�p�X	��=X�!� <y�d5g��U�h�ԆFQq��@�4����4�5��*����ef�o��C8�X	0�t4�AЌ]p�F�ڸ��5YDGc&����A�}gs�֭[��K�옪
]�M�L|��@6Z:70L����yc7�m`s	��H,�����Ģ�1"�1�^f��������Hx��G!�Jݳ��z|��'%���>��.�|P��){��ȡR��-eYI?��?�q}��&0Y�{��؏��P$!q����e*��"���<�E���w�V5)�
�!���x܉�3X7q��;�8�u{�z*@���"ZC��������r{����)z�@J��餖} ]+l֗�ɉ��g����q���,yي���׮3@:A�KU���/^X?=�n���Uz�TF!���7��r�7*�Ӥ��؍th}?P���O5��̬�t��&���(�\Q��K�$�a�W���`��_�Nj]�H�6+Ƥ�M/���[o+̑��~��D7����w�@n��ښ�hYKA&�Hw��]3O���+������o�!����/��R�*�#�A�}S<uf�|$52�n�����.2[@�X���,	_��RZ�
��"�/%w�>|B�u,ˬ��e56^c����җ�d> ��΃�k��P��Y����?�ū�����x�ӟ��0�C*'���o[;�τ	�8!��)C7�)8�d�ZIi�e�)��!f��<u���5����:��V% 
P�AȮ��N<��_�N�bH�P��t�>C�����a�1�i��ZS{�;���
A�旝mzg�a'�Nջ�*����+4�dO�HiĈ��4�Z�B7�"�Q�J�I�ɮ�så�uq>����y�ƒ�**|�嗕��m�D����"Oe�������۷�������xdXl&����Z5��Ʊ����Vm����;���84��?i��_�::_ya%
�U�Z�Fzzt�,}����W4F��U�jkic�N�]��u�����q�����"*m�-��V`�.{՚I�I�^����\C*�V��,���M�E�y�X(U��w5�[.�x�j��k#�B�0��f�R0�sG���>}*b�؈�t�*mbY�|�Mq\�7JA($�ϠI�)�e�c��{�ϱG����ڴ�����9�Sz��D�i�2"��$�A3?*-�m�:�B�re�U���j,��}~=�uF�|�X�:9r�/�g�CG��񭅋�ֈ!�o���Z�勑ʧy;+%%�	�%q��G �����W��} v`4��sXtak#q���IG��2|�/�v)�Ŀ�DuS5�V���9�F�J�Q7��������me�f��%v6�=�L!ig�f3�z˒�[xM[��4����ԍ���(mZ+��q�&G�Fq����'\��C�5v Ƽy!nK�]�q'l�� ��)�-�eId�+���k=�+���ɰY��z�2��[�k�.A<�v1MҼ'-N+��H��p"��e����:�ug���bf�6����bi��U�X�!n���U;��%�UFZ)�6)����'�s(��wvFU��3h�Ԡ,��Cz�C65��9��X�d����h��'���؆���y;�}9_`�V�2ϊ8���S�UO&pd��h Z�޻w������p����U(aIF���\��'Ǹ��/���GO�>��踜�Cw�=a�h��S��>ӭq0���v!�8(��g�-a����gu����;��n�%�ȗb�?�<���4%Z���[��^�Y��x��g�`�nߺ�7��c{@c�?=yz�wL�����c���@T+^ˀ��3���=kC>��G6M]J�JY�ai8������6	huIᑹGp#�[��������]�q��ʼ�������)C#�XVVVev�p�ns��Z��"�1>}��tv���'O��6h2d�|��Ó�'�88��C�+,�H~���k��W��ɋ�嵖��c����8�+<a�M&cc^�{�6+�7d�Tm.|+_���ɸ�E�����z��b3h�/�x�ŧ<�Ϋ��5q�}I�U�' ����Y�L��a�=�^��1� bդ���]k��I�����!F1��F�`b=�a�������[�>��2d��٠d]Ob]�[mW�wpZu����F� r����/E��V��f���q|6;:<�����,��N�j9ʿ��S��3�p���7n�8����O~��K/mMh�K˓��8x��y�	l]��yH�8���qJ�-� ��8}���x�W><�Sux�o�۔�S3�TNf�p*&S佌�U��+�8�H+U,urs?�%e鸨K�QY�v�
sܽc������>N
�P�<���0O��Y��c6&����p��b�F�����[�ֆ�]U��_�����hZ�v�M�NS��u�c%�]S<*�?���.�q���ϫ���S(���|q1?���d�a��o@���s����#�⓱�Ya٥(��r0�Z_�+x��eue�qt�����xjрB[�4jx�!>��K�5�K�V���N���h�Q�j�U�Jl��7!9��Ȏ&e�.WẰA8��޾1Jr��9ه]r�A��'���|8)+����Yd�'Q�<�Mp�C�-�5���l���b~�|g^I�ٚ�Z���+)�$���3o6��r��������c�ͫT�X�Q��\���r�!%��%��Y���0��G�GvZ�c���Rh^0����2#_�T�0D;z@�s����~��d��!%'���4P^É�yYW��b8"-,{���_��
�ݮ�>���K��S#H ��3z}bB��2�u!e �P���O����K�[��T�4.��j������/�ٟ�ٝ۷q�j�y����XJ`�3n୷�B��@W�=&��#+˃�#X�@?��j���q�o��^�|--��n���Y�VՓ�h<S�K��é�v��+�ON�R71�U��������:ceZ9�������9)�`���m={��/�q�3�<��[��.�ַ�0��zD�JuƖ���ى��&<�t:�9`CY�<{��uQ���.�������D]S�7V��h��+qA�|V�������w��*=��ˋ}�q<:dvN���k{� �q1��5 6~�IGf1�7HԳ�Gs����3-t5$�S�|@Υ.�����B�����q��!O�a�G��h�����S�<�
r?���� �иA3�~OVp��xc:�N���Otvr�駟"��Q�Ɓo2�ew�^��I��T�l�P8��װCnq]7J�vƀi<q��l��[ƻ�'"q���o�!x
v-�q�8�!�y����}{m'%��Xק�|��h8��`�	�l�%k�2_��
�ݭ\m�`P,s�*�&�Z-W��av")�f�����Ǧ�O�<�G!����^˕[���� ,�+��"��w�*���G��c�V�f���Vj'˙�M�9�#/: �W�є���Քmj�,����8�Ď%�q_�XFpL�ܹ�S\��� �b{�]��IA�}�-�,�03��%�k�'��>5�vL��'K\g�p�h��zi{����7���CE0Ķ�o)��v ]�/�-T):O1g�~�"Чa�sEa����T�t��_�P򯛑����!�Uc �ޓ����d�u�۞??��h�ꫯBq������ڔ{��Xo͌^b9��&�R05�>�t�|�Ahv3�^�"`�ê�W�/��z�x+��_/�X�@ش2Tx���	�����\37÷]�6�\���3��b�C'[�2�8GRi�%MYr�4��y���d�W(�H��R�y�a�A��A�1yQp�򵉽��.��I�1����ዮ�I�!���IX��L(�*y����oί�<�R�yu񐺖� 71<�����i����6wݺ(���<<<d
���H{�Sp�t/���ҙ�
���:6�T9r���.����@�۳�[sh�z��'���^A��n�E���-I��lf+N\�eK]!$�6�s�b�-�Y�?CD�H�1���
�mo�[���C���C����:�a⏏�����)�l�%��VGG0*I�U��C��G���Z(��ә�$�yjsb*)�.,k
bF�r�28ٙ�,�V�����aQY�)k���\l�J�_�F���B=�ɐ�מn��x��*��G<c~���ۘk�?z&Xd�h���E���ځ��ij�� u''g,�E��i
��l��&��_CҠF����#�p0�|4Os�.�K����<�p�;���E~��j�Pit���Ӛ5�(;>���sq�GF*��	UO��x2��on��	}�م� ��C�U����..��6:r�j*��єk%�L��^��x�{���N��,PW+��X���9�V��_n�[g�i2RϽ���d<��^�������H���z����s߉���:���o.'Z�B�&�?�U�3��E$��y�����H��N�����8k�}i�T����f�2��a,3ug��p��)�AO��@ӫ��	7n9��믿��͛��O�GؽBF���O�XY)x�THl�s�pI�@��0n>!�y��'��w���
�zR���	��f�z�@�q/���� ƣ�8K��l��p^Wɨ5�����W�G?�я<����g�3�<.��r��>}��D�B��#*Ûsn�5��҄֩�X��������x���	<ys�N�i�'X��������OH��<��.��f���P�Fɔ�:H	����B�*㚁<Ȗݚ�3��3�&�b�ւ��s�>�W>�\k�[a��z#"��t���/!Z�Y]���S��}�U<���	�9����tE�{vz*�Wj��U�y�jx�˦���������)���ԟ�b�1�F�nn�X[�k��s��E�[GR��f@ah�c�P(,��%�q<�2���u���ß��׈1k�Z��8"
ͤ�<V�`D�3S�n|e����`�IvJ����?����K=IE��y�o���b+�)�V51򥈐5Rϗ��X���{hO���,7I�.�?">�<<g���{�ZTѾ\P��x�_{�c�w��nb]���wJF98�r02?�1�T�J�TF[��ё�%��$r�)�v��ie0��U����8��nlN!cϟ��{߻��c7ө����/����b���Z�ml_��&ZTU3|�Z~�%͓͡T�)j<�P�ژf틶U�a1XE��Z=�l�mY'���}�����������P6W���>�D�~�2�;��t]p�Zk,Ж)~s�t��g��mBe���5�e��E~��43P����V�'n^yj�>���(l��1g�B�~��g�^z饷�z�6�$�:������[����yt�--5�Lqo�6P�v�\�M��t< ?e@NNN��a-���V(u<�g��ǿ���h���o�`�d�^�G�*)���B��ICt�C�X�3_��u��wb�V7Y������?���7���ꈵ7{�4�'�F��-�+�l�|��g��ۡ g�����}<�R� �ڵ���?� ���+K�$Xc�F�h����� ���^H�)A����!}�p���$3�� �K����J��=9iGO�[�/���7-a������tXJ���<+?��0�!1S�n`��V��z����t�<6JZT'%:� �&�ZNL�j;���c_������q�����*��|���ֺk;�({�mg�:����MG0ϊ�ĝl��,�s9o�^K����T�R�Oq���/�Z��5����;N���h��AA�+��B)c�,�u�g��������'.�8������|kc*�����o>P�������!��X��mc/G�<��$��Fcgz�V�Q���N��+��"�m�D�>�(����<�+����B�f��@����/E����#`��*�����+ԧ���>�"6���_���$�  ��IDAT�
/�Q�������r��I�p{?H���>�	}W�zl�β\e�Lw���+�`��F	��)�.�C�h��$�i@�֭&f��1䝂��<U(���ⵆ�g�WY'E��7�|hHO�W0bpy\��r~1�#G�^�qӕ�������4�Fc�
�m�w��J�Pq����6���XCgD��D�l`�lk��L�/�Ֆ��K��r�M6����,z������@�>��ֆ<S���/������<�h�C9��f#1�hiG�*�
�L�ⶃ��5���ߓ����ab�ԾW�vי��:d�@:��a�'���]��]o7��jc�q���T-�i��K�JE��}E:AW@�S��6;܏IUҖ��eȇD�joB�pw��&��]�h��q�[���|�)[����82�=�����M�Wv��]��=���	���4�	oJ�:���d��� '�:6�qZ�p�K�J��ڜrGBhSMe�ﰲTO���<�����DaC��w}���C������)��4��#f���������������V�����~�ao��j1?%kL��6Fc�%�4�"()�]R�C� ����Z�=�*H��H�EQlY��w�����UX�����d:ٴ$�P���0rxW0���t8pۦ.+RA V�,���#�(�`=;[$�q�&�r5�l�jldȸ�mc�	�F9=�d!v�m��E�_UpU[3+������}/��U�HVB$�U��i�^ٛ
^�\=k�ǒG�醘�Z�̚�!� ��V,�RJZa�nՏ��j���D͠�A�=����0 �V�Ꚋ��� �,�������|��������Q�xL�~2�A�,9�ӦhB��������ײ��m�.U�]4��%�e�RM�9���u׌�K���!D:+6p�����3�V��a��"o]�reV���ϳq:�Lqq#Ȫ]�6�Vaa;��0�t<agЪ\����R.f�����]-?����z�O���3�P�ʺ�9N4�le��S?ښ��*�¥�y���Ӂ��1�;8E�<�9�`��`�����N��;�uc<Y,[��/NP���UC�\��kijD���8�
&�J���Vλ�������]{�?��̚�/.V3���Y=~����l9�(����h�Ѹ�lI�^��P.iT@�UK��/!xYԧG�%i��Ӈg�'����/A�U����2�ᚎrX�퍩��1Y�*'#��m�}�g���||z��3��8?H�zX����c��W]��rQ(��E�9V劵��{�t�'Q�,C�p���1*I���D�] B��7��ރ{�=:�a��X̗\�oݾ~����Y���m�9V-�	��c�	�rg�Wv�j�����X	 ��$���"K3���}Y^tQ�<-���<6����`������7��A ��YN1���WKx��T�c�CU����y���S���Xt�I��F��1(?�+�8�pp�Ӥ����bx���0ھ���!<�r���������k����/��!8ؿ���!j�ÿ��1V�[oݽ}{wgw��ѣ����S�G�L�*w�~���p���$���ɓ��C��9�"�wī]�3rtN���b��/B��p)��a�uK��r�4"㸭�!d2�=.3��t:��-��b1{t�����ٛo���ҧ��������p:�0I!�0.|�'Tn^�s�yr�_~�e�G�jal�?��<�b�Ɉ�ǹ��#�`2)%Ćm�����܂ƴ�#3���K|1QM���ٔ�t~qj@���TL���U�iN�`���i�����y5�r�ja���c�!��R`X|P�n��-*oP�0S����������J�ā���0��F�9��O�1���m9��@@����l�w�u�VQ�]5���>���l|�dD�ALw$�<��Xx��SRL��_J��"-�f�9` �FY�_��jAin\�P8i����ȽM���`f�ow��C%j�|�6��hx1������Ħ��f=��n��rv>?���I䡎�qZ�&ۛ��rv���EYE�`���_=x�byC�����*��H������ŲV"������*$f��+����D�9�R,\�[B��[%L �H`���gp����&l$�! ��۹��+o�����~:_.s&�=�K����m냃c E���X͵Ί|p���[�nq	���������)������8�D������r�ŋ/Rm�hN}��#6bck����O��C;!8ǃ?;�_�+�i�x|F��	B��ͭ͝m�\��o�f	/�<<<����؜l;�P�*/��ٳ����N�.��J+'�1�o$W�����v
z����VX�Ǐ��?���kWq3�e����7��X��)� `M��vꊭ���}�+���>��|��;��Ζ�NUC��q.	�l	A͇��[ױ�����ן>}zxx��@x[�������Cc��4�7Pq%+��;m�66��d-���ّ׊��lC�7�:L%�|�5n�aN=a�������f�f�/�:x~�'���������y3m�������������*�Oc��1i�H#h^uȮ�S���V���O����>iN:��gJ���qNy��t��10�l� "�^YS+'����=91gc��>b�V�� cP$K�>��'g�?��!����v��soUA�yE�Z�Owrrdm[���sʉƃ�ث��h�%I�]��!�j8�m5,rX����ыG�,$X�2�t��b.�����Ҡ�D-uF��}	������g$1�d.!`]��/��A�,(�nϞ=��Hs�|�0hc0�,�dc�u�����@m=�����h��ˠ5��]���UҖ��Lt@a�l�S�9#8���̀r��[$q�R��b�,ǥ�	���T�QB����Y12���P���S��?��8�2����Ϛ��z�������"�T�eE/�M�t�!6#�%G��y%W�A�p��������0@.IGf9۰�%(���\O ��lsj�rD�H��`��mv'��I�6�<N�]z�u P]���2a��GX3H��1�5TGÎ��@�!.tK�%v`kZ T����+{NjO��8g)^#c^ޔ��hU.��Ζr��$@\�e.�Q:��evv��5l,��a�.I]�_�A�D��X����`��V9	�����u�t�u�jE~�lg}P�!]��������唨�z�(����<-�V<|��C�C�i�'^��	<�X?���Tġv!���s��p���+��B��Ǟ�:$@�=\$�3���^W���~�p껽9+(770#�*e��j:�+�d|�g�l�K���7\Ğe<�hJ%�E�%|�M;�Go�I��Ӥ���L�ے��z�r�H[��AFށ�ƈ��\��={W&]w��!��_J8C�̘���PK�����7%�>�i.+�آZFUB�k��.��;�ݸqn������{��Ң�Rc�Iq�E˭�5���R|C���g
��:5�����0J����1J�s&"=�!ɫ.ѐ�Tkq�D��gl<����"�"V��[�>"�:�u������zO�$a�ӗ.�����y�0�~�`�'k@W��7�ݳ�W��Vg�����7�����*Qh��� 00��6�����v$ʱ7kM(V�ˢ�z���RߓE�V�<�;ߔ#� �>����X��/v	����z���#,����L�I/;;��z�:$���Ͼ��h]U�Y#�H<����k0d�rm݄�Ad����i$�*���,|	v=��Ԑ�����6wa:�,�oe%��c|&�X�PD�S(�X�>���M,Ƴ&�N.��ڃ�р��L��;e�EF�����;�^,.���}%\2�������/�jb��0*���� 0�пx��՝kWԾ��=�a8�K�2�I����������k%ANƗ_~�[��b9o�\Z�p����$�ٙI%�.3��҈��=Yq��L�Zkԕ���w��!Z�?��bκ���� ���������@h�Z��}UYM��#hAR? N>:�-Ms��*\�:��I����ڸ�ř�k��_��������g�}~q]��ڦO(�Y[/�@�:��ӶZ��!�Q-�'G�y�w��5jݶC�vpp�T$J�:���Rg��ˡ��������pv�w�z��;�=z���ϧS��9�Y`�J�F�x��ׯvi���3�W�'7�]�$}13�#v
r�+@9�f/l�Z�H�脡#":�*3��=��|c/�MK���nbx�G|L&�p"�6���� �}�(�����9S��@�D} 6�}WV�?�����'�|�)�*�#ne����B�	 w%�3ҫO�~x�n5�f��5�/�!�}�̷j���:,E���ߤي/���e����u�Z8h�g!�:�M|7kH���ǰ�ݣ���Kt��hC�?���K�J>[�H
��԰6K�to"���a�q<��'����*���$���n�.پ?�Ob�CO�~��� <����[�uK�cy��ƻg}ck.�6�r���,�V^������t{�8OLd�Hu}R�N&��R��y'ϖ�*�*!��ֽXW���G�yu�<X���l���&�u�5�@���d�4�Ȱ_���/oܺy��-�y;?}����o����'O���g�������/�]�M�)
�o����^�>�VС��qzJ��(!���q#�8ygPS�x̭���v��Q�_�0(7n^�j!Bh��!6�Rː.ݐ_<��=�|	��/'���L�)�'�����́�g�0�����?���ꫯB�c϶,�$�G-Aο9�����WZ �@�Cc#�/\����"��3Y,��`�����%8#�Y������|S��z�{
3�س"�5U��4Ul�Q�,�0�
�_�j��tc[U1�=��>��?��{P�/��xX�܋�C\��͞V=͔
�Ŵ�a���7$$�y�W=`�)��c��O���e�u�["�<kȉ�/�Z�M5����&?�*��9�>��O���ݿ���T('|��5u������$����;�9��2b%��)I��8s)#ۀ�)_��^i�ߗ���{-��c����n��=lj�l�M�!�L*�=g���x5R��
�E���k���<?�T��`]���n�k�lz3+����������	3K���G��V���Y�C'Ñ6b=�'��̃y~����*�_rU�VKjq�kTGS��e�R.:2u�j-��e9�5������&��#ߓ��Q
!5�G�<!^��F_�Հ3�q}��#85g՘�C��Zئ�O��3��6f.���2����L�K��������t1.٪*I�b�L�Q�,3�%�B�{�\ٱ�`��ߪ$֦*e��m�1�E�6�&R9�,M.�he�^Xe��n��].Z��֓G�0�!�*GTa�� W�K��;��rd�֦~L��:�_>��T���V��i��'��s�Z�{�ꢺe����I�Ù�=��n��ͪ�gM�<�H��M���c��)"Z�t��7xp`22���D��B�~�����ȻK��t�I%.�y��p?�q��e���z�����u��6�ʖ�G8��/�sA�W0����?����=x��ͻ��9�޿*�Җᖆ�&�_�c�
[#b��"���z�������xӕ5+�/������������U��?���?��ώX7��l���3f(���ړ���r�6I�~6;��6�bٜ_��C�>&8�¼Ɋ�3�1|��Rl͋*Ґ@t"��Dݲ����"���Fx�')3�rn�%�O��D5x޶n���g4��K�}�2����*q�k�<KC��H-e��k���&gGA�Ki3<TA ����%]�Z���8p&��^ZCW�H�,��$���1��Mu#'�ٳӍ8���'���7�G�mtq~��f�eT.��������O�
��7����,P;�Q���K����ݾ���oö����կ�yS�%ie�FKK��Wb���xU͵2-��QY׋U����cY7|�"�PIH�|���t'�P�{����isc6<�KczixAi��d���!�H��	l�etz���h:-�e���lV��5��)�Naun��j����y�'?���BV�$�8�v���m���G�0��~��m�r5kc���q�YoŌ��������虵�Xl=sO��>y�[o���꫇���ѐ����-+���PN��(><;�}�)�=��i���1_��ˌ��h8�d �%r��5E�1�����+YV�V<ũZ-!-g
 n޼��R�����7^���~w��ޗ�>'���s�������	i��������Dq�4<6\�0�T�2!>�`�����C�M�\,�F#2.'Cv1���\����e�����0[���?��W^yv��xY7�rA϶\u��X�?!;�rrz<�_P��� ���Ŀ�g��~�dZdNU�u'2Z���g�Xșu��믿e�_��Ϙ���8�i!mC�s��9�"����Ͳ����	��F"Ј`E\ǌ����5���8_��%��,l25q����tja[ݘBK�t%pO�8Hد��+�����e�]7��x`���/��$[������l�'��t��-q�d�u�vPnG`o�Z����W�q1 ����¼Ϣj�Xao���L�w�,�QD�����vR7C�z۸#W�ԃ�Ĝa�)Yq��Wj"��tt��ݦJ���A��R��Ԏa��JfssR=�t���Y����Pg�ȞT{�{��+�$Ԏ�"#����!c�1	k�����f���x2b� �����.fb
�Z���u~<���~塔_����x��.�>SG��*�J}o�<���>�#έ�LL� }RO\�ⵉ�ʭ�Kۧ�WPD)L�'�F}Di��H�҈����.�^�z�X/��O@���/���u�6�c��~o��G�[݅�t�S�Y|Y�e��[X��T�o
�v�lu��w��^�5H��7vw��<m*���|&�_�de�8��O7�o����[���;�V3�eSqn�م��2Ĺg�e�
�sG��S%k����ϧ�������O�w�>����ܹ#�\]o�ɔ_5csq<���i���o"�~��!��_���ϟ+�ٻ�O�� -��������%^��x�&�ey���;��*�jm�r�����r�T'�ɓ'���F9��D��ܼ��^#��ӧ��������]�Z������|%��J�LmP���u�3Swn$K�����Kt�I7>�XT3�ySB��Db�x\�{�po21�B��2x�����]�4����mN�߼���}?�	�i8OIR�_�S��h�[C�x;Ό'�y���b���KT7G8]kT�R�q����^��C�4��D��|��i�c
�]�|v!Rڋ�.��s�>��������^}�N�[q_{�5�	ρ%e^�4H����B�+Gj �oEo�\���wYգ��4^ïh���ր���7��=��p�?��O��/�bwww���y|�_|���T�T�"G���N��f���hy�@u�C���l�U�m�`K�}���Yz~f�����o_7m����80��
�Y�+--2��������=��ŝ�S*?=Ñ�2+dZ������?���MA�|�*)���
魮��C��}�~�����f	�cg-��zZ�+������y�r�x]���X�3�ʜH��51�P8�!֗�jn��y���k����(-�4R����{2��e��w��h	^��KU��&8^�y��;	|:R �"�rg���MK�8��~�R!��d�v�K1�����.�>?�(�pG*�9,
&Š��^��퉔�W�^���7��E��eNG;��N����<Tfb�zFg$�����f�dp,��*ϕxl`���у���Āا�"7�݉c��G-�8�׉]�6�Q]�Q�d����1���W�j،�������5fHd4��*$��-�k��z�6}�r�}��)����uz�fmu�P�#���>e1[g )�.�8��Z��g۹v<ݛ�w}imm��9�g�������B�Y1J��P��ֱA��3�F�F�f)�������?#� ���u@��� E>��X�;պ"�=�y�`�QPK�K.�F˛��-�~||�!&�ݝ������[���#Mť�6��us�ŵk׶w^���B"Z��%a�	�QG����6���a�u�G4�]�GE<�;�1E�,oX�YH
lH�9�i|Y9��(ՠbz3K�oGc6�nn�Jcʇ�?Eml�Rk� �1�KE/R.�'�����n���,�?�����JJ�CIwk:��Cɣ�'!��⿰'�V�8_8�$1@d2���Z��4��r�qiU�RG@���T��I�L{	�����0%��&��ǌ�{�����kw�߿O�t0	�[��j��ۮ4"�	�ł�x{sKy���%�(N7ݐGk�&_3sss�9(���5�$<��`|�8�)%JDEF�#��Y���$94>��I
�����[��l����7���`ĳ3��.E��w�5Nn�G�x3~H�y�$R�����}�	�ig���y�x!�����!��,� �1�F����+x#N�/~�>jo޼ig��l��ڈ/��p��t�2'��!j��+�u�Jj��^��1�K}�|9�7l�:�a�RR��� B��o#\���ઊ�_��GAb?��U�����~��^y啿���Y��\���J�2�����2�]S_����ln*�A]-K��J����hD��:�X�>�S&���}�����GI��&�u0��+�S�RkE�t���Df[~G�x�r�����p���D�M��L��}��ٳ� �J�(�4�9:�<��0��ɞ��pc���_���JJ�ɀVFPE�	����h�K+$ub@Nj��j)+��I�*��Q+�Ce�dv���6��#��Hj`�h���1�P�&>CjK1��Uoo���+NZ���K"�-+��OS�%���Qzas���gG�����sB[��TC?��9��܊�ڸ8�#�/眩��n��K<�r9p:j�~�� S|.�<�Be�sW��y������#�b�#R��d �����tT݃�.�r��mb$��X.{*�K�L��e�O�t�r�'�%dbp�ȅ��)G_��Vb�y�g�5�(���t̊ޜ�dh쫶�����~x��g8�o����}��gx���ޏ��jp��e%$����!��N,ϺK���'7��oܸq~6/��[����������4�ED�����䗖��ŉ���>���vnb��]♲e|�a��t��/#?`M��)ƣqg�n�NR \���M�Kt���[�;���^����*3�/�ɲ!V�1
�3� �k�����O{��w���I������W!�~�:>����/��/�^��W����/��w���_��W�����x��21��9Ԏ�������#(ȝ��?����_'��ݻ
"��կa�X�b�ϑ�0�x~����(�r%�h9G�ƍ�9ô�5H�Ƚ��i��B�%�r�M|]AсTt�޲�wb��P�)8��(���.��	{q�l4U#���v����*e��	�!ݼb1?�=�I�c�OI�>���L����u�V����x��w���}짯��d,��n��'�a�:N��u�zƛK��p����O���������x? ǧ'���ޗ��K/�D��t>�)g��$D���{?=C��*�,Z�Ć�`��?�7B��-�P���
e�ėj%�ʎ�."������������WK�p���@+F�c��=�'�tx�{���"өq"��m��㺍߈a]��g-%�����ꆸ~��n��&:Jg�:�Y~�!s�]vO
��+�	Q�G��&�+�O&�|�X��ݩV%����op�����fc�-Dҝ���hD�+��:x��<b�B&8�v�9�¹K��l(g�Dn#�0T��6��w�۰��P!�$�r�kqz�q��8eO�<�Z�`�Y���͡��{��0I�p0rIC}�M_t��m��'�,����B� �,Z{ͣ�,�e��ji�Fvk��yk�"���;?�$�yHUž��%���Ģx�R��6�Ȼ�K�V��0u�f�~"���b��t�ZBq�O�	%�b?�E��29ݛ)}�B���gi�o��L6R�\$��ڸ������ gq�Z�:U�K�]�f���,Y�T���ǐ�8�z�X�<�4�]7"�d-,;?�X*���;Y%n�υR�6w)0K)�&���lrS�Mn��T[�.�ޗ��U!�R��x�3�O�x�1��<{�#��*����)b3?ys��J38�+���N�� �_c�IB=JR΀t@���d>���Y~�I��r�Tj�r�ɮô�Ge�>R����U�y�r��z`{?D��Y����S�#Wf�G�W/	^W�]�:T���/��j�#ÄW��A�/]�q�6)l��S������㍍�=�4��p��'�ЄGq�x7�{+�㴽X��ݺ���7_G\���e;X
WV�w���bV�3=�M��",�4B��-�+�t4����A�����i�T����l�8q(�m2@R�����L4�L!t籢����W h��]-���X�FG�,I�W�]�U��0�M:�|���OT��V�_s��bFRc֘�  a���:��U���i�%��>h7��>�@��"�i"�1���ҋ��F_��i�X��S�X�w�6�}{7�x��F������/t�K��l{�26ǧg��3��B�)GR]g����DY��HG\m�yJB1�ۤs
� 	W?��t�!�+l�ݷ_�uFC���>zq�����!��ɱ�&����H���z��kx���99z��oN&c\����Ν;���-؜�m��y��meg��
tew��i��6�x��If���m,|��S#6u��j��6ԉ��ϫ��svzqtxO��r(U�V?󍄩o'�[�7�g�*I&�5N7��qڠͶ�q�J>}�8+[;�����6Y��K�
ݔ��$�e.9=p"�\jggQ4>�Sf��`_�N����{{{�~���=����7��="1HS��x������}v������r�̗���l<fj��M�;W�*����n]��l�����69���+���L�}g�a� ��41#��;�"0��w�~vʤ^���#_V֙SUV�9c�H���"�7�NN��_�#>��E�e���3����W� ��S�r^���X��&��ON�)2�fz{uz���zX�p!�IT1�?fU�o��j����.�K�:����D�b��=��+j���*�n�lmmq����\fʔ+��]��f��#�Jy��둟�pD*�|p|ƵzqL�V[������fv:[J�o���]_�����Qn[��1$��ء_B��hs
-}�!��,v�YqO.�z5��1!�W�	����H݀�~qx
���deSe��c�:�/�`;��4 �SM6]�TLdMs�p[�͸��h��
	!��\���~��̢�V����J=���7BnQ�r��{�I`@�֍Te����A�(46B}U��,�`�dy*�IB��U�K8�`>Z,�D��ԏ)'J@�a�\�A�
`_�S׾a9��)[�'�k�X���[���3�D�@[�T�%2��$���υߴ�&�=�>�ƞ4��[2לV�**���Mp���Mu`p�z�ٓY��L�\}{�6!���u�$�$�_.ϼ@��"�����M�����r-"��j����B�)�˕��8���F�k�g��+�>�/�	��P���.�OO��Ul����@&R��h��%��B̢\|�q4�~���џ���KI��������BZ���/U{���#Yƍ���h�������'����>6I���P#����`��SY���_ǣ��~[^��'D���'����
٠H��]hm[)�f��e &���=Nn��:��:osuqN}5�>��NX��<S��K21�:�� 5sh�
I���j�k�K[W�����#t!�J_���_B+~<L�j��A��[Ӎ��\�^,���n�\��6�u�����x�Ų�l,�U�JgyT�(# R���� \�6C�c!�©�膬���c��
�`z��)�7�I�֚����tE@N�����??~���/�|��ٟ�ɟ����X-X���͞�}%{��&d4Z�:"M�ܪ�c�t��I����@��.��ԋ�Hש��S�g��B�Xߨ+�VH���_������\R������[ ��C�(x5�5��t:&�yIQ���A�M��k��	��d|5���^��r�|��[Or��W�����'cqVd:�Zv���g��rJ�ٳ0Sd.�F�9إ��R˛gd�^.ٺ�1Ջ������o�H]��l�V�3�q{�=��Ө&e;AJO���g���h�x'��S���nfn*t��)���h�s?�ծ�HH.�pZ���PN)�9/��J���}�{,�@z�4�.�"�G�g��s����+���N���z���ٵn@�7 I���ב��Z-�M�bMƚ&��]��,�������Cv�:`���(��e��Յn/xw��=��I���g�(d�B�O���>n�t6� bm.����S��EBfmx�<wｊF7jkyњF)����F���8TN�[c���}��Z�]�O5a��eG :靵�%��Y_�=aP����O|~K�=���JJƾ�<TC���~�����g��"�}��d���%Ժ��n@�z�u9�G"D�z^�_ɨ�qxpQ�ȗU�;�;���א��_�1���M�Ll<5;9��!VDD��c\Y_dc���Y		3��|ukUV-{ݮ'0>� �*V�^��&c�ݍ�DE*���
$��fk���+!%����jS*X����իWao��]߻}���&�>�̜xr~A�����pg��m-nx��4c�^"7]Ԧ�]\g弴�rk����n4�ȉ���Si�����:�L�j֏�u��B�N?�ʢ��SQ�Fq�G�$��Z'W��K
J���K�N|]_����@�d�L'"�@I�U<�8`�� 3~�_=┌6 �;Cׇ�5,���@�I�Z��8(~���X`x�uH�Q�R��SӰ������V��g��ׯ+�����'},����������B�Xpy�����5�V\<<](;+M��T�F	���������tsv��������sZ�,uOG��3�&����S�PE��r].-�E������>)'g�ul�4�n#V�[{�����<%~N�y�|	'X6<��N���r> �x�#Vj�2yt$fC%�e������$h�2Ǟ+��C�o.T'�\-��{P�y�]�2*,�ix�;��t~�=��b���6��+n�|v~l��Ʌ��ׯk����M������2���}�b��1�r2�3fJ����Ǳ�Cn���ʤ7%S�������]]X.r�@� 9=�A�9�a�)f��o�g*�rq)�'�g�~�r��>��՞�7߹s�?�$j�ĳg�'�v�(�����C.���,����kYMR��3kQ�Krr�Jc߻�U�(�,���|�E���)��(i�m�����zG'L�$��*9��w��)���������::a�(/�X���`�t/ܬ7���|.��>��/��`TG!ٶ�qL�Xo��%f��sjH�7.����ƍ��ؾ{�XV����3��憎��,,mR��h����p2�+�ec�g3�ɫ���w�)"��c��|�s�X.�xD�%��B�Y��_H�G$���oe�(KŬ��`�$*Pע�@PJ/�����UH�)�n���C�;���w��0�u�c�F�b�����٬�����މE����u4����Y�
L5Tj{�qR���Z@I������O���k�ߖ6�J������K��]M\	>��E�"�W��t��n��.��R�%8�x�+����V����&~�9�2�뿔�Q�K)?����[mB��z6%ɕR��`h��]�=�����q�_Ճ�J^��qܺ�1�S�6�!r9�Υ����Ĳ�T�7`^�w���I�%���s�:.�H<TJ��n�S'�Zm��<���:��9��	g(����������[o������_|q�^���_~��o}�O>7/��}2G�	����|?g^VLU��}����<�1�Q���fR濬Ih�Bp���Z��\��D��T�X� ��Z..�CZ{O\�M ��w��,&�޷�����X��YFA��H"=th�$`Pj�>Ȇ�T�g�g����y������Nu�����v�8�J�Cl�0+�U�j�|��-�XCF4J��1l�u�4J��N������g�m��gW廚~���6�Ix�Kw��R�ѿ�PǣcbSJ�<y���!�ݻw������J�9�mXA׶*��}�'nx��p���^�#��p��>��Q��0��R鸲��9�H����hAK���O�U������H�a<,��|����Zbp���x�������ÍGfR7�;-~�rx��Cu�������������CV)�)�O��|�ɓGO?��s��-ԥ��U��Ʉ`�z����ؘ���t��Q�@,[���g����&�UM�������Ek�&-c��D��W^K���g|8�,0U9��K��*�K����������g5`��w��B��ex{{�|Zz�+�i��;�]�:�V�2?.Y���ղi.�ԩ�O<�|=
��i�2�Oj��J0��i� Bi'�
~Wk�bu�`��D���ga���v��0���!	�)��c-�Ł����G[_����y�
�.\�ˢ�M�Rް.�����۰�T�i>�_U����h8���D#�F�F}�^�� 5�Τ��!�DYאƦX��[#3^�	SLb������5�|\TC���q�����'�z��-�=�/�����Q�;�P�F(�p�F�償��lB�98�(�>T�BX�9��fc:���:_b���6x�Z[ޭ�-R����jS2��2��6>C�E�=�[Q
(9�1��cGI?`�0���
���$��4�,��Qh�^��L�Q��%��Z�/(�u��\(��Ո�uY�Sn1�������4��=}�6P����&!��O �c:b����iS��"�;�{Z��^�~�W�������m�}�olo@~��"eb}<ae�蘘�ɈzvU���op�	�q&M,��=6<ɠZ��I=��ZnJ޳0�ZZ_^��N Z����{������1�(�[��M�k�s��*$bwo�Gn9��nk<������fE�P0�����
^��ÑGLw�\��lSO����C8�E4 �ǁ*~�~mvw:2J�fI�����F�J8�Q䩣�P�#���r4�G���H�i�EC�F�<^n���Cբ��.��=�Ŭ��	����-�%�QD��10vP.AԒ�k:��B!"�_�Tn�?SYG}Z�}�/J��"_B
��i���=���8���\�"������G5���#�P F�<T8ۧgǧ�'�*�nM�'���;�)��{��L6*�.ލٿ���F�S�Uv⨸��Hm�\���+�7;��<���� �M�۞�2�6|�ƁսM��򞝕��Y[��"�l��b93��|cs2�rP��S7"��"�K֡��O;�QnI�^��u�5*q�hy䓍)�K=�C�1 ��Y-W���:r�
�0����7��Ǉʭ��O�
ۛ�\�~�-�/Ñ����sg��R�3FZ�ȵ��3=�,���rV��w��W���ꭶQ7KAW�>[Wk�*
�[�xG1	��p���������ɦ�K���D�U�p�॑O�(�x��|�;x���&^l������K�w�G��m�������V,`�S=$\�����=�Cy�oZ,�z'����y�����*;�/����P�²oia�'g�F��&Tң�ݫD�5���k���*nW�nq�q>��ߘ�(須Eh2:g53&��dʶ��e�ŕ+Wmj'v��(W���nG^<G0�Z-�֯�\��?D$�x��'�?�۶��<;�Y�P�Ob����jsVɷ\U˲^�WrYu�fw���T��8(˭�3ޘn95~���3|׳g��·fr�`Mb0d�ups:���]�!�'�&R��X���*$�C�>A_���`��b�V�P��ڏ�}�W����O�!z�މ'œ�E9�����k���D�ޔ��}ն3���*CnB)�h}�����P+.oYc���KO-��RīLJ�����!H���B_�cLD�\@p8�"�w��f|0�-8�[Y���ުΩ��V|֧-W�!y��o.J�k;l��q��d���&�E�!��a�������c�Y������*��������Ζ�(I*Ѫ=��)}cü)��e�J�1Ld;؋�ϊ-���zsk��]���`b�����xD��_��d��Fa8��?%(�vխE������v��r^�uЇ���~��>z�����FTL��.�mG�K�bO^���������?���;[�O�>}��<�o�۶�$|�G�A�:��s��sTC,V��Ū� �1\��n��\m�����n�?9�ʙu6K42��A��Ǵ�y�������NS����[^��3�7��q�����T�V�@U;�@�@��J-�=����co=F!�FS?)K�l�Jq�_�R��EPAR�AU�SϾ����"����ۻ7oބ�a�"|�����6��j�^�+���T~P�^p �X��
-�|>̕,�d��
{i�z�#�.N�l��T�(ChO*/7Ur�ϛ8���	\.˓�3�b��Qg�{6����3�{rDt�|�?��*k�b�0��,�]N�u��*ɥ�(/���J}��b4\6������A]۰�FM3�����^�4!Tė�ޙy޴�~��X�?�W������O�ݻ�3'-$e�"�w���ٝ;w�]���g��)�I�J�nd�]��&+�k�4������Ȟ�"UԂ���{��?����k��距eH�&F�����$���X�sǟ��"ٔA�r�X~>�ȡ�D8�����-q��0�����mc-�q������Z��ERiL�5��Z�T%�e��21nH�G��#�ҳ�6�[K�!���k��,�.���TMwrv�����Μ�5l<���w�1?p!��ξ����P�K�L�$��)|�]�!�_�Z�L ������� �g��f�%~F�F7�f4
����^-c�*�b�tΚ�(s��pE�"���	R�����	?~"�*IR;!W2Z�'�k�_�U{^&�:���,@��I$K��ϟ;���ٴHp���U���R9>�����5��/��$���x��<���8�������;�[������lX�8rʪ:���kאz�oA�=c��f؀�[�!g���RT*����{�|w}�9Sc7Ov����<�z=�7˪�Ad�!�i��&���o�7֝j�����-̲��ȳ�q�E)�Y��JV\��QR��n� Ɂ�l�����8���S�G��NYǗ�����!�%ݚs%��p�^���Q��AQL�I�����	5D8�z��H3���Tɇ��+v��m��'//�=v9#�J�'O���y��w���ͭ	����ȪmnTKg}����$o�#ڵ��]Q�#�%B��2��A��z4�e�eE�&\2U��`�l�1E�����ONG��%�HWVx#�B�ϲ�㜛�OuWK6����ܐ-�詋�����F�ĩ�H�&9tMԏv�����7�K��B����-s���8P!��N��$ˢ�A鞜��#�V�<�ؾ!�q0���g�l����Yl���l�_�AZ�0N�«[�Q�s����*��r؍�.C3I	�
g���-�� $�"���������zS��F�&�=l�����3[��B���֤��Ȉ1^�%��T��2���:%M��T2���ʥ�H\��rUM3S��_���s+s6\m31	��r+})2<��rdm>�s5ʥ��k��,i91A]����h?�4��9�OMB./3�Gd��/���N'����kh+>�ht��� ��R�*�<�m3�M�ˍ��b#g�Q�LA����o���j�c�'e��#�d���B%�'�bB��d � Fc8��9���=Nj>�rL���ĺ�?s\�$ c�`iC�:���+W�,�gl�DTY��0n�4��;җ�\��%��>� 	��
(�Ѩ^�����E����.Oh*��#?p��l����,/fs-f�	OƦ]���!ԥʂ��oo���ɗ_~	a�z�O�p���L@$<�Z�����B���.m�����������4��^�:�^ݠ=��'�pw���g������g?�٣�}���|zva�@*��%$������
(�9���z�ˮ�\p��9gUk �,�4R�`�R_-ò�Y��/h�_�р��F�փ�,K�$J�H��*֜����:"�q�($�2��g�b���|�{��!{�À	b�2rFЮ����/�@��q�Y+�;����v�3�C3s�%�z�?�A���x ����H �@K�rz��4c��ކ��[�W.-;���/t��y�Y�z6����i�R��aa鮂	��AEh=�����Kl	��y����@�	��Rr�z�DW�������z(aZ*�~|�>�'O�  ��c�%��At� �IW�;G�(�3�'�G���Ooݺ�ֽ�aJ��Ç1p��S'�(��/�d��7�\׆5�
�(v��+@<��4�ϼk�������1�A�-l�K��&�RFN�8ρYғ,^,�6�'�qF�ee*�r���~�wy����� ���&/R�od�)n��� �|�44J��}x�R��U��Z�x�p+VT�pWHx�5�������H>g_����~����'��x��x"�0��N�!\b�Ɛ�����c�e�W&���0$��Й��!�d]����`��i�K*���cPՖ��Y 	DYu���vi $����i|�m�^4�:�ꤊk3ߕ�p:1@�ȹ�l�ex��ά��ۨp4L��#�8�v���fzj�y�J��_]M��� Ѓ�(�O���Zpt��ar��l�BI��@P#�T:��� ; ��ޙn��C����R�@&�f4"�w����~���*_���7o�_�����Mк���@��S0)]�v�hԍ��&V��Ǐ�	��F? ����G���,I8�v����+u>BW�+��rU��G?���}(=H��!��L��t�0E���{&f$8:���i2�Ej���S�s��N(�[ϝg���aڹ�������N��2N��'�K��)�j��e9ke����R'e�Ne���=c
p]��l�
�R0���	��;4�4g�L^m���+���2GX��)�0;�F��h:Ҟ<�8k&��{(uH/�4���#�DwG)�i�&A&�W��.>_.D�L[<E/n
�W ��Ð�ᧈ��d%�D�,��20�R�ڥ´L�kZ�%Yz"���ʱ]�d�I�7��.��ßU�@j��iM�r���{�uxG�LS�z'�F�N�@Ё@ �w��|�?�+�"h��A����}�t�\���p�||"�\�_�(�H�i�dRA���Uu!Bq,ˑ$�BhR��fީ�n�XU7p=y3%Y�����FG�X��4��m��>��w�����9���{-ǩ��,���㿈� �i�w��gKk��h��K�>�i��h�^�66�Z¦��5X�Y}X��`���&�k�yf)b�o���Z�G3�8��I^�͖��3V+�4�f9٦�_�v�q"�G%�W��C��=  <��������@�?ӳ@����ً�#�x&��q�L�E���R:��E!s$RQvl�W
 �%	y������V�{��ϸ{��7����}�k�;�++ �8��\\�Խ��9������j���jڽ���]��h��?���d��ʭ7>�kNN�im�rN����AbM['�ͬLq��(+
a�.&L^,{�"�Q,�z(|E2�4�s�C�d�_�h�	����P�%�J���(
��t��@��8�;x1pq6�c^���%:�#�2���yT�V��]������Ø�:��7�U�Xͽ�D($_v�y�o��^�YE�2t��:I�q��Hne�*�aDm'1gv�b���B�?����XQ�w;o/�K�hS#��J��,�#����{a�#C0����E��׵��U2 �^F��F�Zp����8�*���u�En��<xp�V��%�ipZ�I���䲟��8����;7o߾�9��.��p�_V`ԞOe5���$oK�E�6��ɋ鄽�|З9s	9�3� O��Jq]��-��8/qM�}�������䮑�]GQ��s��֪f����K���ѡB�S����SV,�[�, ����.dh��">�5�5�ߌ���g�i#T�Tus7g��9	�h�9�bg�QMůYήH��v��i9_L�W�d�J��s�t?�"���E���v��F�-{�﬌�V?ιU@�&��Ck��ɧ>��#nb���h���a��rŽYv��N;pZ�䄾_��|{���pD~-�/z����L���}�ѪX �8r)rg<Z,&���<84�H�X#�M�b��_�gK���hܕK��vuQ���=x
���x��<raD]@���YNe ��i�0�H&�K�q��f��S@��R������u��3��3�vrY�������g�j~zr<���Ѡ�*���*����Q�}���Llk�e,fݵ�����`؟�'����"0COe��KZrdz����:�W\e�g|��o}�����?���˿��?���'�EG�<��>yy|5��^.���ώ�o����w;Fli�>wMe�<*�`(xX�{6����A~��gS��H8���`��Em�&P�8,v�ڶ2u�]��^��H�����]@��p�\���峫YN%�E\�U�a�F�)��B���gX�?(��DH��6��:����?�P+����i-��>2,�y��1��=֡�X^�AF���8 ��Cc@�y}D�h9�L14a6v^&�����u���$A�
��&n�8��d���e9"6�^�x6�9��GHC�0k+���@�\S��
9�	��WFȷB� cB��Ie���3'
�j8ei��P�[)ڒ=I*�d�H��x�I�[������;��Aڌ�����4Nz�Qt~qE�}�t^��j�Z������ǟ|J����}6_�`wQ����T!ʂx@l���X�9�~s||��+���^�U{�#���k��Ʒ�O�>��o~�����M�=�~�!���qm�s�_ی���
D`�͂e������gO���JK���AfAm� �%J��E�]���b�����s9��0�`�sa
�۷�強R2�	i}}|�������>x� 5����+�˶�`V�)��X'L� &�R���Eb�������A�:�,��E��/����}�^��R�˂�3s4tT��Ƚ;f�NDG�9�{���V�0\�,8e�?��V��ӓ�vLp���,2�i�.*�UT�Y	*�,+=T�c��3_�-$��ز����ҫ�~US?{��v�^�����N�}��YO�<�?ϱF�X��b	��	, �������@g�$�D�>��n�3����Ny�:b&��v]����>�J|��$=�[��jO�<�:m�H�BJ��B���B��+G7o�d,[�S,���u�3Ky>����|�G��ǖb�:��^&K�ᶑ��x�0�<��Gf��"XX�(
��՟-I���q��ޝ��rK��Y��"O�<mv|����b�9��ϰ��p;�⮍�h�Y� 	>�q �@�qi$I�,ob�T�L��6S`�so�N����x�d�X��7�z��,�^�G/#����~T���R��}F:@��GG��
�3��)?���(��ҚNKP�p`2j:��4�
��n*&�"��/cO<��k��d �)|[yY=6I�ґ�w�)!	��	D߀|�C�����R5�RP�sAkuB�A�M��Q���装	f��d���C�"59�u�n�n���i!�̊�ŷ��`eV�`� 8��m~�^
��S���w��z l#�����׀>����Rm*�V��n`�7Qo�N2�Ѵ��j�_i`�X�9���hZ�Q��Z��6:J�5�e��-a��Rto��Ƥv����-�hY?�y�_I��z^�rfK�Ȋ?`S�ͤ��p`���:����^|0u.�$G#z7�5	�Z�:�T`�0M/<�WP)�Ƈ��Pكp��f���34�N>�,`�{Q�F,�5�jV�|��o�'_�9	�ko�Cְ�, rn��˿�˿����s�~2����}��`9�oZζ��9S�}��]��vv�޽������eb��^.�F��3`�Կ�v�cO�Y8Y����g�.X0n��$cp�p�\����c��.
-ޭ���N����^8���%PB�zx�!����J�����QKΞԼ�!�+�ېq�g89�v�Wn�r����)\K/g�V�m 2,���X��3�
��Jt��(t����L�F*m���I��2�*�,|��ѣ�S�7eDrH��06L\�:�)1��,֟y?LT$���\����HU΃5$�D���D���#/��9��خ��4	V8Wn&�"C��q��S��R���1y���ԯ@;�p��)�9/Q���ʞd�:�}�儧�,�|j����a@N6�C��߰_bv��#�8���W����������_���e��8|�����=��m�G�z@���H���/�ՙ���xĤ����nA<5�δ����5�6*�06a>�X�L?���.�bXʩ?;?��@��u(@\��5$#��bU/o�/O8��x��@�Q�I�ȗ�.0�
�Dޱ����M�������(ə��4����>�=r�I_���-���ɜ����[�; �5���a���`�p���nE�3�#GjRX�����F-陝���"W,3�m��5r�YS�n�޻{�*fH|̈́H�YU6	<^���׳ˡ��ZK��5����.h~�����;�����t�a&]h��3�g�P�e=,S���ّk��RKH�����<��	7�S �<�qTCKqx���⷟��'��������ؒ�=��W��,us�q'<�pB��Ů���®�F�����o�o���x`ZONN�֕Ŝ�N�'��~�EI���[j����#e� �衩��6"} Q��XQ�b��W��Z�
@-�:�g
`\,C�WC $������ϟ"13tO�<*�� ��@Xt�S}�uB��47�k��2Vr'P�J�-�Yy_�p�hyd��;�\�2��`+�qW����C��Z�>`����_{�58���Q�������������
L��z�H�)<�i2W#�`�Hwʓ�O��s@�V�����i`�	�����Gā/�~O����3Rw�&���r.3u�lVV����<$o�����/��Y1]���p�˗/_�x�M��7�D��I�6�ς�c'�t+3�؉������0���7�� �3�t���7Ft�ޭ[��Ղ��ݾ��;�bA�� 
_���Bٖ)v��QB��^B��6��$���0ċp��rK��\�pV%�;dC�\�r^��}$k`�2!8� �=Z���0�lgi-iml����/h͞>}����?��!��k�BPf��ӼF��i��k� ����V)D�Ƙ��-�eHΎ	��m8==��߳\O����Tb2(�L�FȲ�ݡu�IV��heL5F��C��+�;\k�HG�#�B�6
���nQ�H�,\l��$Y<`�D
�B���G��z��E.|��N�?4�n޼I�@�`r��͐7�@���8� ��g`Ҟl� }�
�����y\�K�x�1�ʢ�(�Sz}�>?��������:��g�J��S�VUt�tC�X�^ʞ^��U��L�MjA}�{�D�{�� �Dj��2p�_6�'����߹6���O�c�4M,����f�+��7�~�q�	��V�	D]|xދ8��Xvh{�Q1}P%�E�HK"�#�HH�G�-�-�{}>��[@�7���y�'����3섉Tz+�I���L�(%�I�Zc�W�1������.�bF�T�Q���#�r����n��밂V\e�|�Q���u>�+D&�NS�1�ջ�Ne����=�2]*K�ĳ��ڲ
L�@P�"C�w`pR� s�+Ϧ�r�Cs�{��U�E�}.��-|	I�st\�`dz�Hg�վ�)���t�����傮I�i{�D;��%.�3rZ��6\|���u���g��eys���\��f��Lն�i΁�n��FKҙ���Q�hu���4���?�BƤѩ�N���y"^��i�>
)vlp��Nl_����u ���iE&��G-=h�v����~1�)m���=+�,��Q*�?��x�F��$c'Ct+͎�<�d���
�<�*;�wP�z`��A
���JZF8�[��[JC����`q�D�	 K��ҭ���,�{��������y�p[o��uY��]��1�B�ʆ���k׎�_�A�=����X������ųL�� ��I�(-�'���y�,��8���/��A����(��;�"K(��Gul.Jp��X��~G\h�g\��2=�U��
�S�p�']f��\|g+�zp4b���|&����m�����GKĆ9�fZ�Œ�A#��JZ�h�aLe�3���Y��<@����kʺ���_}��<k�����$�j1�.N�$]��..gt��[l 7�C
@�m]�P�?@��1#��V��r)��s��.�b������8R4M��G �d�O�lJ�W��6P=�<T�F0;��`���BCG'h=t"�$G�ġ�P �`�,��1AnB��=�� �m����3AaS�A����Ѫ��+*�0�g
R�N3��q���W�G�;�jzЏ��yC,+��d^���U���K/���0N$�H_TeMvQPչ��������I�/)�6����e[sm�le����:$t�P� �c�����Ͽ���"�x5���*��ݵ��N&Q�2��.�\0�Y��<9��f�W�pN��X,�[��Y,V�%
�耲�������s�c>��1!��k�����cx��*9Ο�9�����p8���i�(�]����"�$}����r��Q�7�.��l.^WH�!𦧈jU�FZ�q3�\^��
���$Ƀ�W&���Esf$�}��������r)-�Rﹺ�x��G�s��؏���V�J&i&�`xl\��ՠ�(����b�$�eQ����g|�����Eɨ�<�\M����@��쒄<�|�y.e���n�����|��׻�3"��shWi�}RĝL��螟����<_?����O�p�]������hՂ �>
A��S�,/��Gx5�ұ[�̣�����?y��Q�s~W@'�*/�T�?j˨�"m����н��*���u�#A㍆e$}0��2����,�h���f�,y��L�dz8�h�֒M�
7�����cwn�괙#R�q(��h�(����T��d;�ULh	�EvQܰ0qŢb��F[��G��V��:�
6.�`����^�5��L�f�Ѳ�l:[��k�d��P�̂HJ|��ý�m�2? {��S��w��:��4���cݔ�P�DB�*,���2���j��E^�҂�y���(��d��9o��gǿ��w������V�����O��������W����׏n��eyWw�?-������bvzvQ��tv�����tL�劑m.����Ʀ�w�!���a���,j��i���L�'��O?�{��O��a�''g�����������n��{�dq(��@r���#+���wMd\O�Z1�[+��-w��qZr�5&�%��۽w�]V�dV��XRF�h�=��Z��-(㞎��[a� �{�<��n���u5���|&��߿vJ��u���ɓ'��_.W�Ŝ'��um7�
��D��F:�;a��R��
,��2�y��R�8e��t�b�}t&�ɇ����e��ɳ�]�7]��ä� �\����Zan�fT0IgV��x�eH��Sv�>Ic����|k��$ �4lI6��Sϝr�+P�G
��� �Yu���8���#����-Wȋ�fX[U��d6�~�m����w�y����>���͛hb��WӉ!c �X�(tm{���3�t��f2�#g�4�-�{��^_�"��{�i
/ƺY�����_����~����N��>;��tZpr��Q<z��*��e��(g��>��ฏ�@N.i6q���*��d
G#pZ":5>$9�0�K;��bYqD+� ����T7����B�����봍�ɥ���u���x��|?��3��3�'�Bpq`jb��Ia��h��&f�4��u:C���^��你Ĝrnb2�唒������J+m�ԗ��g�������9������
�^�k:�q_�~G�F"T���j�,����S�i�D�F:�+QtK�s���ZN�񉚃��H��vX쯴GdI�/��ӄ"��'�?���=�'�����ɘ6,Ha��4k8O(M�.�2��lecM9B�״�ΒB�+���R !;(=�GC�G�D܈��R����tx��HsPO�8���g�-u��:s�Ul��]�9� �p�Ph�;��ځ�$Q�g�)(��BIM�ąa�<�T���m$:}�sJ��OkQ�4i�#���R�1���v:�h�o�7�pc%@�u����z <�Rdn�@C����le;��֚�z�y��Q2l;������r�4�#�o��*Q�#�8�uk��a+E��y����V!�d�yog�".���Eխ���p�ecpugQEa�e��̱ �=8�Xc.l����*a��lP�rttD��:���Ռ�D�<�IFD��D��<��xs�̈́���p@1�r~A���u��S|uĘ/�R���o����5䏐WE�,L����Q��=�|���>U��K���}^�wa��5.�@�
�@�T�^�bT��_��uȘӲ?����ڣ|�$��\�{	���VWRa,���ޠg*GxK�[���X �pMp�޵�$(�'��5��/��-%#�41����s����j��� �a(Wd�n�&yEV��<��Q��h6��r�{��l Pϕ,U��@��4��C��{��!�ҭ�ٻ�P�Fܹ��خDmPPl�,�X���/� �Ov�I*�"]�;�Ip�Dc¢��&9��d*Y{�xy�$�[a_FU#K��9�3�<�A ����h����J���mQ\mA��7���o` �h=��6����=����O���g����Bo��u���8?�	�W��V��t:�FJ�mj���{�v5��{�GL�cZ���{ѽ�r-����?{~�]�#n=���h��];}�,�V/3I�}���=S^�>��@:��TQI��G_�p�HE*��l�B�qO����r%tB>p��XV�UZsjuA	B�E�$_��򙕳IW���907��r��C�͙h�\��e>b=��z��|b��G����n_�����x�d�����,9��|t�WrFB������j6�3E� ����y�77-��0t��o4=��@"x�]Ho�H�~��������O��98���Ō-Əv���:���~��+jƉT��J�0�c07���C�>}*�Z�N�2�S؋l%���o�0 ����R m�@�@G!݆�kk���mh/h�7�|�t��{�j1�:�`�W���������D��"���c��,[/��0�N�`�����h�G	o�1��Pv+;��L\�V[��=)� ��("�K:�!6�OK<�jW��_5JJcz������<@k@a?��ҎH򽆖x��9]�~���������J�����)��$K盩���x�I� �e��L�ה�ۀ�A�Z�c����?��#mD�����e1�������
h&z���ٓ'O�w�o��v�1ҽ��Hj��ݻqY8`.�F����oQlv�v|�s3�h�cFn!]��쌾�y��>v��.:�7n��ӱ�K�^�v-L��{����Ǿ��o�z���/y�e�.Z;1�4���[�w���\#�41/m�d,�>p�+G�0$tJ�i��	���Hf:����#��5[.$ka��q讠�?��g���7+~P𖂷�s�&k��Tl��ä���	���8h�}*h�Z�ʬ�}��њܾ}�~yu9�ba��C�]��5t��Ӑz���&@Y�K(���ƅ:ʅ1��7*�����1�N�{����^���3���`���H�U��Gn��boo�R<V?X�� �Cɐ��&�V�u���j)����!����@/�m�@�|�E����`��݌�JaS@��?M��~����0�_�u��%�,i`�"�D�(�Xh����?�o�����j�2��PZˑ�s����k��F�N&�|�)/��8)rb��:t�$�)�@W���O/~�ߘم*��e'������-^V�(4�{��P-F\C����{w���l��ŋ󋳿������m�0�Q�0��z��}�NX«	�����d�L��H$(,E$�R�tp9�j�=U`��4ɋ���r�9�S1����j��SH}")����V��A��$~�!XsT,��.��#�k��`60��\�reښ[뀙E��cr���LM�_��PD�$�������kgF��ˇ��p������E�O8�U����Ho���|�h(��$��!��6iᨴ�9���]�	f��,�!(2�1aR�i�y��h<�����5�K	����
a%�O:[�̓�4���<J�~�KM���W!|^�h��F�����f��I�h��7�I�h�!�����FB�z���Z!#�Ќu&�=��y(��Z�3ymlD�s�˥����2[���!�l�)n�)(��1W�i���b�rd6J�/N�3��=M!�,=�����9t���b�,c
�j��N���z��I${h=���y��	�M����:�_s>Zm͆��
���) �$n 9��[����N���|gg���O�s�'�͆���竲r�!iҭy�5��G>����h@&�k,Y���/yBb&�Ժ������y�c:%r.�;ۇ�<+V݃��^�5m�����qg3���t�wi�v��
�۴���`��j�+��x��K93����\��Y>h;��iĠ60��l�U�'�o",�H��b6m�1	LJZ:����W�{�Tr$��-7h���B�U*��
�}�طU�䀵
ݲ�
!���C�%��HNP�4B6�wl#w�����+�w��v.�Z��J�Y��Ò��LOʭ[臭���$�e�Ц���</��9�:_w�k���^ҧ,
�*���1OZǥ=�VdU���.�l9�MQ�UKV�kC� ��Xl!�Nbq0�P���^]^�r�)$r�ƚE�;9	n����
t�X,���$�����
%�1s�HL�0���������)|�іC�]�N��ZG�F-�2ÃtG���uP˙t����sۭV���%��x�@ZQPI�y�}
���P�]mAa�V�.�XzX�K}�F�am��H#�g|���f�@V�_�Q

J��B5/�|1�ES��G�.�a��&�X!� �#a���l�!I��^B>��0��ԥt��t)�+�L�����qH�CB�르��F� I9|j����lѺ�&�#	�)�SCC_�9<��L��y����E�ј�4c�N~�Ah����6N%���w	�@z���7��?x�����m�,� u��	�93�D1�R����s�����P�
ɀD�dEYe�#I�xg���%o;>_�6�,�ǒ���X$e�$�%;�ˋ�͖��b�;���[��
�@l2�26s����♜W�{�>�xpȶ,�eBb5+��q��8�n�s6K@�Q!�,v�:���!�"O���g/������xry������P��Ǒh=�wE��H�7�cXWdܓ��u����ڍ?}��g�3c�"9�0�+}w̒�ԅ�\���p�&pj3Q��,F)y�U�\E�K�5ކG1'�yU��py���q��7]h�Õ���:c��\y�I �p��{�t�.:�t�3�a�|����*0Ĺ *��8��U�C9,A���9B��u2��թkX"�O�C�Њ�V�h�r[� h#��7hsav+�74���^G�
̔tB�]�.T�R%��jG%����i�`%a�M$'#��EF�xqq�����[�U��1��f�ˊ�{\����$us_vGG��Ɇ�d�j�4X�·x�0q���)o���̲�xHܶ�;k�����Z:[�G,+Ɇt�3@wC����T��$�zc�����iOO�>��7��?��ڥ%H��\0�F�s���jJz>����[㝝�����)}4:��_;�S�v~~�՗���6�F;G7nR����Y��;�	h��x404�?!�����aG"V�hQ���򗿤�O�4ۧ������J��B��D����k���-~��wIם���߄x /Fǁ�����	����m�`,�LC����ȵ�h1���
珈��n�W\���H�ip�u8�,��b�@�����=~���A?��� ׎^3���Q^�"M|ہ���=.$�C@'7�cI���o-��a��$Lz�7nܺu�~s�?�>�[��V-��`8������1���}V_8��M�}�g�i������
�ȓ�EO����`z9V�ۘ��;7���,,;�Ǥ��GH'����{���7i�/&W������"�R���`�n$�Ip����>���_��͛75/�գG��� ;����0m2o��Fg[�U40�BN&�X;�$ds �񉗱�p�eQX�����jۿ�կh�������+��ٓ/���ųg�p��G�c���P���/��Ǥ�r��n)�Y�.b�6��	�"Z�HG&��ӧO//'�US3�f�lg��>9kc�k�h��!��0)G쪢f+J:(��b�������o>tYKQj�5�c����]$��=������	�,6�%�2�y����R��t�Mts�5<��o�t�B�P\K�l��%��J�Yt�(���ד�I�:�ra~ı�|���N��:N�W�2�&H�����"RʵT�����:�g��9��m�;6FR7�K�T��r�V���ʮ��=0%c9�]�q�"��nR���Hh^8(���6V�	Ql���������OQ�@�(���x�AB�j��S�k�'�E�{��	I2}"X����_O@_�^������ݛi,�+���?�ѶY3�.�V�Bd~'l �%3����E��\ݐ�л2�5O������r��L�;�f��&l�7����A�v��[+M��3�2k�Ib_�!+���@!kh��h㺥Y�ˮ�f-1�y�*D#���f�(L�D,$	54~�.��#Ez��#[(�mW��ϕ�;M��c��%�(�-	Y?�Gb&-�6���y/��oDOG�Z�}������T Y�7ߺwttD���C8Opa�3F��ģ�ۡ3��x�����(�e(v��ӑf�Z���t��ա����u6LS�:e�L��eB��X����}���A��NU���vR��(�C�c"$� ��\ 6"�T��[��#RvO@��J��$:%�#�����h�J�A2����!LEL+�P�5 Yqj���D^m�h, �� ��`���,��mI��G�"E
��IR~\�Dċ�L�����}��.�p��e���@h�v��J��O����i5�zT�!� +%v�0��G\7>���(T�ⱕ��`-D1�ۮ	p�LGnY%��IjXa�؀���C�=�ѳ`��Ք��;��X���O�����o;-3�w��6���v��T������)V!����u2�=�'�)�h��P`JfW�u�B�1�F��i���qKo�2L'���&�a�D�%Ǔ��>POH��8X��%������=�E/ ��Za5H��A	w%�P���Y�?~����n���*U}���	"+����vb4KFx�����������~��R�.¡06���rtmE���~ ��+��F4�ܤ�Ը��o��x	;���i��P�(����������|:a��@��$�dM�AT�*{��zܷ%�pq���;ߑ������Cn�M"��`�L�>E#�]�􏟁,���ʊ�2��e�U��4L[R�F4�UD
AR�B��_u��'j�Qh�r���V�2&©�����r��3w:�^	������H��(���Ԡ����L�n"�mt�D��?�P�Tb�:Ю�a��,�i��Ʉ���m�#j����rF��4��^k�V��
����ۄ�Q��$<���{H��xvZxɂ���l4�� ք��(�� �C�e�2�>Π�!͑��%2�m�V�x@��p
|�Y �o��[��E�9����[�V_���'���S��Ӳ7��|�J�d�yBV����t���'#Y2a�����8��l�����H3��ٳF���)v�޺~��x8�ַ�u������?�;w>��ڰ�I��C���u�	6$���t�����O~���K*PXJ�t�:g���y�n!`$�<���-C�o�Z���rK��'v�I�k8��k�! ���m
�m���V�y2�m_K?����p��S���|�����'�d�%���<R�̍����Ԉ�L2����M:��q��W�z4b?�v\H�C�Q�{'#v�ֺ��{
.��Q�R4�9����ҳtM�ȋ� ��I�8&���3��؈�ɥ<�. fk#!Ș�g��X�g� �� uH��6����_��͛7�+����z��N���Y��w�;&�o�bz��G�z������)�Rs5:Bӂ4�4��l�?���W���be�Y0��BV���V�bC�x{����_�<y�]��٥_��u�#�meJ�F�!�y:�"���w�E�kkt�����l�W&���!FtY!X!j&�O7���3	�LK*��zҺ�f���'GZ}�o��,W�#�1D��������e�k^�-�^}v�c�tk��t����d�4���RH�D�7L�wf�cM��8KrY���.G��ڴq�(p��M#�������������91i1�,��k� ��6�`���Ny����M͌� v�;orX��5Y�p%�e���M��nT+R�;�ܳL�o�fb88"l�9���C��=Ux@�4�6:2�s���\k�&��azͨ����礄��;)�Ft''ǒ�"�
8���a~��I|����g�@Sd0���Zԭ�+�WB5�aE��-h�iԶ	�|��X���d�7X*���Wv�)*��L�Xp3x3$���D1��K��N�]���E��g�[$R��t`�-�׆�y�l��S�#�T#����&x@��W�R�w�d2[�.�a�!��<��S2r�خ�R���V ��yi,��ӎѴ���TH� �<8CDړ�����ё4Xy[IKm�5�ϵ�eփ'�s�%C�A��q�%�����{����'��szEҠNF_�<�����o��@z���jww�����^�+dDg��蹐%ӓ���q\Ym�Z�t>���<[���,
��{7�L���%ߑ6a���s�L�95�z��}��Ҳ�"ZK��= ��<���\��T�jY0+�r9�Ǖ��q}7�NZ �*Q�
kϡHb9_�`n��E�b�#���ȅ�w!4N��ȣ����2Ƈܾ��G������^.ı��9G�cj}Fk���7��;�'漍�ʳ�Jp�dk*����:OZ��k}|'��g�p��Z��0G����!���Y�)��Ƞ���I��6dl�J��S*1y������{�4��zSab�I�)(����7�D8?��n�ߨ�d=N�dJ��:�$��;��8ѵ�2�[��U'(*R�شd1�mG�>1�&z�`�h��N�������	}(�=�KZGb��|�v����b>_�<&�.�I%�s.�֑��ꑔ&_��<���7U��_��K!0!`n/�AS݈�eu{\�̨�{�YT���(�],,Q�db8ט%��hL�I[@Ƒ3�]-^BiL�tj6��A�e���-�*_B���\Nx�@��ɝ� F�?`�eɏ��tvm�ZҩIv��U�|�M>���t��l/�Z����[aL���v��ב��c����9����Nk;w��W������ �`# �
$<(tA�"��#p a�I�\),1l1�Jț�⮗��%�ɞ���e�MmS�iq��P]��.����ʢ�D&�'B�,�k%�*���0u��y;�suQ.V%����D�h�	⍝/y:
�3�$tҋ-y�N�L9�
9�@�2��&'�[�UQ1�h��G������?x|��������4'^�`����#��í^�����?;=}v|�5>�#������ӧ�Oa&φɢH7e<�!f����ĳ�4�>�"��ݸq������[�cL�Ceiv�0A�ׇ�e a�+�(Υ(J_s����>��js`�F�2�8��iԍ��N�� K��duݺ� 9��M�P%�g5�l��E#XF+�A�Q>�(���1Z��	��y,�E����N܉�v�|eԊ����͔*C�R_l��H�Bx#oRb��1d=>Nz���� ᩡb( OQ�*�z�T�r1!�=:�����������U�zI,��2��I��P6K��n�Z�+��&��"K��N[��
n�i	��mv��
q��"xz�:�gȳt ��t�p�cJ_��]{~yA�C��|P��dU�*�ɂ�/���}u��r�n����F�ދ/���e)�(�t��f�h��ظT:'
��='
DH7���e���h�F�Gk���������}҂9�eI��z������vHo5��.tP��mO��`���*k���ϒ�ƭ�Y�x�N*�׏e�g�⳼/H|��J��y�<i�`]\�\U$��P��h������䓦�e����ď�Q]�ӂ�&�V�BJHxu��)�jK���ۿ}����R�;�'''H��'�����������Oئ�`��9��,�5l�Y)�=9�>n�%�:Ӥ�#���^�|yvv����/�?�Ғg�D�p�ʘ�c�
��W%�:�����xM�F��)�P��<�y�dr�9>�@��wx�e�ba�0��R�N��a&�c��Ŋg��R�H�H�6����_VJ��7Ɔ �n�W NA�`!��\p,��Zf�������T��� �G�HC�k�3�~��'��'�ÿ��D�fo��N��<(V�I��.O_<;��Nf����6UҞ�kL^L71#���!�t����+��r��2y�N��_}�է���n�骘�B&u�P��F��U��d��q��Ǣ��d�G�̋���W�i'ɨ�\7XU;�ۀ=�!�<�[�vB5!�F���z����F9�zȉ���%��9Cԝ�ݖ��/e�{q]u�ܐgӗ�S�`ڮfSrPQ�|v
a��넝	Ʀ��iy�_�j�6�vO�<h�V��F�=W@��ɍ�9j~��Y��c�Ȍ�C��i�П)s#Vԇ*l���`�↓�聨�[\�۠��|8�,`�����1�Iq@�2f���V5��e`TN�ͳ�H�'��%in[�H�I�
�J`���	�i7s�4��7��<$˭Z�qm4	mi�?��B�Z�V�R�F��"ޢ��L6�Sc����K�a=�m0&
�s��§X`����6��c-�K���t9�b��K�bc��LIj�Yp�r� �4A�y>�)5T6�+K"ciRu �z&�0;��*�-�"�������NX���e��l�Æ���7o���_}�����)Z���6� !��)	L4�9�a<�}"������G���?�яHe�գ��������_~�?���#s��LYM�`�`������|�	<�8����M>�tqU�b���D��9�=�Z "�p�c��N|W@)X�ϲ�b��n�����l��q�i�%`���F�rER�#B�*�Gz<;�l��
�B�a�ga����N�q�ѱ=�o��f��po-�i���SN;M����)��*$6��]rx�C*��0��`�σ7�B�Gn9��\L� ��jl��b�u�0w��B#6�[��[�29����H� ,ٙ&96��^�;C5u6L�3g��x> ͨ˦����I-�!L���`8��� ���! v[Er��hj�!�,����B�-���:_%:���7<�t�s,�*� �"H��zI�ख़�+#�0Ph�2U���Ϩ-+��N��S̹�$,��f�WWW6^&Wf"��Юt}�%�ϊ`X�8V�Y� ���)NM2��b��`p�`KG��O�D:D�&`��C#S��o �nI.��C�œއ��i'�0��c񍈍���p����;�mȄ���j.�~z�3���3z^0�-W�������n`gk��҅�K�+^�t���v������U�µv���V�G�;�:��p�Eȶ�������ý}��r���tz�l�h%H�eƜ�9����
�1�JaT���G9���$S�W8��Ĕ�u�	i�Jy�Vf[52�7
��1R]L�(Usr�$N��_���\�T�M).��Z ;���V��r�=B�t��S�����k׮��X��+�'� ���ێ~C�J҅<��LރOɟދM�IH���zqQU#���^�5P�y� �#��bƜ���ʙ?TLLYH��Ќ��v��d�8��^��f�&�L�L72%��l�����bc�EZ�6д�Ѻjf:2FvJ�����|!��<͐�6�_Tr�p��g[�1Sn{3�f(A��갂 �rX�ٴLa��}H���{�	.yZE੽P_y��d:'���~���t��Ly~+�秥�G���'G2��E�R���X�9_V8���X#���޻wo1�d��o��O��O/_r��rUH	��gO����*��X@!��6�T��nM�i��^�IM\��N�T�%�,�M����X���G(�쿑M�?�u=�?�qϴ/_�<���އ��׋�S�_��+�.�����X���_x����������E��%�:�e��J���R�1@3���r_���s�����~�;:GtĂl��c��ʦ��Yi�X����m���p�!smY�VA[�L�H$Q �ȟh���Z��g��a�ɗ_��>�"�� h��QR�䘸sp����Y�n��~�bPɂ�����G��=~�駟|�	�$-��'O���f�-?�
� ?�*ua�#I�\z��ې�Hݮ�������8����WWS���w,>�~��k�Ҧ�2	���U\��$x��/���ɷr�k�����Ig�1and� o[�۔H
�ہWEf�'H�����s��|�NR�P'''�:`k��iOSb�	�����O���N2�ĭ�;�S7�ZcE�BT2%�l6� �� ���?��e���U��"G������ �a#�vwq��G}Ĺ�G�Wwi0 �Pl�!teƏ2W�|2����=�<�r|��'=�G��d�P���p��2�Tv˵Z�n�U��~�儋L3���(��e�P��
ڻF���y�I����"�88��rSKu8w]���a��J���z��y�Ye�Q��\Pc��<��CC ��6������N���4�ENrٙ6>Z���x����,�f�]��Y��?���2.�K��j�&��(�*f��#cᔾ[f�Y@��h#�I4�x.f���#��G�����7bX���&!�І��*����h< i�3�i�kޛ��{1��xy<�O_��`����>��U��̦�نñofuQc��]G�H?��w��fe�C�m��=���<�nI�&m��e������O3%�LuL��'N�L��U���s�s9�P*M�k�*"P���7�#�F�6�,���V,�	�T�%���ĉ�S�K`2v.��I�Ճ_����uH$�w�%B:���hsX�˖��u4O�-E��C����\�6��m����ˋc�`�ж�j����~A٭q��������M��u7��׽$�5�����W-��ݼycgwL��֭[��U��ּ=Lm����r�8�����Uӭd�I��j�J��he�a���d)Y���u���~���o\���>��#�}آ#��o?I����?��A/��ۧu�~���?n�}�����W����US}~D����\϶��8�OV@lE�=�ϚM�V�^���3$����װGPt8C�8�,�&�ˢQfSm���0U
w�-8w<��J�n8h�qGɪ�&3X��.2�B��kz�7np� �A�V��Y�� �:������X$)▨��mß�<啇D��4M%�d�
��:��D�SI�,!B�F|���R�.���������P�|"o~mo�nU^|yq1;>����A@*���aU�@�)�t5��������R��-�ӆZ4��y4!%W+�
�`�s]o1o-h�a��������wܪ��/�/���t؀[����&���G�>k{8F���4��X�6�� �����a-O�o$�b,�'S�X3�4�
ك��"ZM�O���:���bA����/xV#�Y(/�>��Z�xUu �d�8�v�������_M9�̓ޘ�/!m0�O�.��O�#Vɨ%�������d�ޮ�h���/�%!�ikk@�3��ȓ�
��Ǚ�n���=�-gof:[zGG$��W���V�T���j%�b3��Ŏ����<��O��\U;���j���D�ruz�����pgw��>���!�Gq�U�v��o�A�Grܦyڦ[�0� 5X��d�|�$�<
M���"p^�Nڴ�c����X��P���_��t*w1*���w�`RpT��+�#͝h���FO�z�NfSȳ��(.it,��Iɉ͘��I�y�~1C"�q�]"L������
�⢎˪�xx��I~*��ը:��Й��E�*���ɠ���)+�i+�߶~�;�	�����{:(6&�E�I�+�\�#������f>�'��]�Z���Z��ur|rvz�渦�ϙ����\�u< ͑���-�l�����D�A���^?~��L�9���Ѫ�7-�&�w�}���d�J�x0��fV]�u�3��b f�<!G&��./��ae�t��mM�2;��"{���)!������+���'HO�_�/C��x��y-cq>��\��2QȐ{���@p����$��j9r�A��^�����'�n��HI����"zfOd-�	l-���>�t(�@��n����.�θ���}��p�J���2�!z%��&=����V�a�n��|y7H2/�ػo�>������?��G�(��_���I��И,�,!��.���Y�U\����>�)�QU��?[�U+S� �yZ*E"���h�N�(��2/ے�v�4O� �q�����e�ӱ�ܓ�Z���	�*8�ZE��/y<������U��d���4��#�(g��'��~k����}��ѷ�y�j6�7%�"�����Ƹq��Ksf1u.$���@� <�Ƭ[�22���A6�ʏ?���~��_\�v��"K
����T� 9�N�Q���jY����M�,.'��M�B?�b�-x��;��9B�
[�mr�)F.�W65��+�!V6�`W�9 ���uNNOI�I���������_0w
�abG�B�x�p:Hy��!�C)L�Y��c��a�a�	ӭ
Zd�T���.�_��{�b9���������_��}׍TZ�\����#l�RT�5\���a�����o{Ý1�����p�Q��/����'67JIMcA�^�&>�$T�ċbk��(F_2%Eړ�D��,5r�%sE-�B�KrdhKvx"�QXݮ�I�)Y�YQ.C�8}���bVN���6��A߉�̇#��@2�����4?�����[o:�N���c�;�.���M�	��#��ζ��-b��%~���k !E�Lm,����CI�
LV��"��BS�"�x�x��W��'���T�͛7�:�_��wp��ѣ+��eIQ[$�*kԦm��2^.��)~����ݻ��p��G�e<ޥ�(���܍�憦8���9��1�oEc3I:ݒ�u�,C����C��V�$j�穕=�0�7�zLgv������fuM�~L���p��{���ӧ�1��C��Z�]"�sc��b�(��B���N����,��Z����������7R��Tп8���S&Y���X�M���)�t���6 ���l�'y�W�b�s��\o�/N���]\\�=�s4��Ѻ.��O�@�2�X�'�j�w[��������g�s~c�p�� ���d��Zq��sI�|+,)�l�xEqEN2(̔���9�3���qQܒՖ0�!tډ��&��,$��
\FI�`|%������1v/d9�6�!��:O����H���(O{����W0��t�z���Dp�����>}Nմ�*j�X �O8�Gjƍ��v�w�°��	u8ڑv��lD���M��`�D��E3#�9i�Cm���� p�]��_.���6��Bc{�gr�kii�#�1DA�BΫ�|1	�@�Ղ��]TIH�F��Dۜ[%��Z��9��Ȇ��V�����q"��"�C���~#F�,�8��ڧD:,&� 3Z�<� �F��:��V�u�/_H ����H��N9��V���`ް��*I��l֙b�S��W^y��7^=::��#�K7���txN� "dL�iY�xf`V�`�q���m�qX��������^��k� ��>�!(E"mTal���'O^�x��GҔ��J� ���QEڐ�Xd:��Zb��؎���^���"@�+M�<�t�|HS~��j	�g�5=�v��8n\�W������h��4`�X���� ���$ �@$��V2��]'�q#�	t'�#�hD<8�m�:g$S�V�[�;œ2�Hʶ����tz44=AB�_@�G��Imp4���C��fO��e��ʁ�w���I@<j��3֬	3Cly�Z�b'��e:���HR�N'����Gz�#���'� J�T�mN�:�!7
-�6��3���X��>� �#���,�2�Һ��-&36��C�bG,�!�$����@���*`����ò�7����G|�(;o,��붳p�SrX�e�	�lHt��� *('�P+ʌ<d�Eb;��3p��m<�*ܔ0̥��)���Pס`Ș$�%�<3,��gNY�(L��5k��f�3�o�RV,<�S�k��H7�<R2S�1V>��)�����[!lb�]H��4!�9�����_�%ҦB+}��a�v�F�V6n���<�DismV	�A��#��)|��I�ƹ��a�st�'G��{��5�į�O+=��h)�ܹ�-_������i�% m�M�ׯ_��	���c���ȉ��In�'�,yg��G��)�}���K֖/_����H�b��5�����%w��1�m����&�2u/�#D'���a���y'�
���P�M��AJA��*���-�m"v�r�pb*D]f��E��&���Ԙf`#@!�!Ҏ�@��5����,�me ��"�����6��(DAՀ��S�9<�>p�!��*�VB�_V���S/5��`G��dk�����ۦ��C}���_����|�M�>�.@i[�aoo�֭[Œw|���ɧ9�I�$�x���2-]�Zpt���(�u��A�6���D�)�)l�x.�Qz>Yˊĸ7ز#_7aN ���Jb��gg��x�:
�wG��-03U&kZ�O?��.{���V�y�,f�����4_ݐ��k~�	D�B�������Z���g�}��|�]�ܻw���۬���p�%�!I����3n�i�y���F~�In�k��P<-������_P ��,	��PM�b߁7 �����ѣ��c��cǽ�,w`'�o����4�V���FS'��W����>���|��K��H����?Vf�8���e��j4��
�bk�ʀfz�\<���gϞ���� �h��"D�=�K����_2�m����t�
������؇��߀�A��IJ���X˪Qn���ϟ?��)�}�t��5�^ϭ�.�{o��4]�	�"�X���o.1�����!�!��WC[��bkb�$Yd�6H��5�u�� �i�`�͞xK�����d���k��nyw^����	F?�{\��θ��!
�hU?��c:��t�!�ܹ��'���f�(�.f���<�K��]�ʙ�hy7��y�N`M;�\�a�&�;x�h�j�zQ^&�^E�g\��dVg݂�,ح�N�t]�5�%�^���}F�3���i��u�ݱ.(6(	S�$��xFE�R�(�D#W1���@O�	�E�'�g�{ V� ^�J�|H���o@;z�޶:^������ŝ2�q׊:��٧��L���0���=��(�r��l��"k���a����t�IQGGG�Lr�iO�>�^�ج�[;8nX+�����sa�'�!�.��7F�D:�<eK˔�e��c�y���l�XU2t���\��j����,#�*[�xE���N�0:�/�Y*p3���L��'s����ㄘ\��Oi\c'/JbS���g;*O؊��:���`���-�otcK6w 	3�0���.Ӫ�S�T9��>o�b�S����d�R�5M�f��~�6@������6���?�rUZ��"�X i@��-�bbj�}���d�֣K%]bOz��2���w�����\?:`פ]��i�UFH�A�#$��RP֭�����G�B>:�)��BG��=8pR�pi߅t�Ȭ�����x0$#J~ �<I��R�6�y�W��Ӣ*�����r�H*�D'�,+6t�����H�#���F>�Bb1�C����e�(�����Y덋R	b&/ K�� .��f(�O��
�;��G�u�[o�D����5�'K{�8����*��������r!�c�4�+�y�!�`1{���=�;��O�CD�τ�	��ayv9ĵ?���T�Kȶ �B/@B��'�l ������t�;���$+BN���@��1�>�N\	���m�n/�ڹ�8��3���x��xkg{��U�P;1C�wD�$1�Di��6��%0cl&]InYB*�t�ރ��}e!+Ѷ���jmhn�!�� �A�� ��b%,Ѥ�]�&,�<�Z�p����Y��A���yђ����^]N����R�Wt���e,����L�kf+����w$ɇ��Hog����;�%8�:p�|\��bY$���Х�j���33�K8�/�\j���Z6��r���`C��r]����7���2�ZR���1$м�^/��R�b�u{i�L^4���})}��'���������a��b�p��Cܡ��;���G��ϋ�yَ��]���G��S&�bB�a�p!��Rcm()��Zs��8#��ɎD(
�n�ȥ�cu�Ɏ�1�z�˃���4u�B �FU��G�F�5uq1]������b����21(yE�>����]�Z��N1zh�Ií�P&����nĝ�	��gd����4��<S�rA1]�.B�+`IR�0�����M�E��q� �_�#����5�A�"yz�l��1�H�O���S�# $__ԅ��Q(8I+P[���g}����M�,c�(��Qţ�g��'��D�7���[6btY�k+����N|���䔁��kiF$R�|-�z�$H���Uދ��� ��š�;e�Fp%�~[8�?eo�c�y\���9��X�"%��mA�5��W��͏~�Os����m��D�!�MI���b�Ȫ̬����{����ܔ�T)��9{�b\���j�ܚ���N���������t��}E7�<��Q~ܑ�@f�H�牜�ԥ�����y1g�Q��9�;�u�f����� ��@�QT�Dw��(ˁ=��*c�-y �-�f�<� �I�kG�]�!�xc�u)��L��N@��������W^yE�'N%���~�鼃��}�ѝ���b��)t�vY�4`Jco����tЬ��&�ԟ�-������$)�'#�ZKHDPTe]�P'�V��`98?�:��)��r����q-�
/$��gJ�ǋ�ȦB� �8��s�w!D����f~�7p�/^H%�z�t�r�
�_�iժT4	2�t�N�:*������^\}n��Z�B�;d<���`��F%���}nH������l���.�f��`��J,�,���R��sA[�G��Q����nX}.������ǌZz�q�����?�L�_�md����鹟�*0���4�?3"�)���(T7í��h��������E������j�`؎��+��\H��ϕ�=z��Cڽ*�,�kL�t,���_|���/olJ�,���_�z_EA˖�ݫԚA���..f����{0B;D7v�ؐ{sx��D�<йv`��l-(��.�8�?|���ڵ+��� �Ɖz��v���hإբZ,}�������-�2�4�||��~�p<���G���&@��`�S�O{d�.l��+=���s���$� ��Q���ܽm-nYug�&첂�����7)�1�[�n@dA��Y��[ӧT�&�;���>]c4�x<ͭlVF��*p��-���b�J�������K������ִ�1}5C=�Cv�a>�ʑ���r�9�Lf�W���HTR:L-s/����"'�"��)K�7ꉠ+C�s�:R�#�yFA�>���4(]ق�cF\gL)2Z�����2üo�HE6iL(y�"�`d�zb9�V�$��kb�����+�_��gmy��{��)D��B_���C�4d����Yޯ��ÄT�BJ�˾7�"�]gmX"�Jw��u��;R@�5�ڣAg�-��՘opqꡪ���U�`�Z��tR���<����aW�Fd볃c��4Qꁪ�p�L����I��PF*�bh�q��0VV].<G�Q�F3,;5������u�!��;!9�,JXM%Y6��63Rg��x��e�S�>�`�z���:�q�y�*D�k}�����O����n,�������<p٫��Qr�����c���uڣB������~�Q�OƃZC�D��QX�qb���T|ܢ?l8�J�i:������X������9-�L�/bf%�4T8^�'ք��}��;D,�X�К���T�%�u���(�cC{��yF�O�Q�X�G{�Sڏ�Ia�5Ҳ��e#��X6�~�&�Ը�(f·��|XX���Z��Z��c*�d��d麵ɩ�X��)�̑GtoH��`:�҇���x�D�D��XnQ�Sx�W�qp�������㬊�RJ|~���*&�g�N)�2���)��p*'��?�Uo���Ff�O���<�% %��B%�e�Jv~>�nX��E�>�d�q�{��vGu<Tb�N.��^c�p���ދ���j���Y'�q�C�$�Tl�	Rc��f�F.�^�&7�]t�1�d��+���,D�1����#����o��^N�ik��\���/POk�*�'��n.�.���*���"�7�I�6���J#sc�q��mٙ��y�ǵ!麱�.�s N�2c���fk8���e�y8��ʸ����~v�g�k�e�'���ѷV?�j���[3�E8�%�o@y'��>�C�#�no�����$� Z�q���f2���#G	��,�1��<q0����-D�ةk������O�0K���̯EYܺun'��X�
8�d2*�w*��E^3z#�7�]~�D������ˬf�;�̗��0�������Q%y˲S~�� ��m�y����-���>��u����1��`�&2�C�c��ņ�rړ�J"C�:,2��؈�\���m��W�9�� n_���X���"�̺�%�
�r+%6�fg|Q�*�L�E�����Rl)W*�����Ԙ,���4x�+�߸I�q������'G�nG��X1�.����5 !N	Ӆ�)|:�>\�\u'''Y����߂���ݑ
��mf�}ĸT����I"&{�")�ݦ%Ɩ29�#�&����B�L��)�<ytt4�x
lQ%P��-*�u܅rDX?�!r�������3m$ޚ�w��9�8������Jc��������7|������O~򓓣�D1Mܷ�%��^�o�"��灢��&2�?�������/��{�.Ql��y�^�e;N�������I����3�=��a�_�x��%\z�o8L�ӧOي�M5qqz��~��g�]	܂ǜ@�]f����*|N�a�$(I��t�e�}Q*�E�#c��)6���y^�?+�*�!���Ɣ!c��{���c/��.EG�2F~�H��s�ZS���W�z��]��0M��DLK�r��#B��Jd��hb96�F�5�PӃP2�`x4
���`�Q��2,�G�$��HX�Z���ɑ���_�yx�pR�t\k�f��i�T���%
���/~����曬�������F��͛7��_��7�FNcUA�%ZJ#���r��Ur���&L�/����V;��MY�8�Р���lH��'85�0x��m���/"(��Sy��K��kY��jc�9�#�Yw��г5��<Ԕ�Dݴ}��9��N�Kϳ��r���W^d<Ș�7�����-q�fg�<�3+d�e��TS!��t�\�ivgc|/�hJ4��OFl�EuLIw]�6jE����F-˜��X������!g:�Aypu��kd@���IE�9�wu�Ը���k2��Gk��.j����5%U[ٖ�R�Z�v� 0z��dn����r���5b�����ѷ!�xz��2{��5�NB�?vm�e���/������	=[�?�(g� ��H.Q����P��!:��"y66B(P69�恅A4���m�X���`��n0d��B�K�����mm�H*KC��b���Р�'�H��G�~:�j�$S�T�v�]=42��<�,xё��d�p�òb-���L��^᮳�����W�nD�)��Z�!S6������x�c�i���G¾!�wR�-��Ѕ���d�����;�U�����N����>D��-C�M���yd:cf�pǛۗJȍ�oA�����n.��m���'�����~_�-�"d�@�:�K�v�Z��� ^ty�VuS
�<�<pmڊ��y����R�E@���c,}�H-M9Q��"�ME�W���PA煰,�d?L��K�&/�8]|�|U��o�1�JZ��GLE��Q�E��p �*R�W��d�$BrY�l�<
�_��d�zU�k�s�FQ�%$���+�&j`�G)\��Z��'Y2���b.��ԩ�pLhcI<��!���s�8甞�qc�^j��[J��#����|k�Դ5�n^�T�8ggV(s6�tѤ=�h0�[(=��f%S6(�4AĤЀ['Q�8ϒ��]���o���F��s����w�q����M,��H�XX�DP�Ä́�E-�C�("�m��M�Z�Vy�[$��GQ')�J��ra�����i�3p}|�'�1v!ޥ��$�������@�k��� IU&�������heH�v�+0U������0s�`��R��ĝI�c+�%%�'4|�>��@���斘�q�)h�R,�TI�P���㈰s��2y�٤�����Ғ2������`�2w���	3iP�t#1Ó�Jii%1J��Xڂ�O*US��x��V�:&��J��MU���(��v�&[;��〹���K�����#�Љ�.L�V��"i��Ԗ>�𢼪�zU
6V���X�;W�r�b�ilIH��}�v�~I�Pz��ʘ�P����n���m-�%�Mc��͋�[�U��9c���p�Q���L�X;s�gX�!,��Fơ��p�É�lA�pb�}�.��,F���z�y�PFDiR}���t�H��}3���w�,�/�ǣ�d�����x�$���!���xsckX�^{�5�0$A�{t�r#��ՁH���/��E:�v8��|���z}��E��V�A�r�����f9?�����P�R6fb eZ�'j���b	�z���	� ܄[F�+eӷv|�h����Fd%��p�T%|�G�4��^n$�6����	�QZ�i� 6t�U�#W����)�D��a��ꇢ��B�n�D�(�-f$�l�3y#Daͥ�4��|X�X2Bl(�(~�p+e�u)�*�c�a;ϼ2:�k��B��7_�-�w��+���)�]��� t��	|������a�P<���nnN!J��q��#�>��kG�1�r�A��ʓ��ի���[q/	�Xg'\v6g[�v�]����D���nB�B���KVoBn/ii8x��쟴#f�b��̸�a�67�E>�l�KiMؔ*qx���QN��*B��Z�y+����/oܸq���HY��\�e�~��W^y�g?�����-m%2^p�V���d\���l����]��3j��V>v~>gS��|�;ZK����gjA��A��XPzC̏2��2��R�����@��WZ}!֬�A~�)�t��˽���ϟ�^c ��b8ى�� 2�Bb�<V�uoCY�'��xd�S"���L��I�裏^�{K멫κ�`���Ý;w�y睃��gϞ�֘1I���h��淒�0M��%~��Z�Ӟv0��Z�O�=R{�ւ U �bp��/��Pr��f�M�!k�y%@$�Q�)��K�֩�5�Zj��Uh�ؒ͋� ����6�p�+�/�7��;[��	f�J9�*ք�8Ҍ�\�	����u�؇~譟q���f����7���_��[�nNF0�;��Bb=-S��r�+,M�� Ebm���(�r�Om@y�F�o�JT��G���̋W���dc��²JBh%����k��WgZ��[=H���O?���������,}'����_��>���*�|}g^sclw~*��v�VY�$��}�ڵ,s�*�����L8F����{U�h7�л�xx�?���cXO���&���F�8b�-���/c30yπ��گ���v��R!Ļ(Ӫ܇tL���lQi�R
����/4W1�X�����X�ݫؕz�;2�BBF��k�t�6
�)��LH��l�>�����4B��Q#,m��:ԉ}��n��W���e�cn �Fn���
��e�.�q�~l**1�7�nnoA���J���}ax����O���t�����qxx��'��/J�����3��[;��4��4$�k">�Q3�Ui�J�-��qe�)Ú�.&E7R�m��FbjD��'c��8�8��d��"�Y�L��%������(z��X��˝�
OTjh|�QB�Z���5��=�&�lX������`�4A+�����3�Ba��}�(�v׭�}x��L��s��Gd�G~>��b�n��i-~�yf�U��p��	f%��4�"ˠ҄R��ă�.p"���ڊ��_�p��at������m��N�t���=%�'�1s�e�>Cn�bg�ׂ�-���{���fPɞ�P2|)E4����ё����͛�[􀬛w4�<�C�{4�ϓ�'�����~��%�4�c|J)�<��'�С�S7"1�����q<���h�~_@�Ã�>�~/��2��!y�=�U�{�G�lŔ�_��E�ڐ�Y�ȴ<{�Qj��M[�N|BP�H��P*@j�!�}�S��A�5���(�޲��{�u���[���0S.U�8s_�a�1F1�� ��&�}-ز����=���S,VK���eZ��{,6���ͻcڙ�rB=O��p�̭ۉ:�]�Ck��1�৉���i�,v�kw����x�<�r��Y�6��e����bb��k^�2�8NWl�̰�a�2���'�� �ìg�WeN����jM��ɜ0��E^�1��G�(�խǡz"����C��ň97�$�kn��@cO)X&K�݉)�^j�"�5���UHT�ö8=��X`c{�,�ΏQ�q�v����!$���ħ�bj�ߒ���F��/��v�J�ZApt]<!�:�,�R?kϝ�&ͣ�+Ϭt���h�\�#���j�H<պ"��(�Y�+�����Nګ����K/]�y+��!�5RD���z��@0|��e��
�C�ܽ��/^|����b�0�ֹ���@��H,ybLdM`O�u���r��YP���]�ζV�#�(|n�Sӯ\2��v�`e�@x:p�qݺU���o��f��*+�q��k���x�Ҹ�(g(�d_�ϩ<�V:��YV�u]/?��u�E�^Ն��=�km�D��s�-oD����z�V��Fok����`�:�RD��GMS�H�Ԣ3����Jё��>�8�G1�-�<y��Ϟ=c��I��SR+�A������$vu�5�q�sȧ`���Ӿ��L:c�tS��)��iL�[}k��%�P�^8��Z���c�S�1N�����S�H�B��G��$j�^���������W ^y��������������¼��z���=2���"�h�=\�2��:�`�x���5?�c�q����c������}?n��:�_\�'e({T64h�OQ-r��ֹQ�
�L�^�7�pp�hΥ�.��W�d�O�Y�?;�he�+"Q�B�yBZEY9T���;３��7����|߻w߅���}���ů>��E}�E����4 J���]	��W�!��y|�Ҽ����3v4���oQ/\��'5vlWsҸj�`�$?T3�1XSe/��uvF�c䕰�����R�Y#�X�>u�]m�07#�C�4�IV|��W�_~�e���2�҈�����(�|�m2-�u#�}U���f�q���w��.�)	�Q�I���Gj��jJ&��/�����ƻ���ӝ;w�xsHb>i4{�yǀ��^�~�V�7Mb�]p -�M/���_z��l+�������Uh#˝�y�З�̅��� E.�)�՚�a�"x�2�q!��{,j����ȓ`W��/A<P����(��(A!��vȝ;/��l��6�;��/z��k�.��L��VKP�xL��A06r!\��x�¬Pw�dY"��y�L:nf��j��"�+��8��`�e��&*0��~�%�������=�4�/K�#)|%#��h^Ƭ�y%W~���ّ�����%��S�+Q���˯�����E^�Z�f�%��=���X����wv46�n420j�;ȃG/޷���� ��:�;.�DZ�FY`�D���5�¸�doLX�-�i�%�//��k�0�R�.�j{��( 
E�*�L$��rNb���V�]�n�Kei�B�6�:r�a�`�m�e��긼�pIi%�nJẑ�[(�S&�G�^�W�6���Ŋ��ǔ���8��x��(z�"=��V����m'W�#��JI>P�f�)���( ϓ��ԥ���C��|w���֘��:m������=*�;�q�=L[r�M1��ב�1�D[3(dib�o�Y��W
KV�*a��2[Eݎp�ō�O.KA�^���hP4!� ��[�G�VU ��M��d)�Ak�"�n'*��:�h��Vp�Vk}(�L��������.FrkPXa��m��[��PCT4R��-�#�G}�ǖ{Xc��rn��2�l_��p�AWGn|�"nK/4�ɹj��li���+J�o方���`Ӛ���C]��Мƀw��r��=II�+��a�
�	5t�2�$FH��4+�6� �#U��`:����t{犈� {�
��v�C�T���%�Q��R�фz"Is��c9�~� �J�Dn�$#3��<"�b0���􂴌����W;�vQ ��T2BeW�N�<}ʥ�uU�l���N�eg!��!t�q��-V�`mc��=3�l�	�=��f��B��4Vs�/�/W���!eU7!�rv1s�f-���R�ym�:L�`NZ�@�0JH�&�1.�h�}�E�5-��1�T2�k[9�ڋ�3�~��լ�;�']V���O#�8kв��Ŝ!�jL�"J��4J�Y��х�L'b�ĊIN�.Ү�+-���fy!�H�͘���3�K߶8Y�����9fq��k8A���\�bV��W��b���ݮ'O��N/��$M�Y�bi}������N&b��^�b*�et/QR6I�G�*�� l72
eZ�����$�;f��l��GڵD2<��ə������899c�A�$���zUj�8�8�u�Ί,̞B��.��K�TZis�G[(&�	dj.�x>��I�f�T���K���tc2ep}z���f�'�h+/G�o�67���ڵk�n�z��q�+W�D�a@Q�	�v$���5Ǜy1ژN���7��0�Y���@��{O�'�����]����I����xR�ƃ����p�@ Č�B��*1bSy1�����2�T/.�d�*�p���~Q%�K�gb|Y���-�ZS��w�����,T�K��^"�ψ_�����~�$��^_�Žn������oS��vu�2�UE�a�D���������0&ȦF�,���h�ձU��'c��ê�12|��i���ը���*��sV���+t����5P��YK�~o�H��B�9�i��Z��8M�5���.}flƽ���������o���������ϰ����D���O���u��7$[	-���z
���molÈ��,�,��'}p�o֬��*�P�����)��(�&ps�+�2G��1�ǋ�%6���
+��쎸.�墵d9S�v��ܚ`�z�������W�w�1�JY��l�g�����9����?�����^}�U�A���O�>y�$W2%��S���CB�U�Q�u���[y�Ž���Йe��|��1�	��Ν;	�f~o��ڨ�`�{��
���<G+{���a�q&��u�n+��@Q*n|l��{iK��u�eߓ�&�����p�������6�Nl!�¼Ԓ�2�T�&tԅHa�A�[S�W�������n߾�y`�
���?��>mo�%*>`�@�q�4^�ɊZv�cP]6�-�	��t�fqe�ҝP�	i��#�G�$ Y�='���HzՅ>�z<�V_��-���@�B�<n�]��RBXi_c_Br�\���������	�������)�|�5F�"c���e5| S����{�k��F�/�A%Z�M�ݬ��N>�ҭe�"�{��#h���q�F�?�Nر66�\�܎�]Z��'�|r���/^�����]�Ӌ[e��C��_\ms[�0E�/��<Aʒ4�DbF?V,cp����98Tf��h�A-*8ړ�4#�Z����������ￏ�|��E4?�i��ϻ$~~�bcsw�Z4�stz�^*�%}D>Ht�!Y̕�-j�F:��}���$�������7����d����j�u_���z�<u0:�WdI.�-�|~�kM�'q��Z�p��+Y�������`gӶ���O�N��u�&4���������Eq$��8M�Q��EM�a���5=�2�F������Q@Y�ܯ��]��H�.|�Xb��΍?���I�*@:�ۃT��b�%����'ST$i�����TR,����`.$8�Q��՚�L��p,�X�"O[�r�z��[�^h���7��`��3�r�`.�YjM <8�%ϸB�4�B�S�(��@�K��.�<>pɽe-3���ધ�	���.�~���Y�^"�/��Ɛמ[*�w2^�Ԫnc+&bR����΀T�ř�?T~�ܸ3<F�-XBz;7�M�R/V� �pB</�yZx�� F`K�N�ڶ�7��Ul1)�Zc<Q�/�p�΂�PF�R�D��D�M�����簥^�{�?�����U���Ҡ��RUī��2�V��N[�?�yyH�j�c�RdL�<u\#~ѷDaT�To�G��M�j̷��W<қ��ĒB�����8�{;�ĥ���+(g��+��
��桱._��cl켮�#��Ƞ�O�F���������-J�J��x�\7GV8���[aΟ={�j�'���[л���x>�9��I�Zd�����G������h�I�/Vj<<#��p�\��(��g�r��5t*܍��X~�M��>�PR��]٫�E"A�y�t�h����Ӝ%���k,� ���泴�x��޽�+��٫�-X�|�p�����t�12��>oЊ����t��O�Ą���w��"�">);��]�J3�4�B�AxĚ^}�_����,���5�8�IAr\�����/��%[�Ŷ�ʲ�8��^��B�I���Ղ��j�-��C��<�il�� #L�rQ˳�a����͛7q���ۿ�_�������m��ZV�*�re'5���]������������Bp��ٜʑ���6�^�ƙ��/:-�v��Y"U���dcS��!a���[�nq���D����"��bI2u�7��T�(뭷
- ����6�ثG'�� .��E�΂0n��݋7���;����{x�r������u�$���]�ۆ��{ܓ
=Q�?Trq!�H|���o\����o�Qʙ#m�	�"�?
aM�D�hM.�;I�9�8�GG���
��9���og_��wJ4��י�e�i�y�A���S�Y��º4`��2K����๤���qW�yt�_��c��z�'24��tz�&1xod�=�(:��O3�d��06�ƚ	v=
*u*�v�-t��J:��F�Z�r�@�q��+*^w&V��jD�o�G�3%F߀q%�eX�|�nC��dٝ�O���<DBu�o�=RW�hn]Wp�+z���V�0�~���gp5��q �_��~3��Si,���č�?�q��M�k�:?=���|&�*Pz��H�B��J���Z⁭�I�8i��,�e�qqH���=	��M�`��:�,r�5��C�����^պ��66�*�W���>���O1����/c����o�':9;��-��kc��<?AQ�]�H=���r_B�<s�֔��3�w�fP*�W�^=99����F�K�"g�oD�E�s����0�R�y��c����*���Y8r*JZ>��3`{���~�����x�q�ihq�K��ʇ�%�gr�Ȟ�+:����ƿ�ۿ=x�������*B��.�v�P���3��PxM�}�:u�(�
�Q�;A�/m�����:I.��癦ZH˗RE�M�qz�(�Ӏd␪��8�"޳�t����څN�}��k7�f#�e�+c�bL��	U?d>	��4�:+P�KF�(͈��tG����}��i`<�U�p�6��z�:@��4�q��R��ׇ�/ �����q� ՔC����)�y�)CZ�F~�k+��*lz��Y��(sZ���]յ��Ҹ�y^*+�H��jW�C]||\��?�4���M�AmH��-*�ג�E�B��5q��B���pH>^Bɂ�����5'Ϟ=����*�d0Lu�4(ц.1�l�@�ck��n8U�g�=,{��t*�Z\���υŻeE.q�՘��3ӆ|ծX��1�E?�u�]��W�v%UI�E:Ks*w��y��I�n�{>7�)�ۋ�n�$��'<4_���U��͈[W=�����lJB��|�5���4����h�ĉ���A8��_2�/����6vK�I��/Wm���T��@�H�;p�8�F���b@����&B���u�L/�KJ�����D�DJ�1Z�����a��T2i�1��d�e�cu��NeSXһ����D'q/��e���R<��<�z���r#���k��M
�mJ�^�������Q��X�#k B1���%]H ���@�ě��ʺ& �\c��ny����%r���2�=�Uc,����9H{�Ͼ��b�3����QA^��!/�I��!f�ŋ㪜����!�εq��D���B׮����Pt�6Ԁ8��*����du''��+b��1;<,R�!=z�݋qO�X�k�urwB`�m�T;V��\r�����˲u-L�e�f��4:��wcv��D�[���z)|=��V�F$N�ry΋0_��(GE{�Io=���پq�,H��c27"���F�:�ʁ�� G7�3�����Fd��ƽ`�"g3R4�x^��0���6�Zpf�\�|����w!d�|�ԧHܕ�2/Z���Y�}������'PF���|��d돴�K�p��4e�qw��5@5O���Vs�8����1,�]����|a�cwF� �ggc�Z�ߦқ��4ҷ�7�M4|Jq6��%�/���=O��O�I�{�?�7ς`s}�� i	�#]�.Ě^.9�<z)���~#����vtt���x��^�^�?��@&�y��b�*M���(ᳮ`cH������T;�I�^]����8<�4�����-$��
c4������|������wp��c�}�%^�L��{{G�g>]0�2�6��lX�'{O�^��ƺ�T����'X2�ջ� >k�8f3���石���O~�{ߓ[k����������������պ��ߦ������\�j�s\-�fZ�D(��h8�/�ϝ�۶��L��g��sz�e�TM���]�
�!�o�;sh����a|��͍��"��S�#�F>4F��8omA#Ԥ0�z�Dk1�bxTt+������bv~v~��̓K���p��H�����3sq�[���ozh��l���L�r�)���y�(RC<���aT]8�r���ǥ��Q]I��ի�6w��2{1QN���?>x�'b����+�����6�ʨ��wV�����7�|���5��(�B�g�'0_z���y�і�P&��r�	y9�땄�W��� 	���Bw,>O�Wd*�_gg��x�9���U"p�.S�\*-�e(�c
���4�ԽZz	<�qƦ�mRc^�ӱ��Fl;n�t�Bqmd�F�L�j�����5������e�����jg�Em���U0�Ŷ,��1v8�����%fϐ�[K�B��<�FUt��6��?H-?C,��~����C��#����Z4u�i�1O�00�X*���j��H�#p���?�L��I�#�p��Y#X���Wf�?������H2j����� o\���l�@�-���u)r#�B4)����V{0̓��kҹ1.�E-k���-|Us~%�$ ��f���>D��U����Ȳ=ʦ�;z
���,��$YRi��cm�U0�H�~�>D�dT�V2,ފ,��6&磏>����?��?�������A��y�}�78�f�d�F����}�^�6�~rc:˭C`fD1�a3���h����c�0�$<ۘL=��h�+y��X�VwQ��p�Ő���F�g����i蕞��aPL�7�ǩRNL���l�D���$	�Z�t�!t��z�L�j�V��]i���q8�����V
�N��$��ds�fa��w>==x���>��|l4�0Iڣ��H@�n�@��a)����ĶlQNc��'�Å�3+���L�`/��Z�1�A��R�zjqVa��Z=@�&�CA[�c
��8E�#�2W�CW ����@�F����YZ2�<��v�:Y���O|4&�K��������q��R��Ɓ��g���h8w��Q�:��K?W
�r�)�"��f�s��>==����S�c�u���|㫯��4��WW+�)��`�s{�v�� �@��X�Sn��t��uY1�V��m$Z�!��zYdJ�X��� �P��Ѱ�&�֎��7m9�|	���mԍ������j�����s-ʅ�r�ɪ�cR��CaZ\����f������_��� ��������u�������4��l��fd���t
W��&��Y�9��M��kYZtm�0�-�)���D�1eY�"|`�T�:���Ed ���'"=��p9��K܍�[���� mZ2⑥��љ��2�-��<���!$�3g��E�OZ��h�#��a$s	��_�s��W_��Gi�5�4�+d�~1;���|��C���"T*���h2�nO��
G,��`�'�YRC��Q�ɿy������\{+`wnO'�u�sP[ӈ$�.;�r�X��ٳs�Qj�~��Ѿ��\��B�y<�cF��c�'K��Wm� =u���=Dޮ�\���om��rӶ��hU���3�s�o~b��B�����.�cZ�����i3��*'�#3�/�S�r7�e/����q�V��I�I@TBG%%��3A����R���fs�?+m�t�|ppp���K/���WĨRΚz-���˞�� ���$�t�.�P�)�[dpRw�ʩy���xh^L���r劧C%W�Z���*r��"��6�O�I6+�6�WLp�W��*��S�8�֬��~�0�+��>.�s�1��@dS����XE���txGjG
5�^����/�đ����Ȳ�D��(uzlm��ӧO!���ca
����a�(��Wq���.�Yzn�n!uC�z��I��$�Z�OݗNOO��F������Ɠq��0K��.�G�ǚ><5n�/����ep��e��Ms?��;���a$�Q�=&�^id�W���$w	f�[��y�� ꘖ�\pt-�����B+s&�3&?M2|��A���b[=֜����P�A��@d�-������
.�%jI�-�&�ɡ^S>�2�||�	=�����B�k~�eej��J�F>On�����\��b+���Z	��xfZXD�qR��:CX��J�ϳ�g���$
q	ݞSdQ��8��=Bޣ�c���"���ʎ��yk�nE��k4�Y�w����{��>�L�=e�(��-bN]���$�B�F�a�-h�c۸� ׋Rt-\Z���.@c��-�Yi{���q�X�A�k���KUW>dT�AO
JW�F��I~����u8��X}
%�ʭ�.G�+�8�=Fƃ�[���q&�lɰ#��s�D�p���&Q�|foooS���X+�0�()>�iqiV�$?����hJB������O^N�, �kׯ�׹��+b�dy�^1=C�])��ts����~�iQvE�Fgl;��z�����^h]�!�#��2<1���C�[L�D��yXL���ƿum����W[�cH�����m*Zñ���i{�;�'�&��u����5����HW�Z�����ʒ`��_��!Td���x'�/���n�q�Quf��HvhhhQ���~���'�FQ��k�Y�[h��qfV���k�
���k�Ly�ޠ�Q"R�p�A��ac`]؏/�ʄ"k�
��*ו�����n���8R�V�Z��&�4,	����z�0�:d�oZ%�iZ����y'��,��.���Dx����$OG���Ҕ���v�`z��ef�+c�}4�H�y�9�4����;/�~�����׵���O��gϞ�q���Akj��L[b=^��RQ�����NQƾ�re0����T����P5V���jA<���.�Pw��R�q��cth�PI�`�N�� ���:6dkk����Jk��?�������qo�5Wgd��%N:Ɔx�y�GӄS6���6�����1e���ذ��^���'�sJ��H��u��,���L��_��	�P�>g��\��.u�!j��~�Da˸Xj��5��ț�ޫ�	�h>�K]D��v�Fb�?��@]RE�t��n�5�,s�B��-Y�C���/��ˇ��ί�%&[�����l
�Ca!�ĘP�Ѐdxj��T�lHM�}�8�x�֝X�qnnHRv��Ey�D,��2tMq�����=���'�+�|ڇW��{$�e��tx��N�[Wm�B0�0l�<�"(b9��35�*��SUK�����n����N4�>�V�/������߷]���8T6�~�;Xŗ]������d�� 7�mJQ�n!l�TX�j=��M�5��!�6F�X�a�2EQ �ʌ�:��W��Ӄ��U�j�ׅ�M_/Yp3��>s�Z�U�S׈ە�/{Q�x&i�^[c �Ad�$�뎺&��L�>WZ)o�d�>���dyc]@iD�=��c���~�`ª��H��9WY
�-�xd�h� ^�h
�{T��$n���Cua���֌��8�q���w|g�<�q�2�K�Z�?`s�w���!��E�S���"��;������x\f��ZR�c�}{��tq���In��z���b��{�Tn<����:Y�������Oll����/���^l�>�`O������1�S�[�q����{��qMV)���ƌ[ǚ���,������u�ABL��;�W狓����G��F�`�g��0O��źo�]\q��|E� �Mm�+�@Ԕi�^U�/MJ���)C@&�K����e��:wwn>}�Vv6�t��E�k����^��[�WE68=:���k�n����lZJ�^�Mi\�+i�-�+��[��h�ޯ�Pˋ�r���U\2����ug�Hj����9��眨%�
�Y��M�p,�����mi��D�a5Y�*N���ų�sO�W|q2��3G/$���%p���¸�ت`t��W���
w�]̗$j��؈p�X2F3�/��3����QZ��8�����������ĪH,�*!�f�����Xh8����l<�ߓ�ʳ���-�o���@��O^q��p�`
d�)�'����gJ���������!F��Ж�|PĪ21$�g�$������q���h�����\�֭[�S��A�Ƭ{i���
�b���F���ə$	r8ck��d)�c{��s@��U)����t#�0�)���ƪ�������	4m;�^,V��B='��X9S�	�;;�	k�+�����
�]C�A����9���<�H�~�;�N�+����sm~��,�m�|���1��>#�͓`f4�$d�P���O�<a<��@YǇI�Z7n�&Zd���R��:���:o�/_{�F�0�Ϟ#t�v��
��P�|�5n���=Ǽ9����12�Bi��N]Q����������i�:�� 9�b���]�P����u����OI)�:'��ώ��v[�+w�d��\��>���?���q"���|�拴��_��������Xv�?������o�-L�b&4a� xV\}Z]S�ޏ������X���$�F����.r�p|{~v�H�`FWy<���J�'���L�ص+W	=>=>Y��%���s�Ȅ9�ac�6���:�����O����~���]n�$XQ�N������̺Ȓ�BZ��� �$��͛7h8M���^/�R�%�Xg������&�SQ��������V��!U�������x8ZJX�n�d�1�����u�v��SQIк,��#�/&�|Ԥ6��XI	�~���=(�M��s]�(pk�n��f�1���^gX�=X.='7�ܡ⍺�e�72.��J��&��Jj��li�d�!�n������8��*�h
�ˤ䏰C�^٦W�kmnM��S��%�B�9�4U�Z����Vv��lo'��w��&�PW��e6^�	���<��4�/W�'X���>�n�FQH��E��(�^�e�[*U[Z�[�m�1�1�:�ⓓ����~��7n~�o��?����"ꕕ�j�̦�]uS�m�Z�s)��F��j���Zb�6R$Bהk�� 0�ji�#؊�͇
;�X�����ʕ+�rM�;X���-�Bq�V���F�|��v7�F�J#F�h`��>����i�[��G���?�t{{����Gá�'���?��ߗR/��$��V�-�c�0�V�¿z�3�,�L�+5�ֆ��K��)��Y�@���ɹ�9�P<2�[C��uǂ<���\�ǲ
��=#H�Tg�E��*ԡ���پ�5C�(p������xzL*10Je�ۙU�gVs��IC�����A�K��C�LKнgY�/9�\gp�#f�^�i��,�ӎsI^�������}-����CY/��Uq(��Pjb 	���?�R$��et,��E��'ӰQo\��M{F���t�bR�E}��)�F�\�����p�<�E�ZY��3Hu�Dl���g.��C�x�&5h=�԰�ܢm�v-�z�|d��Q�y<�{&�{E=n%nr~�Fq���J�^�'O�L�����7o޼w�>C����nmiuBY^�j-b|8��JҨ��P���]m|8���#���P;�v-{j��Z�2��1��X�M�.x�O�	�:|�������ħ3]	UR71����=�Vy�Ƞp�4(�4�uuՎ&�[��@I��Zݻwo8����~��/��ҽ{w�t��ߏ���0c�T.x��8�z�X=�lL��ͩ͒�9���d$XwW��㳵FTy�,��@LA�`]6R.���6 �����D@�q7^R�tq����<��|���1�	�쫶rA�+*��G�}*�+B�C���Kv�{�Q!p�J�N�M�����*�O�_��(&����B��e(�d�/�J;�V��Fu��"��������Ǝ�X'��4D�2n��l��D�}
f��óF谥[�iu��&�������/\6�8���{!*w���3������$��##��z>Oe�IuL�_��/��]�ˇ��tkD~�l=�Y���
��&���}5�"Wl.�BD�����QŨ��]��ڑD��WtkϭaN�R5�i�gl,�O�Z5�O��_C*�ဤ���.u��*�
S�J�1�ۊ�9ȋ��)_}��7n��݄[~�l{�U�qĵF��e�t�yT
5����4b�"x��H�z�����p�%�{{{�l5�B��	,��P�N2���s�����I�I�d�8\��-Hp�m��d���W��(�Д��C��|g�� 5�}ꅆg�*%atf�����v���Ƌ�"�v�
{W���/#�G��W�|�9Ql�*���A[����!��;Bx����Xi}�Ơ%<z��T9�g�⫯��#X�`�A�*?����iJ-��<����3� c"�����Ǐq�������'�|�>��֞�����Z��z��a�c �H�19S���pLk�0��ݻؐ��r)�U;=����_ ��G+���<�mra�lS�&5��1�/��s�!�:�Q8GZ1�
\ܗL4�q͵�v�$1/C/����C���w���/��j+���%�SCk��j�yg	a��J�t�!&x:�4��\	�j�&62 μrۗ���3��,@#��QlN>lq��ք�8�ftm�i�Ť��?�v����bl�5�ƕ?��c�{��U�13��ׯ_�����<����	���~H����j�0�?n���h�3�~�ܮ$FT2�Z��"�8{��L�cN�4���E�9	1���gD�pH��[�fKd����*=p����}��g�F⻤�x���Z� GE7G��Y��Uȴ.W�0ǐ_�����Ɉ��ǁ�³c�`ct�֗�V!G�V�j!��~�
�!' �:wΏ~��B_x�_���3�����2� {?*�\�����4���;���]<�m�"L��Q�l�5޺/¹�[F��Ud�;gR�����@����0��^+����`	�f��6��C�S���b�����]Ţ`����IZ&��k�"8�}w�4�5�"�\�����-�:� �I�z�k^���݁L�K�����v�(�sAR��T�{���c%�`�#��
�̔e	��cK`ѯ]����௷n��C��@�">�٦��_�^�+�%�ƕ�+x��ǃ���� X��e�+�}l7*b��R1��35�5%ʥ))�K�ţ�".�ܹ��������><�ZO���He]ƑQ��C��:�!���{݄���z^@'�WD����7��MX�2��g�4s�~y뭷f�sx��@$H�L5���$�ٚL�]�(���`�Z��>g�61
]A�������~������������^{�������j>�L ��Upf�|�f�G�2�N��KܐՀj  ��IDAT%�:s<A�����L�5V�c���a��ʪ�^��z���>Z���Ꝺgd7�{MMQ4y`��-[F�Ϻ�X�\�K��Y�܁u��sM�	>F^`.��?��4J�*pV`�P��ಋpc� ��=�e�I���o�?���?�Bd�9\,R<;Kg�p��Q�h��uWLM�
����Xb�x|�,���)U����������bO4��Ċ-Ƈ7�#ލ���5$A�.?Z����<�����-{}{��������5$�[�t�Og�Ǒ�=��|�����h,Q�x�"&x>:<��t-�b'�/���|�;�"�����c&lP��Z���T�`p<����0�V�si�������)�}y�������R�5_�L
�
Ët��V'Y�2Ie�NT�%��qLo�	MG�õ�������')��~����;�j�C�̈́mü���_����l����w���Rw�����O0!�;xk����+�a{$=�`�q��Hle;�!�.��E[��g��f`���!޵���4K<մ��ظ��RUv	9�/RG�%u,V�2+�����9>]E�*�0���Q%��&

���u�J�5YԦmw�t���4� ��8�%�o�D����8;�_)�%�g�d��bR]�Ɯ��cx|�X�w몤�4M��!\��=��%>��M��`k�8nMO._h�%Ƭ�
�ϒ߫�>*[���q�ѿ�U'��Ox``���@��z��*#k.э���o���7A�kT��\k�6!BlԒiz�.njC��1��q��[s^�3l/+��&
�=k�:� �PIA��`��q!O&E1�ٹ"dj��ۮ]ݾs����Im]�qK�:£�2lh��/wܠ�	ŀ2<,xb����.֚�d:ݼh.p���5�j��iy�r�767uc���sቖ����_M�Jn����l٨������ִ�b��l���'K�U�Es�Q�N� ;0�SVe��dę�ͥ���z���rz�T҆��Kl�XFϽ췝�]�pze��M��t��ʫ�3e�c���F��8�Qb]��c����1����#��D�C1�&�~��,�.f�����;�N�&@N��F�Ȗ��	Q���j���c���0�T�yhܨ���䉔����v��uY,Ž{�nݺ�?�ǿ��R *�̝�c���+ɽk���pkS{h�IZ�ӫ�mI�K�K��\dE&��"ƭx*�:@39��!'�ǖ���1�8�Z�a���=��7�x�c1���a2	�|ׇE�X6Gp�0ox|"ؙv�8��h>|��%��X�%�Wm����4F��V��C����p�$��D�����Zw!WT%D�A[��z]t������쵝�j���C�c����ӑeر��9�zP񇇇����3H/����d/r��v�`�I���	'�������Y�0�d�'p�i�p�p#*������0�t~���>�����p�7:�?<;m66�����h�w�z�,��W�N�f�щ�:?�&x\�:�õ�E�F��֧D17Mh�ǰ`*Ԝ�;�#<�@)ON$N]5�ř�^����2B$ӂ��\U��l�F���f�v�a�h>o�y4���I!C������@�0��h8�v�,GY��u[�����G��$5D;�_ǧ'M+�U���ij���y��m\6�b���$Q��N�)��y�C�jV�]��)1?ǜ�����-��+�BOA�\		����O�z�$^�����\��������Ț �J��K�0BM��b}��hP$�b����d|��M�њ�W������{o�?�Ï����R����)ޙ_H��(-PbC��lmW�rs�)���4�����/���o�q��]%�<jڐ��̫7֝�}�������韚�8?>���x��u�
*���^P>p�)F8'<�4�XKGw*<n� �"��K�2���'@�Z�`D���M�I��!�(�A�j	N4��k�x�}*��^�*am��nTk��$ϒ�j��ɳ[�n�f�7���K���z��A�T�9%$�0/:�Q-��y�%��d,U�/�t�0��
�e���-���g8;���ӚŹ��F�
�E�y�+O��h��ښ�Ȃ"v�X����G2Q�F�?��\]Rb�!'��ۍ��r�H�$��m�^.���������?ǚ~��ߘ/N}��x����X���O��%U<V�z�)�DRZ_5q�\l��3:�DAUmtɭ�	�x [���������G�5�N��?!<?��#�BY�s`��]7���0���q�. ����HY�#/C�2Y�孔�J_K�d�/*�D���󱶊���>6'N�?��?CAӭ����:�k�b���z��'V^�s�ٹXA�7o����1]D0/�O�����%7�cr���sR����Y�R_0FF�ȳ�l1�r����L�h RrB�RnBo��[�l'�Ez�����s���t�S|�_��D�a���k�~�TW�$�y4/Hi]^v0h"Qn�T��u��~�T�P���j�pk���a{�a-f����q���L�2���X��W�8Y���n�eΐ��"b���jKHz,�b1;::�E���Z9v3+�nj�h�[q�\�H��H}�]s� 2ޘ��a�#��W�#V��]c�Z0�Q%��YIF�%��U���P��e�h��Vbś��V��᏾�B��U >��o>x�^L҅X�zL����{k{ks̖�a�0����x�0?�T"7]����R$��Ȍ��nm��'D2���m���Ӊ��̸9w�̌@�B�����/D�������h�@VC�����BW���ʵ��o}�	�� d����[�P�V��i:�p�J&��-�J��D~�t�Ҩ�b0�k?HɈWm�D���`�B�q�F�",Tj���Ұ�K�&,O��G��1"N~*zvH����f�j,�i=��"{�ޫ�hc��r�
�
���[#*�о��i�u3�[b�d�95��1�����hN`2!ߘ�7U�g���Ɔ0n�I!���'1Kp%`u��{8	�t�Pq�J����5L7!���k�R�
��{�~�Q�����3�6Z����,u�b���FW��$�����uş���ǽ`j?�YP��r�,C��w2����3\��7����C{�8Zp���ab]�y�O��(H�^�x����Lϲ˒m�p�k�A�@ِYCd��~"�&B�bd���f^hJ+��VԤ�0��u%
l�Bi}���g�/�4��qAVZ(9Hy_7�N�K�-[������;�o~� ������f��4���w�L�Cz��hyƸj@���H��*��N�FuRR������9�u���	�s�:$�ap�/} [`��ƧNY��Th�Y�)�lc�<;�L�)��K���O?��dd�Y��1��z(ھC+D�	�����TK+����̴��Cs���q����f���=�?��˦�[k�J�=,�W_}E�4@����d��\%S��F3%ῷ�Æ(ǿ��ar��_��O�SlO*�Ƨ��H�;��6ƩO `ȃ΂B��]�-hh-�xF�b-�ˌG�/̻�Hl��8�c�P��������#���H/��0WE��XC����i����SY/#w�6I�4��_����E�?��'�Ә&'�N_�ģ1�L+�x��8�cKgym{ޣ���9 ��v3�1R�b���UU2���_�~����~��ߋ@N�)~��z�
;G��l#���жVّj?".1�	�v��;�I��ӧN�u����x7"�69׋�i�@�i�Y�Q�����Є�.
IU�B�m[���)/4��7�\=.�5�x0i� � �Ӧ�^yۃ�x�ZZ���n޼N,awYV��[K��'7��� ���eI��ҚD���@*S�)����k+3/���I*5�
XJ!�-��H2�G�I&8Z�b�Y��֒�������Ǐ;�������G�ľZ.�v%|U5�H��D����>�췒��"<8?mu���|@X��F\�f) ��0�޻y�(
8% �|�ִ������� ʦo���?��/�ZQb�[R?��.ۃ�v�ݘ^rt�֝@��k���p��[XSfd��cj z ��	͍��MD�&6�$iH7�ڨMJ0"Y+J(6F��@.��YyVٱK��x	5J��E��|�P�i�Z�-vr�Bf%禢}(g�l����9ZY�<�Œ��tsN��[�r�M�nK����?`rpq��T8�'�R�����u��'��Տ�
d5�����qSX��	� ��������޽{+!�x1�<���eh���'ww%�z:�%2ۛ=:��P�_ ˨�HX�C�h�.Y�@��^}��˟��g?��a$��/�˃�.��#;c�H���(�jps4�A-��]�`����D��FGG�����(��������o< ��O~�,.��1q�F�ǅ��ѯ\�) ��\o���-o�ƒT��g50"���+GS
#�<G�`j�����[��ú�Z���I����b�^+11���ga{���:``"Ҕ�J	a�|�w��j�32�h݉�{=��)�?e��1���V�����(�]�-�M�,��U��9 �M��H3�z�^	��mYF��r���z%q�v�~Qh�)E�������>�xN��X#Hu,���@+��;{{{����➾&/�����:�Uk�hK��Z��Ȝ�F�h���8�ܨ|s米^�bm\�}T
��`l��֊����PՆm�ʦ�[���r�a��5����r؜U���smD� o�ì�|��ݻw��#�t�b��7�R>������kQJ��7-��L�G;X��_^'�ȈGA[ o�{�L���H��ugf
g£�R��AԸ�#%�r��m��D��ZMd-Ժ=�7	ޫ�|C�wc2$I4Ņ�N�^5�[���%���5|�
݄���(DW�t\��	h�����:�=!B�6��:o���@{�ҊФE�:cL���{]ک�|���N��(��"u����k�#OCQ�&�RTI�n���gSb�&�x�J��  y#�F-g[�I"�U��ƇS$��j����z�X1�c���K|C���d�/�~W���Ue-H��Pe)
[Ni)}���������zt�����?�d]�D�#��oR�l��U�%z���D�����n;��^Ɖ(8t�5~#���H�t-	5���0Ve�#��]�ҀL��V���i�#���j!�R������ͧ�'�����^�|C]HXuf�rK%J��j˭�d��l2��=0Ვ�3�gq:�6&�Q\tC��-����=��)6�_��nh����B�c�pv������p)W�by6�\�8�����]��⚦��K��������DE��J}�Z�U�(_*�{%��>��#�j�YPKc�b4oL�A�|��&Rqg�B�I�e�0�v��MrS4�ä��B�YC�>1R&m���3E.+�2i�·͒�x8)WU$�eDV�wiU�yZ���
K��=�0jX9���v����Z��Ry���J��q�u��_S�ǆx��ր�1F�h�Q��AK����aQ�(T���Ky�I,����O�6y�1˲��MZ�?��l���_7D�E���l~v1S���N7��~lWmKa�X����b<�>7?DLlL<���i�3�'�'�7˸?i  �Y�QcL���h<���4���ԨtSI!OR=�v1-i!ꒋg:]k͌E;;�� o��b��t�J<�����4{�ꫧ0_�8懕����͛�n�VN��md�*~֐V��seggk`�A10�J��ݝ+!-<F��0�}��w�Ź���L�;C���_�!���",�+W��vϟ?��q�۷o��
o1v�Vg�~g�A���4��2O�Z�=0cp�`�)����c��A��O����7�N�q����l�Ϗ�76&��9>@��A�a��n3�"��v�6�,��nƐ��`�}���^3�A��(���!H�ɆT���o���ő��eT��Џ����G��ޕ�5N�nc؁p7b�=�УM��/�\I��BS�#�z�'59�K؈Zoc[D�gG��t�[Ӫ�0 ����\\�M��1|W�~��vab�$Z��.W��r��k�h0��D���[�;�G�Dr y��^n�p	�7�b�aw�8ai������7��뼮�|�8��"Y%Q25X�-�R�s�C#�� �yJ󚿣���HA#y�Cw��!��۱S�h�"%��8�"�5�����^gu�<u_t���s�����q�������q�t�M胅+���lS箜>yF��֑#G�t�?��Hv�spͺ]NM-���NKM%<k����9��s�Yݽ�5I���`<ju;U���l�h߻wox��uM�4���î�8�z���������J��ףř��
�{���R��vt��A��0Ϟ>�{=I*y���v<���<?���Z\�f��~��}:{�6�y�نDZ����]�����΁�ɋ�5�]�]��eJ�e7����,GD� ������	1��#p�������,s٨W
�;�L*â'���dR3N��<0"f8�DՏ'��We;i���#GN`y���'��C�m(�(m��&�QU��T����[����i�nj�ڼ}�6]��0#O7W:�)�ZF�,�6F#0x�M3HAõ�.�^7c*��xt	Ev����;wp=�H�d��"&_\\��&{^�5���/��;N:��ɵ��woC� CA�T�$*+^�;�����/�aڼ~��� �U�X��Z��@�^�{��1������u �X��h���s�S�N���&�y��'O\���/�o~�KK��y�����j�N��y��%KZ6������3˕�{˴�	��"Q:HV`�,���+W����Y��׾�ƫ�q�6~�g	�Z�9o�r�3B�������Lb�;w�^8{�,l聃=��trm���zyy��#LN��Ȇ��YWdu�3�����<Mx=�o���hu�i�9��L ��-�Pqkkkp2�޽{�Ν4��c�Vj�H\4BȊ�<6���a��35@i�鮨PZ'�s!d�M;�Oa&sI\v�8R@/?��q��_�7�W[&�z�eJN�Jp���@q�5J�S�kqc8i�U��р�����k'�]^����={*�2Ӣ��"SN�;�/p��s��~�����lA(���2�!{Dh�Ck�M�,ۅ��r��}���嬬*I�>K���XU�(��g��YʕE�Ks�T�gH\��%�K�@��>t>|aP!H/<޷�~{���_|q~��6#�ܰ�j
�����^d&%�C�M���q�N��V"�Ź�KI*�j�L*�Ps)l�r"�/��'#j�����T_/O�9���V�K���c.��ԥrX�h�K�Q{;C���B��7��sP����666p\|wo/��<���[.첁��N�Y=��)X��2������:�D��T�� ��*z/(�z�e�y+f�WT�`��^[j�%X[1�8�y�Eb�~��XF�CGv��+xt��dn넦+=zuzQ�p٬��7Z���R�r��uI���;�.c%���5'��f�Ƴ�_AJ%��*���$����0D���r�E6=չB�l0�԰�]�i��	�u�ӵ��+�9�l���K��-�.ͺ��1Pz�F�g!+�ge&�G@��,Q�^3&�D�ozeU��m�+���2�WR��'��`����mLY�@�I1ui�*��.�����2����<2�JpiX��+���3!͉	�C�:X��FW?��< te��u*��O����b�3��Ϙ4�й�)��!;(|ic(�[F����xf@6g*
�^Byr�~����שޔ�M��`n"�8��̔~�ν����3i:��7,�'���Q��C�[���o�#����0\
N=��Δ����߇��������=��cTC�Z��d(�<-Xk�l鏎�[*(T�l{���:v��)��F/�F�y4J�Mve����ǌv\�J�Va��$}N�u?�ELl��Ǐ�r~.dy�J���	���/����æ&e�����}[\��6�qD�8���2�������p���&��y]�J�>���i�*�{��P4���ȁBh@�Oޜ�����D�Bωb��]`$Aܠ�f����{��O7����©g��І �]�/�.� /TF��A��k��a��~��g짦��7Cb]d�+#��wN�*:�<��t����[ݲ[~?���3/\�<,&s(|(���b��/ŕq@�޻���E^�}��ɓx�BK��jF �ƃkB9wy4��u�s�?��Ћj�ތ ����I�#��_�
:[3k����C�����bf_o�r2L���d��\[
6�S�8%�%�LF�i%��Z���Ա�|~~QϚd��̪�Y �TSLL;���јR�`O0�B���Ұ�����KbG���/,E�̍�w"�EUۋ7l��~�L^`�W��Pd{ii���������W��ό#ӹ	��_t�+�Sr#��p�*�'��#�-\[f����t�҆/SSI�����k�~��`=�髭�I�J]!����͔,_�f�����.�Ǫ�q#T�~���u�p\���`�����Kv��8�h	z�@�qW�j`)����~��:1y�x��G���2�25�{�;չ!����p0�4�n݂Z�<f_��Kko8����W[X< �5ͫr���8{�Ձ�Euxv�hV\~�!�kN�	�����e&���5�ɝ��]v��ì9��yhNa6=IW���-�D�Y6�K�J�::^�O��O�&���zJg�O>�K
���.��իW�6���Eg��b��Z�
8=�9��쥒O���j����Ϟ=������O��hwb�\��(]�Ȍ�<"P`O���Ό���n�>��A�e�<>�6�b��I"d�P: X���v_Q�SQp�q�c+ǯ\���I��y[-�h9��F��Q�Ex��'�iɶ�(30�
�}��[o��֫����s�ڵ_���$�";�k�n޼9����8���ƌE�g�7���{���G}t���&�d�������9̎�h��{��n��s���mp�vY�-���~�i��w���oRO��|�t�%�#�R��A޷º_��4C*VWW/^�H�2�&밅�1��Ȃ��?��3.+x���}d"0fp)H�>E��I3\���w���,�~���/�9Jfa�*~��]hQ������_�|Y���"�Nh# XHp�&j���·�(��W�絺�ϭ���V#4���8I��-�\U�7�,���
�ɤ�NU"ؼ���:�荓Ge2܅��G�3E������Y�2BN�8�$�b�:��D�N�³�8߿�w�w�)w�&��t̴`a\^ �\yC�(�X;�B##r�̵b�BH]a�*)?�pr�c+~דH���x6��g������0�jt
:�`d�dl�.
���XFhr������EW��vE�'��~`Qg�E��\�L	��~)m����ے�c�*Ϸ�T����QdY��8G·F��s�.2k����rS�u\�F#�$������{)�2�̉���t0�ŉ��4�<f�y~��<>�c�M���E�nW�Wi \g��ư{~DtE����>����0H��<�Sh��ss=ߤ������C�
M.�z�0�gˬno���hD��3���`�t!�ע�0��ez������5�������8��qM�T� {��/�,���5��+��9����"�nP�?_ԙa���9�`!�{�<�e}���jOS��dy�h�>�s�cW�R�g����u�V���KC?S�OƂ��}b��!�)���ǆE�V�^z��9��d*V	�8���p_YHu�<YSD$U��dѮ2��ǗvZ�X�\:p�8zyQB�+�UJ��H'ayA�Uז{�DB��Ԑ+��s��B��<��<.}ڑPD�3��`��X��XPRiD��*���W���ͷ9k�X�
bIJO��#������Wa����?s�SF\� ���@jSU��X~�m�[�4�gq�ۮ�#�* �촦��lS���y=a�>\X�5��hAK�Х��Cq)��-K��ai�ܖ�%͚I���I��z�!Q��P��ĳ2����5��N�Y��n<����nl��/�~{`����2�M)���}��E����AD�����S��d8�F{U�:U�n���y�	�9��
�T��]�{2�����O��9'�!v����`����.�|3G0�M��r&���Lj�ޔ����VQ:�ٴLG�H��D^�������T�j�3Ҿ�A�6��e���5-fY�# ���^�����h+�:NM��2Um�\�(�4�ȿ�%���`0u������hZT��s��L ��x,@E�	��0��فV�Ը9Ū˶j�^J��,�823���[	_YQ$E(�6F�! ��l����ʔ��5�0Cy����+N!�ੇ:���짖C7�ʹ�p����h^�A��_'Ϸw�ܹ��g��?{�>��h8`�C����"�m�7�	����,ޮQZ��8E׼���sM����}�m8�F¿I�ñE��*��6c=wv&8�q����픾w]�s�,ۧ�]�t��c�J��=���adX���c%�w:<]+~\p�a@�Q�Lb�:$Vb2�6U?~��G��J�vw�;���SOD1O��=���1�;�h�I�F�א�J ߒӽ�0��SWp�f
�[�҈D�T�S��I�9�l�m<9����vW��eSכ�+R��z�V��G����$�ml��_�/_��V�妖C^�HH�v�Z��!t��qZ���|�U�ki�aE�Fu��ݮFO�$q�5��rX_	�aHL��gT�vz�0�v1	[-3w���3$c�*^�����C�N���ͱLy��R�:u�;����K�t��1�nh�ᖜ��4]�[<�tP��[�ۙ&�q���������[��C���2v^���m߫����5X}c�YcXr�*����V���yT�:d�K�FKbmb�N+u͒���1����vF�o����#�O�Tf.I�M�ʕ>�>�(�A�*:�$� i-,.x��y�2����{�Q��}/���Z�hK�ȧ����w���ǖ��m�p��X�� ���om&E~��G;����NBC����^zU�ہ9��#<o�v4��Q�mu�r�O��~��f�p�~��:Et`~���GW?�t6�8q�����o��g_<|��Ï�޻wO�s���},B��ǿ���C�
ٗ:q+�}�A�`�?m:ˍ���6�T�Q5��m�i#f6p�J}Ea�jԫ�G��A=L�߬�zF�Aig�
A6c�v�S�Jf�k�OU\n�d���E4���x�|��7��s/�=��K�廪`��	��R	=V���C�BlΞ={��-	NTS�R�M�j#Z���m���p�����B�� �7����͛7��c=�#�ΝÍ]9Y�$�$Bz�9*D�������xd�ُ?���P�������⋸���ǿ����/������/�.p�կ|	��gy�W�N�+W�\���X�^8�=%r?������@Z��v5�����
.��[o����AE���S8#��D�7>�ϕ�B��������޸qc{ ��n_h1¶lk>�.���/�p���Cs_y3���ZmWcK�����y	����R �q���[���Η_{������U/]�:���7����mrhp�*�F�Yc��
;5I|V��v���0&��
����<'�p4���g����g�~������.�̲��u��$]���t:-�.���A5^|��_��V�u����e��%��v���R	��VR}>�괓�N�Z%M��J53�ť�(5�!��<�S	�"5H�t��9*f�jdr��i�@�,�lwYX(�~'�N��l��z\|�Ņ���/_~嵋7>�����)�:��f�_�u�XR���^��LGc�Fi�� �(�6���A���7oI�x8ҳÃ�`���dl%!���	sV ?=�G*�v~)R&�f�˔�e/�A��KB]�s�&P�}�����ZRMX
r%������5��0\'�C��v/]�e��9~l�+��d4�ݖ6�,ͥ{R��C�Ij���a��W���ܛ�9w6�T2fG���<�o�H�$������Dr�%���+��2�٨.��l�_�Ǝ�N2�&��7�L>]ݥ0�?�N&]>�0J���#Y�w�~��,�g�eud�}{���{��D�Q�sI�m����]�Y6�`�_eY���'0i.�j�*H��|#�]X�Дa�!�������֬L�����;���:pb���Vd���Z���e������*�;�-���`XM��D��&��Ǐ��:b�F�{�n=��JRD5�^8g�b9��a��aU(��� �|�;�/C�Q�OYч�g(�?x���")jCS!C�p%�B
 �%Be��|"n�&��ᇧ�l��QHV>�[;�q�B�#,e)�ʋN�5MѤ]�p�g)b[]vZ�*RMyE=�@.8�R6hw��I2�N�:��Q ����pU�q��D+�^�� ��~M�&l?�����U����,j�oM�r~�_�� �����8i'^`��L��D�s�H�>K�r"Ď��ۓt*D�N��W�FU�X>$頧�\���	�ߡU��L؃Xo2+�֥݊^I~?�4U~�V�
h�0�J���y:"�u�TP'�����.�J�֯�=\r�I��kY�.����7<�t�ha#��3.�)��ѼQk����������Y�k)�2�J-���{�ڑ�S-�R�"6���Ȧp8��~o�P+�[ͦ�ǰ��ޒ�*22�?)�̊r6���U<Ԣ��(9O�ik�Sg:�y��V�g@�7��)��-�Sc<qop���/�)�m��o/ƙ��Lm�������B}qr-W
�ç�2ҟq0�8O� ��{�~��p��omA'.̵	�ƿ[[���R:?�s��P�~��#�By�܋d.��[����}���<k���6��#���DG��H��i]i�F�1 �z��'xD�JK���1ba�N�"��%�qj6\
af���!��F�
�Cr����������/�� ��r��E���� ��{���5Z��cBP��� ��Ѧ���eJ4�5�`W���KY�+2R�e��N]��  �g?LX�/<&A�Rʶe�)��|m�!H�=l�o�Y~���ݻ���^#����qZ�Y��a���|�: �g�%�����Sg,�������+b��`ݨ8��������m�s��q�ԥ�x�)�|��xH�*".l�o�[D�a�>�g!ɟ�9��؆@�H�/��ťutF���+�+\�s8(��$�iÈ����Vli4x˵�Y�8#�v�������*��ZF�.��,w䶭ņSO%PHT��9V�Z]a���@��N1v�%3��\�u�%��������H�]Of'T��^?��V�	��̹˔C'�I/!J��Il.$��r�!iͳo�ɕ�s���Z�?��m%�ŷ)U4F���)Ϯ�������V���x%���'D�2��f7�6��e�\�M�w�v�w�X� 9�uh�����`1L>6�trP.//s���8	ڷF'ܼ�ځZL��9`Kl��x�=z��	N{���+�����ە�h#�}�v�{չs�֟n*>��TP�����iac6}� ���xT�XBu-�D��T�xa���z�@{CA¾���}A�g^x��K�^�rbU2M�����/�K��qT��H��	<��ps.^�}��@�l�%�L�VhBSqw���p����W�?q:�۝ـ]��lt`j��TΤ R`/� �Xns�b%Jc��K_��k��v���F����s�����=x22#8Gۛd�ÿy����@R��D�\:�Eyx�89s���T@�ÑB>E��\�t	_�������ܹ���pQ=��I-<7s"��E���y�'n�������W_}����#2����曪rc:âʫ��ŋ'��*�$b��C��E;�!�7�O�q@�'O�8sF�x0O#���*�/�;��������G�T�������ͻ��A���a%���?��W����,]P�g��ql�4�x׺&��7n��hx�Q}=|��i_���֪/�@�3ׇ�0z)�|�M|�k��z���^���8����[����ͯ��]�|�=%���(m��L�
B����+��.v�	�Ӣ��3?hB�>Ys���,t:��Aj��Lo8l�	9;T�M��'e��['�ƷAeL��Y�I�1�m�ײ"a4v�t������e�p��xh�twq@���:�2��e�/k١*p>mX3�GO=��Y�@��F4���&���ǕQ�'��&C��2<�QG�"�< >I0�N*�:pAkl�4������\��U1)
���{��'Ob�N�>����,�м�Z���
��2��E8���ׁ9��o��5�ȸ��?�8W�љ�3���MDt�42�j`�,�m��&'���)�"�	3Co��c��C�'5�_�W��*���e6:VM���T�:��fŗ���W�k;E�χ���Q``U��kv^�<���c����mi�u M�#z��7XeW�ˀcC��4�����zX!&~�����������x*�s%��4M9�������#B�0��Ɠi���( ~�?�!�Ae�\N�)9N<B�_��ru�a�<0 �{�e���l/��cܹ�}��l��rs)�=$��B#"��sk`�e#P��d�=fC��a�����b����\0NѪ]�J�\sqq���f����I��1��q�X��[u���N�43c\I@i�V���T�q��c���ܹP��CNx�j�5U��]jN�c�J��LqQ%�-������F�X�Ȳ�>E�G���³���s��0�ɰ�@�$�j^J�P��4�b*b��b5!��5�230#�.�rgzWu�$Nm/�o�gy%S�����/U��$6_��p�	��Z�_�����f����F���U�J����&Y��y�u;�4H��k�Q�.������VnR.#)Y��Cꢣt�b�b��!�/�����CvSj��(�Ql�������M?�{.�s��[��^�0�Q��O�6X:�+��+�����q���&���n�>��
U�>��/R>��d8��u��ʳ�JR ;�<��H��q�v�UD;?|$=Sw�<������8�[tJ��ڽӧ��j�(��(k4��޻�z�T����Yl�7k}[|���b�5��"����es��2KiE��@�%��L|:��1��ei3Z�����ZMl�m`\�s'��\~]iL���Yc ��J)�ꁪ��4O�����U�u$3�K�NwѢ;��5f�xa��aνvj�h�&d;�κ��.�JT�*�&j >j	����%W������%��8��`I�,�u�H�#��֒\�83�H�N%O���:�rhI�z͚��D��}�o%���Q��.��Ԧ���1�{֣Č��S�`�x
� � ��b"<�۝�H/�2<:Gߙ�Mb�Rp7x9��%���^�o�dw����X?���`��N���n�/��N�X�}�������@�%����SV�]��i0�4O�]��L~�(æG:���\y���ia=DrM�t���c�\H@o���皶9��I�T���g�/�"�íB�<x���i��d����`���0>e��U�}mQ�VV�
s磻�a�(h+|LB�vL��{��^�Y��iN��;�]��X��=L��,�g��*��Y���!t�����W�aEV,���qΩ�rfؓ�nD��9�H9$i�dyZ�I�%S��yB�3�vی�=�R���=��T���R�Q�:�jWU�	�{�p'G��U�;}����4紁lVQ�����rLS��KKK��(�q�k�c��=4�V���LR	��I/3�9�_$�!��Ѳ��Y�`,�1�^��PPYE-_�p2�T~*��R"
< ~���ޕ��6�=F��n�>����o�����	��_F8}�ۿ��{qO"�*'��xAZ�*��1�c|%��q]i���cmD}X���!,,���Uu)��6̭�308!�F���5S��¤5 �/��$��J/����mQ,�/��⫯�Z�9}=}�t��6cwo�4j��oܸ�o?s��l2j��*!R�'OVt��O��9*Z���^�"�2|jr~�Вx�B�JU'����_y�sgN���C����pA`і���wv�9LF���mD)ҫ����X@�y�ZY^���ە"s_�N��N?�v*�Y�I҆\��
t4��3�������U��޽���}��SX/��g��M��19��nYt���p�4�N�O�J'~���i�z�K2�5��o�v���?t���Ȭ�ِ��4���O>�� ��w�=q�8��d:���s�Dtn�	�#R�Q�a/�/�����c���:.���^hg:��o)��J�e�"KC�īs�Y]s.������u%":�w���Q����UI%��{�y��]8�HG��ד�jmm������祊	�@�'t0 r����'�c�\��4���_WV�]X���� Nm�65}����6ﵥ���o���^b5��X83�Q�
S�\A�����p?��<����������'�|�����?��#鋺Wj<�z�kF�Dj��
f���� ..�"特��L۳\��lze�R���t=k>sV������ej��hz
k��l�吵^_�Ry����Z�����4�������~weee4�[9zB%����A�m���߂K��'?y�w^x��\�~�._� t8+��~��O�gV|3�������u�����f6���>��F��c?�>a�McM	dӀsB�:�mXnmˑ�-�1�I%E�ݱ�ɬ3G���BG�A�0��s�Y.�
'0�ºW�]6s�B�n�E�q�pb�n��|d���������nЖ�_��V���R�d����ӗ8��lG�K����S���E8��b�{�q>��K�B?%���,�����u2�o��P��Kۆ0!����VTt$%dչ�4�H��������Ӿ	t$� ���*\  ��ە$�4=���<+"�(���ly�8a�w�Ϟl���
O��`&��ئ�9���?q�yY�<	ݣ�)Sxs�*�������� U�+N:�/�uK�(�|U��S0aN˹ع��iРkp�?*�c(�u��7��r�ɏ��:7�0I'x7Li�׆3F�T�l5�h���m��!ffc�<�)�2M��⇱m�2��azw���p,7ߩ�N	��J?P�������rE����N>�F5蚒��4��4�-.\��D�MM��w1^eFdV�|e��n�T��>�6��������.'B8����f��7 Dzo8$�ˏ�{<l�i;���ca�[��Ln�݊>��wh�s�0��pK��QsbQf���7T`n�)pt�30TڄP^��=�yXDr�[z:��W�ٴ\bzY��fu��yo���g@ ��<�0
���~Q���S��!��.� ����Ӈ�9�r�ڵ�/\�� />|�4h�._���c��.f��f�p�+�8Ϟ=�څ*�N�?��v�%�Dz'N��S�I����g��0j���v���<#�n�SXs�4�Ø�2��&2M�i�Bm9?����M�o@0O���e�����@�;QVD�#&�5W�Y�׈4r~XS}TV9(�rj���TVF����;N\�H��Y���8��r)�*�3ޏs�xr#'�{�Ճ`�����a� !��#��t5\�X4h.�������07�Md�ݗ�����j;�ťk]��H1;�i��yF9w�&�tlV������]I�n���E6K�Y���������;�H�6i����t�Xmf�RV/O�6n�FͩM��_���z��@�e-<)]j�>�WR��5��c�8y��́H�X1�N�8��"Z� L�s�o��0��HyX�&�3��� ̪ss����J=�4n�=u�I�w��9��p�V��C�����)͌�E{ݵz�.��s�`e�'
k��f�TZ1�0(+�n%a�T���u]�7�nO��cb����Ƚ#�c�hg�e����H%�����5��Fֱ�&	M���q��5.�K�Y-�vn]8�{p��]3�9H䣫��F�ɔ%���B� �+�i1PF±����#Ԣ���/��{<ݚ���G"�N]RvJz}�稕x�>ɍv=�a=*-gl�eΨ�J;Ba�zl,M��T���&ٽX"�Ǐ���-��+�7��P���Ģ��]��aV2��'�G�C�|p��VR�1R0�HZ'o�ǃ.Af�ȸ��q���8ϔ𥲑ʤ,��_X]��|��r�����T��a(ޑQ�
�����T�/j8/��2�^�|_*����( �;~Bz��hYZ��l�⑱�O?>r�Tg�0K�[R�i6K r����ߗ��tz��B��0�J��¢�2`��9	�9W�U�����aoC�S�N�no޼��w�y'se��	�oN�>݈���ŋ8�UΥZs��>�����R��g$��/����ジ�8.,�*E�B&HEX
e�:HgF�~�{���t�x�❻?����`��8t�5:P�3iH������ﮮ����;ׯ}Br�Ǐ�L�֑�G\
�x���ƶ@t_�u\���?���r��dq�)]Q�[��(���B��Չ�������/��/"eB�?�ݹ|�2��L)M=�;ƺ9����=�={����m!�+�ڮ���5V+�L��*�Aa|�W�|��r�HF�c��4�jޘ��:���mBsCVn����,���n�jG���(Oz������N�����!$�@������A���U� �$�m^;����(�X�>��MJt?�>��ڽ�����G�Ԩ3E�-ln�CQ��[K��l���L���q������Зp����]d�c���"AkB�X��ʠ�я~�#�z�(��*�d&J:?�.�8��pY���ۿ��~�3Q�	<���p�z���d�\{M3���seo�3d�)��n�ܙr�^��ճ������.�݇�/��>���ݞ:�@I����\R��<|�_���D���rQ�W6����R�o&�^��=��߲��1��Fz=�B!0!�J�>���O7�mc�H�P���GCX�����@��7�����er6�?�U�
ؑ���'ШQI�x驧#�+e�I��`�²O��ޫW}��<A%��హ�NV#��6)�<ˢ
�ܝ�*�O*�k��eT\lR�cl�ȯ�tq]E��?��?�j7k!�;!��DC�{�h�Oߜ%�<�/��u�ry�N�
�!���֍ ��+�;�T �)9ɬj��;���O[�QY�O�v�\w'�.!�Tt+ܧ|#EMu�d:R/=ti.x�.�[��?z�Hl\CA=�AkU5x��<��E�,ƍo��LS��n}�ҥ�<�'j��,O���ٸ���6�O JeQ]7Å�\ŦD.m_T��+1�'��s�cX�*����Le5+g�_`bW��s�V�Cp�k;�7�A�Bk6s*�Ԓؙ�>
tj':t�'��Q˒�+� M�:���Sr([$�������-�I|^�s|�0�X��H1�܂5�F)Ӿ0(�K�)��đ�� y� Z��=b4[Y{�c|��W��\u��=�K����N���^;���9�1�����NQ�t��g����}���ƩΥ��aM!3��{FqQy��>5*��'����7��q�(����d��; �*�����"�.T�����X�k�o��������� ��.ڳ�»�K*z<���N{4�<y�%�$�J�c"����b�fm/=~(_Q2��Á�s�k�O]���8U�XL��w�~�\��1� W
	���H.X����7��a��p�����)�9�آk嶏u?mk�B�C�0/4F�ַ�z���p3<�m�Bh]��~Y˒��yM�Oa�i�q�uk�Z��d��/�Oy2�QL���LW�f)ɀ$�n��7I�kVHk�x��XNu�H��:�llS���&�&ٲJFU����13t������6����H��vMF�Y��%a�?�Q��qY^�=˰�7�b�|��~#L``� Ua|e/+�dr�'�2M��2��� �tT�WH�c�m|:����e�-yp�RJSX9M�R�'q{�O���'KD�5����'ahe�]#��U�)�������'�g��u�b�Q�&Մ$��!�����;��,��e(�̩/�Ț��c�8\a�;�0�g2r[]�x�^w���`,D���q���Lq�V��!�}�V.��2��FE,�q�_��K�v��Fl"Z��"��Af�]m��SZ�E��8)l� ~L�:�^C:ٌ[r��yuX@X��S�e�������k8�ӽ]f�N����a�K%������v�R��I�z&5���f��]zW�uR_�R<��ѣG�}}+�E���E:��髩L{+\>3b�.��ɦ
WDX�f�s����ҩS'��g���bՊ?���zq�����" �Nן)�~Kl���{aFT�zr[31�:+�'|�z�,U�jw�I[�������ɽ��Z�~��2Oҏ�^��c��0y����{��i���Ɠ�M]OO���Y#U,���� �J�<��i4���U���P)�������[�:Q|Px��.��3POe�0;]m�0���5UՁh����ڲ�=�QZ�ɞF��6�%õ8w�̙۟��{VO��S?��.�c�>}�1��#��GP��@���'�p�ر�w�J�N�P9��EE�?~&���tV�8��C�=r�J�m3׋Ԝ:p�ڣk浳Y�`�ܙ���@[���RP.^+ހ�������2˳�d<���j�#||B�ׂ��zl���_�݁M�{�+�N�������d�(��v4'ɚb�ȗj0�X9q��1�s{g���]?�O�����pw�����'V��������������\[�Y{<ʑtd^�(CH��˗/��n�����ʊ�|����j�*��'#,�slX�%����S��������}2��G���YJȩD��<���~��^�&�K;�[CB�=�����g�}�g�g��z��Y���{�=��3 �.����^x��ˇ�te��Ǐv����0_�ȡa�5�贐>��-�mll0C���j'O��;!H�g�}p6�x^�C���OY�L=G���#|��#q����؟<yR�P��e�R?�|�.����"<LD1�#����^~�������ЗLn�B��ó;�L�hq̬��
�[�◲1��9�� �4�gaH=�����}��"h����%���K?a6�o��t	��z~}��������<�Ѣ�DF��*H���U_�ĞQ��$i�GF��w��~����*�j�jMݶh�C�pA����{��ޑ#G��zH+��|'�+�u���S�S�==���m�u�%�q��I���93��W6^�M�t�|���yc6+7��7�6��[wZ���fss��7��?���o�ʩ:Z�v���G8p��x�6/����?�
�K�T�N��@�2F|g
��޽{;;{� �Ogc� �pVYY�Q�b>D��c�dY������3�ԉ\���'pNΜ9�������y1�U$Á}�Q	�q�^.�~UP�a��ڃH�IvF����v'֨O*@�`���N)�"1��%�]_m��0�ݲGUM�����B��F�
uaq��x$yO��C��'Aĳ�H�v:�����)]�4���&#1�IKr<��Q�E֞�ą�p�Ƽn
�ǒ˞%3ʳj�23�)�>��괽ȗ�3����҈�HR@�֧�Pg#
�;�?~ʥ���D>�a�x��w�.��u�"�ಘ�|:� �[eӛֿ�< ~���[��L��C��T:�Sj���._i�&V���r���&��N(�,�!/u%�0rw*�Y���Zê7Vi����#��[��8�^�9Ae�g�x<�d���]���uf~>�<�fx���J�A�P���<�;�����7��5�,{��m�8ʹ/������J �p�}�P:�}UU�	Jҳ�F�[RF�����F�ﬅ�/��G�+[�8ǽ��u���%\
ճ��,M���-+�U�{S�:��s�Ø���@����aY7���hvOm�AϞ�p��N�[���� ����*�d��
�4ȴh����Ds���.^�]L��Yz���;���6��%R5l�p\T� ��]���_��@�D�����`,*U��<�hx�7�����SX� ',�rњ٢�j��d�mrc�qYGr�r���V�Jc�q�yڧBAU�&��ػ+��,Z���4Xki�'�#+	�=�װ�x��_�
|��F������Z
@(�[O[ۼ��ځP�ie�pf���r���K(̰T��	�&rx�0�3����-�,��RaU�*��Pj�WT�O��p�?�n|��g_��7  ��:"d�v�S��t��LJ���#���0@����6��<��jN��I�&�����\��AǔPd��|3��i	:CD��F��X[�;��j�|IwqZ;�0t���;��k�ȱ*��p��H[���d��#�r!������"���%Miغ�̟��
�kW#�$LA���ǩ"Jh%}#܁�L�u~��)mjje�n�"\~F�<�X7�Ԙ��l�+-F6�@?�*�������g�<o��ꮴ&.ȸet�x !������ـ�i=�:!�˳d�����!��"�x(x� #�f��3�-OA���;����0mMŘڴn\�k���f��*�>�����c��}
C��Z-%���G���	�r��a"�t�S�MSʉ碥�͸1r#��&��l�J�Ď���_z�U/�f����:��gs+5��"�/�<���O4q�/��|D�O��ˍ'����`B��\}�Q�� �D�)#����������Χ�~:J��"�ӧ�PV�du��3J�S29�#k�ɞk��vi��ބkH����Ӄw�F��("�I�A��kؘ��l)�.g�+6�ɀ��кu0��9V�(<�_yymm���zj���Ǐ�-�i��]*$9���0��!TÓ��,C� �b��������i����������L���AʀvjkѨN֧}��pc8�)�6R�*�<��䃻�#���߼y��h�����'� 5�׽�uW�sK�;��\u�9���'[-ݡCK���������,/ԇ����������o���?��?ܼ�9�����<J�\����x|�֭������?�#N)aڋs�Z`���d^��$1��y�W�)��<���f���4��/�(g�K�`	����21��E����!i��?��?��?�c~�k_#��ҥK�84��8�b�m�r��ս��q�X�;w?g������~�@Y2�{^�����o~~�������\�-��L2�јu��݅�<�� v[Ԡ�b%�x�w���^���;ა�;{wd�T���G����"��'<TPH)���e\���D=ݴ26�05LuQ�#�k������4�����M+�⍳�c�=M3��|g3z/45.{�S�Ҧ3�U�����n8�n*g@�����;���	&��('�}hc��-�k���gi�]�e�/eͪ������_��׏�/�>b%�Ua�_�]�+s�K���rǄ��g.��M������)A\�˰�����~YGLmг[O�lW�$�[;?W��נTk���\�S׿�x!H�c.>�|�r�2Q���؀L��:Nh���ϡ�!�>�kZնਆ�xJ�B���,�������"N�n?����ܲ����� f.<��z���H��������bUq"�I�~��LVri�͋VG~�K��oJ��j���a� ˋȯq$L"��xZ�\�~#.~F���Pg�/�h�o�kW5��\��\��IEᘞ�������a���e��p�	�ީ��̷td3�F'{.��:���.X�om�QK�F'��:�����p���9㰙M۷��'sZ�z��O�]�X��y�C�θ4�I@ϝ]��e���O>�d�#��C��T��Ϟ�J���f�f
��//��V�,,궾�:����H�8yV:'�yZ\-������x�,p�������F����I�ɴ2��rt��c@�be�~60|M�".�P4���_#ɇCe}��u�SD�����C�p�-��ndX�A�eT��]�Fl�N�Z�qK�hX�T{Ȣq7�w��Bm�Wiz����G:�{�u9?R����q��DR���0o8�o�ئj`t����X��0_�UD=K`�:>>a�E=F�b�չS�l�#w �,��ƜL�š<���`q� V^,��&{��盻U�u�q�t���/�C�� ��rȣ_�:��7�3�Z�����{ӧ�v:�(��]�L�c�k�,e�������>�V��8+J��n
� i!����x�������R��5m_׻���&����W���5�p&a㤸j��}�5J%��`N��?�m<Ka�w)]������m���V�@.T�|��2cOwm���;A��t[���x��(T�'N'�SB�d4W5�GX�G O.�lﺬǟ�tZY��yW"HʣG��>ڡ��r�u�����J�[,1ɨ/��pw_{�s��F��/�p�����GNk�I�O�I�u~�|�/�����i�(B<��b��l4���ziǖ� ۈ�nt�,�t�״����������q0H�[�^��z���ÞkOt��̟��/,̥��<Vޓ�r���V/�Yrzt5~�?����;��x:p"cuͿO�7��=cr��'���~I�xR�Ps��l2�<+9L纝�I>|4�1����l{�����᪘H"�L�×�;�m\�n.5�
��������nU��Է��|%k��V6�b��GIjW���^�F�rIEkX�߈ۃa����^aLg�v��=Z�,G�
�tG��5eRݘ���LR��L,5A��}6=�ވ�th��0���B�0��-G���DjT�EL�0��:��7���X������o ����A'V� ��׼������XP1�[7�Rn)uL�0�\��.�UM$�8X��z�}��5BI&�sc�����-Z����0����]�Z�:��)��*����>}����F[9���N�d:����V�u8�NZ���%^�`���:�ĥ�z,�x��ݰ&{��{�����¼r�N�2�+Q&2�M������~��ƭ�&�����<�ׯ_���l��t��dJ���^�r����a����?
c���ԁ�/Ԭ��c�Xq�q��¿�9d��9�JScL��sk�q񡋫�'SZ�6}.�,�6��$"�����IVcV�}�u4ȩj�M�tB�D{�����p������E<p��%D���6�Y�EQ�=sJq��a�	�X������?u�$�<'�V��Qt��Y9��eOa���_=�����cGq�&���
m��69�!?.\��l�?��'�)~@8������Ƴ����E�u����ln=�`�����TZ�#������WW^����ɼ��i��	�����ې>��x>IB!x��a�p�z��8[xj~`�q�`����jN	�����[x����q;�_���J{o0<{���+wZ]H8k�r܊2P��_��_�����ɓ!r��UF��jouH�U=:�x�_��/��2�8�����eIJ�8���J�N�7�^���<-� *�>�M�y���7n��/_F�{��{����r�\���wx+���Ο{񅵵����n�=7���قm�L��>^��ф�ώ�Q�J�Z)B�G\O�ۓ�2tg0������Ǐ�C8�@+��{�i���'��c���F��:��鶂����_8}���s�sͱM��<~����H����#/��R��//+��ĉ�KG�Ε�{�7�=���2�^ҕ����V�m� �k�u�C��A��k�Fx�V���ڥ�
�b�t��AwM'��}��.,�X]�JMj�a��Hf�!J���5<|7,&���E�Z�m��d'��xV�'�38�Ϊ8�L�������ֈ��������|��/�+)�ٲ<u��T���{�W#��qZ�2��+���
��<����j����IX��T�KH9n���`Ґ��&]����}�69ĥVu�:K��#]����W���7���8���o:�jV\�r�M2I�0�)��Q6�qvV��깮g�Ll��@���@��e|og<R��E�P>���8�����rX9�Bχ�4q3o���w���v����'O�lW�lo��ܹw�T&�Y*�8�=�<i�$T�T���U�a���?��iG	9�����Ț*�@y��u��+�ZRif�W�O���@sG�T׳.��(-eK�<#�������D����Of���γ簒��� �ry~���y�6c�C�A�^���2������P�E<�U�{iQ�w��i�;_�3���q2�N�,�,a�Qs�F/pР�r�@���*.�CQ`��N+�[�$nc��8W���D�Fgq�4Md�g�Ƴ��9*��ʐ��J�>rr��n�����B3��㨋�K�:�W7�:�]U�k&����rx�b2��_����h�]���劅uP6F˧�T�p��]D�52��&N�������G��Z@&>�o)������`�-����2)p2p)6���pD���V_Y��ٖŋ��ƕ��eh�����Ga5��ߦәӆ�A�F5�d�Y�ٳ�K��a���uO�d�"��ZG���P�\$>��S,t��.��B;1��],�Ig��<]�� 8\�=x���R���ALNA,���S#��L�����'�'>b+�n�N�W���{����Ը�Çe���O�V+��3�xAX�O����Kº	�,��z����e�F]Y��ټ��_�QP�!����<�񌄍a���ꌰ^��']b�3j�JgbG��Җ��:pĺg��]o��_���Rރ;t���3�s՘�h(u�I��Q^�/t8�(�C�2��Z����S�x�;�l�� J�=˥���_� U*\*<�"EE�QqN�S�)ա���7�(pw8�إqy�y��x�z�?���0�� ���A�B:�S\�mC��>���4	g��8���IX7~�+1ğo�:��]N�h*��Fl��-2�J�$����̶P`�����X[M"S̏͹S����
�`6����@�p��iq�q���f�e�X�"�)����R�����~-���Br��h�ল~F�J�<�Τ���3g�য়~�EX__��I�g��t�ڭ:���iwihkY��n��-e2x�3	�a�T!�Ы�Z�:�{������*�k�0}"`ڄHSB!�S8��R#1(3�KIuJ��2VƷH�Y�mc4�5��ܹ����b�Q��3Ż�mS)���݇(�f����O�y�	��;U����(��Jޟ�Z�r�?~,��0pya�M�`q��Ĭ����C$�(]^]��b���v_w�tH� ���ņ.���qVLd����RP5�H�m���έ[�R��Z6���+jO�T*���q͏�^�l��jE�ϟ���<ɴ���X0Jd#�'{��a�v$>t�h2<F����p|��1�*�P`7W#�E���Ωo�(�ѹ�6}��������d�6����������Gݿk�7�x�̮s�W�U�2�ME��f�GF���|�p�T�X!���6���<q�dU��"x��N��\X\�������j�	��j��i��]ŃF���3ywv��⥗^�Y�s�ST3�uƝ@�t@��ƭF�����E�̃�cE��u�ԩS�Ο?/]��7.\��d?/]���o~���W^��?�����FH���A�]K���h����pf�w�}�A|�իW񽈂���.���O�Ka1S�d���e�~��]w�s��T��׉����ܾ37�Vπs�Jc�e-`��q8����?�{���w�����;P��>��^æ�\=�%�:�T��gt�u�SHJS���;�G�B���.�L"HR	��G� '��ǳ)��X�Z5]��'S��=�D6����p۸xIY��U\�y�ũ�E�;r�`��Ft�V%*�����`�WVV>|�f�V���L���%)��+D�=4q�o�j{�FᲷ|�A"�졪�9�Ϊ2|���XbÑ���ئ���$�A��X1�*A�t2�C�L��
��0������K
�d:���řhq����ۤo�	��kׄ��^}�UO1_����:�Q�f�&k1h��x
菅>�`[�/^d�����":y]�������
���xi�����_��`8rP��jP4X��/��$^S?��ahH܉4��
��K���A���2��_���m|vowH�W��PË}N�L�A�-�+&��YJ�c�jN��;uZ�Ыm���~a&@�[��Ӈ��}�L&G�>yZ�]+Q�|p�o8��9�I~)��df31�Oد��['���R��,��c$���}� h��G��\U5c��ZV��<��"_G3���A.�n|X^�9�P��?�(�	�R��%)9��+�^%J�0�t#&��s�^�m4����^5���F.U�D8��B�V!"N�)̵��e{�SM^�دi�*����rm���ʄ3�=�FO��>�����Õ+W�N���ݼyZ����s�{��N��,�����ݖ��uJ�o���;lw�L��Z��Fbo9{���ݖ�;t�f��b������f���F��*�(��4[`�8
�8�ʛ��>�]<�h���&ӧ҅��=�>�)�=	Jkڍ�)dK �=6�p�G탥	�:��$2���:0ύ�
�  &��C�x'ѹ�B����&�8�Jl�P."�GA�~�K��Z~�ו{���+/�[��D4E���ftZp.q��&i����������W��2	�W���j��l�/'ڈwvqR3v9�rF��v]gh�p��Ab��"�5��|ݡ�]��bg�)UL"PYKG��"$����	g�$X��m��H<� 9\"�Etkp)�h1�+����0Y\8H�j���o�y����ܟ�eV`�$U�lso2�W�
����<E�=E-͉$�N�����g�qҎo2Kg��B)�;ρP��h:>�L��(OW`9�,��ʟeB�"����Q�R�́��p��l�̭�Q�F
@-���<�t+$0OG����!��S�Ee��^�[����	��x�V��@ǅ��.�NA[�C�_�+��N�_�w���2��x	���o�Q1I+��;�3|���u�O�Yq0��k5 ����]�W����B�/��I�*dԀs����6n0�%_{m"k1kwu���� ��TL���� ��㇎,��=t��g�}�R�j�m2���sg��P� ��[n���Z�Xh��4����Pj�o����ZY�z�褮�p)�r��SΗd��B��-��H��UY�V}s%��xȄ�����q4Ig�B>��k�	����;�?��� �TE�j�{ň��m��B� Y�{b�s��Ύl+�yρ�@����a��q�_Ƨ�������G���tA�$tB��%�0O�L1�x�u('	�%��8�5U��d����l����o`�<�E#�ړ��G�߫�\p;�hr�MV��;�m�n+qr␿���3�$3������OΞY_F0������'���'prcdj\ή�8��S�٪���4�IW[ �"��w�Ah���n�*�3""��X��z��,��u\Ν^�pF�-_� ���`�:��8�K�mb��2f���!<��3��S�ˠ��(��x@�?S��.��R�E	�7?
�D����8��nܸ~lN�7'aO_�	xb`tY4;�S�����ʳ�k|�=w��C;ꉦKK����$��˃H2���~�d�Ν���q�ڝ��<o��GAZδ�^�������O���>��	.�mwC&�?�Ya����EV�p3���TS�N�"W=sٱ��̌���Ƅ�VV�tib��]~�i�Ry�@F
 t%%����(����}f�YA�J2��n��Ω��h6Ũd5�Ի���<����A�~k?o�,����[�>c8!��Na� ?���N��W&z��o�٩ZC��7�L�O;���ل����>~��	���� � a �ܹs� ��
Ͼ����]�u�)A*\ f�^R�;��+�?~�z�݊W���OB1�r��6e̋�!��k̍�Nd��Lہ�����h�?�������ŗ�m�:Kaq{���%����7�>�v��Z��;_�v����o��������泺s�R\��)����_f��[��������[;�o�n�(��ʨ���~`���<�6}���ƺ}�+_�m�YυC����q]�7���P6_ȳVb�PX� ��$�� J�`>�������w��\n�֎L�>�t�/���ɓ'�=FFj\*�LY�%��>ش��mڎ4�2|c��������Խe�wZm���Lg;�o�fH��\��m�Br��������F�D�*O?�7��Ǘ.]�|,��p��*�tSgڊV���xcvbFzgs���Q���p� !O�lY:�M�@'�
�#%�b�
dQ�ne-��:+��h4�y��qY]�3r��r��G��˫Q�&ƶLs��3V2Ng�F�:6����K ��6��'韸tu��^�;�j~������|�+���/A���l���?�կ~E��3�ҖF��ql���c_z�%�˴~I5�`�|
f(���T,Q2�j�S4�L[x�\F�[l1��� n�Jk�p	��ث\��F.p�e�f�E���ڸdGl�P]���>��U�E�M����Y"zQ���s8ss��`o�PVѯ���G��#P#��9�Ei�XQP��R��(�=�p��k�/:s�����)�L?џgْE���޹uO�,s���;�ե(��)��liD���>�O�{%0��;e�˪I�ͺv�Z�
�v&�j�z@Q������/M����6�)��"���[�xSʩ���I�^%�`k6|g�%��9�8�0�~~&R
!�����+�q�Aj�C`O�hdc�r�Ԏb�<>����G[�sXy5qQkQc�,��6(�8�,�JKF�d���bK��.g�,�r�g@�� �^D���Y��b2���w�?���έ;��6ܸq%�!��Z� ba��V��m���l:�N�|�g?�15e��;��=����&�J��%1�K7��u`F�5��hY�I}~�fh� ���p��������U�椅�b�q��"��1��\��p����x��2��+N4��i�O,�q�g,3.�A��8U����MκAnH�P��5ȭ��*�#�TF�'��i5k�4q5��`��
����.�g���[������w�%4��ZJ�(f=�!ru���ˤo���f�^�;�CNܳ��5+����D��B�_!L����p���$�YX����V�|.u�cee�$���[�j������ß��$��e}f�t�����G�4G��$�x{r΃���<+4��c��T=�W?�����d�	�Кd�l����[��b�.48�E� ʍYCꖺ�$�bnӄC���S�gL�_)������e��~,;��3ޱ���z ���(��I�%YmKNd@�$v���?&ț���?*d�MM�L�%�S�����ꩺ�[w:c����]��� ��U���}����kㇰL�6�w�����=�[�îC�c�iy��<n��$}��=��������Q�+�W�dr	8?wi�_���ݰ�4�x�L��ѩ�%�x�C��Q��}���usx_�d3���L����ca�EO���:|8��љL!|#Ա��Lrc��q;�N�����0�fwe�ҹ+��J�������К���[S�+�$�?|�̑μoe� u�"�o�!kCS��V2q��'u��sF��he6o��Ď��8���s"꙱%{���>�Z���1"ט"�g"��u�΄���uH�r�'�|�I|��͛$�`�w!�z���`����	VG
��dZ]��'u:���y@�~�7�y��y+���������H(4ӎ�3f<���"u�Oҷ�jJ�)�[<*��޽{���_���P��t�:˰}�>ϼXe�)n���N"T�O�5���Σ������*g�5�ϳu^,m$KJE�$�n�Y�"843Rc���3	ޮ���Q�̗��#6�(.un4��Q�Ҏ��`H�?����ҥ����d���*�Ve&+iLR⾋��p�v�`5�Ej�8�<�SCj�f��S�JZ#D���煟��))xZ�*V�e"eoO�M�O�A���P�<yYomm�<�ɴ,��g�1��#=Px�[,y��Pq:��Y%�8�Ջ��w2��s�Gf�xL"�dJ��.$�xT�\��Z�\&FɣJq��U��p1X���P��\KJ������X�9+U
ђ����K�tu5��H���W��c��Cu?���ںO�W��>s��)aO�r.up �9��.�,/��,��`�S���1�y�.����<�3�d������� �Rͳ�����n�8$��F��ٳ�����;w�����������k׮�oAA�����O�KKA/�nE̊�=�~���6n
o�/��/ �����w�1�Ko��wxΥ�e�~���F_��p��}�s؈w�}:��;l*+���F�V�ӟ�4���믿~���ңJ�ǧ�$EiME�U��rSY�"m�'��Ԣ"��y҈G�|�;������A@��D��29�������HZ7�&�m+����j3��N?�d�|���ɝ�}l�
����4,��)G&mĸڂ*s^�E��eTxο����%�����я~-���X@Ǵ}GЋ˫�o��6�([�pe<���
���Ϗ�Z��WI�,b���C��m���8�yӡu00���Gi.��7�{���cq�>2�Lad��q����::�*�� V4������-+�y��9�?2|P;�k2�*����1I���~��:.���/��A���8Y#�LO՗�̦,v�*��!�����w�O=�Z�Ȃ�%3VVwu���ߛ�3W��/�M�l�@㇑I���z�ڤ��( ]c�7Ak��V|	
� =g���e�QhU����n����G�05!��nWxN�e�P��9����=ľ�O41�I=��@H��@��p�i�_��U}��q�M��o�䥍�$� �66$��rkkP���̳��E(�:f�>�-`�����B�wv.<q����8�yR�_BT����a�:L��j��<e�2�8�I��J.1�q�R�:���t��<D�}o�����GZ{�'�$�[sX���#W����&#�6���µ��h�l�w�p��8�'���L6B��xaZ����Z+
 ɃC:6yPBJk��Հ��x����h��h-��K����L���OE$���&)�ihE��*��^qr�Ms��1z�r>�Ҿ+�ܒ�h�;=5����dv�����Ͽ4D���NA����"Cd��૖Y��\x��u5��s�SAQR�/��=b�v�����x^#�W
,��?��;A+ ���O&ii��.ʵ�b{0�E��1w �TWJ�%aXҁ'Td��;��Ȫ,�+DhpM�i��1��zlϬJdӁ�(�-�J҃���Ù���;MIn,�T���<Zn��Z���Q������S��
b�nq�hem�'�v����a�L	�6�3�_M�cZ���u"MW�p;�Ó'�cvwz���x6��Q�Φ#�������-u��g=T����{�RE�u�.�:����i�H����e�L&%�;�Ο��ȴ<�dZ��n���eT��� ��;m�_Z��	����R�3Jcj#��0�]��xv={�5��h©p#+�q7˦}�G��g�z���Nv!��(jaS�3���a�<��iF<\�J_Zֽ�7��E����U30�%à��!l��H��r�����F��8��RuT��D�&���v�������U��A���8̺BG��STp�x�3��1LA�{q%�GMV]R��d!����*ըt��*8�Jb�Ŝ��tm�te��N, G�)�;:̨�hE�a%��l:���T��XX��Y\^^���]��.u�һ�va�qg���xpU29���"Q�5��u�ꘫSR8�zԌ���
���p����H���#��A[��L��Ȗ�a��Ѿ$���I]���йrpi�g�̘���Ʊյc���ҖI�Bk�P#�
+�a'��N�}x\����<��s�2ϖ����������D?Խ�-fjk!y�����v��gB�b�U��d�e�Ig��RDR1�]v�ti��l�'�����~��)���H����19<h�Z��L���Y�������Ȭ�K/}~?i�x�������)����!��ڥ�2�hd%=��Hn�Lv��
7|C�Qԟ�H�B9g��s):�ުUF&��0�7_�v�#���T2��1I������6�ů�i����,s4�G�
��ۣ��յ��h�u����߽��Ъ�4Őf!zI*�-��x�l�'{�:̶���+C|%U��J��^<�����U*�*_[[c���[�2P��cR��u�q�����u���nJ:��Y��}z��}���O�;}���ޠ��B���e��r%o�c9��rt�9�����+�I˂�4ө��Xj��x�%P�18n��AJ�^*6�	?���f*"�I��<8	�T	T���Ni��޿����n~|x M<E��ŉ/��\ڸ55,N�7S��s������ރ�A�������zoo6�����۷Μ9�֯��K=��rL<�f�����.�Hh�o��:N�S��D
���[[xl4�=����W�2/^d��E�S>fs8>s����	�v�-���(ߨ�p#��>T1<���^]�Ãƭ����M�K
�=��>|�?^�ɧ�ʘ�g�i�(u��Y^����NCy,Ľ02�����V ~���])�L����T���8�������l?���q�SI̕����!j_QB���?�����|��ɗ^�/Pt���/8���r�t�����cY�ω�y�7 �82���g�7oޤ���ᩥ���(Kqܤ�=��#X��̉�,�V�ᵀj��L���ի�����}��������:S������kئ@2��e�
!�t<���=7�5�3��'�b˰��>��|�c�������1DJeΊ\�¦!�T��eگ��&ub��`a($c�<���V�W���dH��T,���b���[7o*MP���z}<��O?�3��/�������G/^xbt�?�gu���qX;����E�����6��U
k`�_d3��֌�И
��,oTkeã=b��d�j�r6I��YϦ{��q�Ã=�u!�:R��w�FoO"���&�w�,сl�V�x0��lI�[|��el(�a<%X��$��U�z��N��b	�;���g>�o|�8\6��-*0O��2:�#�L�:p�X�l,�3Lh�t��BP���L�&�~T�O���I��O�i��2�vlY�y�v��#]m)?3�ޤcR���6P@K�0�Ș,Rh����@��f���h)�w4T����J�U��&�؝;wp�+W���Orq�(jf[��GNK��'�bP2��ȧ��N�p7�f^B���VB�d6O��&1^oey��K�KL�Ry-sfe��&��_��%(�Ϛ�FyV�2V"ϵX�0��{K�+��Wgؕ�}<��En�m,����^�q q��!N�da�(d�
���G)`é�+�1M�<gP!���͌n2����ϟ?�*_´(�4�kw����&9i-Ƌ�U�W]�&t5���/�}.Hh��Z@J#���܉+Hk���å������x��3�Cr`ѩm���t��s=
���bX�"sX�aw%L�s~P@�A�
*�l�`-��=rG�gnVqx�禍Jm*A,�����}�kQ�լ��*�}�y�ʦz�:�S�Z`YW+�+N$U��maaC}#kþ�FY�'6$]`8����4"�:Q�f��b�h������M����5��c�W�D޽v�W^��+?�/5C%S�=���NV��m��G�A�C��YHO�һj!Ș�>�m`h�3&���|4�˟�Ա��5���w���� 6������SH�ۻ�&��Sof3Y�Ѩ��w��p�HD��f�+#�t+kR���""��?�W
�T��f�!�d��;;{� ?�yW"�I��cS��¢+둟�vS��h��I3��[�/}��PK�Q�yP��/�A"BV�����gm�`KV�c��imh>4��MF�μ��m<Gb1����E�KHh��K+�뭫��c�ֆ�^\j�4T>U�Ҏ��c�Mb���>"z Q쏖�W)7y�Jm�;3kT�4���C5&I3�ȏ1\(h����K���1Qc�u`9#��;ݔ�������red]!V�k��&D�@���p����}O�>N �~�G�OeVb`��G��s�HjC	kM�*1��ױa]�҅��/t� �Pܬ��=9-��"�p7oAbɇ5\����sJ��{�ƛ���zeu��ҹ�!Qԕ �,����eC"q^f�5W�M�3�\WY*���3�'#�׮#a��ן�2V��a�Y�X3ým����yA���$5�����"#vd��#�hqh�
ڀ�
���#
sЄ`$֞�cR�_�t*���c����:X�c����OQ^fL���H-�.�C�`1�E�^��N�(l53��/U)��k�=���'�<0��Mzu~�Q����n<~�<>���+�L�g��ht����r!P��v�o��Hjx�$U�Kv��SA֪S��ٝ�QV�����a&Bi��ߺu?��\k��y|��0",z�e�c��-K]�W�^}���u������49[ep!<��#g���c�TI������`SI�//�B^n�8ԡMg�Ɔ%�<PI����e)h�K�kYYy��������˦�_���\I��2��=�^�f��$.�*'�~����a�B���`��x�׷���/�9�w�+N��
�.rJ���~��/}���Ci��T���1�?�y���9�7�|��E���D �މ���>>�P��"���ׁ��T��843н� H��������������Ξ={���"|8��H�Bł���N7w���D�/�ۃ��'p������f���k��H���Ν;�<���o�!���#��E�"�mIr����뭷����˫){!DSPy���5H��A����}�6��_�:G�B�וʓoĳI��j���+۾S�"��8=0�Y5�V��w��
|���lnn�&� .�oYPKx�ȧ
L7ҽ��ˏ�Lb���Yz�'p/l�d:�����<zt�āO����ޯ'k�����ܻ�����j"��ݻw�Eݸ��^^��|��G��T��/�����!".��g���� ��8�A�~Ӯ$غ~����K˫Ʌ�:��!��yz�Y��!���=�V_��v
�6����s#Ξ蠟By]%K>m=�N��w�����R��tFς5;n�jbW�%b6����?��_��_=��lG;s��	'�p4q7�z��u��`�th�ӧO�`����`S�x&4՞���h�}��j��<��0r_�>9*�}j���Qǆp�o#��j6]$��!��w!p������~ ����F����㋋2�H�Xh!l��?�yJ�qh|KmT*U{0�c+�<�6���"��%PD6N>���P�饋E%5#�5�����>�2~�v\z�JkuuZ4c�
G���!�@��Õ�>6V�#'�h�BϬ:���\*8"���<��l 7Χ�.�\C�`5^_и�,�i@����\}���2��b:N%W6� �	�!+�˳����QP�2��{�1����
�E�֤=�����7�C;%bY��5��$m�@�Z(*��81�Da�_��C����G���`()��C�ĵk׶n߅�S*gV���Y�_븐G��OuF������1���ww� ��KW\\&_�*P�d�!)��$��0��eM�N]-�F�Ln�����>\�2#t��K��C�{R5C��|��P�6����%Q���iǕ�g�ʮDse����ť杣�7F^��qE�	��s��QnC�%�<��)]��V�f6�?W:�mԆ>'���C[�4�+!J^j��Gx��y��͛7?����?��|t���\���b�R|x�Uq|_mn)CK������N��%$����+���]ywwܕ�'9��f%!�
�ި��*E����V�U!�L��n�$�	���7�#��G;�zNHL�'��,�Uy���yY��ܔs2�|�{����f�U��ױ�j�b3���jVsx��`_���J���%��S#���I���l<�+�[��OO�����r�*blsB	��[�gܔr��$�I�o�~ˌRd�Wh�OO����7U_u+�Қ��б��t��	�}�r�Ul�|��A�h����f�oa��>��@��TFv��z���K�t�6��.�~�ٍ���B��^W���³��L9�yE�� c%dY�U\�~�+,`B�@i��E�<8�SZ��VG�0��&��,>}��J>�t�$�:\b2����:��&NXnNI�������E����j0����<��]�.?L�Q㹙$��p��1�wǕxY���
���IGl¥}r�=I�^i���.�9�@�M�H��־�^�շP�n�F\g�y���ezZY5��U���-Cg�<�{���x"t^#rPУ�+8g�l&�-�g�^�*�o注�p@2�W��H������Nr�u`��Qv��L��ă��:�h�J� KM�8�TlI�����(��4e�)���U��A 'c$R�2A���duu�
��a��`��.~GG[x�25�2>���̊������s�R��E�'3���[�gxX[=����ɕ��A���!~^�Gm�᜻�Z�C����4�Gi$�l�Jl$ͱ�SoX�A�Mv�7�)������� 耺��0|����8;����"�k���!/�i/�5b'n��ߔ��8\ �T����k�z� �������nZ��!MtNEwZ0}�aPGz�d�5)y��H!ar�_�"h���m�1�Ku�� ����"�˪�vM%i ��t��5�	�n�CF�tT�#����HTP"mz
h����P1�t,.��,���K����tB}U�J�5].���qk2�ux�e�����ˊ��ğ��6��q{צ���X��j(N4�������"��Z���Ν���tQ�i,�$]�	����������8�.���lnn�>��O���P��y^|��G�E��u����;���E�1���ojܽo���S�����^��_߸q���@�a�eEUΰD�^�S��̋�ugZ����ho_
$U}x(͞Q���p����z睷Y����?��x�/�f�<���៿������������]1sAX��m�䵭S�N�s(�l0�׏�@⓲���}�7/?}k���G�n�X�k*��@j��!�;ʰ����
^�������?<y��7��M�������Fx*��YYp>� ؔ\�{����/���|�p�7�|��X��:�(�UU���b :�ه�a2I� �EO�j�J�~�2��P|!>�vbUc&a҉�;SN�<�rmo?�5?��&�G�$V�9���ނ~]D�5�u�^�`1�%IU��P*�)�����i^E�t��N�1���rZJ�������� �a�{wkot��kǎϲ�{���D�F�}��GW?����_���|��>9>��saV���o��gfv ����1�֖�ɰD�����5�Q�y(TX�kmUL��%G457��6�y���3�{l�өq��z?㣬��\,��<9v�
��Q5jg��ύ@�5�&Id������b�o���/�������W�\饝�� ���y��r�3�vr�5W/5r@���^{��_�:}�K�.��ǋ��0X�
�ip��Ԕ�x��Z�	�u��l�j��~��b�Y�Ylݵ����fy��syњ�j��XC��x~�\#l}y�(R��v�ԗ�|B����|bS�G����o��WO?u�-��	W��R�qn��S�(��r@`s9��)Y|nL���,T6T'����Q%�X�N��5��u�ye��tR���
~;�M9�9�G�l6,�S����+��:*H��4ᔮ��8<i^��ղ���i��5�N�S�k'���������ch�4���+�������R��S�v�2���r�
^���a5��Դ�c&�g!�Y��0^|��>�����&#\hT5e:�l�F0F��s�>&M��[�i��H����Q���ْ�fӻ�N����U|	�j=���Gá BK	�ǣ���ҝ�wC	{jz��ÿ�e�����v�|%�5	�P��a�Q�L �Xby�a���A�G�!��+�-����/��X#=AY[��TQ-8���]�n�� ��q��Ԧ�I-m���tW�oE�7��g]���ɭ*ZͶVUuC2X�1�3f�?�NCm%z?�U'��Q�<�X�dB�7:�)Ƹ�����o*印Y���a��K�M ���=�5�(x8�,[g?4TP�����O<N��A�冶ul���v�#@�X4��̳��9_�5��TV��߂	u6�Qt��3���tw_l�u�J��-�Ns�ñ�,+U��o�9��Y��9#�kP���AV��ɛ�̠lt�F�������2�.c���.E�0��*[���&B��=�i&}\JC���@j�a=�O�#j�1
��i�����z0�l*�$X�y`6���nR��d�� �M�qI��n$Rk�)��|��N;�B����R�E��@��1ٮ��7R��4� �H@�,o|��)W�q�|����@X���e����G�.ʍ	��h:��Q]2�l�jsk E�:�L��+�e;�̪�k��mBSLf��Xk� �3-%
D��qY/������|6��u.Pd4ml�dk��\C��<�]��6��	o����x#�vu�t�[���<%rX5F�|���ZZ�&������w4�Q�F)h:������4xo���b!�f�DD�/AG�͘|��Ӈ��g�>I �u�!�$�8P���w�vY������5������ }��9���'�acy���G�k��í�-�\
�@�H�F�c��(��y?�x`�{:��1 q�y����-�sW�`���R���cx��xI��Z�\%V����޿�oʹ8k��/���щ�0��ޜ_Ϩ{��I�\��휖Z=&�l6ύa7%����}D�Ú��q�d+S'sa�;`�.ȗ$��M�t�M�VX�q(�p�t{T����K.{O�i���$~�*�ԢH��2������J@~�$#��RCx���+�k�T(�O]�D��B}���D�[�Z���Qnl0z����L�xcibC�SkP8*�Z�'�$�T��A��T`n�^��QCn�0vQl(�b��r荰�dށh ��#_���5�G�v�H�y`>|���Ƒ�I?�?�)D�C��/x����ϥ�A3J0-���%:e2P�1�<Q���#aq�֖��H��(3�t{�֘4d�HF����XKb���/��=$��%���,u�Ŵ�1��;�m�T�;�DH��@R�J��j�����-��=�-PY�L�|n޼y���|.�������\�m�{���o(z���|{�����6�w��9����cT�o���h��O��O�'�����x���.�1�5xv�Z4���J{T����7�/�>�,��0g�����������5Rn�r���ӄEv�����p[�9V�+OSK0'�[+���U�L�'N�;�4��wiy@3��2Ɛ��X+G���F�(�O�����׸��"(3�z/^�r�ʩS����ߥ,t�V`�>tN���Y^�Ù��/�����T��Ι2`�8g��:{�,V���W����}�B1�Q>���@;��,��Za\�.M��*j�dyl�)	�'����C��=s`<�WV�`��x#���x���N�uc��*����-��a���ۦ�����?��?9vS��R���=��s8�&��v`�F̉p�֯�kh��~���?�8�Ǚ3g�<w�ܡ$ֳ���S�2��
ƃ���a�����Or
S��-�qw����Ɔ�sh�wn�;He!�U��G#�(��߷	ٴ,���~���[YY��|&���c�(:�@ΓX:�h�Ν;��lݹ#n�fT<qF�$N�f����r��e��Z)�z%dG:���z$!�u)А�!V{���L[/�������t���7�A�/E8E��=<u�����Ϟ;�{5��D�N��1g�����n���kMm��Y<���UcQQ����6Sntgk�2���yP�#�� ��u���t�W��L�[Y��>'T�Y�Z^[�vM:��&��͛�{[�c��[,p2ӹ�A����q��.̲�q�B���9(�m+5Ob�pH�ֺ]<V�K�ez�u���:����J귾Ls؀^�.���^��&=������:�o+�B9oA�&�R�"�ϩ����>�v ��F<��.1}A�uf<��JH��/>Ɔ�vb��~nlS�1�U¬�kX7-���7�Yk$'�4��3''*�Gmp���t�%u����HR�����bK���%n/�r��0�)�������J�.��&(A?���~{o��&ek�u�*��ncqL`��Ě%y��ӈ��O��}�蟉�J .��|���ix+T�	A���N���`{��Ǿ��3V��Q��O��O&c�C�N���M�7���uTy6�?����u�>��=�'��DB���$Z�q1)V@���UWI���_�qJ}��P ��D�Z��=���郠	��q��b�z8u��ʔ5٭SB{��=$f�h/�`j�y/n"��
^L���'t������&�:,;p�)�nҥ�b����`5��g��4`(貌��XlQQ�>�r.=�0�4ޤ+��y+iWe���"���)ߺ����dkը��+�M��3�儞nK"�Z��>�f�(FP4�0j>,��?��6d�Qw��HXI��{��'�"�}�6��pj2��Q���w�Đ�ŬB&6��P�"����*..���ҰP仳)�1��R���L���ڲ�#tk`��sM��q��#��X�ť�	�y6��z8�?~�����0��+ҟkD*#�G�����J��S�%�|Q�++KJ�%+���p���/�i]�B�!ì�Аp�j�wg�	�!Nl��PgF�M��M�B����Sw��O�C��~^0�.]�\�maԐ���VP���'�)Z<�̛�Ft�E�WR~+u ���{6�Z=�,�!2��@����,k&W1�Z9�^m8��!M�T�(!w�:6ؗ-�eݐ�z��"��j�ƨ[��k,��������64����Tq�"I�a�pp3�x�w=n�×�#
���t�X�A>���֙����r�����"�+Բ>:�z�.�_~�/�(A'98����p����SŮ�Mc8�ak�
��ݎ��8�\ځ�C�f-��x�W�!û��f��"n�|aq��_,��6Hshi,3�xk���g���?}��>�0E%"�)�LH��%Gy��p�³�>���/��/W�]W=��.E� �v����<&$B�����)������Ai�P�/ZU�?i�h+�'��J�f�qԧ?�i��g�L8�H�)�_��9�׍�'�x�,u����Jj�}%�������,fM�AqM�=��m;&��� ���*��f������i-*N�ęy��%]�,|��=}����(v��MX���mZ�����P-�&6e(j0I�R�D��bO ��^���3�N�Y�]zZ�ů�3K�Ґ���!�?��H���������D�D,//޽w���Mg�w>���/v� ��S��������O⠼��u�lp;"�ƪg��R�]:��ߦ�E0�Uu�Ƶ{�����7Ϝ9�}��or4���e�w��SaXx��|�ᇯ�������]�x���>��-�/UGu�g�^��!?O�[��%��?w��}�^����{n:�P����g�Kboݺ��$��Z:ܾ�=O��96b�Szb+����Ԗ���h��hoa�������AQfC�ͫ�W�Q�N�O+,r����:������FY;�hw�ݝ*
fE��?�S,�Ψ�?��cP�����[w�9wn�ͣ�Lx��������zq0<�g��D	(�=�R�G4�Qk�,ߥ�rH��ی�ʆyH��O�1M5q�k��:�����67��&[��'F�a�L��?ǣ!��jb����{)}�y,G�����,PyZ5Ձ�Y��X\���������������}U:�pmy峟�,V �-e�<c�E'�����W։�h���_�?�<�DaT8Ĺ{��� M?��t��C���H�Zd�7�����x��Ln�g-iǙ�b1���ϩ��e�-�S���ެDY�8�� 
A4�:�������
�ҥK'Oo�;�v���̱\���f������hwo����2}x.�SF|h0B�YG�(�BXR%Ϲ}�6���'���������BC`+�C=�H�J�2�&�2P>��Ex��;��q8�q9�����+4����Hz�
Ŀ��)����ݒ��% õvv�_�%�Qm�SY�Y��>���!pd3��p�O�	���I��n�|� z@��L�6�5?�M�4Y����"�����v�M/n�� ��k�o.(��0v���k�� ۨ1������f�?r�Q�|����b^?u$3RJ�i7Sr���B�RA�:D����KwN�YѠ� �Z�������|�5q癢ɹ���+W5w%s!��ߺ��������Ʊ��x:աd�I��E�n���VB���<֖l����X��.j)��R���������$�zu5���FI��(T�c���C����� ,���o2&��s[΄Z�b�o��u�����t*T*����dL�W��F+������F=��S��%nϦ����0P ����p�p���˚��Y"|�T��&�Q�R[ic�Qӏ"C��x���� �2�jdDf��J��Tى��{�:���Ba�akd���v�h�"�F��N V��{a��;TR�`3�F0Z�X
E����[���bO�\���HH5U#v�/�r+����x��(�+Y�ZL�� �4���S�OZt�'�P\
?��/���8n�U�Ќ�W�)0bm��k�E�-u�f~t@`3���N�,WfJkjp3I��b���Kʼ�=?^w���Z�`섧�&|��v;A�<�V���v��l�Ŀ!x�"@��f6��\�C��9�oo��[l��>q|
���H6�8*H}d�$�X��h��
_����%
�Rp�q��)R���5�=�-vm�ed5~�睘;�.��1�P��xInJԂ*'�.��.ieC'(�r��u�2��P����s��y�A�������S�0�	'�Z�	DS�N(��QR8�a�]��D��lD��H5� ������=��;�Fr�'N��.i:�ð��
�[[w9JBϜpzy�e������)`��̸EB�5&�WhZ-L=2k	���.8_����qy�L�}�Ѧ��+S�s�766����z�35�p[����_�W��w>�O���1v�`����:u
���w��
ODF�41kq�]<ڡ�l�o)�z�'�Ʈc�tt%9�]2%�DH�
�����I"BՉ�,R�Y�!:$܀!k``�ب{c�k�F��c˗b$S��(��c�=�?����l^s`�Ş��n2�C`��&0c�H����yǆ,-I���`������5xU���(�Ѿp�!*�򗿌'�Ay埿��o0�T*�q�/P3��A��r�(k��a"����%D�>_��X�%AO�MR�b�uގ�>_$�L�|���C,�����޿�?�O㿏��9�G/� �r�lJI�x�$m�O?��ɓ�,��q����qdAn����/�7hAu�:�WO�ܱ!na��N�T�C�4�:V��q 3�<��J�j5��E��!K��?���kʲ����D~З��O\���K��{ｇ{=���ef=#��E̥����]��-�dGI����?����)x�H�F��F���k:ԥN���ܽ{�~�2`���e�H�o���P��M!c4Re6����e"ON������HVR��ʒ��q` d�I���˧��,<�ڟz�)��aOr�n �_�P�%���ٔt�G��k���r6�����Q�!�0=�;�zk��s�����;��Xv�Y��G,R�~���ַ���O���!��W_ŭ��2�%| %�2~��~��X�g�y����h(�aX��� ���t�
��{>��7�E�f�bi�=��$�[TWԙx�2/d*�r'q����B�Eh.]�+k��'���oY� �$���*8�^�Ii���F��l��N<�T���>�yGv�,W:]k����:/	�;w��ށ$�v���,�tK���`d�4��WW�0��k�U���zYh�##�ab�kモ�X��H�cCK�#p~����_��k��ȟT6�1��(OT��@���˥�E�b���(m`b�7�@�&�ڨP.���4Ǽ��-���+i+u]��7��?��O�$/���6�֗.]߻wo2�2U�[WRGSɳ>��w����s�7BJC�S�1 �����}H�B�i��&ִW([=)2s#I���Aw��V_
�a=8�QҞm�^�0�ͥ�����u3!M9w��@�l0xd����sgϋϯ�&hA��8���R)_Ys��6�=��7W`GY���	˂Cz��5<����/��r�uM�G�v}kQu!
eog���4�_�E��G�@�6����ۃd�1N��;Q@\d'��H䈟�~]�&G�e�tXr�s���-f�������-w�c�z"C�R��e�PN�ɓ'�T�1ad&	�B #k��zu�>*��� Yû�('���=8<.	W�Nm��|5��r�a(<cc�M�pp�U#b�a��#LW#<��:�<�����H����Z3	�in�y!u�^�
������(��qfo~x+CʠT[?Ǉ�T�z��~#O��/_I�Q,:m�b|pX���깒K�A2+罴���O���N�Ow
OS-���f��Q؁2���R�������N��r��yGq�&�dZ��hi{<�5C'2��B\���r�፣J��� �`�G]6��̵[��)IP�`��<�Q�:�:ё�9�{H��p<?*�U҄���	���yB�6Zi���U��LYh�}��l6��țf�2(f��Q��Ez�Õ4��� �,~�WuS����l��,o��\�܇�lЇG5I�1���C��������Ĩ��j<!l�=��6�KDw�Yu&��-'-!q��J+���M���&q�I�����n �	�1��,+5��IdVZ�.�T�[҉ j7�9�I7H:aP������ʞ�m�Q��eߥ�_i�_ ��;�d�U��=X�;E(,��|i	�9��$Y�
Ǵ�C�c���'�Tu�)���L��Н�Jv�����	���"6*��$���,ci�OզB�+�.���X�"�m6H��^G���؈IX�u�E�b�26I�˝��<gg_w�l�M��d��ʰ˺/�,�-�u�@i�h0͔C�#�la��W�Z��x�i%s��C�U�x�$M��a�
B6�
�~2�����AUB�9���������p�ϧ��tm;i'�������PJ����H#������bK!,�o��� �F�d,�%��.î+��K*��8֝n���;iO���lPw���������$��i8�c]!訖�.
T�*����¶pmE�䍤�*�.�No,,�޺���^mt���y���B��	i@��B��$�H�H� V����2!9�p6���<��7E��'Â�ݏ�<��|9�q��0+�����m	�;�&Ϡ���n�l<��n��N�t!��1�4)��NI�@�p���⓽��X�8=�)����-!���e����fao�}傪�vw�q�e2uNs-0a- ��K��*s����ԡ�zN��9yok��7߄�,e�w�M{��������s�jkV5��qƜ�:d�p<88\\ҨC%.�X�"I���˗�^�
�E�[����+roA*h����]�}nI��
c���14+U����A��$uc}�έ��V��B�'�; nU�(\'�5BEJ��Ai-�l���$�*�^���c���q�a�	I4))����������Ǔ�<��gH��ҭ_��_�K�h)�L����	][�&�х�TE1󇇇#5@%K�yNV�Z=����3|�>䍣�Rn�;�'���WV$(�l�l&���g���MY��d	v�q�
�/���ԩ�_~���L���;�r�`t8ka "t������T�9��{�gӇ��`AR�U��Y86��~�O����$�ǝ���֭;�I����l,u�Y<|�����&���U�9n��:{�N|dp����"����*���|h��Y9�`!�K�a*��[��|aa���F]��<���M'�8/�>HVV�����?ԛ��%O�)-��Ⰿp�Ȧ�ݙ�'nݹ	�Kr�����=f�-�t�z]S����OjA�3a�5��٠�	t��gd��L�:�V��?���,�r�c	��`�O:�x��?�|�+��R����?��?��?{�$L<^�ߕ�𞜎��g���JX�N�8���O&B&�P�a(������N""�����P)����2�Y�@;y|mm�5! �@�򲳹���5t�C���ĭ��K૟<u����͓��1t�\)��k+���"�b��E|/�Dse&C*TB"��I�
ZS�ˋ+r��8<���4]Y^\^Z(�kL�*����NڟNŇKڷ��K<\:>\�8�xTN'/���ݻw?��#�wZ��r0�[��߻r�ʽ�JX9���oM��ҥKK�/������_J��p8��W��j�+���Jr�I��~��X�?��?{�g� �6�q���3��P�lzT/0����:���iO=�Խ{�d�����n;r���ܺg9�����ى������lN�gB�s++a*sq!�GeU�q>,�Io�����N?%�H�<I�D�����t�	JWr�q1���;w��:v�|�3���~�֝�0N�0�e�ԩ"�Ӽ��Q�l�-.i����OE����g���_e��p�ѽ;y����/�&p�^w^�b���d����.1tg�i<:�f�a~\��l�r�B��4�}�#(Qfd&��&G�e!w�b�[����;�p��;2��s��%ʹ��4�,�F4���6F��'>'sR�|>��!~����vR����?^Ä.[m 3L��7b#�Ӄ���D�3�V��d_∙�@!������ޮ��駟�ҭ��m�=�?!���(��L��Z�K\�x␾��{��9q���$��$C�@3ݼg\�3pf�-�f����F��uA?D��	,���q',�1&����	[��y)dDK]I���9*�WqP��X\��|Q�dv�w��ކ6���崟v%��B�N�n/9~l�����;������6GI?V���~��`#`Pd"��Ӂ]��R�_]M��.a� �`��ޖL�dt��������.^������K=�e*�Y�s���g7#Ꮄ���}�������A\�b�S%@ե���H�&��#B��#Z��W�ر2;	�qHѠ'�]p�e�F���jbd�&qg��ӡ�)!�
�#q�pN��F��H�k!BO/��N�� �
���H6���� ��g�xi��~lq4:�D9����gySHF�RU�� E�}����
m���J,#1�I��R[^X�.��HH��'�F�#�$)d�m\��4��*�>��։G�ۡq�6)��p%�Dvb���Y��YK
������p؂��oܛ�Q����v��y&(�����Z$��u!�j5=9m�k��\�B�.�v�XƐx��\N�rx�������'��>#�ϱ��xT�	c��P��"�a��Ph�1��hh@�ڦ�Z�m�g�~�b_A�A垽���;J�pE�@��J�0��fN�i��ca�x��(Y�IQ�Ք�j-�E]z"6ju׆ڮť�9���V���e�ux�����V�g��&Y�Z`-�a��V�7�����9!�ϲ'׾�]�O��L��X���ʫ��_� ����1+�����J��Ù�������H*���k^R#�尞Q*~��fn��Z$AT��p�A*���
q�s,�6�6�;����WĄ'�DΦ⑷��&c�M���:l}ѕ�Ng�� 5^�v��Gq	�����mUE`��CR���E�rYl��� �I"GL��DZ�.�� ��O%o�p(�{������Y��LF�N��9�y��.�X��&M���./��3��%S}�B�3M�5��K�s��V�x��K��I���Pݝ��#YDi}E�ar�I�����(�V5%�L�Fx�>\����[�2I����ٳg>�U�P28��}V\a{V���.L0��D]��e݌*�+��^���ppx,$U3)W[ZZ�8s�d��)��������/��x��0�ڸ\���
��4�m�U�,��#��4���xGl��@��P�<i�*�E��vG�Z���.�C�| �^�Ԛ6Q�$΋b�����Cw�5�t���%X*�� !V?����ll�kI`1����D0�Lp[�a��?'S/eǊ����I=��c��GU��R�Րc��~�(o)��T�3��t��vn�,��yɈB*xzxI5U�O.M ��ڵk�O�&���x�C�X	���g����|���˲�Q�D�Q���F�:&٫RV�3�%F��E&v��M~Д��0+/�b=�,�T��1%{X+&����&/�;R��v�/�CG�Q&�X!��=�q�پ����Z޺ug���wI�1�[dm�5���c_�
��|D@�5��
?�D2ts�@@L�"�rq�pB�d�,���mDm���శ�^?vHK��@kߡq8b�!����h�Ȝ�i��Pّ��N�k����,5Ad��A�Ab[��}�*�Ƿ�_؋�,�j�i�����ik�=�ӿ���E�oY����d��_Ͱ;M67�-����Epx+Ey���ˏ<|���T�8��|�S��������"����D���.�
������{�Rk!�y%��3�Su�TH�#Tr	��֟DZ�3����r���M��A'�ܣq8PP�S����)?�</IG�w��C�ɄI&U	�/�O=#GUJ�%�7yfTG3�]���>��.\8w���Ѿ��ݽ�{�ں���%��`��w�ep�����/�.���/��C��a��E��6~����W^��a��U
(ƞ�i-ǃO6b;�2-����^����o�_��O~qa�$�'eil��CK��2�1&�ȝiZc�kNp^祗^"�%Ѻ]g���xA,�i@����tS�U�X�;Oy�x�	K�B���HQKG���ղBm��nnn>��_�������c�IERE�����,N&;��Ϡ^��������l���DR��vr�dm��'���RAD��,�c���$=�\�o`���ZS_��Ҽj�u�[�c�5�L�wĥ�(����M���jw�Y���ae����0�x4n�I*�*mX�{&�����Cf~���a�{�9<éS���Y�|lZ��B�f���d����ʘsR�:Ra�whHj<��u�P�b��>I�H���7B)=�[�l����-H[��z �I���H���Xԕ��{����+4�$������!]Gi�HЂ+�Łr���в��ز �6���\_�l߿��	
^��`?��h�~�7�78�_��W��q��%G&��B&a�_�~��0��c��e<kq4����)������@bb*e|"�B�Op���>nZ��ᇬ��=
�+�@SZ�$;8���>�
4KZ'Ylݣ[��}�@y�����j1��C<�^u,��dLgE�z+�[*��9���=�3����}Mڒ̯v퇂��G�E�Ҵ�+O��6��|����ǘ��{�6��2N�@W��)���tw��_(\gX�#�g�=p����֢��@�RR�j5E;�EVKsV*�me��AU�0В��p"3�UFq>�u�i��#Q�G����u�<D��0J�2��^���2����V���J�v*��J�1�'�B6=Mfee�k"�i��c]�$�K��I��%s�+'��)YPx�J�0�R�fm�:@�d�$'^j2�
d��$�R�	�Q�����R�;�5D���f}#�sj3��4i")�m�>b<�l �F�CS�Wg'��-O�D�>�@��#.�X3�dR����S�b`^M�P����#4F�,��@1�Gen�
."@u2�3�U0�1�p�y=�+��e�+����^fņ�q�vu �����f��]z�Y5JJ'̪>����:�� j=��g�2Zta�4,���w;}��أ���O���;��Cu���<'ֵǲFh�Þ�΍���϶��l�jT�$�W����4\IU5�����q`��RF˥p'�W�M`�%W��X'm�z��ŉ�a�)��deeyi���C�Fo��&H�jU�J!�#σ�-;Q�,��q*5��o��tê�>5�D�yU^�1��]i*�	����P��r��|V�o]��I��tR����(�Zx�
�=@P�h7h"�#%�Ե�]���h1�,�5쵽�����S�/�f�2� �3��}/\M�p� ��P�>�� �[�.�re"d�s���S��g�u�S�<�l?�y������T������o��uꋙ���}&|q.�04��$:�^��*5��K��xN��y��{��R;5*NkuKiD��3A�A��'cƍ�c*ᅎRU׭Γ$2��H��%��!��!b����i��J��I�],�����vB�t�ڔ�
lsyI�w�&J�I��a�m�Vgs��f���5��\�P�J�6X��T�(�.L�bň��%��U�����o��#��u�,>�eIt:��'�9��D{��s���;`����$G�[|���Ʈ|1�ej���WZ��M��R5���ÉA(i��� 
�t����k~�Q
�mjܗT�7i �g̍���{#Ie�����
�ȍ�S�+��iBm��p�W\)=TR�,q�Ը�JQQW��A3�3sC��)/(���%��Ajx�;��G�!��Z�)g��#�z��ɓ'�"<�p�B�W�n��J'��q����29<��a2Ht0>��E	{Ue�3Z
HH�]ۛ��.\������Q]	� �V*��\[Z􄒺>�$!(Ãń��9�H��Ñ,QE������_�4/�'ŔJ�b0�Mo޾E���r��ǲk�
#��BRf��U�"������C�}2��[|U�z�r#=k�)�L���k̀��.��zhJ5Se��u�����^x���������'qj$_?><}����ޗ�--J#��h?�O%��b��2
UT�ғ���CI
c�_\�|A%�b���t�c��oT�?:��pم㷟I�i��������?�-�q3�*(����ߩ���ޣÃ]z $�.������m���x2�;��\R`��r �ұ_ۻ��s����������.�={�C	���e�����u��O�9}����=�~�����x���˷n?J�"�ly�7^z�%l���/�)jX�K/s�
�.߈�������������b/p G�OP?Gu�.��/� 괷�z���}����x������7���Z����ؙ����-���������V�X�h��z����4�>$v6�`M�{�=�q�+~{G��v��P��S>�oQ�������;X��ݺs��3����X���{�ª�7k8X��r9j������q0R��F~:���y�i���d�����VxxX[�{��!��iv�R�?�4��#VK�F3sWi_�d��g�2j���w�6J�c�O���FE�{d<�����T�w/����3��븿���XG�Ǡ�º�[gB�ӈTY,r0�L�� ��'�b��L�Ɨ�w�>��ܹsO>�$K��O��J���C�֕#��5�����7jO,VF)ӈ��
��r�yp�H�۰��f��u*��V�I4O��)�[�}ܣs	�@&"yi�Kd�Ah��e�]��(?'�GI쩢��R	q�d�u>3|�x������~��)��O����ڞ�٩w�J$,]�������������-�pH��̗��HAJ\�k׮��� 'pA'�1�X� 81#A;��[S#��7^[]�A�����3���ݝ����8M��T���--U�L8"�̉��nq�Xݞ4�hx]G�8�7�zް,���^<UZwf�NOTժ9Y�c3�!�p{��>F`�<�7�ۆ��6#MѨ��膭z0��2/rxz�'��k����d1�D�U�x_u�����y��"#h&�WN+�n|/�����b����!��]�e�����N��Nf�H�a`����b4��Ʋ�uz]��˂|Сַ�S�5��s�DS��&5ά���=�� ��N�J{_!�]��G8O�6WD��=����0\^h��h.x�&�Q�)2�*n3z�p�f?�tES���ThD�Q��!�q�O0�����u�}0P���}\QW;�5�����')a#���M�]wmO:���2���%��Z�ڑ��NO��r.1,da9��3�q�9?���ʊ<��)BC��ig��l1_Ԝ�\6���bw�W�w���!uP���lRS�k�XyH��͉�@���n������U���9 �a;\��(O*�	��B��s��3,p�ӈ,�s�Y��1q��y��mD/;ĕ	�Qb����[�-�׆�;���.=�oF5�K�4�7��<J�|튌�x�ʓ2����BO[�D����S��*�j��Rl�N�p�D�ȏF��~4�fos�$��0]��߼)3�����h$���1�s6��Ơ�������,�P=�B��x��[�hYL����pb%4iշ�D�h}�*���W���c�c ��_'H:�(~���D��C�8�c��%U�4p��9��3,�xܔ�$����`
�#o����w�S��n�V���s�p�ѣ�q����9o��F�S=+ޑ��s58X������lfhh3=C� �RdFs�GַE�'F�a|����*�l�-�-#���J[�k˕���g�md?5c3���Z���퇻X�������2Iʇiv�ab�H�Jk1��T�%���I!G�W0��a�骲�N���S7�����НQj��� �>������?���J{O�xJ.�-?��d����x`KL��bnlCT�;�!�%+EW�;g�cri�m�@����	��% -T��J�xn���æ#�y>�W,��7�����n�olC��!KLSa�A��򕩍)!���[h�)��A(�ț�����`>�>�-�a��U��-2#�)��<�a�C�}1����?�ƍk�+ظ��R}�	���a�I���9�"Ӄ{2Ak{{wuu�����J% 7�\�)�+���+Wx�N�t���;��eZ!x�g�:��w>� ��R��T?��J1�N�h$=Pt�hq��B��2k. �8�Q��cwt���($n�N�Jh�5bi��<��Iw��j.X��Pjӥ)��0����!����0^��64"u���Ƭ�F�_��W8qgΜy���U����}Va��Dh��*dmm5�l�dx�dw�
R��˪�� �F���ߗ���ճgϮn+�'�&HtBo@8��C�QV�X��g7a7�S<��������<�m�$��L����Tučv{1w���'
�����Q3Ԍ�Z\��ae:�|��s�D��tq�{����/]��Â+<�����Զ�>I����y�y���[!�;�u߼yr�̋�c��z�)<�#͓�+�^���p0�3��W^y�������/���h2�~�:�H:DnF�I�ZL.cpB��W����?	�)���?W����<�Z�t��a�_�u�Vn�i(�e(��!�{�޽��_=1�ւ灥�I"x����M�� �W�6k�w���`g���xwj��f�:n��(��}��G������8 �B#�3}�M��$Զ��(�`#>��C�|�	�
����5���Cư�RT�9�u|�uҎ���x�<Yۨ_7mek��A�݇iǧ��82ptly���W�Yu�����[��1U!C���g�=����M�=�C��R���'U8�K�U��w�[u����"-���[�kܷc3���r�jު����/��
(m�am`s_��P&���s��l�ˠE�ɭ�M��Iy(Tۀl��oho�*]J^�~�D������H�5�n��D)�ϟ?_͔�?jj�|NlM7�şd�g&ՙ���ν����{�}�3�!N��G�R!H�C�Q�za!R�����`���pj� .P�����_��`�7ˍ����?�����=��/ᢧ�Q�dumچ�nO�3��5^�3�����{��b�2��M?V��,E�Ot�{+äų�ZW�_���p��¾*+4�-�SdSh�c���x��pi��{����]��&S��z�-�lrm��Q�`�Xj���ܪ�o�߈@�� 4�9���6�L5�1����W��p�����<wٱ!?m��u��I����z�(π��<��!�M.oss��I�d�My�2Ī��i�:��Ҡ�e�jO�&��²��0סL̐�:�:J�Ag��CǎJJ�'M\(aYǽ�'< �Q���ƱV��m!E��[�8�L�媸�nQ<%�U-�͞��jK*�z�4�5�M��V�t�O>��XWBYԉ��ԥͥ�X9�'�wWs���h˫*��w��0��l�y`���c]P<�X��]����(y�Q^���C�\������v�9�B��qά�q�ON�>�����}��=x��߁ U��Կ�GO�pr��_T�Uҁ��XƝMZ>�$U/�B�fYa\E�3�T5���c�V��'��<V��j0$i��<�_F�n<��g`��L��KZ��:Jjc�-���S��鴅C�JI�:A:2�P�X�a��{����z�^���<p�����f��*Τ8D�i1�,ےI@90r F����i�.��&$�F�aӱ�����")�C��b�ө3~��Y��k�M���A����}׻�g=+�M��a�4�� F�"[áP��81��ꯍ$����n���:�,֐SX� �P]��$@ЂK�Q�	���\��P��������uIO�A���l`�N�� g�����a֌t݄�z�z�C�a95�+`��:[�,�#]��y%�\R
6ۋj�K�A����5���:�I��q�~A�q��'{j�~�Af'����X�i*�{��#:�q!PAA�K]�?
��Ɏ�f��j#�O�q�=������3��{t4E�0�.�*�OH�+�[p!e]�+t}B9a'n.-����:�x/��Lo35(
���F�ӻw��٪�FC�+A��sP�!i��jt�f�I!L�9��D�uQ�A8aUR�`��2��{B-��~'�C�U�+�¨��9-�)5�j/]KL8��X��z���v�������k�4z�r%����dow����F�N��d��!5�N�� Gc��ϐc�Vd%+곙��9&�G�����ueV�+�Y��ԜO�dm�nl%����I�斐7c�a�)�d��(Ҷ�[g�%��y:���4V�?6��ҡ/(�@L��Uz8yxw��PD>b�M2}y�Ľ�E�~@f���!��l�R0iW�V���)����<;�,����y�@s|l>�+ҹF��|����K���Ȧ���tB��ES�k�-�ű*���5jJ��E�9E��QiT!e����H)WI��s���/���.��#�٪Z��8鎆�Qؕ�Mw�q.�ְ��ǻ�ɴ8�?�u��6�w����[35��˗q�!'��y/WA�@�`aS#�8�V�b4���^x��ͽO?��p�_Օ.Z�6*�����e}m�.��t.]qiȕ	�
r��w��yS��B�<M�qy����1t~I~�-Z��Њ�Ļǂ�Ż�Xr �:]�� ����9P����2E13�
u�&�h�<�0 �������������;﬍�6ܝ2��=<ڽu��R3bL����~W1Ţ�;8���i�\N��&������ހ#_��c�.���ѭOW��w"k��lSѵ`n��>�Lt��]�<���=�
K�rs�)b�t��ˉ�T-�-R���� �7xP�,)]7(g�i��z�t��m<䪾q����=�C��__�_�9sJ�Jc!#pǐ'4� �Q^�0��O�$z��/^��+\S.]ۉ��fx0s���,���������g�}V��Q�j��q��2e�[-	�o���������o���ţ��xG�j�6
3o1��>;3�W��B��^�s����+.���������P�`���J<����,j4Gܴ\𴭭m�>}Vw���dGy"Œ4��F8�*������})X���C�%Q�2���������]��3g�ʇ��`<Z��b�I�턘��}�#�Ƽ�N��<��?��=6��,�SQ���	WVJ��X�?⼧��t�Gm�%��!�)0|�+�ݎ-���R_Z����b�X�5�����8���+T"q�.\�0Ө�c���{��7�~��ͩ��ޤ�"�B�Y�"j�o���_���&K��E��Ä�/,�;<O(�+S��o�z@a@�Ј x_�b�<��$����s�S~�v��52|���}����@`7�ӣ�����Au�R2%�?�]�taS��>\��+�Ʀ� 0�I-Ws��/�R��W�\�-�*ER3{8�酽��xqx�_��\�p	�B�?88s�� �Ȓ9�3SA���NG����f�� ��\
���>�&d�LA���67�����G�y��l`�'�������?yb��3��d3m������i6_��:7�C|�,��4���#GU�
:��7�#����il$*�Ւ�.�oP��iH�H1����r�M6?[�2q_��ʀ���43��O<GO�~���>r�ɺ�M�ҦN?ȅ�O)��߶�p<�z>��XK/S�p�i����2��zu4�3�UJ6Z:����(�2C�W���._�mp��kdA���}I��L��{Q	���rKf �U�]J��ˤ�b)�Y����&A�v�!n��$cG�Ֆ�����\��0p��'z�n�F9��+!A+�Uhz�zSϔ�:��xmA�HePy�9��n��JUNV�q�ruƎ�X�&m�F�:��@ڥ�����Z���W;�J`�[7l�����P}�X�(fk�byE(�Y�vH�6�9�ܾ&�x�\"�+�x�!NdT跿���_=Q�s�@I�N�������}�S#׃�nӰI}�	��t��xN"\5�KƠ!�f*�8kJyY��[�B��=�a�;�%�{��8�!�S�#QH�P�u��Б��#2�ůY�<c��Y�ؒ	��}�x%�\ɫ�V�ĩ�ǔڣߝ��y��8�����R��b�;w&�K�P�BpV�ǡ6��T*l˚R�ꌓy�B^�.�q���K-qC�ab��B�{8\'r!ԉr���̌l�n��`����BE��4��@g_6z���VE^�FC�p7�Oa���j�𲌲z}�.J!���,���
�Ns��&l'�u�}	t��ɕw��eI�[T�K%M�*4�XW8����1X�6�u��up %�G;��&9�+���I�E7�� zx����H�#��B�yX�g5�$�QU�|�_d_'�IԺ�&yL��d�V9�2��˹S�ӉRi]4��I�e�O�I��h�:S��I�� ڎ+ NO]��14nP��Yr�k��=��DN�Z	���W�Y=��Ĭ%JT�,V
^`�'�dlH,m�)>L
�B48�ͦ����3��6A�K�Ě��� ���ІR?:��I��[Xm�Ս7�׿Z
P��"~��)/���Y��t�!���5DT@dP�EW/G3i�9����1Ga�ܜ �>��#�Qn���b��q�yL�������{�3�u�G�"�K�� ���D&�&�*#ob(}e�,��_���*�N�[dP:ӄI20k(��̀�>����f��W�~�F���VV�6�6��2������-�\�d�x�
2�eQ0�*s��b�|<AV���/�?��O|��tAMve�z��na��0v���cA���/\�vMxVtG:���k-GI�F}�&(ʥl3��'B}WJ&�5�;cȇ�L���M��2�����+�� \7<��;��3/���a�器�@S�M�l&5}62+y/�����������q�2�O'�W�^��~��'%�9��՞zꩣ�]ae-&/��}����D�oˌL�zr%n�$dMґ��U�Ӹ/�.(u=-Xb����m>�>|�0oԌ"�J��?��Z�b����v��҉"Len�o4e{�Eq�����2��0�*S��@=�L� �d�[nނ�%*=�,�jw�����?�����o���a_©��wt��)9݁� ���,\�������:}������I�lsgg�	������Ư�Ϳ�7gϞ}�7~�_�iJ,�[�yVvB<ۏ~�#|�K_��s�=�c��� b�K�W��5�0 1O��Qn;Př��m�m2���0Y)2 Q�3�c��׻��OʓL��#�t�SJ<��QR�
����	4��c�#���F+KJ򼄚U�xSxp��^�~�ʕ+�n�"�>���eI:��
1�M�p@����y���!�bzO-*z;�z�^�|�&�[����GC����_?Lۗ۸�vPFEQ�NE`)	����A�+��4��=E"��b�h�X֐�槟~
~<|t�֕���y�=�E����7�7�\�:�ʗ���7���W�*�lu�y��ٖv��4k`���0�+c��Q����}�ug���4���,�Z���)T�B{L��E�3{��#zc=eO��vhhdN��	6Nb_�$���D(+�e�c?��9�����/��ҋ/�(��"!N�Ύ$'G3]sa?�d�a;p�b��`Y!��b�)���p�q#x��E����*�lHn��I3鏹����B�5�������'�Ia^�f{{9{z[�ᔰE�ʊg7uccM�6Y-�,����}l�o�Ir�)TKk��u(�+�v�#4-�,�j=��i_�<#WkQ���w��y��Dъ�Vhl�ABC��;��j��x�X���!�����.{�h�p�U���F8辫�W�X�㭽�(�X�C���5��Yڤ��A�&�c~-�ی6\=z�'�<HАmta�@�QX��Z�V�^'��95�̊ͭh8m�o�{���{s$�/�Q�Kx�����gpﹶ0֍R��L�j6�Mk�'�F��3M.���kȸ%ɖ������Mc��XG3\C�,i_se��E����p,a[+!
tŨ���;�:!�{iү���&�'�2;�s���l:Jo4�ǨCzxM|��Ct���Qj��64c�h��@a� U�+J:%�XJ���-Z�Sd�����Lb-<��kųx���6�SKU�"�҈WP*��Y7�;ɳ��J��E
/��W2j����~]ؑTTX�Ll|����^�«� �S�gQ[8�?R���M)�?YR!���E�'9��^">��	�l��_�<�f�*}��i4�
-ꬴȚ���Q��J�E����]�q�GUAh�J�HV��y|_�"FMǷ�.���faIm�L!k�PJ�s�t���`�^�<t�Hk��[����E6�s����*=QV��Z�=a+Hb�n���@��uX�	���?X��ϟ�:IRF!%Q���[[key~���-����GX>급�R&-����yR�˶:8�B�бˊ�徼��=�̹�t�D����=�tӖ�j�:��H=������HB�I�U�Ȗ���3'�6����,���2���dtC�:�8z���+�
*����)ºAW%t����xL�����)�ZnW˝ǂ����_��oJী�L�S�h�ɂ��b�Ë�<w
)��B�Zp�`�*n:��&�
B�UgF
�<�+���K���;wT���%8W·:�:ݔ�)�nm̤���܂��7��"v=���l"��nD��%�nY�ƅ�b�S�J�c�7��f'Y.3��|����GR�3�xo_&*�M;!}��'Ov�����J��;��̯��߻w!"}�#˃����wBpF:݅y=ov�P1?�s���WS����C���V{A�?�~��?���L��W��Z�/�μ�rf�/s\vmmK�eK͊.j$rv]�Aq
�@�����`@���ʐ�_��4㆟�%Z��¬�J���VFIFq��f���H7�Cq�L���;r`:kH�ۄܲ=��Ϝu�"���Am�� �4m���eN:	����FK�NO�2VQ=b`�b� �]封��ΖuK�W&Ov�����$N�Ϝ���N�7n	��w��<R]�BXW`��"Q��8��͖8�Am"h2����ʋ�?��{���q:?'���T-��d��h������/'G�_��$Ϛ��It���4�
a��'�[�T��l�����8o��S��P�F��0�W]w��w����N�	!�):��Ұ���'L�i)�1itz��듥+M����񀝶*0x�h6����������׆��S���'���M��<8�~�:IrD]��
yW���ĉS�t�H	i��	��w���F���a;J(�"� ��i��M�+��*o�vA�e�/��á�=+=�
� �Dyy����F���*+{^���PeA�V�1���Q��><:`�-�\���*魘!���8�S�*i1?<}�$<���?��+���ω�X������p/�;���r�qGy�L�����ۿ������Û"<���j������ӦI���}��_�����7_x��/b'����k �Ng0GGG������~���~�����_A����B1�4�t�[���S��~��wU�ڼx��<��f��{r�K/?z��׮]��!*����MU};tRFU.SV�B7B�r���4�-�B�Gk���T��I=��f=�>�	R!��XՖ��s#���GG�іIw��J9']�'t���w���1a��9�&�|����g�����$��>	�����1�A� !��R'0)�~z�\v�4ny+�:̓��aP*��WY��j���*m�b`->t�Yڧa��#G���QNt�<��c&S�;Q�'N��t�v,Ѥ5����|W��ThA���nA+�j�UbO������БQ닑&ձ��ng=��2i�9� jq�o�`L����G�:�k#��l} ���<D����r���Mǻ��jk������F�ӂ{��4J�\*N�������Ḋp̅�%	�[n��8u��'���P���!�ν����/���}����\�����@������!t�Ct!X<��U��LP�����ƣn& �A,�p�?�KVY�G��D�r�6#������J���E�������o���ۿz����J�R"��x����>��^�ֆ�T1���c=:d�fH�"G�|v�)�sj�z�`  ��IDAT��b�,	,Q���H�(p@"�0=#F�-<�f�5�%��`�$�`��M���tIE.��82j�H�R(�J� ��������s�Kߡ�Ke��*���ٰ��49�Dz��fR��� |��X�(�4�.�P��E�¥��@Z%K�G�4P�m؉�'rĺu�I�6�Z��@ L.<]\x؏�H���Ç�Á��1f`SD\���[�g�����mK��O�D��S]��P�Z�jH�a��?w.w����2Is1��\�1�m~1_������«������5��
�# <�W]{���-����_-4��� �1��5%ڂ[��L�,���Z�n�B�飅����V�)�	�+a�k���lP?"��e�A��<y��'�<>F��D���-�K-1(Jh��8��Ts}��y�h���{oww�?�@g�u�tZZ  ��l\�xq��AB�[���	�х��	� s%��2����o�B�L灍[��y�ht�A��؀��g�hx��jZ�"'e�S�f�V(��f�d���2����cYi#��Rh���ֆ̱%�R]%�^�<�lzt<�)b����&��6��e�CZ]�������-z*l�H��Bh�t�S/����dr���>X����Լ0�K�;�.+��ȣ��>��^�	n1(�$M+�����)Ii�Va�<eMBu�.�����7���E�B%)j� �&R5(�/Y�RDh+�"Ս��<꠫E-ٸݽ=*@�:<�xԝ��ؘb��M���ӁM�e5��v�D~,iv;�[̰��8Y�S�h,?"R���%���'O�z�9V��.s"-��S|%�����H���@�q���&��C�t���9:�S����rI�`� ��mS$�O�F$ ��O�������Bi@Gy�o���3oll���l���0��1��Z�eq�ǻ;p��n�8I����pK���xYed�,�Mv��IKC�s�2�K���?纂�q�w�(4��8��+j�ܦ2�b@�x��Jh=�̖F�҂�!2���4�e/;�N0'1.ro�C�/nǍ��N���<,Dw�6~���[�M�Hlx=loZz�#KD�(
�J��Qb�����䫼$�b �Z�յ�{������d<�Ո�X�C��=n���ʳg�^� �f{{�N�-c�:�\�h���W������T5���+*_�&�T���<�쳝�ֿ���z��򓟐վ?�o���΁�o�3��ɵ0��f��g�#�g�IIH%J�)	�K���l�U���6��6͆�eT�S�+[�~Vv��?Ek6em3F*���Hm�0u,���r�u� �t�_GH��2&֟Ad4�h�����_��_������#֦�;�n�M���7�߸ŕ+W��{_ş���;�%�~��W��hq��?u���e�V3�j�~�ӟ��My�����������
%���}S�����ںz��0=Yo�SO=u��e<�NQGY���j=�,�	�ݾs��u&�I�
u�'bu��5V/�Gï}�k���V�T?�я�z�-<���?���~�z��#,
�ŋ/��s���$N�����qX��o���Ǐp��!��Bt�j��c�!���3��/ �	�V��I9t�b�7���������?����~�+r���DmOZz����_���^b���O?�R������7I� ������},����~�i���>����C�H5�l�]o��D��Ey�n���m�DL�H��^ �[[�W�}��>ɴ;���9��Mj�n��,�����Ѡ�xY��\�w���ٕ��PxV�?���l:�#���(�&E��B�xň`(�O^G�&����;�xj�+��|!��"�ޏ��&'�������牭5͋���+�m�����f���0m��v�4=��]���X�/��| �a�Y� ���VW,�|��ur�%����C�UM1�ذƆ��'��q;[�Q���h�Ir����G-Fj��5t�ClUtG<�|0O�P�Kc�*[(r߯���Z�J�P��G��6��O��N�������.#\�aO'h�$R�03˧����j��������g�;f*�x/���}�#��g?��/~!b:�Ն������(ũ��(��y$�p@(Ɏ c�g��P[md��n������-$�N9'���I�s|�L��`��~�r%ٕ�B\ʭ7�9#u����pD�y�0'O���K&f�jd���.l�CKǙ����z�r5��F�Qf��,Dl���<O�|��ox���i�����
ދq�CY�0�;Ok�	��{��13�U�(m�)o��U����UB�c���L+	���)Di7;����V���3�&2���J�?5UO����x��V��jy��@װ�18�|P��I�.����g���!\Y�g:�AM�þ_ˆ�r%�H�
8�MU9��~�Y��\���^��}ǣ5R,S�ʢbZB`{#���1]C���
�[8�.��ސK#�+@'����ȉ�e0�"kF6T��掊��t�r#�j��f���&a���C�� �t��X�q���AMs�X+P�Vk�B�&}A�h���l?m���5���{�s���%ī,	�.���%��_�ͨ�J3��q�UӔ*��+ad�1�v?�TWftHP�}�D����ln�$���|�.�\�ֆI'�{�������`���V�5�����UW�U̋i�oO�9}��+*	�狸�j�ӄ�����矽y��*[ P�%
t$P��Ca�~W��RGȡj9���s�u-�j9���T2��c��[�yX�)W�$C�Թ�B�1��0u�9��<��x���t��6�Q�W����G�A����֖��n�I_�:�<(z��?zR]��rzص	����ZR-��kI��j�YT
�Uœ�W:�/^<����48�U��S�i{����հ�hh�64��XY���-��e*s(j��*�,��].��]��Z�ٲ|�\�'C���u�`;�ܘX���Y_����4!�g����N#�(�!<r'I�)dNR'j�XJ�EV�s
�p1�08P:�Z�Z�qS����@ꆼ�PN7���Q^Tx���p}c�L@�u���yx$��$6��uXt��b>�r�*��v��&��&+�YE�D
�U��J�PXi�h��Z=��|6)�L3�<�|&ͭ���T&�b�р*֡���-�+�\�O2���\�F�Z�8L➑6�5��
�QhS��cF�����h�,�����^��+�K#%���2�زI*�>u�"�pY���a�$��2�v��
��J��}�칠��R��d�Q}�mes�s���LUU.�ɖ.(�4j(�	FP��r�`h'�x}�I4٠+��?ux8�裏_ݾ}��=�U<�pLa������J�_�8��7c�@�)ƥ�V�#-2�o�|}��'�\<���C�F9+=9]��f���F�M�0O�$�=���,l2�����TV:B����pc����rc �l�U�
�nv�E�JLC{HY[����T�LNeF�S	��:�e]�������1�!���
�px���y����n����0*`G�Wփ��		E��|���|�<���k/���3O]�C޻��[��檮����$��CC��L�n��f������7zQ����N����~����Z�0k���0oNQ<�����jY
]����������ae&3�lwۅ1KM7�Pr��c���� I���r����=BBC���s#ñu�yё�J���0��MYZ�Z��37��o]mDΈQ�d��T�-T�{ｗ�l�$7�����ܳϋ����W.�;{�U)զ��L&<�2?g��+�zZ�S���f�˗/C ��x�.� �q é!/~�%�$ǣT�*��Η��z����� U�k������?=<
��W���:AŘi�ԩ3x�����H�Ϟ�`sCzbƣ���_~�[G���W^{U
Hiz���g.\���D��oH�sϿ��w��s/lB�O��]��������$Q�)T���~�k,�O���퓧Ϝ��7���\�	�uXj9��
������o}�[��믿�� mj��z_����{��v�+_��s�=G퍃�=�m
޺XI��\��ݽ�}�oֆ��^{��'��R~�����{�X��w"��yr��z�1��=�E0��h���XßC�����)�8��K�����՝��I���h<LH&me3A��w5���'�O����O��--G'�CJ�N�!lg����Ŝx	UV�7W?��*�`�No�If�5fK�P�G���ayE��V
.�ͥ�`l��g*X߈ĦJ��='�n65F;+�&e������,�k��6�264j��Z7c�Y�m�$�������?@�~�Vt�?�˗�Z<����y�E颩�n4s�.�\~���3��6u�Z��.T�ngCC�����ʿ��qf��
����\���ܽ*#\�
��}$��+�Q�E��B5�k8���Pi��]fa��pr4�~�D�J;��r���ʘ�Z�,�T���l*p,9X�s�S�u}��(u����{����������A��{���ֿ��Ly�	7�D�r`K;�5@�^����yLp���	�{
�9F��-�I�I��F�X�̖\dg�����!�8�gYMYCFIW��em<���|���_�A�C�5j��2�-v�	-[��nt��~)H���(�s�.�عr�u�E+�Q�͛�A;�'�3���8o���|_nݮ~�C++j��,��������>O�2R1R�È��$�xrx�b ��r���A���-ؑH��'2c��	�<���Ãi�t�C��vP�5d4I��r��{���h���X��*@�	��[�#-on�!��@)��j]6 MB�%��'NHX8�����ӧ�0�)k'JC-Qu�F`Q�F�2`(�L6J��e�#շ�^���}����
�kl�-�b�z�LYl���f׆�),�Y��q�j��͗i���wM!A��|�|T�\^�	,�M���0�_��(u�K��&u#�r�8�\����V��S{y3��St?����[�p7lyCR�$���a ��\u��q<����& ����_�O<�Net�u���1y��b�؆��`���o~����p�P�Z�A���IB2�r�+�V4*���F�H��vvj+�d�9w�G��4L��gt�F�����;v=��pq�{&a+���7�K��m�T!ʻ�E$�-�P�t��ف���"���{W#k�#Jb8<��v��MY1�v<�:l:s+ͼ�HJ��Ʌ"e)�b8��?�lM7db�a���`��_�^�뫊���U9�����Nm��&�M�)IO,mЀ(
<b�牷�'�#�\W,c+�
�D煹�R-����Ek��U�]�=s1�Ք4=��b����j������k�<&�N�f���<�y��&o�t��0Fօ���9�����g ����KgXUv���ڬ��LQ�U1.˶b���E5���#\�c�ٕ�w�o<�5�)�6�H�0�y����Oj��jh"���`�/w��*`d��EQ&Y^�>��eᾠLqQ�=�����s����ӧ^z��X"N�����2��&�5pΊa����и�o�*�X|<�;$�D��+�n�<�#��T�=�ؔTii��q\>I�!'#���?w���V��F���
�)Y��F�M����2EU[�⬙=\J:��Ɵp�\f�R�g�#�����G���F^���*����\K��<>���c���ĵ���\�x�P>�ub2��ƪ��L;Ž�[��Tu�Rm|hԇ~�U3�Ht#�;Fn�H���/]�M��^�H�Ʃ�:_����%�EpJ���W͘�Ύ��`;�;��?�v]�a�Q�=,�Dn>Io�܅��Ϝn��տ�WP��ލ7D2OuH:�`�����^ݴ�j����亁�B6^~���r�N`�h4����d��qu�a�����+������?׆��O~�?!�4�� ����G[*�>΍ϑ�QV�-ZSЪ�3�<�0�R�]p�;J�A˽�����\�z��K�s��;w�Opks���_��
���|7�T�tDq5N��ZU�h���]\�~��CDz���.���ÇD�t�����;�@���d��Op*�������Q�����SR�YMc���G^0P����:P^���x��Wy/���Q�Ǽ���n���
o�HT�P�[{#���'W���������o}��ٳ�̞0�ǂ�L���ł����߿��`;���/�~��=NNg	�1g����?��?��t��}jH/ϳ�ΕW%#������'B��R��͛79ʓ �<{BOÝ(*���c���T�k_�?5�\jM���:�cڠ7d9�����٥��b�\H��p4xR'#�2F�w׮]�-;��t� q'��5�{�Ӣ�H��tr̧Y�2B�!����Qa-L���WST�K�pqʛhݼѺ�AJ������,�����,�YؘWo<�^[�}`����OY�Re���q%�Y�����*+��4��@y�2�c��nMh<ZR�!4�>�,^�y��7����Tn}x�EKHvA}�!�>�I<MF1#H�l�T[�L~������^�������q��U�|g�ď�`��X)<7ZiS������؄�~��ȳ���ʾ�V�*=4t���ڒ8�E5g�]~����x�>���A��5+�Ze�H��_2%_P�Ã O�� �gN�s9OQ�V�=�$�?��믿����uA��s`{��A�k�ʖ�����=����i��<uj��$�ۣu�b4�Φ+B�i�4]|�+˫����a� �=q�:��@��+�A�\��E���hz����2���Ϳ�w��׿������:�p\��������{(Z�n�������O�@����Eȯ�N�S�cKSYݗ��*�g[<c_�`�ٱ�}i^��3�Vj�
�{�X��s��x�� ��r��#�e�8��4�G��G�:��ޫ�/�b�3�S���N6\ߚ>��`�l@�,�U?�)�E3Ɉ9���ٝ��3��tP@��|4o,c&�(,�:B&�oR��4��\�dٳU�c��P�u���ŜDpl�u�TY����^��u��ATu:�<�&��"��&��NT�tQ��Q�����;_5�=?&&H�O�D�v�D�"�%��k��������HT.S�.U/��5�*��O	�_Pm)�.:�;���K/E2�VY�5��¨-��]C�r�c���E�r���>EA=[�$oϯ�F�^��3y�	_35�ğuI�?��'/_���F�{��[�퐧�d�.r)���,��&h:���t�ɥ�O�����p�Y^SoC�͆}C
2�Ch����[h���*��]I��^sj�G��	߫��U�LU;sr�{��W��drY�%����[jDJ`Bd�ġ&Y�!�M[�o��;��%��5��иinW&L��^y��IJ�]cG��pϯ��b.��j��e�i��1��E8Sek[����N���,�o4�j(�������6� ,�=�b;��*�%!΁��R\�G�2enܹ�`�ڌ�J��<��s�d4я�
B��+J^���nR�eIl&=E������E�*qds��ۓ�kjFOO�ORlkC��k=�HMF�2Eh.�0�v���b�3v��(�	W���z��IZ��\ccMQ��1��׃2
�$��T1��m�d�l_��><{�,G�A�ame������ވBq�����Ϛ�'��5���z��J�>c���L:h,}�^}>�g��ǩ�lM�2��Iprx��B����1_
�Ju��E�Ђ�B�B)u��1_%���B0��ë���{���#U�B�hgg*�6�k��Y��X��ǌ�::rW �O5�Dm�e�q�S�N����IƛB� ����G?��u�7uW�i	lQ���v���:a���v��H�D�*�)B߁�77��l���5���37G�~�gc�Jm_()5\�H�a�dE֘T$k&5%��/+�thZ5�fD}�v��ixשiy!oz�ʤ�m��`R��O����7�kd��bZ�/˪Cm��Y�L�E>T�,{�i��!�����h�k��Ыk��u<��3K��]q�k�0K_�I[��ӣ|�����O�;8���q�A�r
-$��� ?�H�*M_���2�	c��`�� t���	����6}�� g9�b9�دYq�֍�a?�o����~��_�+��޽�	\wm��-�P�x��~�˳gΫ�NuD�:&tN�X�$%s�,�y%1�cEưÕ���۱�6Ж�.���y��?��˗/C%��z�-�^����Z�s�鮌"�s4�u4Ȗ+O��M9���]�D+�#D:x�*�_�t�EO{����x]��ݽ�C��W�}����o�hr��-H�J�y�ٟ��S�L�j�u67���~�)@*Z���}���?�f�<L�rRΖ���L�6{��m>~x09`Z
��������|@3�cUp��i}f�!����/Y6�.�d�ɑ@w{]���K�.e;��> 	�Śg<j�b���{�X��r�t���c�qYj����rR��NT���U/��_��1V�ي��:���`F��W����@�޽{P�o��ƩS'�~�ʣG h�w��0%�YjHʯ��E)���?�����?���?����{�e��H:���s�dY�wE������{��^}�U�2?Zi"++P�x⩰�7�ڲ�?k�� .b���O>��_x��A3׵�����q�ԙ�w���	h#1�k�,��S��>��:j8�y����ѣ�l2]	�h1�lzl��$�h2A+Fy�{�FP#Ѳ�HzQ��P�Ǧ�e6��@F��d�B,�"�k�"�彅��o1<7\g�\G�N&����vj���1<"D����*���)�!��s[^
Z�r��Q7XB֥<�W̓�x��z�}�CmD�J?96L�`�W�;�fb�s���Q�Q����sC?��s�LmrHѢ�c�$7B:ORT�Z�Y�k�nv�МĚ���𜋇�.�N��.Md_�X&�
k/�1ӭC����2�[l��n>gdd�6E��a�!�x�	�,!�R���
߹}���'I�t����*R�wVEH͔m�9�[�u�|��\z����8�&<�|��/a���D�a�I�����;\���tFJ���
�5t=!ˈ�C�F�F�����l.Խ�x�w&p ���;;�X�i�bK��D��,���C��򵢣�7=R��E���g� /a����	���lG�{��M�7��׾*�C�&�F�M����Z!O����)���~�k�7�?i�j$,��g�B�0_-��#��Z�v���=~��EyW��ٛğ�hZl�.:&�����cO)�Bt;�I;k�x�N�]$-��I��D�?�5X�Z�l�Xe�߰�z�� ՠx�Ju�-H��+�8�J�|�ƫ(sV�uS�ľ�6�=M��Q�0<,W�~�_�j�(��D E&��J�]Ty��b���rd6��wj%jj������ֶ�cfÞ��:�5����N-��7@����SM�Y�m��ß���^P�,rt������H��V�T!j=$"�O�ܬؕxlxf٘ZAvq!�-���!�kV����Ω��[���W�Ma�	�$�����pڑi�ū�1ϐ���7V�+g5 y���X�5�Q8��(rx	n����o��p����'�;�����v�|���ܵ#g~���n�-}��uG�*3_�W��d�6�����FEiI��jR��"F|ި��FN���u��ρ�y:�pF�^n�*�ᮦ�����ж.m���#�c��&LY�
�w-F�rz���]a?t-'��݀�����:t��+��t���������$/�r��
�"�Zhx"��E�	�оR*�D��*6 �;���wM9xk�QB�E�1��Y
=e��>��$�q�6���V��<0؋��akJ��]؂#�?�اm�q����欵b0܀k~��tB��������?�λZp_��q�?�����S��
��rF���V}�J�Yf�����5J#���,B��&����aas������-��e�u�|��#ƟȇÎ�"6����q}��tF�M=�V��S+;i;��d
�"@"�E(��K�����d7"��z��:w��b�<u��ٳg9���o~��&�%2�$]��:Ȉ)���I��8;8Rk'���a��1�?}��7�{��G�}bf�x�k͞P����+��p�T��ĵ
�pe3.)rx���}y($∍��O�H�A;[)d��D(4_��+�6"7J�����#0�`ì�)�+������K/y�Pm��T(7��$SUh���(_�ҎXlJj2:� 6�<4"�B��"�
�`�G�e3v4�
6�z�m�_A`��9��'�T&�wz9��h�ϔ��@z'�yE����,2��TX'�PM:@H �<�?x饗�ݿ�w����n��&�
Ӯ���X���H����y$�����zTL�������	���	�������yB��tm����f��9�@a��ҥЃ���_��}g��E;��g�������ɭT[_nooY�9/H��s4,bbC�M��g���$��?$]���a<X�;��͖5mK���2ӹ�s�ē�OA+�
�1t�w'���M�Lv���O��A��O>����,�0 5ل?F�N�1�'Gq}��x*_y���ׯx��Ն��>F9�n����Crd��f/�Ĵ�Ah�u(f�)��M{�,�K�.%u�Ϝ/Y`�N����⇞�]�tp
<A��6��:sF��o���-�XkXs�WΣ����>���������eh�}�k?��k��}��������Ñ�q������������z��C�zB��l�����%Ψ6�[�$�x���`��y~<�W�ކ���DY�W`C���'h}�ך����[7�p�c�ΗA��>ܙ}�{�{��g{�6�΃{�%�����V������	���4)�O �,u�BC�Xp���������$���̵.�(���V��t«�:�]b�M��6��9T��*���0���s��.{��c��x�4a��7]P�����I/cp�T��8 �;�sM�(T��.��ܹs�5 � �ͺ6�?���yd���"ke�RZ��&q�6��ߝ]$5F�����w�mY��I.fdC}A2�SW�0�����H [yWe�X�a}�l��>K1X��.��Q���F�L�iM�)1x��'���v�0�i ��+�Vn*�1?k��H��}��j�i&a�}�x������`����9���������g
ч���cD�s�	������ࠥ��\;2Q�ǂ���8qDl�|����K���Tt����07�w�c2�O9p�j�U�Uv�
\����)P`�dt��Ʋ<H7���z�-���_y���Is���@9���}*�VF���0R��2����\b�6��~6��pτ�-�w�o��n�@кB��~�����M��3�PΏ}爼�x���ĎHA�p)s�������%1f�<f�T+��g�Xh8+��8㓨���k�[k��A��BT�Z�;�o.tx�ȇ+��R��H3�|v���/�sõ�T,P؉��A�&�b&SB�v��h����ᨻhFAS��6���^,!fb]��Ȧ>5�A��fwù�`:�[�5���a�V���#@��`��É���$S݄��Y����M�=*,62X�Ƈ��\X��_���rCX��IV	:Gx��I$E�KY�"��<��c�������KM�z����Ղ��!A�zH��ؔcs׫�|n.fЀYY�Cؗ{*4����*�Em_MB]����p�{p��ݪ_{�B��9U�̖�<ֹ^�q2-�霟L��ѣG�~��M�bӡ4��2�r8�ⵠ��j��O��RM-l�8�z������^��Mf���$����u�^�A)��;��&/�3�1�Lᅭ�!C\�a;~�[2�b�nQs�6�*n��2�f�*h���0Ħ�<����
r���vbNъ� �hYH�$i�9���99�w�B���P�X=��8׌�7��U�/�g�N��n"!�B�����1VC}���D&���!\6:F�|������OB�to�cO����Ah-D��ί�<���
���&��M\�EU
�˸��!��שf�)A&bE��/"�~Q�LMY,���lvt�8��(�K�A��&$&b� (�v�ꙸ�o�q�`b���z�z��B1�A�MÓ�6��.g�3���ol���"�<K>t&�tS�a�����;�,K��`0�<c�GPLM���� ���J�7S����hE��)r�[q.MA�:3(9�K��
���h7�׉�F�%֛5s`�{V�E�`c`�S��+��YPbb8XCx�-�7���Lg�%ދs��-V���6�e��h� 
�s��]�^j������hK����Y�&ṙ�1�8���|=���e<z��t:O�#�c��	/h5	w&��Gg4U��E?�TW��j&+�0�iE�e����DѦ�����|i{D&��	�jcg*E�����MH��e�ʖ:(�,1o5�s�I�X�'O�~��%�FJ��,�i���b&܇��B}k��o?�J�#~X(����P�ql�#�L��ny�Z	�6׊�o�#R�0�W[b��Jj	�D.����@�-à&g�� �U1u]b�%"c����MY���[0��Pʟ}�ΦG�����j������CAF���t���a����pP,9\䫽�]����IwK=EiQ��{��]�|!e����_�mlJ�i:S�'Z��n�����$�t�ڠ����>��;��;㵍/������_��_@���h6�"b�'.���9=Z�n�BР(��k{����(������h��.h�<։y�xF���6kc�1u�N���g�;w�t:�?���&Ջg>�&�ѓ���u�[�\��#�>/���&��t�M��'�O��SOq 	��/8�^������	'��?��S���ڵkGS��\8V��|�������$U�Q���w{�[���������^�[�Q��,cKF��:�T��Rח�2��^O��Ν&�.���p���_}�R����F�.#c�%�h�{�r=���}�Q'OmC��}�=�߃����!��W�M��>KMrE�N������{X
(�P9��ө���?-}��Q9
���xA�qPEx^�8��#��L|�+U)3�����}��W_�tI�tV}����r%�#�ϓN�����q��|�;W�\����Jnj7I�(���R�����������U�o�A�A\�>h�3V���w��l�5ϔ���ؼFBBd��{��<�x]�p���/�5��X�k�8��ps4	�.�>{f�\�@���3�#1��<��/��� �ZR��*�j|������	N!�y����P,��)x�Jz�,� 2��2�jS.�у����'X�������<���斸 ���xi^ήbWoݺy��i1/,�Ր�\y[wldБQ�0=���F���}B���=�z��=!c)-kɼ��1�6����E�^Z%RXК`!�I6X�;+[�!-V�ɣ����X�A�&��2�Te����B�#����4R��(8���0�\�E7T��S�w�|�<�-��+�&��ߑ��ƐN��~�o_���X�bP� >	ۃ�:^O������=�Ō}����*C	�%�{��m�JΤ�*T�S�o�AZ��u���Gd/��{����O:=QP��IG����b��fD�p��_�L��ݯ^�z����y�EjvlP 	p��2�.
*?v��xJJ �-�vrc�ś���
��tW�g����������H�p#���ɈoI^�@�`>��@��bua��j��_�;��K^R�U��璥���W�� z���;.�q�� ���e��P�G���}ah�]j�m'")È���օ�n}��#U�ހҎ=C���E��
�����2q#�`)����T\�:u�6��?�9�&@}$9q�^�)幥t�����}a��B2c��U�f|y��NU�=� "uw��C$�W���i���g$�	>����l<.�I96�#Z>1�����kc��(���Ŋ=��F1�:���Y���KG�곊*�w��S�Fpx$�a�A�5u�8S���+�]���hq�<q�a��C���s����1���q�o�����J=���]�#��Y1fv_6
k?�m�Q~�}Q����]'�lS'�x�ee�&���%s���%;8�^羼̺�+�JF~P�[A���c����x���0Vf�m�]
|�W�í�5o���9�V��,g����O	^T�֚���+:-+�$Y��AC����A�\�O}X	����Ǌh�� 9�&y���G�Bq���g�T��~�{<��D-N����ySO5�Hˎ����縚��;h�g�P���T\q�Y���v;�u"�A���uJ�� 2W��n&�h�
�F1��껫�M��t;����d4�ݫ���nb\6L�v�o�U��Œ0��
h\y.��M��a��k��j���>ׄIm��
GO�5�C`��,�Hŷ	 ��.a,�/nЅ1e)��l&��x��\#9T>�%#�uU��)�h<ܥ�Uv��@w_
�B�ݺ{>#�n������53���@L�i��c=<�f�f5o�F��)�q'���C6gqa�;\�'%8�Ϝ>%���h������H�ui�lUA��wI�`��޽+�	���1T��-ܫ?�����4�t��N#ic�'�y������<�A.�3֠�G�J�a��a���'��B���� �/;�����VNǭϞ9� ��g88���� O#�Ӕ͡N;q�RkN���D��8���
nn9w.��>��)Ʉ2�P��9�)T'4�2�R��5�(�λB�s�8�]7���8����_,��y��(�FF�9CF-�8�=�"'��H��"0-�6U>6ք;�Z�]�������p��l���`l�1'�R���Yl���|1��h�+�����B.��ɠ�y�7W?�^����b�-�����6�y���+l�(OU�����g?��܆�x�'����y;�<.ߣ?���u�{��3�{���1g����d7a�A��Q�2���T�������Dlmm�B�"1�"��V9�a�eޒ��<����] T��2�{枰����ᱏ�?��6�7�$<<���5���7kk�ደY�
�˗/Cw�X	r
��0�3e�g_�x�c͡�$ 'J�o�U3�r�ĝP�T35jW���]F[j���c� ׬��<���ĴhQF�6bOI�����ia>��#�~VZ�V,�����8���x�.�{�b�wi�#�qs}����t/hp}�8���tX�L쭂H{:e��}$�m�"6xH�^���W������۵�=�I���|��7q�?��?�t��7��\�9<�k�K�1���$S!��}��ϵ��G���x,�fr�[X���v��<]>[�~6E_<9����jgΝ����9:�({���8�b|��P��)�4��ᰁ�������/�::Y�L��"��u��%������H���h�Q�u�1r����%���/���[@\�A(RH8�����Z�&�s�M�Q�����ڲK�e�<B�qd�mmࠢi�����&ē׃���RB�_H0�y��ͥ,m���#�kۂDV���!���R�g�ꚶ�`q�:^�!�H�6J��DFyL�Σǰ�2����uQ�%6+���&ش�Gb�Cb�Аr!�F��5��ڛ=.^$�H;p!��%.;eơ��-��� +���}`7Ǒu�P��ก,hu;rx���z^�D�z�jw��s&� ��ҋ���Lx!ֆ�\2^y60+��o�%Y�p�a�l9*:�s"�n-��ٛ/s�H.ٺ�����0��+_��7��2��_���O?��q2�������tBـ���X.q�e��i��6i�E��Q���R��5�A��a��$����T����"��Q?h�(P|ES,U�T:�~��#$<C��4?۴���c�Zi����M�<��-#D��T���y[�x�(,��#�*�����������ڒ�â�irK��R���P���r����c�_{�5u ���ʕ+�de�0��5�n)�VLk�U
��<L��n$�n��|-6�iB�P{�X�*��,a���~�5�u�:��89ּ������w��i��d"�X��.%U�A�������B�lȬ�,�=�a�=��K�^܉�Y9kj�Pp��M鯖�r�����e"�c�uep�$Hٌ�����eL��06c�]��pQ���DM��d��^'���NMW�'V��Ө�P�L9��#�d��u厣a_���ܝKw���~��p����k�LF�m���k�\¨��a	���km�qk$�G}t]c�=�*Jl�a��-��%
7W8��k��q���!�LjIGϡ>r���k��x��.|b_~�/�SA��<��Y���%�\B7n�x��wi���r�����*��$q�pG&G�G���w��2ĭ�5\�t�ΗB" ����Igs�Hi�W~���ŋ����|��N�٪��d�R�-�/!mi�e�~�l�B�f�r��%6����;� #j%��UU{��nּjvS�<祠h�R2��tӡ�J�����K!���*
8,�L������i�l\rt�()C��@L�涒�4���(-털ڤ�:Z�>��N��u���S?��A�)����J�I�yo]Zg���\)��g$�Zm8��ʬ��}��Ni�4x3ʆ�S:bM��چ�/Iuɇ��9�h���u���^e���,JI"˨J�k=�XY,�9��n��A*�4Yz�_��ʼr��ź���Z��U�m���zU��s��J�O��n��t�P�� ����ǻ�n�n�I�ú��C˺,CI'��T��h�U͵pR6<�b�X梪!����;w�ܺuK�,���+�h{s�A}�$��d��TF=K�R\a���\ɸ������5�^�~�c��1�H`����E��Ɲ�a�hf6�$�lbŒ�+��SI��G���{�x���(v��3�4���Բ۱
��th$�px\�u���Dj�_wX(cVb5H���_̀A���c�c��r�S$DNa�	?��K��	�?�@+�ON�͠@!���JbT�%�>ɡ+��F�-�_O�����g�#�X3k�����Y�1���{_"^.�lF�TB�k�|v�Y��k�
�aӡO��tN�&u�	:t'<��m�󭞺����=ޓ��
�y�IM�}/ɶ�UjP�����Pk���:���QS�"�K�K�/��b-�� Fdrx�,�9�Oy�TƑs]���N"�"���\_�t�|W�E���;)�j{{���qPe���^�;�N�N���S�z��g_|��L͎����y�Ѩ��	'��\� �`�c�Q��M$_'�ClS��!f;�fýf�:��@$im5O5�9���~�@��0��!���j���BXp��溎�Yܺu�S��FÓ'O2CJ�<�a��|���/�z8��L,��3�r,��Ӄ#�N�G�6#(�JP�O^�'A<�a���)��� ���� tJ�q},f<�?~<Â�?�B�#A�]N����a�ə�d�֮0K�:�TdiX9� ��[�A8ц"��{������8�66�݁�j9���;;���*is���o��l T�3�l��yitL���E�Ξ:}��e�a���ȍ5��6��|����k��+����O|�_�ƽ������i\�� ���j��曈���o\�|�;�����/�f�H����T-�����W��
�<�̫����S�8�9�6X��:�x}Z.��W�ڞD�a�#,���sQ��y٠��������en�~��3�=+�5���M������g�
���p�x0+��(�Q�.)�����J[�е�4�QA�P�x^����7W�<k������
�Ii}+G9�M	��L��>8�$|�������r��Ex��5~ă&t��g�Z3Y5d!ǣ*O���$4�[�M���#-��m�Aq��`�C^���x���W@��`�L[4�������$b\RBd
���Rܯ4tshX$���Zy���$3��ir�<���l�n<9b�)	�^p���R�xCO��f;�a��;R?c��&D��^���Y)���ک�ʘI�V����;� �B(M<�n�K��J�A�N3�L'������+W򥤮�C���C��ee��X��-�މ�$�Bq���2�l>_�?�Y��E��h^2�������!��o�������ַ���e��"d��DJ�B�R�-/{��`��_ә(:��S�iFU�vp��5��L(��I �69t�7������QI�A̋H�Ť����HC��b!�b�)n�f�E�ÎTyʎ����ƥV��Z*�K��W�l�!�}l�.�����f��G �pk�b)&*��=��_��:�4����j��a��������ca��%S�����h0�� QG���:�vh*�<���;]��>��_|�K_������WNg��:}r�!N�d�2&�D
�l}\����i!�<�Q�$lx.�q�P�W�0֧}�[�i�/ب�C' �vp�����v҆��S�,r>�ww8�q��}ٜ���F݇���@*���d��7!�����A�P��hrw��*7H'�*����l�б�6*�j�y%|w�q�)b�V� {/ x G���H����$���9��:�2����2��a��֎D�$[��dK��S��#�q-i)QD�!PP�?nzg���I�r���:6��OH(e��3i�,3J�m Th}yQtܞ���yh�����ntm$ht���&c�9{��?H�!l�|�|��N�cx��
�׉"�e����jWt*ރ��c���(s���K��t�������U�H�Ze2���R��#i'�L+~=�_%�{�6MTt����I��;�x`=�يFPK�&��O�M#2�[��t3�j14v^W�DАQ��Ï&t����\KR�,�W�9��Q��'�e��eɤ�9�,v�q9�=A��Co�Bx6��IE�%��j/s��t�%=Q�R��t����Jt/B�Ъ����Uqf4M���W��0j`�b�I���#�'��$#��.aJr��@��RK�R��t�pM���p����YI��� Fz�ݟm�|�x�r���[�_g�j�^ش4�Qz�#�%w�51�&�~ZO�Q���4EG�@��*�1���֯>�)�B»2�r.j&�����nwX�̋ح�U�Z|a'��L�c�o~��C��4�2_��!OIE�tӋ�u�7yd����.]�!��������z,��3�3�s�323r��$&I�[�E�˂]�5�_���Ш�Q�G�h�l��.ڰ%ۂ�i[�HqN&�#c��=sk}{�,��ZH#�=����^㷾�Km�FT�8)Ȭ�@��R��A��#(23_���qyM�7X��uML�(�0ģ�(��ț��(ϒ��a�lQ���爪��c}ꐧ�ի�Rȹt�m2�@z.Q�2��x@�D����[��ѷ�����Gxvv&��7��_':S���a@��D���wB���R��א(�ޗ.]j�����V �u�'W��b�5�'o���'{\����E���H��<�)���S�j�L�eF��M2���ф��}狷�8A���<�J�ܮ2��AA��QD���0�mm�8�$��	-�uc���V+�d�J�1<x�8����_X"fx�@zfq4�[���G��0�u�g���:�u����`x-��͛7	����oDHR��k98>�jv��Y3�2��A��u�Cc��h�4�5�ajZ~ʝ�6Q7r�6u��.O%]n1և�#�K�����'��p�4e?C���>��9Ǟ�t�ܛv�e�=h����'I,s�u�hT���l���&�n��
��j)�0_
�i�s����?����/_{�L�\	��k��{�Px�K;���uih[p���s6p$ cޟk��)-�<�uQ�uVFBMu���+Ʌ�8lgS��!����_|Ah޳g��әCv��< lt2��sOGScHŨ�}���5_����Ǚi�A_X�Ij�#�;�}����R��~�༼����ƍJ��{�=�'� �N>-t�.�������~������1��]����{Va]�i�@ǂc��}
�����䃵�w����S`�IK����U�-��j�_�~�ڵkϟ?Ǫz����駟~��_�^�*���$hM�$
��\
�W_}�/:�aMNO B����e̩
����J��ͪ2%��x����!�x�Ç�<�YT&�=U������,���&)��漖�id%�=S)`=!<��%4cDIX��������ΰZ4�G:ؾ��
��lo���.�"�gK�t�f2�K[����2���R�P��Z���QE�v��v�p���K�Ұ���D�j�th�4D��ĸDږ�ŜI\�(sm�-��h�3�3Lv�K���XW�,]�o+�����z�0�Ҏ+!�����b6�W^�|d_�ޑ��e"��5��"W<[&�1o�����Ql*+T�	�
��o�Р�i�a�x'��n�z)���4�YQ�f������X�" P���y4�27�ʗ��Q"��WG<�&���3�zR#]��[@�j\�0�|����?�g����r�۠�b.I�sT����`1�/��[U�}���n�TN���Bـ�D���ŷ	���r)�Bs�ŋՒ��t�|�� �S,>���h (�(0}履ڄE�4nn��c�$L����"���V)��4���~v Y&��G�ǦgΉA`����v'o�e�Z�k�&F��%��nu""���
'Ϛ���oYڨ�����l<þC��\�g���#���}�������K�^�1������x�L��1ο@w͗��6U�'�_)�r�6B|�8�v���b�|����[�Y$$TQ�([D8;�[o����:�� ��)��`�����g��[��RV.��5]�Z{���E�����:ֲ���it8�����,���G�E�4��0��Of*��R��\����'�.��6�	���F��`x~8	O�*h�	���A$Q�f�5>|P?����ui<
=i�5�N,���b5I�eOe���(鍶Ȩ�Z�l�'*+P+a�j]}Va*Ee)DOI7�N������C��Ћ�XQȡ<��@�f��}�4�e�
.m�0�y=��,����!\�������R&6^ݸ4s���v�ж-S�US@ q��n4�q�m��[���/8��"��ⰲ�
^7E��L�&�g�E}��LS%�N���ɑHCs�qd�r�T�=V�	���sF��4���*P~�FӅ&�)�`���suݤ#kp���ә�a�B�]��!��_�R�9`j����c^��x'aq�s�9jR�I\a�W6����I���d�l��g�EY tb�g�e��x[�4�}�tr���O����Q�"��5�$���i��x”�~��
�V�~��]���on��j<�*#�'(,?�pL#)��~[c�]��u�r
�a��^����svIА�4tfI���: 
Nӂ��`Xi�BO��Y���x�CQ��k�iP�yS��~7Ka����A!D����~��4���Je_�#�O'����.�llJ�iU΃��䦇�8���q�Z�@lu\D˯�eL��6E���ħ�cr5>!�=i&�5�$�����Jec88?��a�N�'�m� O\�^"���h>�����{�Ŵۉ�������"q�U�X�8eU[:��k���ޞ�I��B�*��.Z�X�8;�PCK9�S'~�_{~7�B�z�� �T[�N�'��t��Jf�,��"'���D��"�j�eN5U"��n�[q�ȌL��Ҭ�At !1��9j�|1/��А/�����x���0k�phfM��g�0򜽇��fq;����o��̀8�1\��*_���%�p}B��0�uS򞯼|D���G��/�B+A,�F��N��٘J�o�)S�x��e��Ԁ._�/j��U8��4�X�����~��;$��:&�5�K���!�K�z؅ӳS60�2��v��`�=<6��4�>��<I��Dj�}�V�"G ��t�E�	�G,�/m�wv��]_�>8�E]���8K���[^+ܝ,��"^�ٸ��h��&�x���8z��,.�*�G����$��P��ZG��Sخ.�A�Y�뜞O��x{s��v��y^��/(	Ն�b5���gٖ�\����|�b$
MNn[H����UAX��Uo0�����A���P�D���!	�Vǂ�����~y�VJ�0Ly���ܫʦ�V�NbK}<v#f��b-\Mc<~=�bzz��������r��%B�ռ�e]*咀4��:��t1����Ɠ��|އ��ea�a�+5T�����-�Z�w�O�֓��kW�JRcks�m�W^��x~�hh?�˹��T��|Qdi
G.R��^�F0�8��J5�©a����!��`C�ǔ.������[�e.m�\����ty��� 1��m�
��q��a2��#:�k��Qr��c~�7$h6�>x�etu������>}����ON���"����R/��|.�0'W�^��>̰�a��F�9�	G�AyQ����>c9Fe
ۨ�$���Z�V��B��P�L�2��|���� ��Hq���*X�r19qq��W�>yY�g�On _�fbw�]_v~o4�fׯ����NIz[���ڊ��x�R{رi�/��:93���U5���&��H �uє���p���^�/�^
X� �V�ٽ�ww�.A �|�H�T�)%R<��NDS�d2���������6��{�w:��g?�YY�a�<�WZ�^z�_~y��û7o��O�S���5�^�H���G�Cë�����[�o.g��{����C����ǧ�����1�AgIOJ���uoܺ�G��k!OL:]MP�?x������E�	���������^y������h{6bgv���`�x$�����\�O�/8����4왒��Y���ް�}+�:�R'��ŌvPg}A�ʯ�zĜ�x������SH��"��]�Y�2�K����B�D��4�������@5a��_<?|�T
9�U� n�tÄI(6�ő�XҺ�2�0U���/�*�`� "�ę��9L�4�u���<\�.h��#qZ|[SB���u1�0C�e	<�XSW�*�ǕDIM=��ݥ&����4���/g,TF��Y�=/�ƨ���
,�cT�m�95�+2W0�e��*�r%�;H`D��
}��
;��2�	��,���r�1Yw|�}�ډ���g(�20d�����g�-}�b���]�STb!�B([�*�ڵ;ͤ(�D��jT"��Y=erY(�KHhSj!�9��O	'��N�]8�%'
J` +Y�,|h�{4��
י��2�)m��`O7εά��t6ψ9�낋O�c������@�¹ /������/$��*	m�"�5U��k`X_�������������_�����?;8|�젲�β�aY���E��9��/^�@�T��|Yt3�Q/�z�Xz�aGJ��H�[���3|���J���3��m�?	@�,�$#�\�2�u2d+MRK9���h�ڡ�A$yie͵�\�a�Vv�[ću�a	�c)!��E�A <pD�̇/�����&q�\�Z�������<2�����M�o���O��SM��,�k�@�	m�����R陖Nx5��� �� �!	�a��d��O�X-ʦDy�ڵ����㯡?g3�/�\M�j�(�٠3�|c$0�LBx�,VX��
�%�8X)��$N�h2�S^߿zz*�������� lsk�i��\�L��`*�����tsK��bREL�"$�]ȴRP�
=�g��GΦE¸���A̉PAp\�x'Zxg8^@:K|��lZ�7���o[mOO'ҭ\�*$���J�/;��>]������C�lQ3�z�	���S�ϐp��ލ��Y����e>/B�W��V�6�!5i�ۧ�]�)I��kdP�zHX���*E��ذ�@W������J��frd��[9d��}�6���\����m-�;�p��u��x>}��}2�t��p���c�?0�`kT5xDK����
����qK���`>&u�h���B+1���N1��߬�+��K�f"A"���*h�k���,}�����T�K.�Q\I\�e�����@ۈ�g���F��	&g-81tV�Q�,Ų�P0�{=C�*
����tA(;�M�����UFM%m�����w	��,��+�~29?==���/uѝ� "���0����$B�U.�@�����˗���v���9֪.\z��Ȼ���p�f
�`X�x3��dҷ�� ����R�����=�ЊeG<y���_���l{E^,۵В�-N���K�!��`Hw6K.xU(�!U��[M$G�~���;�n2s�+!���l���B�0D�ܻw{!AT�L���J՟��dI.��)~�+WB �1]��|�7�_�B�0�c�MS�zE	)����l5�t)��Jr���\(7?T�lb!3"b����!���}����0H\�H1g�}�:	L@Q�y�(�B[�.C}NWu��q�n6�84�q{υDfI	�Q�:�Ԑ����������7�>�6�ͳ֪FP���c�ȥ���9��ի�ٝ��<~�x.�C �"0Z{�������y�̪�+4��A��L+1�ZW�qց#��	��~}E�_;�E_!ĳ����Y�Z3ܺu��$�����/��_~�%ކߐ����f�,E�i�@^�f]��`Q�����u:]-�Hj���ٜUw�D(��3Ζ+~�c��ov�R�B���-'��.���+=nLd(�zA��u
!��&A4�CI�4mvL<VZ��k��)�M#H&.Ӆ�A:�^ܑ�A���,��1=-�2���X���o�5�,\fV|�\Z��1�����78z�.l�vS�wA��:�;��<�������Bq��"'!�$]D�z��js�܊V�$�<�0Ol&9�=�tk	"j�&�!r����<>��lTr� 6�":�ޅ+���1
��#����{�|�������_�\3|�uz����A����gϞ��_Qt�p�ca��Q��4�s�9��w���g{TO�ҹj,�sj�
<K�G���+	9-0���Wk�(?D�-�,Z���ZCP
�d1�x���x���&�Ñ<����D#�[�lpf�uxР[=�ڀ´�A�Hi�tx����'˫Rd��짱jq�w�y?���[���A��<�{y�^�N�|$6%�����m�4�����6�R-cq&d��������������e�I�9�ԖTT�p�<E��f�4.މ��YƷ@ɳ�j2Y��׿f{���>��cC�Px�w��V�9Yد�> c}����l�6hCx��Rm7�`�Z:3\����{OH�k���m�Ն!.�?Ra`\2c�J(�^���l�	 ��be�Wae>��3����	-���6�s`G��Ѵ��E�D��'*{I��J�Ġ�<�HǨ�t�w8�Ut*�2��� N��̐n> ���i�o��$T�6���Nz���ֹ1�m ���+�͕Fo�=e�H����n�G�n<�8�׳O��[�����ֆ�c(Wq(
��s�ѥ�(ꁝ0I˨�3��#�}��	ϳ�D��'��}Ñ�bLgm��3��:�c[U�-!lk\�m��-� �Tb�|�l�g�K��W��a��lT��ǖ\�)Q�}�6M���ұ�����"!��l��@�׵�p�����/~����?��i+q�0����"�c�w*£?�/Zx�n�����8�텃�+������bK�H����y��b��]�R�[.���<�
m��o{+�z��x�C>�	~,K$v���iDv�����y\:�)�2�a'��ͦ0N�#c��&���|h�j�0��ʦ�ނ�9��ڥ5��,IJk�t���5�<�[�:��b��b��i`��ݹ#& �K��L����[�X�(�86 �$�V�(�p
*1��jN'*P&k߲���(�TCE���QHqe�BJIpʦ�/�/]Z0�~�����*Y�JNN�6����
�m����0M����v2�����Гk�����ҕ+Q�/��õU�5EU��s�0�'��(/�J�|�G��IƬ(��gx��S���*jHڤ�Hܺձะ��S���k�$�?!��=U��s娐&W�k��U�X�'M���);g��Q�t�T��U�S�(sm~��SK�(Z�o�hIyyF����_'�hS�������b0B�6�Ù�"ˉ[Y��x�5�]�~��tf'I�ŷ�^�t3��v3��qꘆ��k��ty��]�����Z&-[��T�c����u��?�5���@���D�T�T�'�Z��\�����UB�y�hT��3�ɻ�v_}����/�o����T���P��/��b珺�6�­R�\��It�Z�e�G666p���Xr+ze�E���Gi����J��Q�jUY6 �YH���D���l�X	�s�U���_#�T����,BB(>H�?;�������g�/�=I;�s>:g�/"��:]����h�Er"�y��)�-������ED������_p����%�udgb0m����r�3�S[�8���J8&�z��]뻽9��ݎ���k7���9�jj�e(]��ʥ˧�1Z]B�B���J<��T<Z88���pNU�N�I�p1�"_���㯒��e�P/$M���>�5�5�mx�\��_>|��͗��&0p��\�9�B���L���S��v��#��}��{5�?\	�S��e>�����$�����|�<9>7WZ�`�8_��B�k'��/��n|3��c�Ͳ<Ը���b�S!]f�c��9<<�N�g�k��ʠ4i`_���{C�B<����!���,�:]�o!\��;�2x�-�]/d������$â�X�_��҂PHm�m��0���a�X䤖F��.�q�lmI�%��x�x<Q�����@��aa��n{�������m'�D�t{IUb1[,�lz&VwC�OW˹Qz��(9��m�A?���it2&pKX�P"�R!��j!@�,{]S�Q�3�ƨsiw���N��8j����N��)��i��E��]ۿ��d)QAs�pнq����!.��5"�:
a1��Dj�mS�ޚ:Z����M��R�S�XxH��-zϰ�7�2��A����t�u�D-��r���ma�>9>�S�Q��ߨn���R)�.��4K�e"�,�:I�uH�O�T�:׏>��ζɊ<G��p��坐���J:��o-�D�8�I� ����P�(%ƞJ2�\����2a ��W��w���Q�}X�߫ꖡP7��z>��x�ϗ�E�����������g'�g���?~����?�����Bؓ�(e�#��*��b٫�`x�Gf�2L	1w�[�e9��]��j�Y�y��,�1/��@�|�P�
9���ޛZ+�)��v߂G��hPk����T��Z
������g?���o��h�>�#��''g�U72}�:PVB�z���y�"��'O�x�o��yU�N���gu}�z�X�� W1g+����Oc��* ��G��?!�=��@�G_��js��;rbr�,��Ĺ5d��Ѣ!����آ��Z��E�����)���2�^sa�A&���]��u+�r���8�<>��Y��W"zRqNŉ���k<����������y�װz���*�������8N��{l8t�O�S\�����\o�����>+�|U��]���|YU�?|��߾s�Nc���c�{a�	n���������hcK��?��̺�ó���N}�{�KSmb��Ƽ��K�P\
?C��5������=}��ѣ����41��\_��c�K�I�hl_<�0�wJ���>$�])�1A#�������7�C0�,*@N������}��ǧ�U�q$�UP�Ç!H�1Ԗ[�v �~�A�;�-]%�b���n�ߺu���6�X�#O��R X5���M�H��L,6�M��!Z�8҆�<�ݕ�4�AȬ�R���Z�$>+5)����px�ͦ����0t����Mg>�Ӻ���b-#z���Yw	-��������+����eFb;fAc%�9�u�	���@�枝=e���v1'3���1�Ed�â�@P	Wk���w��~c1Y�ea�-g���m�X�������t���jmi����#��^.`	ٹ�x<����T����"�&�E����+�J�H����I���5.h���K�V�4��.[@���[۬X����я~��Ex�����\(R9bSjV�f�2��I�p�3������2�̸�w�]��8%�^D��Vz�X��|;�E�g2X�)���8,4��STR�+��x3�l�s�v�Tc�xmpA� ���Nh4���I�Bu�&��f	5��I���;�rJϻ�qW����vb���Y�Z�4�HT&�^c{y��0I�A�e����yh��xA~���0Dl����-\��Z(�/�.?U)7�Z��<WT�pw`��emceO��ԜŬ"�8�S�G�VҞ 0�tRј���
G�25�JՉ�p5�f�5 ���0����ފD�L<�=;�F�*��#���`�qK��9��|�N\��I�3Vw�(%��.KU��}��Hi���@T��k��l������j�%�s�g��������<�٦
K,{��k���|���v��UU�NF!s\g]��3*U󆺌mH:�buM��e�bK�ڬ1F�����벁��v>Pk��E���;�}�.��Q����÷���]�8бw Rr
�"��v��
�b�Na@�kx�$�	���-3�?}E�I0��1㮆3��u�1q���`�\�_f�˻	,o���2zq�Eۯ�ʂ9a�����)f��G��Z�4ݸqC<����̧�#�{ZJeZ�[�����;2a.LY�]�������ǈ[�I��KG��D+@�mllA�]a�<?;Q�%��uS*nb�t�6�J�zH�W�0�y��x����&�:'���AG�d��J�Ժ��L�׍�t˵t���c|7vJ���*��,�3�<扝PՍ�� v<�_|�j�w�������}b�+ΰV'��BCo# ���/u������=i��&�)Ae��I�Ag����W_A�aCX�n��vG��±�zϲO�ϲf´)�$����OR~�/��5h�w�G��т��ڔ�L
� �!u+,@W����]�v��3D�0]�eL'C6ŞDED�y��?u��̫����M��q׮��
�υs��_)�;�z=��M��Y,*�7�H��/�����%�3Đ��(M�.�^�y+��fFjH�BSɕz���u[�gQ�|��	�#�W��$ 	#$�ֱ��8wDAB%�H*U.>]v,�|&l;�O�l���꽕T\�q��&�B�]�QG���;::�K��3m52�B(�pQ1�S�Ћ���m�2{��/��ŷ��r���bpH#���͇��+9�e%�[���4�'`I������Z��T�7ݒTh�� [�7G�W�^��௟}� ���s~R�0uuh�Z�K>�f�Ut�)-Sa�IK?��d���?���������#A�X��%Y��Op5��(�����4������Mz������2�Ue����=�e5W$��9h5E��VK�W{�]�ݳ,�Db�ƚ�9>>~��񃇏>�裶�;��ll`�^��y��ʕHQ������#%����'���S��Mt4�
���4��ŵv@���!2�Q�Cuv�Q�2��Zl���H]���M�4���S!���s��$]��񤩤b��c�ǿ�l�X�gϞ�t�����e�OP��ZR�/!i���b�z�e//nݾ���W���͸*֫|���L,j�i��(�Y*�ڎ7u��	��(��*v���U("�DL�VB�@q��<���z�����i�=�,��*G�ҭ�Q�g�T�#gJ����BO�x]������+�m���k�����q�Ah.z�0�������B��ݻ~��7���ʙ��&zq�z��,T1/�P���^�A����IUI�E`��8��Mq^��/��y���ݻw�f�z���7�˳-#��x���_�|A����I�n?����	�q��|�	���/S�Im�;�2�#VRVpo0������C�¦/͜�Q�:�&W�/��ĺIzW]K5�:׈GoJbWu�(6���QY��������O��D��r��8�T
�I(k�ϳ���5�-�ˡ�vd��;�
>» {��z��������ֶ�V	�s2�+.C��O?z��z��#�+˨�#� �b�l�����;����"J�˴�z�ezp��,�y�3m�Lcw����k����
+Y�A��xڲ�b� �����4TTD9Q1jv�HZc��.Z�v�5Ob��w!�K�1[�Jb����<@eI]��qi/FFN�SiS]� Ɩ��利�;
��,Ǻ3�.-ʂ F%���O���b'͜yv�Ic��\����S*��0�W.0	,��	-ҍ�ʷ���Ncܗ�NDzx	Rs�٤Ӆ�@�֩��Zf��RQqq5�ryF����ل�a�Ϳrg��L�"ZC�g&�Co�~,�<㬱�͆��	���������y�Hb]n�u�M=[F�����J/��������U�oA��bs�xm6���fH�Đ�ʷ�.]��X�g.�L��de'�$v4Ek���bL����ZB[�ҤcO���6,��u�nݺu����1�k�)5Bp+u�]�t� _�X�L��Fk�s�n1�]�gΗ&�����ٌ^�g� kb�La�\j�LR���)�R��I&���'P����,�R�w�@o�	��ʩ���R�++�D�ȸ� 6rCU�,��
v��Hq��e�ds�#^��U���Y6���(�C�bلW��O��Ptp>*�^�m^�ð�����q�5D�;X����f�Y�����d�7��+A�!.%�a$)�0��F��__��c�
?�%��4K�L�eQG���xX�JB��h�9R�盺��M�t�K����g�6�'J'��m'��]�&�ur�f};��*�i1�L��-��y	.|��p���@���i���wuj窄�nX�%o�`bX?�5VN��%(]�1�ک0�r�Cm�]�кk%������?ȝ������A|��)�2bO=������ڶ�C�b�#Pچ��8s+�S��x�rda��h#bۖ�6����o>
䮂�c�=�B\�z�z�w/�@Eʘ�zU`���e��$C�sr<E���1�k#e�;&�y�h�o��<�|:�>bv~��~$}8��i� �U����]zf��
���K��\5B$Ld1�W����X-�hyX?g��=l>fK��H�Łht��O�Rsh�R�gL�N�-�qS�1�n�F����O>���~��㞰��{��,f�Ũ�����Β�W��7���</M��M�ajA%��G*�o��˯��L����c.N<�
�(��PL��e�d=�0�];[[�n�8>:�y2���z:� 0���\,���R�d,N�d<nj�����Ji��,�~')���1����|�m���]�76F�����=���L� M��f�9|Ǣn�I���Vی��Hh%�1)�L��x[��4����~��޶$��?��믟���7o�ы],��#��l�|��U�jY�>�D�;��n\��T	.��k{YO�9�+�:z�fgg6��9k2N�L��1�'.W{���WO����x���b���q��u��@�t��x<C��@G�(X.fG��!ƕ(��l��h����?�� S�����1ՋC�D��rʊ���&V5�*��˗�lm�v�$P��Ȩ;�O������7(�¯�,궑��]�۲�S�ILۇ+Ga0�E��Y��b69;��	�mO �Y��+|�!���mU�R1���H�N�7�BLP�Q;v�s�R;�̴y�+�F��b�%ߝH�߉C�i�q)���Wn߾��K�d����dY0�����AI�Ϧ��%�le��iM��Muh	;w�-��dN��G66�:Bw^�~���p�/�Za<����7�1�E��MǕ_��OT~Y�ӞQՓ�'�N���Q��٣-aF#Y��;⣗��Ϗ_-`!�n\��C�lւpO�ǳE=�/�鿌�~�;�n==x���ɻ��{;��q��s��#u�����2��D3������X��f@�=.��p,ٹɞGW�klѷ��#�
�ٹ�d�a ٮ�t5#Y���sFю��z�B�f|3�um'��f& vd��Lp�V���a��I�F��fx�˕wttr||Z�9�Zz��lƠ+�*������|:9y�D�
c�S�Y`�LK�p	��h4�^��?	��'3Q\b���� �4x���F���U\[ɖؠ(�AFc0셑?�OL�ZF�����@e�-��ƙ��B)	o�G8�B?�$��pꊅ��BfK�;�E�[B�����|�3�.]K_&N�2�������e��|�:_h�(Y��կ~��z����������C���r��A�)��2�w�w��������+<n~�!SEL�2�b	���H�����~��pc��A·���:�N��_����.����[�=�1��Pc��M1L)�@jK��p�!����v--����W^}��ޞ�;�E|3����l�:���gcR#�h\f���+3.���d��*��l��VD۵���l���!3.�h-+�K"�o7�g�v��B�"���K����ǽ]��TP��{Pg޾א���_�+���8��3)�z�����k��.�a�9Jr��PA"T"�Y*���{������la,��G�i�@���c�瓙�����`oy0��R��eX*�:����\~Yu�&��*/LKl�.~d5D���/) L'���ca�Df�����.��1f��%�\�Z���[�ҩ,�C3�v�\s�7��6-W����'��B��Lc�Z�C�_��y��.�|�@*X/�9慖�E�.`�-�bk���~���;����(�(L���%2�P�F�OT8��gS�4�NhKKɥ�[N���#3ȟ�>�`@n6���Ĝ����B A�to���u*{���)/erXk*(^��Y�Pq
�|��/����ԏ$]΢�K�A�����6-I2�耀F�!��%��҈�E%C��Zr^�J��z~�)vEn3U�D+m ��Jȓ�D���B����>�{��h�.d�H���
�6�5�ѵ�*b���:	���� �s�bv�~U){f]Q_���F�:,vg 4P{{{/��ʝ;w�j�/�(H�d?k�"�hk{���w�Nr6�ĳx��w�P�44�
Ȗ��lJ�na����R�B���j�R�UQXւц���
���֥�y¦�e*�8�RA�U��Y������-���T:���Rg�s�<�m��������u�o�tƳM�Դ�E#7k��A\/Dv�fe�9��ۂc)�)r/n?��z6.��.猷����"P<w�yf��iR�(����d旂?9�����5+�7=�"u
�\S�F��#��h���[0��4en��S&��$.9�'�-\η L�4�#�h��}�M�;��g��*\#qp俞M���޳�	���ߨ!(��̃�~l��lbc���M�;�_��#��g+筙�Zۜ��#;Z]U3.�J�*�5����>q-�SÂ�*Pݗ������%�X��ώ��Rr�vV�sj�A�W���
�ώu��b�F�}��!��"�劍��Xh�р�km�.���"�������ř�Ne�FS�)�9��|�z����*��{�S���ꙅ=9�$�������p��]�g�/�����V��H�͂�ҝS5�-<N��h@(�@p��N�6z�#,���v��K������j6�KR2��	/}w[���� ��\�o#�4��O'�+˄Wn��I�5�K��-R]�2�7����z�c�:����`}�������g�\O1`�! ��� �z�X {��X;���E��u��ƍ��<�����m�4v���;j#��H\�����d�V �"�`|f�_)�"c�S%~0��rK����-E#x�l>'�����'fD�R��6oݺ������B'�]���n�����n>~"�NHu�BQ���Dd���lKvq&,fO� nQ2�v:"�\g:�*�J,��{
a�����?^W'H4�X
��ᮭ��#_���{�u R��&����6��<�c⮰S��M���CP�x��ԁ���c�W�g)�Wƛ�Z;8���eUSF�����:��%K/���A�͍�(CS��o���5I��)�2x�Pر�Žd�����,�T<$��4:7��uؼ��^�/_f�O����o�>� �D���E}2�:xe��������`��7Bz�"5��s��ߋ�D�j��t��D��-�A�s��e%C�(�Š�M�RmGh�t
i �JMSK�"��m���CyQ��:9=���X8�����d����|ԐI�y��
�X�Wp�� jŪh��V�</l<d_*c3���ټ��y΍tICZ.�5ܞ��ێL�:B&�;Y��V���GU�`�]�~��}��3+!|��=����;�x)�	K���	�x�h�+3�65��K�;'������,��KL�gI�`(�N�x��S�]�8�S4wm�θ���,�%�Q`��4j�5�«}K�"�����&oy.XT#���%�t��0m�]W�l��������"��vpB��s]��I�������-�����e�������W^!u)֜��[��/�k����'������z��7�$�˄.s�Z�P��2�@��y�\�[������(���B/�Tձ�ɼ?���o߾}��|Qi	
!3Ҋqt������
\�,I6(	.���5K���<fi�kП!��u�M)�
�·�/��]�s(�-O�k�d0 CBl�f�>P��[
3���s�`2�a����K,~����&��f��r��1ݶ����f�̷��m�7n�K"5V~4�*[��"��&I��3"���HHM�[���bg���T�S�M�Ѷ޻w����A�,@�ҋ�"iW���F�����&SG;��l@�.�,b.UYd'&����ڲ�Ɏ�CꅖX!�&� �pWހ��5�ӹ��M��eKt�-'��ZC�Sԍerȗb�ȔJ�;_�J����pk�J��"Iɭ���3��)�a�r�<:!�e��J��׫³�	.X�ɠ3��|�������52���m�S|.���E��N���P�S*���Iq��tlR"��� �Xnt�ia�	N�0Ե��%I�;� ��D�t.C�N�7�u�����Y�D��O?���Ls�����@ǹ�`���_��� U��\�����'��.M�ecgI��IhKrU.2n�&�}ϲ���Y垝�@&k�ZUˤ���_��..��O	Ёf�+�2�]�$&�x�Ѭ�k�"^�
A��(��V�!�9mmQ����	+4������Atʹ|\<-N�7rI��~����ܺyO1?�?�7Ѵ�BAu�ä��.�`���L50�[.����)W{�T�3R����Է�ø�e�a�I�	3������/�b�n�kO��L�p�%��0T��]��K����\��5f��#��P=3��JF���J-�6���AI�$1
,�L���R��ZDt�ɑ�<kd���[�H$���=���Ul}������sG(��o2����i@Y*ס��g=)|��Z�B�
�~�A�����\z��M�T8΄uR��#>h]�����ą&�a�X&��!���j�l�s�ή���s�bbgNY�~1Y���v�咰|Ci�*x��ֳ���r���h;���-�[F�m_�]�@U����W�U����4o|��CK��67߶��up՚e��Y�6קo����]ò������@�O9���XV��B���<-*nv߻샫FR#����)#���f��\��*�Zr�5�(�Ø�e�,/m@�K;2�&��K�鄦8ʒ4KŃ�W�8<:9��Hڴ,]�2�����lY�����f��`��
ՌB[����(q�Z'~��{2n�(�����O����O����7w�ޥ
��{��@�ؖ��M�)J��L]肅�����ܦ<�I�K�I��i׹�>�R�z{`a���о��?::���/�?�^������:te5�y�\�:��6�f�U�x�C{�I�{y/��q.1V�Rd���\�X$��ѧ,mW�S<��J=�ڛN�_}���i�m�஺u�B� ��A��+�,�Q7K�Õ˗!3^�X�a �ܤ8�`�:i��ك�B�N�����B�8)�6�U^[J�l�"�ï�J�F������P(6�����&V�H������ʦ.^�k�O��V�v���f�ӃI�yrʷ���ϟ={����&� ��.� ip�)��bA�vBb�-�GgE>�J��z^z���hx ��@	��u��l>��#z�4_�~@�ȼ��&h�[Y��U�ס�S��h���V������
u;�������|v��l�|-F!_	�:��@x3� ĉ�t|��ΰӁnIZ�R�nlux^��B5�s�-���,�Z�uJ__��L��և���R��=m3�LөWWq�u���I6����捫������h����iP�Kv��\3D��c�mi�����BY�D9[��~��;����T:Ԅ�11���B��bѦ�ŋ��G����Tz��f�:�w�PUK�'2�='����L\�S_׻�,_�8������r�M�lc�>.����1���U�V��]#ꥮckm���j����M�h���@�)���_#d��i`��E�m?~\�%\V8��W51�*;{>�����h��K8�s�3g/��9⡓�D�Bk�r����̋�l�;�&��z%%���l��{GF�U�����@�˂�-��Yb0ȳ`��I�8zҍ��3��x����Z���j1���$�{sd�ͤ���07ہ&�7����E�W-K,TH%H�b-Dd��M�u%c�[>}��֭[���1��"�\B�����R�����O�
�GH�z�[}ƺ2Q���-��+}�P�����tx�ޖ�ic��	K�\jk�s�X}�bF����o�-qY�B�H�tұjO��3<NB7
Q�P�ƺ���1���Hh���H��
�C#YAB�: *+�f>�y�b��:( ��&��[�+�O 0��֒�1X�=�[`����P��������x��?���b�S'���j�X����������^��ۿ���z�
��!pq��t1��O���)&��~=|��^���0%��{�P���#D��:j8E,	����;;[̫R���E��̦|�0_���6�7jo,M˞J����x�[��Y.��	���,&��L���7JC��̬��f�:��nZ�SO�k������<�C���m������ .#�Juc�ҫ';$�J̔�ڒA%�_������aB8���+H�*�aa�WA��(���!�$Gs��a�r
7v�^}��W_yE�~'�x��D���GU�����ONY�Q����֊���ׯ�z�В8E~������2j6�s
3W�m��"/W�N8�aP�*$�� �TQ�2�Z�^t��}�w=Pb�lr:��k�B�d4�J�S���h	!��j�j ���9�fvVU�$Y"X5|Ӕ�rK�+�E��4s���*RT� fJM����m=����L�س�
�|ƶz��G��TK|��gr[q�<�>�~;��Z�.t���y���-iʞ-3a	&R�����iY"���;"����!��-=
jc��\P�.�r�O�On�#����ja-���4���`��ay)s
%K�g�
��������~��'�z�z�*���I/�E��(��������V�����y2��m�-�\+A9hKVm� \�`��9/=�L� ����Hyrі���˕ j�k�/~ b^x��v§��ļx�β(�]GmX�]ܶV��9���/"��b�=�������`�v�t2H2,��}��:}�_7�j�d���7v}|p��t�ӿ���w�w lR�WTSe�|m���	�|�La��e`#�B�V�Yx5�$�!��������x�ʶ5���POY���o>��N�'1�Ll8/� �j�,t��#��~���%������)`�9ѳs��u�$QF��6�j�yrς
]�KS�>&�7f�7���z>^�I�0s����I��ټ�6y��,�5����%uIw��I��M�h��7�:ׇ��d�Z��^!�j󇾅�y�+m]7�t�����,0���7J;��m�+D�e�jdYI#�^3�),�%�������-�o!o�Owۮ|��!�8c"��\'ǉ� ��zV��j��ʧ,�Wx�.�~���x���lnn��Ov)�:qT�Q7t����k�n��e]ݣ�*�K����ujtu�,����Ը�8۱d��ᠻ������>bI[��&�����W�j.���4څ�] ]��)�G��(w�/#�[��1�ig������i��vN���j�oK��x���9�0�D*�!�{��j��!7�,3�RR���k���SJQ�\6da�-`���k���9�S+���<_���h�O����L:z]����#�כM1�\��M�L���4������e�"�g�����cbK���KQp�˯��J@1=��aK8�ׅ�<�E�R�+����gr��	��&�+�w��"����J���r�t\$w?�#}d=��
��Q�Pc���"6#��g:���da����7o�}3՚���.b���~�>�l"��K�"I���]A릲�{�B��&M�g�/�|����ݹsG|���O����Dk��;���"���B�̙wJR)�A�U5�	�gJ�Xjlv�ލ���ooo�lj�ܡꖋ\[Gц�X ��������B�Ţ{}���a��w|���P[����P�U@�x`��3jz.c�YK�����ϑ������4���W���qI-ϫ������/�����j�:a��6�I�h(�/jh�#�D����F!��r�&�yi���9�PI-��v������"
/�	��Wʅ�E�eS#��i���6�޶3:|�1k��;t��XJ�*\6\���)��$���r��֧��O!R��nI��?	|n� p�S����;;����i���_:���t2�h��3|��<+�" "�F�]��^Q�;����c�Ƣ��V꩸�hsx�9
@��o����O��_�f�B��LGjxgb\a����e���rR���"��<���iղ��5����Z��[�Բ��N�� dj\Y��m
��d�"L�8�)����;v]��.�c�)n��x� p}m�e���|�+/E9[���6ϲo�q¬�me���&Ɛ���v��okZ|:'��=| z,��v4�~k9^�륿_�9�@lqNEA��	5���rֆ�)E�v,���.����88���2!#U
uH�1e��
�@���1��F���o����}�1ڸ}�6.��g�QƸM�ŒQ=�B��z�y�|�?���{��'�L�6ɹ(*�U"0�H�t�<��7��v����ޛo�In>N��F�ؠ���T�V��Zo�d�ȡQa�����Yψ�2߹�/D� No���ފ�>�Ȓ��*N�Xn56o2�N�oБ�ǧ�TY�Ւ�'����ǊHCf��u�i\���x?8����>}J3��'��zm�sb'�Rll3�'�K�S�9׍7��xv��
���_����l�u�ǡ�\����z[�YٖEb.�m/%��K�Ŀ���)r�*b�q�Y�Z,m=�a���/^�����"�������N֣^��lnm�i�q�dq��o�X�7*�?��e.Q���	���Μ���&=�NGj�/ye�fb)��)V�'x�5~��V�\���St#��M��/��6Q�<�fm���Yc9�JK�r�4��L��k�V����{U�Sh)��%'�-�y60���%�ܥJ;���]��),�Kҹ��;ATbܬ֎�#��e�(Ɂ���A���:� ��&F�A���BPB|����BF;V��<	|iC��%�)T��ݞ&[{�~�O�����Tu�'O��r~����c<�gUT �а�Lt�����!'�&@4�T<>���9�����oY0��BRd�	�+�&�鮽��#�!\��#�Z�|��M,����ﯿ��h�ǹ;;>�at�'��Fs���ᦃ5By�m}eb�g����mL���,�n�	8G#Sk�Ʉ����Ǝ׈<�"����+��������K{0+�f��VLVV���l[�M�"�1+�0�is� �*<�ύ �7��ۉ�&MT)���A;#�w��x��97���������&��򰹞�����ύ��ǔ�m?�Ha��+�{��l:��(S���k����K�`ä[H�
[�adB��ϖo���ы�[��|�|�8^@�h���j�K���Nҩ�R3p$��dA -^�6�n��U[s���/���r�ܘ��6lT��|�m���l<��F�t�ŦN�=K|�=)"�+�"(E(���E]���EŌI��`�m�b%�[�5̮g�Bۣ�@���A��.�����r:�[k�sp#Q�ǖ�5����	,fْ�Y"��[��nm�Z���Tt��œ�DI������)5�$/�皃P��<y&�g�M�?H��M��4[��2aW��qq�M���k:1\�򛄸�=��=��E��r��\�gYԶJ�{�v)E��ԕQ�6xήT�𛰪Mkb���>M'�/>j�8�H����\�b&����jU�^��:���n�vV2�+����A�D��E����� �䉊��ܐI����+���l^,WA���Çk0�ק4l�.,�Qm��S�*��Bi<��ig@9tF���)R�G��E�'�V8�Q�Q����ɯ~�k��[����A���:�<�Z���[�dD�2_-V˲��&�
��ළ�ʇ�L p��źs�Z��Y�ߝMs�JEz�HFË1Εf�[-�{ݡ�(U�ԍ�������!�Q�[Ђ��k]��<_�\�:�nm{;[��#����|u��=��j%�EL���ǽt:��W�)$��(^h��n�z����M��{|x$�!��lz�o�~�����	w��)XJ�%�4�31#�(��S.� P�����Dص뗷���m<F�&k�3�o�$��0�3]�z���ǿ~�},���pc��3J���)�'B��]���aS_~��X���[�A�uQ�O���$�*ʕ��a�%	\�pi>�'4��x��_}���eXO'o�o���j��X���'�B��������ml�ߊ�#�G��:��"��#.,~�p�t��hi}
+�ᡓtkS����6�e)�1���t1����s8"��r
km�c�6FW.��"�To��@��:p�R����zQ��붵a}�ub_�+V��r��9Ηu�w�ʰ'<Y�n'�p�
�,n!�¡��B�*Q��;{:k�����"�K��L�sծZ6_�8u{�F���/P��Nb��$B�\�(�w�7��<VL(;3#�(u�hl����������5�k�'�&*�DX�HX���M&����ߌ���(+���1E�WI�@k�˽p(@E�e��;���G/^`#��O�.��	 w�Ƀ/Ew�:��y4.�v�������(��t�Fh��0��z���x>���%)�J<��&h����a:Kn����	<�����^z)���x�u-��O�>e���
�zډ�a����~�)|�+.��#;Ҕ�9���f(�X�$13����i�,�]���'����[o��'�'�61�����,�k�M�S�ݻw���o�ߜ�	�t��{�D'�S{��������阴DrWq���"7���0n�i�\����2J*�.��Q��%^l2.d��x�'G>�r>��JU�:���-�V`�RJτa$�3{W����2�B���Dk
m�CKmI�)��$��M��K�ܯ���Lr5`G��\��Ԓz�����\��Z�����?��\��k',��9�d�`���h7���&�<y��u�~��0-�N��'��!豪:;?�o���;�������o�����O����-m1%иj��N0�?�я����޽{��~�_@*<�����<�m�T�-LJ�-�1�% �[� V�+<��5��x����D,��*��_z�||B=K5�4ߺ��o|�������L,�H�I|O3�x��C���c��hy+U�TP8�j<&߯����yk��ċS�R�F&���ӚX:�Т}�ΕQ�"�'/C���[QP��ѵ!���^�r啗^�䣏��c����ژV�%{����WL�����i���ty�w�-*���1�ݎ$��N��l�!>��9�����+���lܞL���IVL�3�*��)+����C
uПM��>�¶��Z �~����{�wpF *�1���`I�+N$�q�ӂL
8W
�����K���)�b>Nb�ҥK]͉��ٺaā3�C��2����6�����V�~�{��%7�����ܟi�%^D#��J����T�����q 5~�P���2��v�
�Ӓ<Zc x.9��ڔl�k�l�?��*�{|�c��[�b�����B�Y�Q�Q!�K�K�O�4G��<z�Ա�D^)%��sY�M ��^��+��t-��l��E*ס?��2˓.�Ō?# �W.<vh�_�:�5�o<�ʆ[	�F�����pæ�JA�p3*x��/�Y���%�.ܕ��R�)��<�I@0��]�}��l7l!Y��E�Y֒|��p�Z���Д������/^Z��R��WO��әw�������˯܁+��(8�����aC��P�z��&0@���� ����6�$�^�線;�=)<˺-����p@�����6�i�2��,���+�l��D?����,{�6�d
c�[;��W�w��]�����K�o���v�@���a\�e`i�#���*�ic��T�uA�7
����)�vGԺ_�NH������e�5�tMOf��09��-�	�yEv޹�Og����^�q��V��Ms8�}�^��@\�$��.�{i4	�ڈ{�+%�h�P�Ěg����D���h�����04]���<J�4)13_�SlP�W�囦n]��?�mE ��\�$msUt�R�w��[^�
�B�)��K�RCe{-��C;�2��I���u�w1#쯍�u%��N4^ϯq7+��Q�A��>�>wM���6����i�4��w��(�B��`��q+ɪ��s?�ӱ��1:��o6}=-��"��j�f4�����"��mDJ:9�j8֤�����nn�m��\��6�;��8~9_�O�H�@�Ӥ4c1*�~��4��#Ԫ(9ߊ)�$�V�z<G� \� ��XB�6����8ik��%��횂Od���ƣ�����D~S�>��3(V>��1ZM"���ًQN<[����b�[��r�ö�]��79F)��mh���0��c��U��J���x�b3NN���w��� rx����c^d��ޢ'M~M����"� [�n�|�},��T��^�L)X"����X�vJ���<�-1�lP�r}�!��gͩHaE._��E�6���!��-P��,�����Y�!�>��gŲ7�*��q;�m)�g2?�g��Z�*E`��x�Cz�|�k&�r���Li���_)/:�l����cI$�ׂ����llw	�g�/+*�+	?�P�V�#�3��#�#Bַ#}�]-�UlGx㯐�E֡:�,'�i������ׯX@^��C�����y: �׮]C�%}�]3+@�oX���ƺk�2���G��η�G�OS����VL��V��tz���ސ%�'�
V��[�)n�6�u�:O���G�ZW��w���wXc%�ZK���%�Վ'�3��A��1��N���9v63!Pj��YNg�څ�JQ�$��Z�t�I��
o�|��Yd�9��n��6�D¬0�� ��xg�B�F$�sZ.��:	�#��nn�����ZȆ�����1��@�:q����~>[�P�X:�����ԣ>��$әN1��ډi2_��+Π'vl�R�K���L�D@�L>e�*Ln�+(� �t*�C���eh��p���tD�*`	"M�ȮU��Hy |��,�=�����\���@\`���G�̭�Y��)?Ö�Ad�]���~�����jv��u��f7d��F��ߖ���m���=yvї��T8xF��L���u��@���GO����!:�$P�[j�	,�6���jh�]�W&8��{֏�xx-���08"~փ*trH����&�QK�\�wz�R�L�|p-I��� �{L�y`�JT��=9~Jh!���Lcݸ&���L�V�Z�k�#��������r�����q?��;�s��mvhB,Eꉠ��m/~�:�ٟ�>�[��,}�駰�y��\F�a���ӳ������?�����߻w�
���D9���p��jK����D����S�ۥ����H�7O��ެW��:�g�s�9��X�XY�"���m>H�,h�نe�?������@�a�� -J�@Q"�"i�@Ң8YSVee�T�y�1���Z���FQ@w+PȺy3��9{���o}��=؋s/ i�b���L	_⒪��FiO�����W`z��5����p�A�侫a����H#^��ٺ�I��{�>�P2��+�JO���z)N�sj\����C?�X�>C�U����_�n����(_��IÓ��SOݺu�k�F5^��zY8��\@j��y[۪_�{߃r�I&��YkCg�
Db��J�x�ʯ��G��R����z�-���0��L'�o�	/��g��;���rp	 �`+JQn+�۠�������q�?~z:�ln,����,Wr�6�Ϳ�
t�9�F����a<K�J�:b�p�;�:�EY�u$����IIX�,	�T�T��(�!�\wC�@1�Axy�J�KD}ȫ�k���ڈK�_�pz���W�S��L��S��*�q�֪8Zao>�u'e��f�|���4����1�Ly�#t�����<*�C��5�E+�2��\�X��҉u�f�dack����	5-.Mݒ�c�������"xe&-4�~��^_.�@�6�
ZD���?J��|��0���� �N5	��d�h�Qv�2���TU¦�Q�@�/^�e;��j&մ���l:!z�v#��5ΘH��+�#���ى1j�O��'!�F� .O��TzLE+��i����:����j�s>����`��Uꖜ�՞zc�6��nX�O��7����H�YG�I�	�+�`;`Cǉ�Ҙ��#�e\XÉT�Cr���ʶ���Ē�y�8j�E�l��u�f�ԭ`
+�0�О#�(T�4�.O��S1�v�mU;���)m"=�F��Qod�)���뼯��� �u���L�ɼ�`��7
�~/���ȅ�$�,�(�8��A؆^1�Nv����M0�Y�IF��\_+&�jN���qSM����8��Q�!��B��U'v=P��%t	�н|>�qԂ�.o㚅cǀ�n��5ɶuo�fieTW�a��,A�ҧ��N�n �Ћ�z0����ˌ�_'ǧ�4�Ֆ�֋��YhG�B�oU�
�}j�Y��2�3}>�D�˂$��-���]���]���Ѳu�Z�{�2����#� �2�5��gCE_$)\�%�(J��UA�����	.���x8�l�l�ó,4�� �H$�t�8�!Q�F���f8���o^�������vҴ���tz��0�ܺ�P�.�Ц���$��bq^;qU��6nl��'�����-QFn3��
�R	ZE���'f��{�.�ֺ�T�l;�Y̗''R ���TڅZ��V���wG�@	M���d"�@�L#m#q�p=ɉ��Qb��r5��q���$nR(Rx;8+�����dz:?�K\�/�������*� z�N���l�i���I�W��G�>HL��B�FPe��e�6��������jK"�ۑ7�Ae������ˣ]o:�*	'â����4�b.xIA��|�Z}�Lu5��M;>K��?88��T�������뛗ۤ �cǢZ.ds։SU�Bu�M���VG����S�q�U����Q8��d�F�S�J���|t����G�D�b6�hL*�5�D���:�r6�iT/̦d>�Թ����?���9ᆅ������ks����|*�{Ӱ�K��m�?�Ә%���"_�	�>Q���Ɓ�/V���|کT�r�Mk�K�v0K��ɀ���˰�ɗ�ӴV�!�É̲���
Ԃ-�o������^O���p��(��5��Ү�T�2��i.�4N���;�H2��H%���~Hz�����<>���3*4�U/�+�1Ќ�F��T��`�a2B��"�m�/W��.E(y�m(��IP���|��IAYfC;j����q�xc�d�����,P)5�hc�V���x^��̚7j�.�1�R��`)�SG&�w����Ix�p�nݺEݥ���+�9�*�5��2�p|rr*�խ������)!u��8`ٰ�|K ���:� Z���^���R�%ðө��fww���n��C��6K���$�Ԣ�ĭ'F��նg$���1���n��z.�I�p�Ʉ�^f[���6fQ���b!��;v
���W_�W���7��c�F��jZ0�����ի����5^y6A%����~�Z��$�9NZ���������T)������a>d�Z��=�W�41Yt���׋�ԙ�ex��
Y�ą�9�2�u���be~�xD3���L������%�l�o0�eǇ���֚+�}	-�p�I^��wS�ޫHWr�^�@��T5%6I���W�hk��ߧ����	c�1������si1�pἂ����ʥ;� ��c-;��`����&=X�~�X鈪w�y����}��_��}��nܸUI��We�	�Q��?�s<����?���3�KF�	���ė�D��ד���Ǐ���/cI_z�?��?�}�6K�7CX.&���r��]�F��Ұ��)�1	��6�у��y���TE��3v�1K�:r��
�X0��yv����Ç���c����.�u�5�ԉ��V�!� �{����wx�S���ý�h|���{��E�2���������ޯ����Ц�$�X6�e<��`���%3�>�dف�̅s�In���$b�ON����Y�H`mI�9kH>v��.���fgg��?|cc�}�ʕ͍Q�e+�ypx kx���дd�#��d_p8b���o6;U��V�+�؇�����q&��'�q+M���cq������>C����?���/�˯}�kӓ���ا���!�����^|�E�����.~����̦R���f����%~8��=	qN���w���������c<F�l��!*(�������Z��<Y��D�lz�������<CUT������M&��m]���s/	�x��ha^�@Bb|4��V�9��${UK/��虠�Aj��R<����,��%{�i8�eߏ�q���;
�]��M��̃��~ǚE��٪�ڐ��C���ň�V��c�u]jA�!� ���� �;	m�H���r�1�m�FM	^����<�'镩Z]1(
�2JhF��>�$^�*�����Mc`GgY�3%��m숧��9���hߪ����V-2�L=��g^��u8]p�/�x�-v.+ �����ʼt�k#����)#�k�$pgr�g�ZG� j�.�
�R��D��;n�mu�	�jD�ݞ��t4)�j��
�/|!�+7f�Z5�E��&h�~v����_x��T��Y�x�?޸�>�rq�*��J�s����-+�t��VQ�ʠ�C]�ք�ʭu�p+eJEK�+Y�B�"f��h�����>�5,�z*�K���O�xi6n��3O�JH=q$"�{c�,��k���
A�jW�j�w�:�nL���)�0]�zQۂ~��%��M����3�v˒}��%k�i���I6�p��^�Ha�����w��a>�ٶ~���i>ξ׺�qÂCGÜ:»�����������m*t��h� ��=��qm��k�JdV�0���7�E�L1�+U9Y���0r����N����K�$�NQe���������Z��&yԘn��!y�|ǹ�L��qӸ�-�I讕n�<=Z��u��E�?�I�F����`L�M�xrʙ:��7v  ?%���A,�m�q���=���s2��dz��_�`;T�l(Q�~�z��7��c��U��#��&��ɲ&6���J+�6f�=7�)�����F�J��W�z�=h�#��Z:κ�׏^�8�~�ȁ����`eһk�ٖ�eƥ!����ܰ��Lz�x����^��6ɿL㈽��Y�������'����y�x%���P�����X8�p㤛�(�k֍|����A�EV��$X^���?#7^��Oue9���ǂ3}| �����(��#��(�֍���e�|6���cH
<������M�̵��`_�)����>��B����4��1���-����-��MH��^8|x��:`�ٺ�r�82V�L�"�>[l��r�k՝,�r�9l�(E����I�ck��EzH6��J/4�L<�!M%�eZ��
ۑ�:����	ʘ7�FN,m,a"�M�֬�U��(�^�������l�k���RD< �Jc�,d#
:xX)�/^Z���}Z�hIEa��2�F*	r��\���B*�_�<���[��;x�}<��j�t��^K�R ��6�Xo@E�Ø�NZڑ����}D����yͪ�<���vP�*ũŉ�)!'�Z�i��6����pr����7*��apm��[2ཁ.�֬/�ەtg�����~���^��y�/}�K� R%�ǁ�S;�
9���9;�i �����X��y�"p����#<��y���oÕ�9h.���TV�|��w������W_�~�:����������m�������g������_���pp������a��:ǻq"�izlg/P��̤�l�}�;
�����K��n�~"�'ѬL���3q�!��L������<���2�C{�j�0���gZ��l�Yt)ҡCNљ���*��\�AN҈�|�@�C�����vV�IE�Y!��pҧ�'��4Z9�A�nl��|���{��=�,ϛo��o|�W �D����[��}n]�M�4LFV��	�r��e��t��:�:p��vd4��\����H��>��'�|g��ի�=��=�KQ	/d��~Y�h�6Y4Y'��&�TԺ�>�"����0:{{{�%�g��M��=T����z\�����J���N�����u���ρ�q�۟~�I�����1�MX�a0�nnn��8v|�pT���ZG�P��I����R�'�4 rB0�:l��]k�Y 2Q�-B�� 8׋��Ε�J��y�p!�$+׆兄��,l�r&�7����\*I�.����p|n޼y������
�a�p����:���{�=%���j8ǒ)��|)�\�������&��f�wx|�'T���k�'����w��O~�!��rY3t"(^��� ?�=�IRR'����*nݺ��G�*���L�a�_~�e�9g��G~��c����#���P��P)9O�V�m�[[�,ϣU)�Z����)��t*�y!5U�N�`ٔ��ۑ�3��y_�gc���>ze��w[�&�ڍ�q�|ңv��.h,���}~E�6Ǉ*�K�M2������0}]�ֳh\;ϲw�< ��G�˸�8~�VP��8��}�Y��^d���e]v^V2�+�ꕸ��q�I]1�O��<'��tjF�����Qs/]�Y&�&v����T!h���K濵W�\�n_��a��^{�2���HA�O
A�j��3��2ǰu��Q�be��6.]��C��$�W�ZyR�XHO���10a >0��36�ܸ��T����簵���,U/�C,Z���^7�������9dYwQ-�;\qW�?X����\�a��ǰ?��f�ILu��7�����tJP%�4���%�qu�/�rAk���4� 1�$x1���Dܕ��4�T��
WG�-+S���4-���3J&J5wޞMU7�T4�6f�0bD!�ڭ��S(�+�IUUY6q3g��J�M#$'P�K!gC�J�NԄ�bӪ_�J�>�Q�c���w�y��3p/�:��dWد���X��F$_��v\[��y��qw�V|6�	,�	��IȄ �N�[I벞��&�۽���B���R�+���uH:��xC�gG�����y������8+�z`�ϱre;���Y�ժ�L�"�;��n�R�j����c�M=]�D�窘&۱�C�JF��y�0�9��f�Ѹll������#��v����+g�*�[*y�yrrį��@%��Џ0���i�����{X, �[�р}���	��O�/X�9ޖ����N��PVA6�������Ⱥ�G��raC�ؑ�Fo\�QLBh����AŎ�֮�{���1�.S�2N�{,��r��k
��\iUC
Ld���ng�/I�,V�纑y�0�¨�]�''b��PCq���@�s�����;�'���k0�V�|��� .�����|e�\�]|�ɮd
��C����:��A`�Ly�2_UqԴ�,4%Ⱒ����h���w&��aߴ�k�����������=U�ä@��R��Y��5��4�,M�l���$��I�+]?�� /���ˤ��5�媪3F���P�)p?`�X��y �2�`GZs�BI*R�u��<_��]�\��\`A��6~��9��E2��@rQ/��q+S��8�`�^�F2��G��,�!����*"�@g��ҪݧI�W���u��%'�v6?R�ڰ+,��Zb��쫛"�M���-�z=鋁��F����G��R&�+�c���eM<�C��.���b���9_�6�Uө��~?��n+9���e�^���6�����	M�l����A)5�8�ap���
S��<z�t���Y�ƕ��pJ���Y����s�S�q�I�h�Z�媩�,��(�?�6�~��:�U�+�M�q\�������~�HdI���D�{���v gAZP�8��e��V���㣶�B�2��-�W�^Än�;=uz>6��pQ�4���s�mLK�8�]�M�3D���$��'K]V�U�$�A �If���� MpOk�ɓi���ۇ�ϦS#v_쬵�x:'i �'���R�[��U�����y��������7�|[�n�,�8��o�|�Vע�׋���l�y�!��c�����ѩP=�z8	J2y!|O�X_|����]�^��ϡ��٩hD��;��&��c�M�����w���}�{��ۿ��?��X�?��?x��q[������
a���O"f>==!u�|��E��+W.��2 �)��
����J���R�r
�QcQ*�4о��f�tf��8�D�ZF��ⱕ�dF�ͅ�FO�ymGr�s�/�ϲ�n��-,#�d��b�Yw�&�iiפ�2�{\��ܟ͇
�g��6����H��
,ά׏�߻w��i�F!���F�p��Q�h�V�� ]��[���7��g�}��ŋ���o�a1��`��u�<x��������s?�s���
�~�!s�r��6-���ʼc����;;;W�\�޸~�:N���Ч�!nb���YF\[6��lm���ڕ8��1-HX8�߹};t�B��ַ�7N����Q�С���M揸��R��\��k��.���|���d2�e�����aޭ�]���ܹsL$�{t:NG1�=X
	
r�<�Uf$B�1%���jB��	��L��,�7Cd�����q����w�0����P�P *�2Ogt��F4/�( =pv@�u�������?��Uh	B�p�w�ܿw���˗�a�ҥK���d{�Ν{��0<�@��;�M�c�D�ED+�.���#��_"���4���w�$q���O1��ࣻ
E��Ç�f����c-}����?|��'�^�tic2J���6����dw{�O�m��E���弩��֕a��h����q7K���W��g�m/��=�1�'���Fv�5r�3�����0����%6YΎ��wv�$ϻi��PHg�-�H���B�UJ�eb�x�⧟��Xj�5�:qºN",��~E��kfp�hY�o5���>kH��9��5/V�r,/C���(Q��|*Ч/�2�fC1�F@���ӥ��$T��^�J�k���"��
�Sօ����24c[�)b�^D~�� ��c5�D�Z��C��A�q��?�wԺl-��j0��؎C������J�rS���e��+�<�{{k�ڕ�x�����0�l���*S�O��o&��T$��`����A�HR��>u�N�� ��~B='i5:�J�4bS�����uge&�`����f��b3�Ł0��t�OG�YkU`5L&xVӜ��;[
A�k�}����|9O�`c8<^.V�L*Ɵ-�䎣@��c�֯����|tj�H�e�G#�_ai�J,Q�q�p���i�s�Ch��i\��r7c�u�,������d���yO��,q�qR�c�w�&!\Ů�g�*ǯ�A�����Bތ���;*=^�]��y�S�1���W��}!��h u�K�j�y#W���2��rIRε��Y��}�� ��j]��{8�Z7�u ���󝻩v�U���ˡql�@�UC��:/���lc�j�"�,auF���V�ێ�짨��-T|Qr(���+��F�^�u���OZ
Z�Z1bn���)����\:z621��쵪IC�{)l����J�@��_L[R��q饝�ia. h��Qhm$�a�;�R��r��G&���dQȟP�2�4
�t�5��1l9M��q��8�E.`�G���ܡqxC��8�X4W���'��{ �%��9�YO�l8WGڊ�!�Q�'��Dx�t�5NnHY�r�f�w�gi)��Z��T+�q�[P��/�H/���Y���J�~�ȓ�����:~��D�#�=t��r��\�r��f���� �[B�8��|^3'b���`���j/�R���n3�&�@�
~$ݲ\���-OgԆ�U'p�O������hE8�Ǳ���_�pA���}��ʭ��{��=Q�؅��$�ԕ�d
�ؠ�保e =�]jD1��ѽ��If޸�T挈(����r���{�:<U6�,��������
G� 8C5	�!���!�3�x!���G�����ڲ��`���A(��=�m��R�@�!D1 ��
�^���&�������ﱬ�NPm��֩����сv��1��s.x@.��r>{�h��t�=o������D�`O����G	[�i$��� 9���w��hT��Ă�i��z�<��c�Cl�����õ$L8ua4.����C��x{�:Jb�����9���[G�S���"�K#�m��)�c*�݄�d��9V�hkO�	%A�X�Q�4O��nG��#RZ���k�/	���,��*~� ���o��o6:�Q��g$������t�DL���ׂ��  %HQT|�(��|DD�z)��C��&!P��	�0����A;� �o����Ф��t!�FWg��zR�E�g�ӟ���~���_�p�~�$0��G�T�ȡ���[*!q�X�W^~�Ν;O?}���u�W��嬤�'��~��y:�Jz�GP�3���t�mf
��~4y�K[3��茙lR{�g±V�f����ʉ|��X�<���pv�N���j�2�C��Z��
�u>I�(���;���I�O�ҽ���R>	�Y�_�ܢ(Ϧ"����+ˇT�Z��e�B2S��B'\�^|�E|�����7���"6��E�EN��җ�T)�����	�}�6	݈(Z������կ~J��W�$E1p]S��Ti+e6���}���/�AW>c>�3�^��<�[�e=ĩZ�D�=O��->&A!֟ ����oW��NJ@&�
ߺu�7�x��gײ���ƶ~��\�ikV�D*o�7ҍG�~��J|�H!������)L�3t�{�.�"�NMYEʓ�u���nr�W[~7��
�ﳋY��J߸������x�k{�ƍ���'�|�'���"����>d	kH������>�ė1���`����7C8�1���ˁ����������O�$qDOb�����ã�����೟�,o�)\_�'�4F��P��<x���ÇJ�{[�?�Ǩ�R�G�g(�k׮��
^9}�q��喾�8Z�����ކKE��QI�8�C!X�7��=9=������%OPF�'�q'[�
P�ט���Ǆa��&B�x�v�g-��+��n�$\���WF!���_�>j6���e��>�q�}��X���4��2���ͱ�zCa`K͌G��_�<��Q5�2�n�hhi���p��=W��M��x�%�m�Ma���/��<�>�P�q1am���5���9>�U^�$e|T~��g~��ex���g�4��Z��\>J�[��T��X�	&�!���ي��#1�=�,ɧ���ĩo���(��%������PcO,=vI�W�^m+q��y���{�ҎZ���c=%U���![�$�n���(��϶�I�ؾ��E�D�Xl5��!=��SKZ��5�V�Y�t}A�g��b�w������Y��"H��s�q�6�� <`)0�O�ip�C%�c�:hJ	�@%l�o�ϑ�������U��^��gM�-ry�V�1�D����B�]E�tp�̸����ȃeHv5���F�3KB0PZjV�v�O�\���<�:�Xa�r����X��F��ݸw72ظ�%�]�'����k��_�Ի~��[�ˣ����b� �>���%^oV��OAL�5.�K���Eˇ
̑h���g��k8mQ�U��=��6g���������8v�>��a�{�A��ܡtӐ�A�N��j�M툊�Tzc*n��-�;>�0�\�M����~ծ	ȸB��Mr�-䪨���č��nOMNA�B����Xдù�)1�U�f����,�p�[�qF��,3�l9����yQ̗�~n�AYY��J��1�ڡ���fڰ�=��p�hm�g&��$�8p�C	��]z��1|a��Ь����¦��h�}�9v<^Vg�c� �6��W�i��i2�+��¾�p�b8���@u=bD�Uq�ჩP���"������e!*���\Y�nwXW��|�3��@�2��|5�q��d��d��'QS)�	[����zf�Xt6?�:�n'z�O�H�W�I��GU����r)�B�'�v.B]V����[��%���6��|�1���x�jQ��W�-4�5/%�6N:���a��s۪��9�&���<�J�n�3�ڧ����NN(�0R�
�B��Y�-ɦ,X�3j������l9�a��\ɝM�t-%�S�nvzzR�EP��%�C�����is8�{;[��#[b���"��U���lM.���\����|1���=�$I$iǍ��5�JU��
Sz��(Lb�d�S�i�F�[ޚ(�����,�����X�$���n�r)��XuvVP܍23T+�#�%qo944� ��d��n���֦�!""�RG�J����%��NR*ApX�+��[��ڨ+!L:r������橧�bl<�NLf�[K!�ې�و�S)��|���Y��tQ�U'ɰ2x��dfz�*�|35>9����� �#e�
�T#*^��Lʳƃ�D|���`�B��)�B4$P��{|��/���ɝ��� �NZ��`$��ᘖB�*ϳ\s��i���9���\��p���dz�*������������_��_�w�&��ZJ� �b�Ns|��-J�+	�wo���/��/^�{aoo��҈�	e'�Ѭb��=�¸x�O];v�?>��j�/a����H�Y&�0��`�=�.�8&��Z}9���������J�����~���Uw��Pw6;�9��h�]�s<]�z�����ކ���B�5�Q&��;2���$���!XB�(����ɠu�8�C��m1�����z��H�f4��Iw�tB�Y�E8��-�Y홻�T���e�$퇐��d��O)�G������"K�glϑ�iL�����A_F�Ј�l���M>�r�C%�nĄqy"F�I�x/�^W�v�t��EP*�8���c^�ӟ�4���!��n|5ݼ��T�!�_��W�k���'^|�EV�~�ӟ����O�Ŏ)�_����.8O~�3��:���ņ:�6�ƅ��q�7��޵�fOpq>��"���N�i���Z����E�K*ˠ�*E�d�O�̧ޘ��I�����?���q�s�N��sXc�=ƽ��.�.���$���yƒ���uį�g`n�*�H�K5�>ժ]k�aƾdh˂��Ny@x||]�v�I6ϥ��<+�@�!y�l���q���������W�+�u��}DU�>x���F�?�t�C���|�!��K��ꢞ'>\�=��pa�VJ%��˗/ay#����{Zo�w<MONO�O���&��^*����Ç[���ܢ�K���n�@pA���޹۷o˰����O���͛B��I'�܊N��lW̥L�z�?�������3���ϧ�A��7ÞNl�l38ZZ��&����˜ȣG�4��� 8lr�Q������s�돇��ׯw�#��������:��Y�"��hN�9-���;iW�}��A��r�#��荙XO�S��(�"�y$���Rd>�h,��8~�_�M��0#����Yrf�ön�H�hj|"�g��u�<���T�X��_},IH%��V��-!f����g?�Ylh���0����rZ3l,�>O;�O׊2��n/!�74^��d�u�"7@f���H)S	L��e.�Vn���@a�&�h���$�T{���ő�����rU����t4I���,�Q�6Nm&�:N�y����� �$���ED�2��|1����/�I�pi�*�j����B4�jU��ie.L�-E���$�z�K�� b�f?���ۙ�moM>���d����$�*�C���'^
/ȋ4O�L����6^>���~W�nwK��t��4�	��9�B	�p�1E�B���r�v�ڑ��{Ҽ9np�v�����w��P�2��ܧ��a�7�sƵ������eR�+7�'p(B�V�h�Y�O��[�34y�5�C~c��ur?��Z��+S<��?�<US�ͺ��sa���e�?#R�W��#�3�~-�f�خ��Ǝ�Ч�|���"��	���C�pg!��ZCkk{�S5�31�K'Ҭ�k��c�k]�ul5�[�j������	ZJm3���+���x�=噳����PJM^�)��,�����>����L��p�r�/�L"�"��f�?����8�&(q�\�@K�\7J�OO�k-ϔ��R�ZP�<qB���W0:���V��C���#I�L�77��^8�N��`���΋%ϵda��T#}D:O�{y�U�qơ����1~�j�f�V�Y�q`�3�YH�uЛ�8#�[�ZB]�3׺�d\v~:3����+=bk�ꇎ�#VlA��9u�ja��X��Ď�,�:B��F�r�y<�t`��\X��R����+a^�q`]����1;��%����7�VYJ�Ek<�q�5w����Үd���7k�h�L�Bq%U=�>("�b9_p�T���[�����NP�	�$c���z���h�:�s��e��2�gL@�X�p��[��e�_C<r���ʲt�kB��N[�e�{Hx��Ȗ��)&:�k��&5��H�8�cϠ�oz����_"� in����+�?|�:jH�{ꩧ�v6��	2˃�`��h[\��7�DE��RoYX�T2	.LGm0d�7��u+7���l,K#�(�[�Vݬ�۝�;wn�ѡ���O�Pq�����'��0���P{�Rl�8�m4����*��㱀8�'��2?"�Gk�K9q:;����k��_�?��e�,9�R\.pBh�ؑY�6A�Y#O4�e��Jc*ۮ[��"��,�x�"~]�Oy0i�(B��\s6٤Қ���lj��E�a�J��rv�o$��Z�X���~�1���+h�p�'��\u�?�|<�Md��V�m�2lj���Zv,��Lu��GGp����:��g����q�Ǝ�~�7~�������^�z�f�����$1�%�!,���[o���g�w�&��Z���<��z�:���cE���DP3�$���V�!�G.�4=*^�V�A��
?^�ق��+�|a�e���c^����?���b>��ه������	�2����hWq˕h�>�	D����cѺ�j��4o�S�P����I3u4�����n#"�R�
�?��A��r�5�B{!�k<ƺ,f���R�u�)�v�m���:sj��[�ً�G���MN��G4	���6vw���`^��^�����b���w�E.���A��f�$.m�D��L�&}��]}�30M��Әb��Hڋ�Ç���o�=��������~�#��Q&�;��-T�w����?���������?��3���?~�(�TI�1*�b��+s6=��*�2)0T,�h�6p�9��^���4%}�}���H�ܸ���<R]�s9��q�8�n� �ePJ��VP6*�+��؝�M�	�ay�7 �%t9�>���6x���SJ���,3�V����A��|K�F�l&E�^P�c�|��;w>��WC��!c\`����%��y�bQ�z���Y�{㰺���5�_qw�n�34���X��5�}F'�K���嗿�eX�������&�ҥK�r}D�B�(EA]�|�c9r�����~�	�Xp�3�Sk���_�Kfp�Na�Ⱶ����S�.�V
Z�\�C�K�v4��y��!�( �o����/�L�J�Axy|f�n��C3�o�Ǳ0��j�&�en��40U�(�DoB�hR�]p$q�x����l��ϸ�*8�w;WaA�R����I�Y��%
}\2���d��N�؊�H�0��~�*������!`���W��~z��'����]��� &^xMތ�,�W�>�-R�V�9��7	y[̤]����3*X��g>�-�>N|Ī�)�z &�d����>�s��Og�<�+�3?j��^o����O?�H�p���۪ǣ�H�9YrR��%�?h�����1nF)t\U�s$V�e�7��:��Z6	�M�~�0r��[J�(�p�HEk��~Wr��2;�\?�Xq	tb,t�d{��{��K�#g�_W��ZӃ��:�b0��<v[WOu��h�E���Z�*��+��F�X����kUF��Z&�	�V��z�(�}|s�up7^��`�KŴ}�R;�BI��A�95E��v4�áR���� mƭ)qKI�H�z6o�{
7���7�@Zv�B/�U[�C���5��ĝ���i	tZ�;�*H�ӈ�� ׺�Tf���c��0d���aj�KB_a֒1s��3�1S!��$X,������r�5	L�^�
��(J�ĥ����V�|I�f��g����ʒ�7$vH��L��2},'X��Ў2��T�2�G\{x�FA%�ɔ&�ي��0��[W~�?gOYG�P#�����M+�#�2��Veїʝ���,c�5Ǩn� �J��K�r+c���m��;��A���h~��(�eI����&i��*��:�T�-��M�'j��
�y��c�{�i$*XY'6�h�x+,���T'��fI��nV��ċ|!��<W
m�|!ܕAw8�u*ߪ*;A�R�/�u�yMQ[s�_���Rk��Q^�i��ߪI�^���`ф��X̥[��ۺ�iG�υ�k�-Esa�<(D�gI$A@�5�����O&����&H<���ؤ՝�>D����	Y��d�0K��Fnyr�x"����V����gݠi��
�/5I�f"��U,�U�AOyH+�ZS-� �L3�w�~��bz"Ӗ˕�r����K��t��f:a }��oؚ��>88m���2�R&�N&æ*]�k#�Ȳ(�PhX�8ɪ�,�����#��M�B+Q�
螲XV�Z5dC�}!ĭWE������m�:i�����^����ǳ6��索���HF@N����hz�d��_IX���;�;�mU�;et���ر	�E)NB/E��5��Z�6�*c�t]T�иe#��*e��Ph6;P��9��4K����-��T��	L��u҉���I7k��r����_��e�I�̆D�C\87��v��.�|�9n���	��(�<l���t~<K��\���$q+�r�j�c!�<�h]DA�r6`���L��bMW7a���m�@���#����}�+ǽ���[��N�j~:�����#,)�������2��3K���요�4E7�{}�$��*�;#(&��)�-�f}�������̚��xd�qV����^'���7�u�U��d8����:>/�C%D����1Y2u~Qu�K_@"�rV,\I�i�	o���ΡV��G��3�:J��z���âȉ����u5�̫�`�}��-� ؾch��Gb��*�����?y#IE�����͗�B��nڇ+�y1Kj�l
��5���[�s��₈�&���p��5�e��E�p��TZ��X�x|o���C��	�|����Q��W�U�w<ŋ/|R�1¤�sss���(�:�����ݭ!w�tI��ũd5;�u'�n`Q�������ǳo����tY4ӹ$=>>���
�W��2�����O��Z����ŋ��5F�lnAH��R�/粓dX��$��o�'�h���/���/����@�e�T�e� rt
�aW��9L_X��D�����GC����%�L�����]�uP��	Z�w���BFz̐�ֺQB�kx=�Ϛh��l���B%3��"Ch��hW�w�SS�߿U����s�=w���A^$��)�̛E�4E�C���K/}��{oB�B����ϖ��(���a%�I�����D�2N�]6�>x0��>I�	���6I�	�0� �F��E���	e6�1��Ĺ��*YJ���,�>�Y�Y�J�p^5q�U�g���h���|���Zk-7�c��R�<�RjDao2��2�e�s=�מ�����z���[��b�7��.aI;Y�c�qo�c�)�ܛ����Z��2*C8G�x|+r�Rp��T:z������o��A��)�!��|����|�
�@����_�җp�_|��;ϵB�K�БɋA���7�ѣ,�<~�؇��f�ߚk%�P��$���oB�Qf!�| i�@)�%�".���V���'�/�#�!*ҨA#8�Y���{d۶Bf�?��O~��R��������o��G�/�3�}v�d`������(� zN��N?>�c͚ ���%)��D�M{|xP�9ȁ#�adQ�a9p�d`n��@�1�6�k���0|�d�8�ì��Rx_5�ZQ"���N�I5m����T�����T�%^3����Af�H�N�����L��$��A�}�����ɔp���&q��
2�I���_��r(��P�eRm��[o�q�G[��GQ���=�1S'�ĩpqW�-Z���Q+�#�-LU��_0#�y�h?�ۤ:��aT����:ƃ.����-��(�u6�7��ө�t',�&�F��x��Z�W/_˺����JK�x��`8Ks9���B���Nt�vg<4y�7�89<�����A[������Jݺ�Vf`)Bʣ=�_��;�����b��穡�p$���$9 0�aP��������w��駯�����,ʏ��~���d4.��d.�z�Y.��ld {���Q�mI0��K,�\͘4�`����yj�dpa��֐��O�ƕ�d����&U�V!��kҤF2����X��=a0UW��6mA��ِ�-�|��Z�8���Nm��4���������!<v��8%Dt�*�gE�8��\:r g�Z~�!� ��@�ʥKO>q�P̏/��1Z��p�e
�)�N��Y�HR~[Y�
���G��+��ӯß]i��a_�"���:]ꍵ�bR�m��eC. L%�7�v�y.gP20.�w�,����;/T08xG#�eJC�weUҐ5a�Dy'���|���j!���S"�mY)��ƴk�X�#�,�gsF�&��e�؎��NI�7�xk�ёt0��š��3e���{qM��Ӽ\���x6����Uw��m���c"b&	���j��;��Ad�����Xg�!\�+��� �HH(���&R}nn��Hj�Xw�9ZM��3A4��>d��]�����]��8$�ϵ�ɣ�F�Q�^��_��%�*�%+�	s�����?��	�`���M��,���n�.15<����j?��S9��l�-�ܭ�ن>B�	+�V*�2�ic�0
��nX����
n�h^����|���
p=z�x`&�^[yu.7ⰲ-]d��#ؙ���zLXk(��S��(#���A���+�ͷ��譪f���(q=��F�R�[�I�3�����#��[��7���R�^�{��;k�0�
�|��X��&�xX�d+}��Y�ف��i�R3��w�C�b�X���2t�\���qF�d�9uc�=̇�IX�㪊áe��A/)�,-� ����g��S1��]��e���"�3�8r�N>1���#;���
��h㋗��J&��� d��;��(�Mlͮ$�/�����$ cr��5[)�ִ��}N^��Y�H�$���N���#nߘ,�S{���n4��ϥJI;���N:��(Ay�s*<��:�|��xxvUm;�����ݬ���w�H:ڵ�ڑŮ��Q�-ߥ��	W��!bZ�H�<����M �;��6ɐy�,���8c��V��sj�D����h뱒w�� �Bq�'Yi����Q$쇣�zW�Z��0MIo�!����U|a�����=5�-�D�X)�Vu����=P']�Fh~��s� �/t'��cmsP+�ɭ2,u#�| 8�Gx��3@������_�8w��%qI[���m��L	�τ70��Xy����#�c�����9�҄eX�C5>lH�#��M���q,<c �X	q�oX���$�޷Sheet����_ۗ��(X���n'H$tc��v��+*E9MK!,?�5,�)����-e�;wz��#�Cm��������L�n��鼗ͭ1�{W����oOz�;?8<d"���c�Q���ާ��xɏ��	ۈ�����&� �.<|(s9qeQMs�QG|E�V�_2��m�L5���W���[�U�S�FoyB`K���D+����p���U@�v���B"�}���*�(Nʭ[�pK7�}��~���_������_�����҉�|i�W���T�(�$��������)p���9�gl�u��ԥ�9��u�#Ԑ|��<t��|%8�ΏN���QJ�)��==>&�'p,�,Oɹ�G�����>�������޻w��L�2����M���{�^��7H���ő�s�6t�hF���P�yZ��,��E�c�p 5c���X��[х��lk�rb�.juKYMӥ�+���	
-���Q6�'ޏE��q$�d

#� ��|�)�q�u�p���:G��<Om�;�1�ԧ>u�����SF-rҵY31O���2;5�$橊����|�L�8B-�߄  ��IDAT�±=��Vx�7����K/���� ��я~�!׵�J� ��_�".���|�s������_�$T��0���U�X�x"׿�]��`�k����B2����QJ��(�5٪ ������̴k�#���M�:tz�D�ٱ��Yx0��/[�<��?��?޿�z�F�֜�𰛲�������K��X����1�*�H�-��0��+�f�R�ܮ�[G׎������_�g�����/��k]C"'��v�ʕK�.�G�����Bi���nfq�n.�H�X�)?~L��6`� ��Bd8���͋�ǩ�h�loܧ�$f+)c쾪�*gJ^�C������1\
o����S����L��gtH����&�a���m�#hx�f��֢��E.^�XC�28Â\[.h���d!'VF�Lr��t��T͕�B���|�2�U:?p<�K�Io޼ɭǧH�!�WDQQ����������ѩ���&�ʅ���Dr���L��?���A�珪D�.W�v�6��
Z��:�)�W=����@��⵽�@O��������ȇol8И��ͪ�#ڄ;���Z72��J'�$�D�2�b�MU��=s��{\xw��P�xW�y�DqbO�&8�t��;�[�"!Y>�����._�_����By��ֶ*�<�DJ����aa�D���2���J�p�
��7g�3�k^���SW��)�K����3�+}�JQ�2��<���i!)�� �q3*]s�~i0���·�+�{k�~��4|��,V�'��X7:��'?���#��(����Oa�:�=�b����1��*)��Z�n�dҡ���PV��+]S�� g��(�V�U�g�^Fq�G�+E;ֶ�NJbf���ι�& �b`�?�}�� 8���Yr${�l\�V�G��"�Z�{�dB3��HB	1}q'��d&yKQ�Hy�� �Zf��:�%(jw�g,x��A�(�xV[�H�Y�ce2zZ9�_���b'ы�G�O�Y�X�>g��Մ�x��#�ӯV�l��P�fQ[;+�|�ZB���9n�&�;�zY˕�\�7��0���Y��@���q!�.i�܉�_@��s7:��W��8]1��0����c� ?X�i���ļ�S���i;)m��k)@'���,n'e'�p?_��,�9�}���|�TO�a�{���B��̢�`U�72�|p�a�+�s#�.e�zR�`Te��v����|�UQ����/��D�t 3s���D�]�aI�K5i�:�R��7)�n��l&)�0��C����9V��&9�����Z#Ml������^'��X��b����Ƌ|I��҅u��Z������N���9������?��pxxhڲ��w�,�VG�ڧ'��9�	0M�^7�a�I�/f�.��Y.���9M].��ƣ�-�:�8����,4�LG�Ku��o�0Y.fM+�l������Q�g3�@%��q�á 9E vU�Ӧ+�.t��s�͹��z���p�iz�k,��s���/�r��#5��h4h�=Ige�'���.?��UJ黈~k�G�u�8��8�ȄA��)1��U7��U3�ՏO},�(�y��#|��:3_�a�����m,�,��)d՟k�+�=�7���JT�s�q.�k��6r�߆��V�o�`ڂz��k)W���fu��T���#���qo���)F!���4�8����N����g����k]ꘜn��4z@nY��Bֵ#|#Iȷ��z]ږ[d)��a�A��M|�THZ��#��i����Ӫ6�*���T��r^օ����om��V��J	��������`��4sQ�y_�����,�78���_O��2Xf󩺶"�iW\o\U�N��r5g��Q\㡬�`(^����1�'W�mLS�<��]3�϶�:�'N�����[r�@2˙~!h]I��a����׾�+�����-K{{{����lmn��f�+p<����恀���%Ǻ�jm��Bh̸Y=>9��ӂ��z$��T�S�>�S��@�2�6_I>k�SA����wc
�x�rݧQ<�ި�K�0��$M����w;�s�=�?�w����ş��&M�v:⌗��F�O0�BĜ�l���҈��:Ƿ)p�$�a��6�|ˍs�͆тo��i5��u�rخ�M��CfO�����x�S&���bƽ{�vvvv�Y"�C��t�,�)U6䙦'3!���*�7p��2��9b}@=}�&[�% ^��Cg�3k�#�����:�pm���v�X/�V��ʱ�Dn�m�c)U,���.�+9��O�8gO4��;��5��ci�i��l�����|x�Za�f"�W�r��9�N��:4����&zd�R!`�S�n-�FYq��u� R,�:m��*�d=�G`���G^�	~��7����S�B(ˬ/n&�nD�������W����K/���+������:��d5a�M�&:�Lt�8�	S�n��ǈ�.r��WGn&�.{�Cbz�X�$�]�q:|��N��f���!]�m��"׼�&t�9�Ǚ߁s�ǁ�<z� &@[�1��S�K���rܷ:Q�[�1h6p �3]�p��1W�q2����6�n^pkq�r�'\L��ƍ�_�$/��B�+=��'���c*�T>�r�����g_��o~x[�#H�`4f�Nt~�/5��4rJЮ/�?�����{r����WY�]![�W��Z���G��O|��ѰG?䃼�ev;��c�^�P�6�s��^�|ᩧ����`�����tS4�i(O�!��{�h2W�eɗ�]AM�p�L�&��B�N5,��?^ҩY*�Ύ����X���ڎ;���m5"}��{d���&��JQF�;����k׮]É���q4��30SV��FE)��p�U�,$Ds�����x���:�D(���0�.��*I˂���R�&x�]�ve]�9I�]��$�Y%�h��SB6�U�KSUP��۟���j79�kb�P�z��������[�b��ptj���o�ƢY���|���v�ʮ@��ڢ������"&�(��5,���"CN.\��.�Q!<��_�e|�(LC�b{zz,���D�l�V�qӭ�	$�\�uh�bu:mW��i��vM�@�c�`ԛlp6�E��F�$���0�K� v��$�z�y��2��>Uz��	Y�� �2=9=9އp���@	����	ۏ''#��賁���I�Q�ե��a�/կP:Lg��G:���i���ƅ�
1�0����0�������h_����'?��ޛѨ
�	nv�*RM@ p�E�S�-�㺄��»�e\�+A'��NVBd�5����7�������uV��bk�"�^�k���q���ʍ�y3.=Č/C���V�v3@i�|z��<��g 7��p۳����3����W�R[�0#�eخ�Bz�u�5���1d;?I��#�|>���a��g�\��cKZ�B"��|��3(����6Y��S��h2и�IB�-U��>��v��٠"_����M����X��}��Ո��3*�ƕ�[炄��:pR�
[���*G�g�)U5a��qya�(�l����2[!E�����+����b�;�O�y�8�j�ʬ/���h�-ʯ|��-�s=[��۠UaM�O����1#�)���a��8B98�H����13��=� O�C'����:|D�|
<�纞�AZxa;CU{b�{}����'���{w?�@8N:�cU����M�BG�P`<���5�y��V��/�[��sf���.cl���;L:�Z�s�'�M}����<]@|{?�� ��>��'�:X;:G\��ꫯ�ݾ}A����6�{��!-c�����Tb@-?�?V�dPÉ|�r�~:C�Gh@G��!؁Ւ��oƑ%���ܖ�tT��s�$�
C�[%J�ȄH���x^
C��iE�i��v�!�j���׭��YՄVH�Jf��q�cr=�+�F���{C�U�^����T��$��d��;��ټd��YhZ��g��K��hj{����]�AnZ7�ew{��Rr�6���Ja�<�Us*OQ��R��+K]%t<:�d�����n��lt���T��dt�{�zc��:=L70K�U�dϩ�ڄ`c�'V!�Y�,�7���#93���4��H���͠#.*�R.�P�r�g�mEGBW�iC-
�j+��l���#T�W���d��%o��
��$��0QpyӖE�N��NbZ�ʕ+JP�z��[��[c֓�x�(N�mc�DĎ�#�,<�ة����j���y�#D�v}>oCNܶu��gL��Ҿ|�
¡�/2��p|/bihܣ�����L�n���f:�H"7�ps�咋�]�ā���%��yN�W�7LF�q�<B��\��Z1@��8r�P���)`��cf���Q���W��U������?��?�w��[������5T����ٴV+�|�z���AA#���)-ﭩ�����sJ����*������h�=x��߿!tï�� �&�X����f�(��T��ZI�7n`I!��=�u�s����9,�������v��#ܲp�z8�;�#�x�ӯ]���������ZҠ�n�f�0�V�ӭu}�X��ǌm��#��y�RB���{k��-'����o��5�^����1�s�W�Y�DXp�b:�&7x4��ݽ{j����;�.!W�������OY��mn��.��@<����>��da���|�
����z
A,��޽{LX�,̄����7�����W�^����|���fj�kH�j��-q������/_�v������x�Za��8ebǛ*p�X��k���CN+�	s|ML����v��n]b?����3���Wk/4�].�>�1u>�7~��5��ﾻZ-��������Q���+�Ӫ'�Jf�
0ib�Jч������>?�9e�������k)k��8>>�}���?�ŷ��$�R

�_��_�����������v.H�p���^��C<�Q����
Q��;R��$ �����7߄,���;X�؍Q�+��>	�C��?�k�[㦓���BDU����3~��"���M&w01un;�"�I��ĭݘ�+n߻K�9�1�Վ�Zn�C`K,�b�l����I�FQ����c�S�f�k�2�#W�;�g���YN�L����б���G��O<A	��str�3�%��Z�rũ�QC8��z|��9�O�fl����xc�N��'���P�s�u���s%�lt����j�vbzSB�ӓ�`���������c7�t��ı"U��1����fT#^��I(ne���(o��]2�Ʉ����8ĕ��yk[~l�M��d��a�"mGm%��c�c�0��GP�Ĭ��d�Z["�'/.����"6��YP�n!��yKA�K�atL!��A��4>��X�,�#|���dwMR�|+��Rv�DppvH����r#���NO`�?������z�t���C;�Z� A�Wo�]�z���6G��W���Ҡ
L�*�;�|8�v��饃���Sv!\���n�`��0.�<�,Nt6�Q(���E*8ݫ�㶨���1(�R�[�u�Z���-Ȍʄ��:�j%qV�.<z��O�d��tk5�5��p�i��3���l��Nc2IW+���Ot�wk8����mG
�+eU���T���Hd�+���W߸©7�>���<��5{�&օ�E��/�\�m^ԡ�)gԌ����j���X�f+dAjM�'�R������CIz�1BTHE�GL���ꅪ�Q��Ymh��o��D�-^w|C?Q�Q	��\��6��kӄ&��t��7'�1�5,!5#�,�B�4'��E2��q����K�z�lf�'_!�@���?��u�vۘF�^m���J��j�(*K��P|��4c� sO�PQ���L?�®Ø�y꩖v�3��a;+�9�����%��qC�`��bRo���`�O�'�[=m�<Q$pM�eh�0�����^:�5Q �b�X*icV7e�noo��f�9>�����Dٯ!�:X9p"�~@�Ʀ�^��bV�Ű?�ҭ8����&�0(�,��o��L��V�Q��l�`�X(���N��g246������0M4n��tEԣ^����8_q��.�0������;��8�ʒ�o-�A��f�4�d@ރ�NjF�~d�
 �2<$�d��c�����9{�ɮ�\p�1�3k$�,ř�yeI�dе2���0��qm����~h��r�a@��mH6=¾�$��dQ�Xb�5W��1��׷��v�R?�U$"+3��9{���o}k�T�Tcr��P[�1]<�p��u�lƧ�G����J�K�XfMg��۰|��4��ߣ�J�M❜�y��9Xy�+��F�br���9d�E���K���D�:q92�K��0�y�#J
?�T�=��߸�-#�|��0KϦ�.�U�h��>iF5��pvz�;�)�Z�jj9J���b>�S���ؾ�o0��r�'�A��C�0��W�hGCZ�C�l�z�8qnV�3��*�%����lD�|����6P%j�ٜj
I��i]�i��p�����2�FC�� �.�p Y��hsC�B����-ۀ��|�*.FY,t��:�`�rt�6_>����m� ��t�6Ό#��?N����0�gsս%|���s6�\G��>r���_����Ϊ(S�9��H���Dw� d[Vf>�;��t �Oɲ�b����8כ�K���Z����tF�&�P��+?;99c0�z;�f�Ҥ-',Kp�,���5�"'Vf�N��DJ���Ҝ�3N��a6'��[��X΅\\nR����~���=&w{��m	-�:"�{{�^��Í:�khH���[�������7��/J~ӿ�S^xJ�����T#1��H��P�0��u@-3>9e\��a2ey��c8��Ý;���_~���{��������;��:c	��y`sj�e�U�%Otm�J�UA�sp!]���ǧ���Rd�Jgu��5��Q{T��Z=71���ʫ˼p��铏�	�'��9=IM���,�T+,�;w�v��g�{�=�۷��������2�n�,�T��omS��3�e:5dj����J����Ԙ�X|"ⲱ����ҵ f>��Fs�֫E�K��j�F��:ij����TmnZ�>C����AHl%Ɛ#����[�iDs���:����;�o	&�\�v��]��k׮m�`��rm_@�7e���G�M$`�\�����lv�3�<}�W^yeK�(<8��f���o�E>��O�j`�z��y�Y+.�<��*H�����}����?���q �l��o���<Ζ�K�u=�n	Z�n����o����h/�h��,�1�&_*z���$F���'��ћ�Ɉ���� ]1(N��qLd��:�_�z�3���Л�/vo{G|��ᨲa͸�zU����~����Y�a�<��߈0�H�h�[T&D��$�9j5D"������XS8OX�Ń}u�#?x�Ë/����HLL�1W��U�:d�8� N2���Ľ�v�P5����w��޺g�Ӵ&�Sq�q`u�@�iJj��F�����Vn1�򟭭Mg,J_E�m��1�2	�$�hm���.F��:Et|tR�EY����G�n�BDo<{��_�~��������鱈��?|��j��q*	���W�J�!�YB9�cU*e��Nd��Y~��Oa>��G���p{�Dm�����?���4r��<�W��u�	����(�$��������BՐ�-SE�^xݩ�����d�r�*"����r~	`�1��u��(s��D�g�h�MIs���fB���E?>|89���U��4��͐��C�o@ц������S?]$<j�"`+��xв��:�����kUe��+_ð��� �f����E>/]<Дw���N�69�������!�7(����;wh�� �h�{;"�r'����=���>a�V]���}�>�B�%�q/������/�N7��R_��m�x>�e�Գ������h#�0�^>�r̓�=���?sx��"��ţAM�T%oIU�i��*�s��l�&&��RnO�|A�}��;��_�O���}��$�:Cw6u@�%%H��y��@���H�z�9#.J�b탌T�D�/]����q����������KV,��UT��d�_(Γ��Y
͚�W���$`����O9K�� H��"տ�d�@�A/RK�4� 1d,�e�D&Gc�|!�^ӂ�9��NQY���x��w���q8T�>H��Ⱦg޵�G�VQѵJ�<6��y����'+���A��g�"GΖscm��'��w�۟r"˂�Ɣ��O*�Z'r4��3_���B�i�Kj{t�z�V}8�B�f�N<¢4���:���E�� 6,o�*��,�l0l�Q�6���?�M�~l�j��U#���X��O|����}['r��d�*0�Eq���',�Vm�������!��1R���`1[��y�c�Դ^�{�Q���u�3.G��2�aB0�99npu2iH'��w�a��Y��YW�>qd�����4��k��z�M[~m!��5`��Jb�`s���)��ޤ8�j��T����-I���C�ԣ�J��Nd9��0��]L��З3|����1D�1W���&�c+ِ����6�Y�,�ܸ�q�A+�ؠǏ�29F���q�����¦5���˗ex|�ߟ�'�qr|RՖM�`�������t�QS�WC9Ŝ������I����'ye�g��nx�<8�R�U�Gn!��}�70���1Q�u<1�"�"��E͎$�bg+a�)0I	g�σ�j��1sYlC-�i�#��b��s�A7jAZ�CG�|My�4@��im�[FI�!\B�8�R���\��`�,�Z�?��9���,�w~QQi��zg	�k�Iq�0I*S}
��,��7١�A�`Y6�!r(`(��8p�9N��PN�c��`c���a��`�(x�;�lT��P*�T�S�*��/kb�4AOmP�)�z��,��js�I���i޼й���р�l:�E&�%�_�y�����M����iO��v�\MqT�X��C�i8]�!����E�;\m�%��{�ԋȠ�I�W�5-�쵄d�|�� �{
=s6�޻w��6�&F�QB��&f܅����7�@.�g�[�n3��J�{p�O��%��<������K�3��p�J����\�f�:r�Tk������ҥX.T�kyhz%�� =�reӐaP↉<�k�Ğ�QH�y||���������s�������~�?����������!����u�՟;��ض/�]p̋hϠ���E�� f��|.�F�<�!�"xV�a�青Ք��h��f V��E�LX�Bք}jtW�7b��߹/��(�Ǐ��ݾ}{{���c���G𹋕�V�^Ι��Ҝwq��cΎ��ړ�a�<�%x��Qd�QVn<�!ދ�]�&�4~���p��92n歹V�r�y����,�8\������ͻ��xj6|�C*�9�)�+�v�b=�s0o<>>���"'��_�����X�20�SO=��k��1P��bhdk��FOL~���~W���O��ŋ�}
�[�"�(�? ����GGG_����Լ�������U~��7��P����g���i�S#�������߉[0��xg��K����J���R[�#�*>G���s�������"���<899��*�p���m���wd�%����w��ݞ�#ȡ~W�F��Q����,$`�v�lBX����@l=d�8g�U~]0R�A.���Sy|ٔ���{��J���+�7|�{��q'�9��2��`#��!��E�:��N�(0>����S�R�^���v6>�q��`����N��e�8g��R�>g�K&! -����wi��uJ�
.B��]}��{���ty�	3>z"!��V�&Ì�\�T7O	�Dm[3�}M�̵�$�U.~�Q>;�i�����&J��n��'�~�:9[��!��>CT#��Mu�t@>���:Q�0|���f��UI�2P� 2L d&&T���χҲ��5 �h�
yc�-���� ��Ǉ���O� _������h�	;�I��Q�q�hv�4�����Ġ��8
���P��� U:e�^tf�7���+���J>T�D��i��ك,8\�z�<pUT"p�`(��U����V�:b�Q��kW(�1i��v��~(QL�RK`׺ޣ���|�h�Ʋ����� ��V"������B�f�S��������G���S���1k�w�����rZf��!Uby*����"���[M�˷|���+�G;�^:h���+h��U�X�DN��yR@�WW�\8FF�� e#�"�?���G�M�2q;=�2q頗�Tqfy3�Xm�4/CځMc�b�!{�%~�|a4HٶU(�B����@�*/3N=z�!��u�=��,����J�⑇Z��G@�&���b�UV����f�]���)gU�4�M��N�xgi(�%ON��D�C�CYk�o�񖦎�)[�(!���t��/nP���B+E8PG;!�[�Ղlhȃ�t��w�?�/�E��T��]�V��w��;m$gO�y���	2�{I����le�����\��hM�V�zA�D}d)������9(���x�J!]��o���z�}��1�y� n��jX�����z�e��ȠnPI��B�F�#�&���2�R)0�4���S!2�'����O���`Bp1_����tm	&6`Rm�}�=ec4AB\����D!��ȭ+�g�Xf�"3{����ZNA`�ל@��� �2����Js�Nh��RIFu����2� ���c�����O�+��f&�����ʻ2�9f��U����|yg��H�?k��"�c��q���� �ZQ1�=k'.Z<�`&.P Q�I�l�wD�zynȤ�������H$7��k8���D���+˫��$0>::���dQ���l9�Vkmؤp�7�0��z��е}6��iv��fu�#��L@�j�+�n�X<(�<|����x�
j� �dec�=��'���K�F�xw;�����`|�A��5W������v��Y�K<��i���7F[�7k�tL3����y�)�M�?�P��
������y�D���I~�����xr�f�[�\�$#7{f���i@> �aW�+� 9er����x��!�����%�౱ueY��_�9����*{�2����(�A�ѐ���X'f�E��0��{X���r�D��F�B���Z��$&�17�rS�k�ޘ��S��%�B6��̺`&]n���˲/��zr���9{E�� �! H"p#x��	ǁR�0�X錹
ib9�&��Nn���T�f�:R}˓%��;E��v�%R9�K*~�x<Y�ĳ�/�E�X��+��S��
/����)����E.�0'rCڣ���k?.��y��ӥ����t��}�N�)�K��3uں3�w�KP�e|��d��1�vM��,�ݻw77�x�dݞ�re0�W����p3N;Q�9�M-F$�{�&VN�N@�X"	(�r0/pX�	�u(P�5�5	+#�;�c�,��UE�����rm>�9�I�2�(��P�d8\�z2i8�Lo޼�g�g��{���O}��_��/��7��?�S���ݝR��ߒ���t�E�����oZ%��*���I�x�(�{��Ő!�{(��4"�PEz������g%��T�|ߜ������J��HNP\���(J��t�jA4�[VW.]% 1�,�f�4���
6�ƈ�����6OR9K���x�pEi�!�ak�1�)dW���!8Nay�ѼPg�&<:s5+#��W�����zy��$6�O-6���f֥��beIf���ĚԜv�p >�~���O>�d��/\��s?��r�n?x����6!W(>X�K�tD����f�E+���K׮]�o�C*�"G.��H�'��śZ{��������<��$Lx���&����tN�0��R�v>_ݻw�O��O����7ސ�Y���?��ʜ�;��0$�]%@C�N�&����h��D�vۛ�P�l���0��
9�y�.^�zuct~���$�Wa�' �~29�w�����u�iz�[eUh�e3�Oyl�oS?�TM�/0$ڑP{�O@?��0�N�X�QX}��ɡoB�tCư�S���"i��N�f��
e�+N��^;k������(aR����
Q��O��+���{>[���?���y-�Rs�����".fE)���:q�
������>����� ��_��K�t�r_,n�1|"p��l>���J���c�W��/���l����a8X
����?��E�y ?P��v��y�ߏ��|���8Ϻ��,W����|�B�7�Q�)�l�{� p��ӓ��t*������[��\AN���c��H�0L��G�ų�A� '��ۣ������	3G(��<��<���N�;xk ���l\�����`+߯*_1Q�R�CG���,��K�,�{r:�S� mZ�jNc�/��h�+��,��?�#	�Qm�W�*Ñ�\{k�
����,�Z�����EV k_V±$v��U����h(�0����`k�/4���k/� �������+�,/>V�I���k|1#\�J�xH����L;�֋� �l�F��x��e�s�>;R�O%e3�h6 ����[�?�/Z��ɣn'(�X���,	�Y�ԫ����?���8x�uI�N����x�5:�	���j_��i��$,1��(���/�m�Y(��[�׌W�G��֏�P�}��}�;���U�ꈱ�ur
��n_b�u�����$T�Yd�o<���[��^}�%��VȀKx��t?N����TC������:�92+=�^.�	�s��p�պ�t�<Ni�BI��]��O��3���Nh`�t��E�E�R�q�ӂ%����\XO�����uk'd�j�Q2B^)���`b�QT�M�=�M�
>hlЉ`��Yi��<�Wd���
�� m�n�W���ظ�Zch5?.t���pV}���2Ǐ��#[�SDlͤvE�D_�;�ZJ�����HoUL��-aC�)� ��Ag8����oK봲�}b�Jb��G�T�+5 a0��Z�����4|�#g�M^C]�B��|j�ηr�Z�����S��g�gxUd1�}Qa0w�E����sa�!�?<<��e��V��5�/�a\\1�{W���ǄP	�<wUm���l�R�SH677T	z牰��x^��7�<�}䋖im$��M�
iG���,�fX��<qQ�;�
��Q�n�p���BN��$��Nj��_\�z����6K�z��<Jg	/�hn�s��zF�����Y�'?awZ��C����&̃��p�"��vv�
ce^��	w���uD�����L�s|���_�җĪݿ��+jN�i�PP!�����ȭ>|b2���{O��O^�%�&;ӱ�솋�H��'�ʺ�3M�=��ܣ�h��G$�!R�H�H[��>�u[����S啨��|8�&$�2�x�@kV�x��7�e=y���T��L��{�=�K�6eF�O�J+���УG���PSv�B�D�Բ��B��0g�Jfi�]]}��_���1J,�˹MK�Mҕ�`剓6D&�E�����SO=��1
1*S��>0�0��2 ����ػx�1hq��e;�	I&���c��c�%V��)%I��Ԡ���zX1W�Q䗋�Վ{`+��W�~��/_�R=lԐ9FP�T�p�����W���[y<>#˞�?�;8]L�]m0������|����VWr���Mv\"�����cV�` -Q)���~��i�G�+��b}����?�T4b̺�5�-��A�pUwu�)i��G�Y�	ŝL��Р֫%��읨�۷o��>�+�N�?���yx1av:R:f.bEC�KZ�ǪT�$,��1���ȍ�^��ecW{���Fl���ԩ�	�N��'{�aU^�-1s7o���׿�ۿ��/������{|���`
�d��7��&A�le�sj���f��2G�k�C҅���4�a����F�\��q���b�9���-���	N,�o��\K��N�jX:����ɍR'r5�N�]Z?V���lG��8ȹ��b�\� �q�;�z25���5�gB�\�T��.��\
�!\�����f+���X��
�Էލ����[G7�ɚ���*f�/�n��kJYg@r:ޞ,ſ�˿������?���_���� k��I�1�C��X��\�)9>�ZN	��}�-�v��Z��ݻ��ǀY��Ν;��7n�l����"B�Y�qF�(���uYa�{��������D�M�^<|�PL<<��|�p;�g�	� �۵������H�>�T��+*�k���>�t���>���K�.]�r�c�嗢�x.\�&���G���)j���huy���6qj�����X�BD�C���-�%���D�eoo_�����.9p��Nb�����ݬ�s,pf�]�ىO�l�|#ӋQVF�!K�6Sܐ�)ҝ���x�^��[����<�l"O^�c�����V�,%�&�#+�:ʥZ�����b�\,��LN���5'�'�Vd���2m�O	���%Shrmy%��`7�:�#@%��E�*�-��	ʙ����?8��d��q��&�(?>�@'D.�a���G����>�Z}^���Yr����>�ty@MÞ�_�$�I��<������Lͩ��0�B�]���R��9���v`��%@((��z��Ҕ���u���*�bh;��R�t���OT���D~��/�o6B'������1d�kM'�-��[Ѻl�A?�wD�^���?�3��l�p�2f-ji�֕�{�ׅۣ(ʢ�ʋ�-:6��SqZ件wP�M(N���v�V�$�3^A�>Ѯt����9�S�:]���ސђa#M-�jr�jt�
'=O;��^n�6D�d��~�mQJ�n�R�/)y%�RԢJD�X�Z專,�7��kk5��D��A5����Ü�R�0�!�|#(�%��=-��#��FsD%�o*"�\w�A�ķ��v0�dۃ=�����ml�s�3M-!҈���F]ߖo|���Tm��i�~t2֞]x����������]�x�YR�&��G��|���4�2>K���a�Dq�T*~lJp��0�)=yj��%�Xt�;�����0�"	�^Ӫ"֭&��;R�����9 ��r� %D_^^}~�_��MMT<� �	~E�P������ı��46�25�[ƱO�ŋW�F�|U��K��f��D6��'����U�z���y/�ї�[8�r�6�O�6"�P�����f��	b�����m{��j�T���"��vC�8�B4�l������6�w��Ԕ�I����l4ȩ���B�Z��Y��@c��Ӌ	bb�P��;(�K�0S�t�c��
aͧh��I_�������a&�W$�{4�բA|ҙ����e�LK2��\1�n��	��	�ۊ�,�:���(O�fY�E�i�y!n��-z#�F���2��n�b�G�ٺX�3%i����R��n�R�o�Ƭ�z"�G�N��(��:�`����sL��w������B�J�k�����S����Gc�jcow����5�*��꼮�-�i�SM��H$:V��!B꜈ٷ8�v����TfUVb���"8��#�V��ސc�W���p�67�W����
2ؠ OǓ�ӱh����ٲ�]7�[	�y<�IS�*�z����V`V[��Z�s���MB�Ҧ�uw��ѱ0�a�1I��UD��x��O>��ѭ;
�_qJib]�T��������ehd~ ��O?��SW0)u�����E�Q�.Isy��d*W�u�+/ȝbc#���S����v�K�04�Q.�?��x��#�ݝ��K\[d�.
E+ �*�t<w�9*�a��P�P������r�cXd�*Rݧ���̟z��g�lR����l6] m�Hmd��H$y�����c��C�Yd{��t��α�o�M�~���`h�����:=�T�$�Wu�>��h�Ҵ�����T7����qX[3Z,�ny��Xd�3&��h/�[�U����X̟�������,$n\�`���ܿ����=ŉ�5�ڿ9W�6�l�f�e6��m����H�ɳ����6�퍉���R3�]��ƙf�$�b2�<����E�ó&O4� ��[h�{�6$ڠ7��{1�R'&����Pta2B����1[��Б��
YI�v�,�9���<]b���.������¤Gb�M�ʘ�`�%+&���e>[��^�.�4+�EEH��2r�9� 0j����l99��g˦�d%k��8� ���>���/����]�y�w�~[λ\��p��!	�F:���>xk��Y�	��y��l�4�i,Om�\��;�X��Fe�>֢B�Ay`�6����
��i�6>G:���*�;D�X��&��,5������'�ܜ��������\�G�mq��<n֑�e�&��+��3Of�Q�O&F��=��sZ�]� ��ey�n��\�?����Xj#v�F6�,j��s��m�a=������ZD䁇�� FJg)�<�bi�/r/�ۛM�9>>�z�*r%F�u�z����gy��n<���}�მ7o⃱C7��T��;���$�'�|";+�Y�-���y���D������h���߹{�����|��_}饗D��_��L)�u#�*����\1�N���?�ӯ|�+�?��|��.`d��6����/N��cE�d��r�)$�����E-���$����W�\a"��T��r�<���L�������7�KAT=?�[(���) �K��z�)1���w���	e5���ZA�E!���_����죏>�p]���?)��:�ر��$D.���HO����C&���r�
�˩�i ��DN�+ܼh�LrP}B�	l�Q���`��r:��	P�M�!F�s������7kz�6q!{!zOd�?����ʱ����h�\�s�xs}h�泅h�ޠ_�$\��T��������Ǒ����`0bbʭ;�v�1X�$h��� �#ۃ�!��$IT��O�rZK��=: �1���S��xҲ"���^����ZS�Q�ܺ���	��U�&z���3��.W����j�2Bڢ�&���4pM���/�Tx�
q�/��=Vrsy����}_�y�����b�:
�?{�q��<%�Fʙ3U²앙�o�r-W�]@�$؋�`��fDDF��1�ta�vM���x��p��-�q�ΪG���oS%�A�WceN��;$�Kce��lP�n!�ėǚ���L��&w���oiZp�9�증͡�/qUT���x�2�1G�+i���$��&��},V`F�b�A��l��a�)F ��ȳvsR�%��;�v�T��C-���AO$_vjpao�`w���-�Yo���rRT8�
�������
�j.Z���jy�3#^Uj=+�����{6�l9��'��.-����ƫg|�y֍�p](]��(�拲p�Z��w6/�4�z��Ǔ��������&ej�K1�pf�:p�K�K���¥�����7d_�C�����So �$'�{o���\5UQ����/�e�\\��SD���/K���e�.:�85��'��Ou�v����2A�p�ʷ�#�#`,�A�����*`!��ƚQbn���2�_ܚ�v�Y��3��;��	Y9��J���%���mfߝs!�����S6"4�V�-hX�uZ�k�ߡ��&ޮo�N��6�-v@�}�(ܞ#C1�Y)��V|6�k�ZgeQ��S��5Ңv�y��ޗĨ ��);��.��dxq��d(�W�v����)R�[m5geހ
$�Mp7Î7-�u&���m��u&|�n呭^q��LI����u�d���%O���3,	��P����?���"�DLfy���W6�?��X�|�3�����;��/ZGx3O�CΦo_5�^�	7N��qƱ.B�q���y��wYt��%�	u�E�
��cJ"�k֊v1�c��GK[�q>*��%q���£�VZ,-Zz&��wK�h�8i�.d�[��*+WM:�mu�X�!'�7Bk8���EM�sԻu�����c�Z`�SWe�S�X��V�vx�[Z�V�l+�
�N�m��.+�������3ݒ���Z⥶6�؇��X��Mv����m+�W��+"�J�0fO�>1�!Έ�)x�#��Z��h���ݤ���p�|2��i�Ь�Y���2x���*	Q��!�m��'U>�Pz�}�!f#*�3��F��m,9b��, �	��)&j/!k�kd�77��I?~x/x��`Gj=u-\&�/��K�.2p�
(��X w�JI�["d��#�_�������:@w�ޕ�����ӄ��i~>^ �mb���q�FZ��ћ��,�Ç�e�N'�}Y Rk��Tb�Ţ�x[&/�**���PM�R�f�#b�Ȟ�W-<�RI�(�L�"M�u �|��X�SS�����l�����f��볐h`�,��4���Mh�
ejCdhsBt��X�v��nC����#����yx�gB�����Z9O�p��tY�ݽ�&҆��׬�ҡ�Ȉ?�2=��snǕ�'�Hz$���A���������s��[l�@�\9D���=�ˉ�ۀyY,���I��/���>��o��o~�[ߒ8m���I�%�9R������QR�u[ \��}H)&��Oqm���x�Bf0��Q?G�9�6V{磯P��5�L4P�G����3��|�S����o��bŲs�̳WD���.`���׭S��X=��gU�H�oHm.apuh�w0�e���4qy�J�+s��6�.nQ��X��]p�f��ƋtOb��j�W���Wjx�/Ձ3�Y-	��+RG���ߡ��'ҡ
m���7~�WU������Q�ѫ�c��=�<�N���:Bd��D��Ν;,��p���=S�E�嗯����+Wb�w��o�uDF��˳�~~��7�P��shÏ�c9>㳉j�<0���l)�<��]��Dy
�P cꩵ�m��D��oܸ!q���.��s����;��T� ���/f�{���(��
!���^�z�NE��'_Ĭ+��Bd@`J�|��='j����֭[�����~�m�Y(VJ�:S"����Z������_dp�xR���r�b̲*H���3TJ�Xr������I��x�Ti��������6�R��G���}��&jO��1H���ud�ev��s+�&��n�������`�V���2�:�h�t�!ucm��?��I+�w� �b�-$�[�K�ä	k�茾x�2Y�K��$C:l�Rd��D�����C��!�Ζ+�w�}�ڵk�.fѐe�Q	32��Q��]`�¶�<�U�j��I�q�{����^�|��HtHaz���͛7_{��b���y̕���GI�/U�՟�s���8��~��&ͼy�FA��X�\b"���1S�g�ibc���!�87D٫b��8�?N�4�qHP�C�Y��=��k��g)Ʃ�h�#�":��P5��S������!��`xe�wĞ�Z7��H_N�N�.���ѵf��P����8+I����$0��$D}�"�W�^����ӌ�H���^��	K���8�)q���V��l��ka-��p6��T���z��|�%��[�5���Ԫ��y�[9��YJ@�(��Z�N'�Vz|xR[ӺЧ7 WU1_n��5`�r�m٬��.<�+��_.EϤQ,{z6��p,J�`��W+4)1�O�ہi�l��l\F��.�tt&����l�.Ĵ�M�Hl܇3>���#˩���>$�h>c�e�"�
��~ε��|!�q;���Y�1�|c���C�w�GC/n0qA_�3��,_�>�$&:Y|yźg�x���˟}���f<����J�=9�Y~��C�+ 7#�o�91j���5�#��I�r�{e��|F� *ۑ&��7���6O�w0׳6����nA�|:�T��G� PW�V��l�
�!�e�������.~f|`��QX�
�v�lN��	������Ԩ�����&\�*0M ;&�
�#�64uRg����ٍ�K��m�M�Xy/ĩC�
-$*O"�H��s3t���� b�S~Oǩ�8;����B���-��)�,Yi�X�	�5X�H�G1�	SqΏ�S��T��1r���kR�+�5������aYi�1]f� �;�ke�+��$|\�Sn^�ρ�*ֿ�W�%!*�}��0�`b�Ml��ӺZ7���/2#P3��k��$�0�^�J̎SBz4q� �;�hS�����'L㷏�g "��/�]n�gk�67���~I�%ق�1����@7rt�e�}e�3�y�\�OeO�Dl��4r^|��g�Q�h��-н����$��ب��A5�ȭ�g��}��C[e�@$*�L�����e�ȴ頲!n1ƴ7��XF�=p�WD�g�V;@P�t��YX���L�7����~:'M�T@^�����ƘDL�x��b%7��İ'럝,�������t��ƭ���ϓ I1 t[)5�:�b>G���T�7=�/6�H!��~�D�SP��]�#-G!��;O=<���W��S��i!~���ú���8;�΢%|]L�(�Ӛ�y�3r��"	{�k0Eq�.����"�?%���7����ZtN�g���`��L�RWe�#�"q�y.-K����:�'� ��I�ɣ�
����}����C�,DE�y���t4�����h�%[yx8�i��q�ɾ
��ʃA�</�Y���J���t?꺵�.1�+�N�p��mg�&��m0SL�'+��$И��3���GÁ*󄖽������Y\�u��7�ʢ�7?��ܽ|�r�&ݮ-�����Vg�g��ѓ��ev��>΄p5yi��)���J��F2u�. |@�H[�U]	+
��E�N�N�z�Z�k�?�:�;x���o�������\�p�_��_��_���{HC�A���KT�:]��PL
~��n��]sV1�9-�L�q�E,^-$���2;Rl�����r��;XY	�6�H��ǯPLn_�~	��=��S"c��^߽{7�K=��u��]���ݪ�5;=|�)�5Xh��T�Q��O��!���](+����B�$�f_�ݪ��ny����?n���4��1�S��C���$c� U��($N�����Ȋd��b��sp�#�)�uU��on�C��,U>ne�C�(���������?/��v0V�ZR����P���w<��@�rZ*��/���&����A����{{{����n޼����=�D���{�'�����~��^z饗_~��DΏn�Z�d�Kn�'X$�Z��yG*�^B;�������>��/�p�F<?�G}�6�"�4��8)�x�W*=ъ�������j�y�8�b6����b�Cyc��ODA�{;���aϓ�� 汔T>�V�(���x���2F��?:�Eق �6~�����XL�D�Pf�RHwbA��g�U�J�1|�X�Ş'BW�����E��l���u'��c>��~��<��6;���b�|K��mmmTE��ѥH\��Q'���OM��Y2�"�&Ow��UM�Գ�\�80(Cd6�]�b8�Q��qmIT���%~�����B��d�q�s��c��c��X{�����nmn����uɂ%� Hu�g�JQ]�&9����<��]�~��5�'#�){+{z��=ؑG�E{��gC*<R:9�j��7y�F��i�D5�zdFb�j�*��O�#r��U��t*��'?�	0���1Vmmm�G�޿���<�h�����H�����O��ʕ+(��}�IE�o�[<�L9ap�<N�r�RM�C��r[w]c����F2�9�؈(B���jP@|���X� ��9�����Ʈf[�<ݠ�i�bcП���z�>�*K����x�$��˙��X��nҠ0VLgh{W\K�oΚ*9��i�y� ���m����Q���0y�D��;�g�\��)M�YIƹHtR�x�2y/�F�������r0�>�hy�����-��KL`�w��8K�#/ƧǪ�q�Y,
�仪4(���i�K4�¢i�Q�XWDF�f�ھ��\@{E��?}KJS�S�4T)��;�E�q�8�bǳA�m���M]�b���u�����dskz6�m�했s�b��%�<�,���f���$N�ǆ�UTgF#��l��Oh�^�޵�r�ŕ�\��b��#�:�c��`"3�����D�I Ð��\�!����q�Z�"x��%�r�I���K�U�\����lLF��m�RY:�1�X�07�m�Qg�Rb��V�|�'�y3|�p�+k����� ��m��������]cGv_}�7&磍c��5�1�v���CNt��<G�L�dz�h٪�l�m�_x@;uqim��D-���;u��������=��0�ZYݐp̌����+�ٜ�P��[h�KC���Ћ�b黓k�.��:�i��O�EBw�)#���j����]C߈W��P�Q����� F�,Fz�Y����_\W=}k��IX������(�CSr:U���&sU��q�9)��tR�S�}�,5(na���rf]K�p~��F�fM�4��jOu��&���X���kZ�Rjr'g'�uRÄ�ZdH��`��3�7����0��w�����C�
���JѴu�9#vU�h��� �*�ܪ��H}9<��֦�(�#U\�h���9Vۊ���w�B<���ym
7��AO�a�$v��y}�sMT(Sx��!.T�'qa�hT�[Z<a�
sw�{�!�Xy�)�x�|?Y3|EK�P��S�VwI∡���9+�z����(����*(�X�UZj���3j5�LQ���Z�X�O�HB����gby-G���f�FF�����uc�֠]���~ꩧ._���lJ��엍���F�T�x���C�:���`C�sb�|̬Zs��<�d2��q�]o�elDQr� �{��Z�P�X��������&�'BՎ�e�Ii� �9&�86S��=�
5��b
�����~�
�r���D��0��ȳ\���Ox�ڧ��a@�� V\W5!�	����o�٪��JY���C�.��|���w��=��)6��:�r�3�+E��FO@'���h0���{T�r�yo\Xy�J�P~�=p�}��'�����Kb%X�C'K���%��(E_��d
�S�s,G-��;4��ȑ�)��������Q���~U�S��$c&�ǜ�eY�'k %[�w�w_��/_�,����#ĺSq"BlS�|����� 3!V�W 9X��^ۄl'xkΰl!���}��m�u>����`�i���5�)�X_����^��=�����oߖ�8Rh�G����4z5� ^M�u��j�T�\����\����cH��E#a>;����hZ��7�d����8�-F�`|C�I�'{�Qj��t-�Ѻ���er�7�4V�Ӏ��$+j5�UF�+r�ƍA�����7�h��!������1�/�@� ��	&�p(��JT >`��y�|:g�^ޞ<Λo��[��[��O����y[�+8�8*���zK���+����K8�Y����5y܂ pm�V
X�Ä)�>�űȘ\P�ub�^����X�
��U�kj����5n�s���D���'+C�Q(�Lv�D)l�GL'��+N�}������������|p||�7�7~�!�c��B�Vl�M�"6p	�:D�q�p�����%r��ߋ~(�}��$�L���1<��T�_�ОB{���R8�bya�����
 K!��0T5gH��kF4�g��P�.�E�Ϛ�3���u��(���B�k��M!���x��C?��6���NϏ���e ~��壬ȁ(EN�ӳ���l�\v���m�o�X=}��p(���pZ:���Ç@$)ۦ< ����������q �q�(xr����T��(	)�
�]��ZdW~����������ln��r��M$�w��=#Ct��	{�{�=Y�_��_����y�
`����Y�xm�g_樐�v���Ӫ5U)�v���H��h�0�����@���Ã��,�2d�/�?8�0�o.LVb��^\�F�o.u����Cx�#5ث1�s*fCl�qW;�PHu�/�h���fsVFCLg��g��*�`[�Q���e�uS<�xyf���o���7�x�_��2�vB��r��xU]%5j%C�,h��g�����Z;�r|'̴8+����=X���&g�7��VW8A/�A)�J�%��׮]�����[�qx*������r��(u�^Y���>B��v��#Q&���&���frx�]a����x��{�1H�c�F�$����jN�%%�i#�q���&���X�"�j����*�Yv�'���7:�����qd,McF��i�A��,$�W7�yM)dRJ�uf:!Sr[�:��Hl�j�(9�۱���X��k��<���i����\���9�V!������)�͓07J��X̋��p�.G�6���h�����e!B-�2l%�k���fth�f�"3�R���?�o,��Cc4��w��O��t5��ٜw�ƍ`��ׇ�RG��7-��}�U������7�'g�bYD6� �R	�u	
=1(+�TS�~�E�XE��2ȒVe�`/Dc�/{'�Z��䚢�<a���\��[���H8'�_.�#�4�%F�"%�b��X���85��jKuw�T�����<�����6��Q�4M���+������"�h�p�����������G:+-P�h�Ⱦ�X�	�+���+�����>0KRF��ш:�����r�I]_d���`����E���iSY���JX�yX�4(<>���"vlƜl�G}ĕ���H{�t���4/���敨�)#vYg(��c�raƝ�u�(���U�RD�,���k��B�#&����S��GHt�#�����[��A\��\����m�7q2�s�� �:Hz#q1:�l:���o�����9��ߡ�Â�|��Q<���nw��좘���`�l��h��i��?�w���ZM_�SzYkOq�K[ ���%��
`�b&��*.�I�4Np0�2�[�wv����G�z���e�c�^�����mpқ	J���4���^w ǧ0�q�=}�eWK���d"�@� �k-�?E!G�y����˗�S�N4T�T��"a:�%"��d��ܝ��$�b�a���@�F����#��gf���	4�mlt����y�ӱ��r��u��8O2���j���������*��Љd�����Q>��f���Ĺ���'"�y-�\DB�b]:�j�9qA�R���E��"��߯JjN8m� *�䶬|MjGg/����,Y.��*�������X��|��իW�}ćG�p ��s�!в�ý���_6;�.��|�|����g9k\\J�t���0�]6��Ig����r͎B�f����ռ��qZT���"c�hcx��8���g� ]�����H������Xc���w�0{�!�!6�Bn�ԉ@�_~������Y.�e����t����zb�j�Md��Ԙ�Û��Pܞ�psLC���ȡQ�� !qA��Zl�fm�*�T�-n�NKc�Y�T�ÎҤR�=��������`_�*�'gM�Uu��G�����u�Q>�Α>�����jjP^wR��:�
�۷�A�)2�bm�'��~�2z��Fl;x�<��\o9Vb6�y�(���T����ٌW�rW�t�U-��z�B��(9� W�x���ś��ৡA1�:6��h?s-��������x���B���hf5R%#'}��MZ�*�0<B��|r�td M2vŘ}q��_��W^|�E֊^z�%�R1l�q��ӭ������-&oܸ��
h�Y�OL R�P�5{1DLlVfi�I�!xdDJ�yS��0�8�HY���3���1�?Su��0��r���1ɖ�cW���w�B1>��1�$6/�16��,������33� &��^U������{ov�#k􁷦��
ӳe�Bo0�V���WKx�bnk�r�t�'��vvx�e��+y�r2���$O��������1�c}p�4g��$��j���l�O�V��Y�X��в^�,�%F9�� ��C�P���m���Z��ƴ�goPQ��@��5.���d,���lk(H��ҫ�sYd�FP�,ĉB۠#%�؃ٜ}Kr��	<�/��%?oo�/S��g��є�������&Z@�~���~���rU���)����1��.��Ȟ��6r�,5��&B"�q���k#�ɔ��5D'*��=����߭Ѷ�Ǜ7o˒�a�2�Y.��P�t��p4����"Y1�r��$*�`��"g�T|��O���\�"�h?���Ӣ���bj� �6D�\��z���pBz�0���n�վPT{.ݐ@�X��qfb��Y��U��W�4�V ԄX����-eد��	�E��܈�����d��\�$�V<4N������a�[�W�gq8=s����!#Rh��O�XRMg��
.���g��`�&��2p"�y�8YR��wOv��|p�ҥg�{���Hs���̳q���h*	QŊ9 �#?a#��_�b��-}8صgCm_�E�E���Yf#���\'����(����_�ZW��L<My�N�)���x�k&X{aݺ߽���?nrš$��>=?n��ȣ�l)A�|8w�����ݻ[�b��]�+�Ï=�m���ѣ�=Q/����]G���Ş��-Tz�	�M&HOK����Dc����1���i'bBZ����P
V��k�,�93R���ˌ),�N���I�e9N���w�tUp����	i�ķ���p�]d�k+�ֆ.L�Q�;^x�II�Zgt��p�c�(d1aHl%O���ㄐ�i�*U�s����i�.�Yj�ը�rA+EV�~sc=�����?��?�JĽ�
-��e̝��1���c%J?��`��v^�j!�y��`��>(���j�c��0�����	��jE�gxe�9Ôݕ������0���9��$�Z_������z3x:.��<�*�g�Œ7�wa��ףQo8b/�z*��� Ž��n�����6�9'�NO����w�9���zե�/�G�Q�|��y���Y�3�UcN5[\p�i���� TJ��G�-��Qy�#�~ʃXt��C��4�݀����BiZ��{�mg�2��]�>��ҦL�"Ŧ�ހxb,���.��۷����ӳ5b!O�B5���\=`�H1�Ƨ�k���5J=N��,�5Ɨ�g~��C�6�P�&�
bN�ʊ{��$�j�=��k�Oj�P�\Z76��K�m)��Ơ�F)E(Gf����]�ku���+2� .�ّ�,��=Iy�ߕpA~*1$G.r�J��$��V_n�N�;Y�m�{�m�.��Z|�G�k�='�;������Z�� $,�g)����]���_ޙ(�4q1T��>زt:!Q]�Ă�9��
r������^�1B��c^b������L�g��{A����Ƹ� E!ٜTA��<k�y>J��?|4�6�����)���0Y�O�<����l��bD�5J�ϲS&�=��%�>U��k2�e]J�|vk�+�<s�u�&D�pP/0,=?RE�%2�~�'GӎWG�[$�uf�Ľ������g������o}�[���w�~��W��Q�������O��y��ܡ��abcocS�K�6ٵ+�<-.ݵ�0�����6�B�sTbm��jMv!��e=764׀�0��a6J��Z�9D�b�&�=c{Mg�h��	Ij�R΃@���o~��}^�~�W~�W����0
�s����]��&�)��������/ּ�چ��[b�3�!�x`y��O�`T;�%��"��4V!8����}E�[����K/Q��p�^�+R�����S��4�H�k�a��<�'�+��y��0#��-�V>�ʷ>�׾fcYZ���P��{����UvƷ�l���=o�>{�!�lLm@�$�3�Sv066�j=E~�j�B��e�	�5�&��.��mNOO	l�4���C�-1R�����mv��i�K�!�.�o��oEf>��ϋu{��g�Pݾ}��g�[@��vr	����J���~���tȗ~�{��p��҃��*�녏+J�.�h�7n0���RͼK����;{(�Čg֋��1p0p�Q����X �V�x<GlYx�Z�A/l�%�3Q(��Ѱn�U,J/���c���W��y�b���2�T�_+â�Oa�o�~�A�Z'W�r�ҤfD�<58��`#�~�xϴ�r��A^[�Dv�E���6�����<
R1� gU�f�.^�x��%��`y"?߹u���8Z�V.�|��_y��������sT�e`��ty��
��Y��q����)��t{DN64!(?��8�*Z1��Xmq�FC�A1 �b��n��S~`G��O�����;�#$n�!���&�BjS�XQC��oȱlo�B��k1��=x�����b̺�$��
�t���w�g��R��~������|@Y��7o^�p��=�v@�8�0�%T�+Q/��������M��������>9%�Oa�T��#�s��1���� ��p�a���;TD�Dt���"�/���ϊӠހ��r�PJ�>����$�dp��*��_�Fh�oDI8=�h�#b����bEs����m1X�F��̖�&|���𤾪WjA ��Ǉ1�PK ��ek��fv[�|��E�9gt֛Q�_��7F�Z�4D�T}�Q�k�m���,4_�tc/X[��L#?*�J�j�wx�=M�����Ť>E.Wg���Z+�t��m�o��b���M��"�t��|��- b��g>�kV�tC)�C�:�?��y䭨B�LO�a);��ޫ�3}�����Ԧd�0�5E�D�q5�b���56'���t5�9{4BT��s]���eF�(�#Þ�6K��������	7Y
Wv Gs~�q�$�Hc�o`�0�Ϟ�CL�;:���ƣ����}��c�W��ՠw��:�4�mu�j�rY��ũ��Z^$�~lI����5�mfBm���P糤�t�OJ��*>�\��gHR|�����'U[_qs��#�hq�dw��&U��ϖ
䋷�C��j:#�yh<Q?ϱ���X�x��G.�Ʈfi!糧O�V��U����윎�I
�sK���$����cdPbU&�(�Rw8ȑ>�u�	�#.�k/~�Z����e�9���P΀:緱����y��18��>U�u����f����y魬ż�,�	a[e/Tghy��c(�e�F4+�w6��BI���p�����d|2�{�>%ЂQ &_���uk�����q���l�ܕ?9V���]�� ?I�Y��4S_@WR�,^B�p��^��|W{
����M�=t�:�j?#��X�R��E6�,��v�2!�Rakk��]*� v���=�[��͌�u{{���N�t��MD9�������@�ZĀ.NR`ڵ�8�9U�|v�"�~|�c�H��!��E��,`v�T�����~���16.�{�N69�HSِ��&��?��
�-�Y�-ʥ�Q1���JR��|v�/
��)z���F��6������s����f�ym<���n/O�H]`2"�!�u�pG�[��U hvpa���γ䱏�5��Z3����*����t������k>չu�.N��|�oY��*0-V�%�L�)�Rӻ\<��@O��
�z}�T��\)	ts �7F=�=�4����z�c%2q��t��g�#������Ǎ���;���Oj'���z��,�%]��U����U�k�HA*gy:���Q;OS ���=��!��SW�|�_�R��흭�b�	�t���rQ���O|�.�����Gw|����a���o�D���4�Vq�m+����C�BU�n�8�˗/ǩ��@�!.��!�I�.u�Hr�`y��N��~"%T��ݨ����~��
�,ǣ��SO=%���;�\�A�ѾHV��y�/��������߾ʹ8��rvJ#�*�b�S>,�R�p�yFf�u��
���M�6R9`4*�eݑ���}��&���a1Z9O����O��˺9'ӧք�8�(W���<��4͘��'�k�"/��O[���㈵���ID��f���K�B|�N�9�x����G~0�4���0W�ԛU�<�K�o�Jq{��7Pk�"�WT%��T%�bq�I dG��bY�=�ѸX�k�ᚹ	+`�n�B�1O�Xd��Y�P]�:�
��x�XǪ�#�1��F����d�ȹH��+W�v�]�~]�t�ڵ��~[$�)-Rl���}��[o�%?����c���r5:�ٓ�8�;V�J8(����W���/�ѓ�Og_��n&?��k5��(��rLv�Bɒa�+�IG��駟��G�[,q�ݑG��K?bZ��*.&E.�	'6�]��Ϳ$��+"�Xf��a:�|�s�=G^}
�J������׭����p]H5��Q��[s(��tln1E}��������b<��(��/ɟ�gf��_e�� ;Ÿi�&:�9*V��[C�aX�P��wyj��"��ߍ�����x�$m-��.`����hfjkg[>{�ҥ_��_@"Cd�1��?z@J"��K���\y0B!P������� _�җ����j�O>�D�R4���n�����>��cp�\>���+7n�� 3���/����ԏ�Ab����u�Ħr��^{��0����{b�G�O%�b������D-�Wb�E�y��[�;�{��{�&��uf��(~,W��+��T���W^~y N����x��W��߾�H�yp�Q���p������Ӯ$�{�|�����}��o�_f�r�q�pTx>���Ȟ�C-��ͅ���xCA�*(�N���ܫ�x�P�U.:6�t��3*�x�_6�	12ϔ�0-K`0�+/Ow�iHc�xv6V�Yk�QL����-Gq�B櫥_.54�U�\	�����+��x�
.Ւ��T~y������-�h�$�t��;�6$"��{|�P���t�����"������������XWӳ��S�E�!�	�5���`���I��w;�L�_j-�T��}ϥF��	l2��N}2�qXXeXug-ndK������{��.��߁e�<Ւ��bM�*]�����>f]��%ś�S�d�Hȯ�x\�U�Ԫ��&�)	鑪m4��>tͪX�YW��$ޛK�<�л*(�\=���.u�R?m���H��y�z�:�5�F�|��Px�5Ҫe�)���N������İE��z��1����N���6��<o�M�����g�u�9]ާ3\p;�駠�2w�)���칦��lB��3H�O��]��gXU�)���l6���p�*�`�N���nj
�Z�J+�z�D`�U1�O�>o�f*���Ø����L1�i�7[5;�m������"cH��2��QD�qǑ�(�7m%R�~П��~zCbp�@#M����$�sZ�|��%�A�49e��Ƀc}"�u���,=�ϔ�1M�B%-��!>��F0C�Wb��!������(�ӣ]W<s+0��=D�b9׼0q|X��:i��_���vԁ�;仓�9>�({����D�lݝ�v�]`�����״C�����|2�W#�K0���܂�'V_��*,5��q�߮���tq��O�$1X�.^�0���L��l�H=h��c����d�D�U�=��M��t0 V��ٵڰ�H�M%�:��l�,�\X�n=I�T[3��V�{��-cB�|v���`^[�Et2xAͷzU̬e �ʷ��?��V� %��n�n�/1��P6`l�Gc���'���g���Ή���E��\�ք&���B��C��Y�L6�/�����=��_"�#ֹ^�+z�fs�G�>Dk����h+��x�j�d�d"�����8��p��Dpc�_rY��[F���
��ī�8����PT~D�>�pL\��^~��kK�����w6]�ǐ ù`{i�C7�G���T�Γ$���ÌB"�7���ٝƁD���m��YF�OnUG���%�k_�=r����4��u]�M�1�r�C=|�1^�������k-b��*�6.��$������r
{Cg����J����/W�V�[�~���G?~씥���\D��sR/1�d�Sl��M�H����K�����<j�z�8�����l�켮�N>7v @ @H���]$��U*�.VI�?�������*Z�T�X�$��� � ��ӹ�擽�^�~���E�-Ԡ����<�	;���J'�aI���P���	&z1�15"b��XB.�v\t��&B=潞 g�3����`�8��+Q��j�ʬ^?����3����������訴�b�{���hF����<(!Jx��jE�[����q�4������ ~��C���OΣ���t�ӌ����KqYz ���������Çt-���^������/j�JL���H���	j<��N��w�t�������B�k��B�upp@Y͘>I�=����XC����3��'O���n����u_�q�L)È�g_�Nh�cN	``�2�F���vb��^���SV\E7m�p7��������%{a7��2�;���9����Noo$�N��H{�	+��O��o��~�^z��K/��M�������i�jk!�@�޽{R^����o��w�}�]Jcʫ���w�d�K1�� n߾Qp�Ν7�|�rzv�ӟ�"���ٓ'Jo*�ũ+H�c�[�	9�!PۃA5�'b�a��5�o���[�����fM�9vz����N%g��g��D�A�D���Ϻ��*@J�C��/����o���_��_��Ur���6j�xlAk��񡮔���*���-vWe�$���t�
o+R���$-~�vww1رա��5t^���j�mi�N�eH���b&<8�Em�1{���g����w�nb=~��Ak��vF�f��al�W^yۯ1OF��}�r�O`���|�����|#����ML���)v#��B�|�4����D�Lb��7��y�ul��lE�K;;dT�$<�;|�嗱������&HBC��+��x&D0�Rӌ�d�52$�l�:�F�Mc+~����W�"�Y|�l?~�oݼys:�q�ȣu2I�4�*m�����ى��%��w��]��f6�KБ'���b�i�����Z�J%	�T���ҟ�v��%��8�+1�:1���E)�C.�����G	��MK����R������k����1N�I�ՠ^��7���q�ލE�J�S�{�U���1�M(³m�q �F��\��\������,3�J����j
C�G?��,t��N�a�ǹ�}�~>??���O�D�|��15'���٪^��0�;s���̧I�b)��Q�,�Ob`��"Fq��Y�lQ��K+��u��Ї��Ѕ�Zm���;^����J񍀂g��@��+m�	�Wv�f(и6kJ��Y��.D
N=��ÖR����u����k?s�$y�
Ai�֕�G�(��R��K�6�e/v���A��d�Q���m�r�h�Rs���r�]eQG��q!b�{��\J��&��؈u�:�!��OB�Q4�ZOJ�Bm�Rh1���s�������n�M���2Ɗ���UV��?�Y�#~R�":�1wv+KM�f�4K�\��	��]r���s�$��*8L����:�%�0�C�'U$ $�t��/r���0d:�y��a�:+z�(�1��߸�c&�N���}��':R�+�J����;�z�N�K��J��:�����X�7��k١���z�_�w�|�)���cT�8�09�)���������z� �Jo�[U���d#��++��b�m���U��A�F�ތ�~&�l���ŲS�I4t��]�Ԟ!0G�	���WaaOE9�����1|�6������: ��JMX�ʩT|5�)q��s��Ea>�Ky�a$���w����F�ako�Z�jGB��; Ȃd9�����mk+˓�\�0��v���qRwr U�a���BF+lb*��~��T��1X7u��a$'��jY�������_]�ze\ᡰ"��O�*I?���%u1F.�Z$��H�θ��O�D�mM�X��4�����Egt�C����$�9�̆X��b9�����I��j!���L��@CBm�r4Hg�ad{��o�t:��6�-��;�Bv#��+�
-e���Bp�F*a`�,q���;j�� n:�،�c[t~�����s�f��NO��9����@���7��C�ڗ�������]c hE��]�K�%����{	�O��.&W�����J4�4z5�I����~O+�;l2Ƽ�5�u^\�e�E�wv.�ʻk���a>�����赕��ql�94�h���óc��DE��	�J���*-�e�sU�4e L������	f��ѩ���!�~}�y�ؙ==��{�;�"Bè^�&E1�ḩ�G��<:�������PP�(���ͪ^���V�$�}��	���	�W�m�������J�6J��I!�ʦ���c-��j:�LȀ0�,M��Rş'Y����3��y�0�:
�VB��d*�	m�3�Y�kȳ�^e�j�i��6��LY�����
�c:;9�g<܄W�%2N�`�%�t�pS��|c�B�K;Œ��n�ϻ°��b[Gq��ltrqO�h��I���� ��Xm���i����,����t�c��	�����â��B�66�///<z"�P�r{s\֘�po*�uM�*f �˿|�K_����y�����S���s6��"�YpVì����d�6b����_^5�\����tc�S\ͮ=:=�A!��i��o���l>�XZq����O�/bO7ŪY���(mc��ӛ�B������+�3��$�=�koS�0���h����g��t�*$l�=�Ь&���Je.��#e#BoXl���?������;:9���6P_�ʗ�~�m�����1-�V{���[�xXͤm�{!�\�>����[��)�E�S*ͺ�P��DwK��n�/�LZ�fZ�.
�<��`SRi��C��ѡż�I%�H�h�0�Z������@��L�|��߿���Ţ�+����N�%�=9;�g� 1v��!|0*�����sZ8>��i��s͞򰹖u.f.��$<�<K��YP3�#��ĝ1���Ԩ�}�&���Q��5m�U�	o����"Q�鴞K���p�����_/��v�����q�(�?��g
���AedDi���������ͭ�D�!&����!��@���Pڒ���iҧ�	����Z)"a'5aCV��V����&R['A���þ1���!��)��%Ԍ��k��4K
�+<}��_��_�W~���_���ፃϾ��| ��zB��e���jr�O����~�w~��/|a����;'''}X�
?���ˊ����+�����w��y����JFG�?��6�<����}c���7�5��͠0��*��ٳg�F�p<5�(m!�&�_M'{�7:a�(dt�=\b(pU�	nz��<~����ǘ4��@3PHx�p����%����_\��ip�r�]K\�¿��t����݁��{�q?�_���ͮe'���wBW/�EۻLB�C]�L[J�*R,���v�M�	l��B�)h�T���b��{�/�Z1G;��@��#�x���K���|P�����ۿ�+2�-i�{qy���G n�&哀�#5{ml�pB�!���`0*g{ov6���|Z¶�?��'?yp�>��`M5r!��A"���������D���O�㝍� ��z,W���	��m�e�߹)��+I7�N���O���^7:==?;��ԼI�2��!�/cZ�Q��Y�*��߅a�/|A�a�0&��9Tw�n�1,�S�:�X]Ɨ�˳�=<��>|ק'�O�/��ɶ6w��{��|��?=9oD�F���J4�И��AQ7;;�U�]Ngܽ'GǸ�X�����|���կ~�;?��ַ�u��=a^Kdڸ�,�Q:��d���bq	���"��������� N�7�5�����"�,�[u� ��j�*�
WC*
�/�%v�E)�]�\_�sc��7�����F�������L�T`u�cj��R��1�W��Q�ScA�����b�A+E:S�����F�A�Z����+�j-׊$P�I�E��Z�*�x�J۴"jh�B'u�'0V�eqq)"7��IZ�g�}2�Uz��M��6��)	-a���*L������)gN͗��&N�ǏU�/������G��,�<����x`���Ue�t�,�E��I���]%�Z(�)�ac���B��ȋ��n�~,��i�����#�����\<���|~Qb �%�8�+���m,M�zu�}(F�|!]A�<{�Ν�H����Ê�K$����qQՄY<z��V�B���?@�jʫr-��M��Ú��[��tc��l;�Y��P�r�dO���װ{�		 �D��f�3t֕�G��EVJK�WSa咟q|]`���z��9A�5n�R8X#���Q�X��B��a�Fy��ȫ�ڍ�^~y�F��oy,��F�ō�x�H�}�:^�+c�g��|ƙ�k�}h9X� ��Ǵ�p�Q�Z�y]�j˲$gSc��z�.��i���a��
uu!�^+k��x=��%���v�*�q'�0`��Y�C۫U�[k� �e �՝cYZ���p�z��*�^'�R/,3��j��_Nro�є��V��������}h�q�ƈ�*cG���l<\\Iޖ�ϊ�[�\)��b�H�J�2������u�]����1uZa!��R�Ya
�jՒ�`t�|m��C-*L����*�Ek���jd���E�I\�f���ay��Yc\���&�Z.�Ga�c�JQ��=��-��Y^�������^�]铄���fƗ�+יlvdܓ����3���3+�d�3��$����ou������Z�į�c �����x�c�
Gs�_ǽ�_�J����>��!b�ӧwJ��G���}%�˥�n*H�^��)��1�]�R�Z���xQ�Y��2�dv�G���,�W���Xs�rA��W��/��C����woC��yF�P�Oi;9_��I�� ��U�M�ܢH�D�7]KD�3*IBT��Z��^�$?�������n߾��!���_�t�F�"BS�c��1����ʠ�q)1�/�����K}���4���;I�8�Ȥa���MC�%�4��Pg�� <m[�ϥ��
��n�+f�<�S��^K�r�1o�0X?_�<��K8�_ʲ��5���H� ��%��*V���b�H],~�$c��o��v�.��EsKebb�5��zc��+��x�W%�S�BȜ��*���Ae]�(*Ŷ`�+͊@@��W|�b���n�[o�w��xC�6���6n\8Hr͕�	NO�I��_w��d3��h��Ed�"�a�q��V4uQ�JBT]��5��_�;�H#�$�Wr��n��i`�aa�IM��\we}rr��PI�<�;��bsK���l�ْ{���˾r��a��������x�������_����%g��
�
w����?�p>_p{�jTٙqL�C.eug�\ʢР�T�DL�&���Ǔ*"�]C#�-��%��u���=��@5��%�aD����_���ӧOy��sa��V<;�<��K����UTژ:�).\
{#��k�=�����'ƬRiժ(�������B�}
��X��O��>�,y5J�R�TfmT�;��9�W0bH���a�az�F����0b�>��-�,�'�H߆	'�G����^}]*+ş.��!J�D�ƪ�:��o�{���c�_J�ǩ��;2<�7���z�$�O�!������?����7�d8����Cޅ���_�|�x^|�ŗ_~���(�p�q��-Qb��믿�Ʃ��k�b#y��*
�i�6���7�P�KjC��#��v���ƞ�y�&$^���J�b���?��W���#e2�Ĵ5�/~���
���TRx.ܚ1<�4��ʻ�si�ļ�4;?��b�>o\�ϽF,���m��
сQAh|����$C{⯭��	��+j���~��K�q=-!��\�۪#}d�2���ֺ$/�ڌ~1�}�H����ߤB��ĭ��P-��T�Ju�1jg�I^�P��rlV*2����ax�Q�ƍN�SZk�y��=����Z��J�ƍ���rBIK�`	��U�ޛV1d假Rb����;����D�b�e����4�pM(9_J��t{}�Q��V�KOW�B��5�FE�W*{�)� ���}���J��g���
6U�56h�uH���L	@��[h���dU)g����[g�xa��K��rT����[�6ϕU�&����6&��8����r�k�����n`D�.�F�kh����ZCG�f&"T(�@~�����|r���w^�"	H�E�"��3�����V�[5V��d~uC�<�8�`~��{��T���޾��=��,�v����r���tJl�a��&g���ӓS6���ğ�"R�m l��r�[m��1�l?��-���|zI!���.D0�#��O� <�>���.d��<�/X�!k� �>��U��G>�U�~�q�k,H{`(v�*U@o�˧��}A���3;��J���=h*t��g$'#/�BO~���{ߡ�Z�޷���5q>pk�ƞ�v�����:.r�-���hJ@Q�IPnb=5U�H�i��Y�z`���x.hj��cy^��X��:Y��M���n����1ֹ`-�����\����	��0C�X�q��#���Į�Sm8�h��:m�֦����bz�=�y"��E��i�� t��؅/��ʸ4�j�뙉���m���B{%Fj���������޲���cTޤ|��ւK��l�~��>X9y���:m�*PJy���j����
��
SK3P��|V���������7���Ͳ�/�������S�}��	&Ǽ����H���B���I\�D��hc�Kxp�(|�M`��r�,��Z��#�Jz����[O-��z�ղi�ȱUhs�l��u<	[�������vI�rskK��FuOb+�B�P��Z8ؗqF"Y	Z�T��me��k^&�Z�T��j�PF��	����W���M��Ղ�[-Z�T�įAUwX}��\��L#��ے�9�I�[n0葕�zv>Q&���v�� 5���I@��82���Us�`�c5-2��8�����Ga���B��n����]���][#���.�=gOO� FMvM3�84S:+��!1�A�a�::*�1�7Zl+M��Hlջ�ˍG�#-�Y�	\��d��J.�Put+����M��'��0i�ԍ��kk�*�gN�(�@o�����}6�H���^H�,�GXA�����}l�]\�t�xޝǱ�1lo	'4<"^�Q�J��w�ߗ���ۻô��De]ᱺ��֍�	v�d��J�����D&;V���]ܿ���'��ۻR6���4�A$|��P��i��_�ɝ� `eB���� x��E�ǭ��``�S�����v׶�沷�&�����'F9os��&f}��C癬��U�N�G�� ui���­�D��EYM�v+uʚ��V;�k��^��&5�P�?���u�<KKN&�����Z�0`�խ��5e��K]F`�91U8@�	<>9��.� m�ߓ3`��-W2'�Pq��h�Ν;�7p���~�����!���g�ע
�'΅�3Q+���RB�����e~C���
V.m0l95��{�V�,Xr�;�N�5�'�$�`&�틟�?�,��7ƂH�����I#���݋�ɇ~��g����B��'�R:ކǕ�����f��������V���3���`/����[���O����>~�q~��G/��2�[�GR�j�i�"W�j�N�e���|
�kD�c="��b\��=Vj�`-SY�*W�{S�m���Rf�F��Z��q%?�pC�t19=>�F�I��g�K/��ꫯ޼uS��0c�R��J���:�`�7�����,����"�7 IB�#3�<��x0I�H�(�x��omW_\\�ܕ��Ĳ�l�D���M���tW����1�!y��HT������唒!Y�#K���5eVw��\���U��x��٣-Q�,��x{{���#�!�0�TQk�����;�R<�?�1):[kp�Ob�VfN /d㤴7����Ȩ���?��D��@�0K�^X6�aA�Z���1r��/Z�wS�f#��+M����9����D�K��ӓ�������J3Q��G`�L�E_K���w祗0`��~�T^G�KO�>>�8��ƨ~��}A�-<#� Ot<�j�9�ƿ��A���Ƶ���Փ5V؄�뢚��//.>��8��d.г!�%o`l���'�|2���+R�5�����Y��s��@V��[����9T��V���K�U��,����6�&ʅ�x|\/Y��)�6Iհ.�{�W��%�\h$z�t�q&}C����DC��a\����M7F���
k�rnr�̥�?vi�R[�b�a�S��m&5B!�F���tO�Mhy�@���nb������?��ϙfÃD��I"�\di�F�!�Q�<>>��U�3������>ͳD��Nؓ��prv�09�R�Ng���Hdx6�H��`(]צ�+���Gt�����p�ĸ[؛Y�}��zb��=%h&e����\*�|������>q}p:?=Ü���ڂ�7�/���ϑ\���j��B�!�����8�>�vY�|�߃f"c�^w�=�E���cf-#k���N[km��BG[�����Ol1e!� ���SNRhҴu9��0���))t糩bɅ?'�B������7~�^� ��$�|���ɴ��C�M��� H�0���q�Ta'�q�,�_��Q��z�+��#����r9��t������VM�\-����d�� �V/Nq����\A�	�vgi�
��m#������ N9�hYb?�
"�y3C��p�[���FnA=F b�m<���ȼ�K7?���ցn�F{d�l���Z5�h8�e����_{�M� �ۍ�s`�i�&��d�ON�&��PF��>��:mޫ%�W��E�]�����ƕ����%鱒�ٮ=+�lʲP�����|:��
�c]̎۴����Lg���y�����h�Y3������G2ǻ�>���?]��&�����:�������Lx� �>>��������R��S�&��Ֆ;���Y+j��9�nn/v��yn�yco�������>��Y��5�\c<;�!��zk�O���k����Ool@����}���Ѝ5B�"�D��򇐑\�kj�Ǹ��`'�{MT�C�HŨ��/
�ZG��w����T+�t?�HS���H���)���KZ�7�^]~K���V������>���`�İ���a�1��l�Q��<�x��[.�Mg��)�<�ZV�	+�b��ûn{4�w�u��#�ۭ�Se_�q�VS��Z��|��
$�0�q8q�H�Q{�R��F���t���x���_]JQ���Z�ҪB�t��[<&~�L�@Da�L���M�ɉ�l=�(���y�HZ���/�U�s�غA�����.M��%�4�j��=� [y2�:�P�#�B"0����>���&���Z��������U�S�p���29��+O���!Uhm�?�(������p���]f�iV��й\\��9y���H�*0�G���6C{�6�Ţ�����^7.)7җ��Օ����'�zh	��ZfY�v-6�k��*�n��N��{777�~-ĵ��C4U�<�b[<�<{�L�@}���oL�S�ơ�9
�mg85��@�/)ɽuK.9Z�|3�|8�'��S�E ���-�h�g��d���+���-K%���r�*���q[˃(y�KT�/�DC,���R-�j���v�U耷��ei]��JÓ(���?²�n���1�1�	k�Z�R���"��+���ħO����]�O��Wt9ϲvJs�����p�vZ������������������Í��j~WJ3���s���Y+�@�.���胕ږZ��l��P��T� � �τ%��/�I߃M/mCܪ��
����?������[���7�����4&[���߿-�s�v�GO�\a�'�B�9b�cs{�T_8�cl�o}�[_��!d��������_߿n ��S���*C"Z �`�Q�{�������F셶HfC@pQ<����X͇'�cE-#�^*��t�X�ėR�kW
 .
��p�R ^KC�7�xc�1`s<�ҕd(�	�Xr+Q�a����*�V+O�Ձ�ߺIH���Z���^�O�j�~��7��L��/�x�6t�\�/
C�(��E��gl]u��D��,s |=�n�=J�gg4�>�|��|��'ʨ�MJh���'7�ܜ�mg������"2� '�O���C�|�8kV�l������x��W_��o�+V�#c@��3��26�G}D�D-��R�c̐<4���4o}���	�WK���[�FԎ���4�D;�>�0����������{����]�����4f��W_WB>��	YA�.������"���+p0\��g0Q�%4&(�͞Nd8}���{����ׄ_�����s\�ɓg�~��g?���1e����^�w�w{��衉�!��az�B�7Q�o��3r�(�<H�ލ�����B��pb76����b��;9��I�}�*�ȑq���ݻ/�r�+��C��HdKȹ"0)�������:~��d*
C�Z��5��UFU�B�_єj�ݽ�O�H�m/c߱��C�X�HI~ʌ �i��#dSq$�f��������^h}���$r�r=�UGG��EF��!-Q֊����(B�\\�� x@&6�d�8�ў>}*k1_Pur��K�Y�)�]F��#yLX�RO}�j�\@'T ;n��ɴ̧�ʚ6����DC՚�������af���Ļhf�0�������n�@�ӛ�	�X�<c���vkMG�e��:��b�oml�l� >߾ΎҒ�+4_���O���B���&����i�Kpǃ<f؊T�~��������l6�>���43*������U�,1ĝ*2Y3���&�]ǰ8���l˶���Ήhy,#m�G�m��S�W�����յ�3�����S�K	�е~�u[���[�����3��;ϑ�<��y���'J�2a�S�fg�*C9�8#���K�S�t:&V�z� �`߄۞Qo�5�6��.3�E!���pQ���!K�4�X�Rf�Ƌs��`#Iʷ�4]�/ʸ���H
�2Q�u�m9C���5��.�� 3������s��"$�L@I3���i1x�_��r��,��F^������Ldh���ōѦ�c�Xoo��5\���O��A���}H�Ǟ��5������R~,2@"i������y�6�m<
:�[�O��e5���[�WӰ�"�ny�?=��{��,�!�ϷW��^�� ��1%7�Wě2�K� sN&O�n�v�G��'��5�ҳ�f/�eZ��;��VRp�i��S��K�1
X*����"t>q�4qn�*�ajM�k{�k�W��} :2�qe����к��IAt7�okU3�%&9�i%���_]��*�i%�@�(��)J���Z}!�se5Ūbck��8�0��&n3h��d���;���Q� ��E�F��� �9�X�~��޴|)S�(�=��$�rۅN�keh��߆Q�0���E	K�I~8,B���8�V`qv~�������G��Ae{KSO=^G�ix�� �k6R�R�&��f}ݤ�ĺS�gg�Zv2[J�3�7�P:-��`k4f$U�v���]���-e*Iֺlj��(�p5�N
n�E�pzU۱�h_{,��riR�t[D�W+��2��r��c�lnn�X宭y�!Z9D��J��Ƭj�'��=])W���Ǟ��"�hX�Z�m�[�g˪lVB/�-��
H�����K%s��	FB�Xw�'���������L�r^����} ���.��E��&ݳg��<�Ӛ�Y�/c�-=bS��*�qooG�R�fZa-Q�,��6� ��H�;d�j�&�P�mA�����,f��������4��YKC�l�h�E�V��a6�z�UJ(��qXR<V܅q�Q#��@On�m�`�����9�d*'�0v��h�\]]M%"��tMl-wX�#)<I�.�b���nZY�~�,'�x}�J܌�r�X���֎-DԬ�|2n-3���2�W�i�+�)i{�OMq~y�!ᇷna|�޽�J��⑇=e?��
{����Oo�&y�p��.+>U���+ �Y�ʭ��H��5��U^/!�䝑�2N:�
|]}���^�U!,B������XN��FZq'F�<\.��0
�xYVW�R�S%t���┣2DR������� j�br5�pQ�hwA��z�!0�byq��n1�7�p2��y�b$��b~yq4�W�n�*���{w�&)<XH�.ě;����
[2R��VY�{����b]��_����?�����o���������{b�j>\w~�n�b⤐�_kXk,F�3�ԯ����h�4F~$0��he�g#KQ3�C�=C~��rQ���ҋ��=�/�.P�)q���t�A��&�HF�a�Za*�m`x�-���w�����ALo-sb#A�_�Y��&9����Vp�Z�����*G^D��7��r��4�x�Y�Miw�arle%m�����9�ɥ����s�x�}�k�
J�q���v�G�a��3�@�+���#������z�t�(���-�YY/,���~9>��?�1�lt֟��+ R���;u�u�?-1|�'?�	�7n�����=|��䄔,>I�cvڱt#�:J��>c�)x����K���9G�e-q���bzuVW�~��L���:C1s���~��Z�����/���������c3�C>8�qtt����4O�3�X0o��qE�*&:�*�<Q<x�؜�ͯN�%5솼���������nc\��[���*�C�
)�e(�x~.�sgk��?==�DI�j%��0s��o�J�)�;K�ѿ��a�/�u%מ)���y�\ ��j�� V��||z��j3����Ӂ��������h������
Ҭ�X�V���^Q���9&beјd>�U�f謻&e���2���ę�f�E�T�t�T*��[V���k�NH�^��-��6CX��m��,Q�\$C�EG	ބ�=R�ye���?=;��#<t@u�w8a�tR��J���(�$}�?)��Vc��t:�l��7��B��$���8�,Q�ݹ��e���΂�4�h���kCz���}��l�I�iA����*�J1�M���p��9��ʢ>ZI�e!>B�
c,Āl�"��%�슶��-2D%e��L�Kx�N��I���+z��`��i4�~��	G����$Y�D|t3q.��$�'5Fy2�^fQۈ<�dX-p���Sg3�8($'0�t4��b1����_��T9<;����w~�o?������=~��l������C]^�I0:���<���5BM����]��dX�~�V�VW��npz�4PN>]^���XݹsC�|�ר���lzu~q%�u��<��f)d�m���3؆u�I
B�b8nRGG��p2�0y&�ߒhog��\..S�5�Y�v�m4��E嚕3ѩ�p�ZLS�i��\04:9}�:�*+�(=��s�o8��ܵ�h�Fڠ�UD5'��Ȩ��8�Tͪ�za��ѓ�#�a���p�8!���� |͟:.R�V��"����ت����֒�3�TL`������V�������r����P�e�k�?�֚�{����|�/Z���c�Y�Tb��Ե�Uj&�I^�)A�gT�p5��1jv=��(E��(([�n�{��E����.;J	{��O�g�޻6�C�[2��W�'��qzS+R�%g��I�ˬ�K�~�k���
��5n=5�e�>@f�N)���쥗^�1��x��1������3�D��0�P0�.!���A��>��X����+[�@z����V?�Z I�-g����E�U���ۃW��"��㝄����!���ӎ�.[�4I���PQ*�nAA&�E|ت���h<�d9�6�Ֆa�p��{Z�h�@E�0���0Yk5w�!��#v��Kn���x�Jվ��[����I)�,rأ��݃��xc[X�F�}-�8�*j=�Zmj|�D�/�j�&��ӼG�Y�Z'JÊ�Et8�R��n�䇹�$��;Wӹ�0�O�WG��x���QAh�ώOJkc��.�ዘ2#��̽�Xv�b�dR��9��,p���h���s</��!C**o���el������ґPr!G��N��Xs���_��+�%�^n��M!xx_��*5�/��b��P�
�g�E[�3��j�QOP]��n�Y`������lи�3{���[����b��R/��#�\{�[l$G?�r	��� �C~(N).��V�r?���a����섎�4�����F�E��V�Y�ְ0�Z#���L�^�N%q[(>#1�f YT+�$(�6��t�Q�:�T���5���L��V���X9C��^��|L�u�ەki�Y��(n�'%��h3�֙����-��a���e%J�v�9iOvY�����ٶ(P̋�V�ɤ��ΔF�<J�t�=�*f��Ek�Q\}��h�_�!�vX�@��w�"�+�S�������?Z���'Q��e&(^��� }�[�Xd�.&�5tB�1�ȍ��o�_����/j&_�g�+�'�`�N�FBNƂK�"�f��/��������Ǐ�/��_��?��������;?��p��4'Zp����ޖx�b6������_�;8��׾������O�:.ZW�ԐNޣ�x����
������1xG[(1}���li=�֫�p#��
,��/zԞ���:a���1
hf�`6�yC6���b���_�UH�n9�V�"��d��1FL�!ӂ_��y���T'���>��9�E�/�J���X���bP�P�fi��/>ͳ�1����B����թ��P`n�h]X34$u��K�a�Mt���f!ה!�8T�޸j��:Xt��ě��5�F&��f{����[���f��Hdx�x��_���?����z��ݻ��'�|�Y�;2,!��@̓8�N$�j�'�Vx��#D̗*V�b�Y76M��ł+ܼ)U�Dy/5)�kb��"G..� ��z�vOS��=���Ky��Rc抒������.�[|��_�ؐ�_�؏~���.rcr)���sQg؜�����d��,��Ԇ�h<Qj���;[�Bé��z���F��|��QxqC�tJq�,��|����K��X�$>{�
T!ؖ��O"��cA��Ա��ܼuH��ťL��(�1Z$�j�$�&��a�>�O��� G\2�҄;qo�H�M�N���A�F���3�E����Z�B»ƈ/��G3R��67���h)^( �����ȩ��C�:�5�x�ٙ��I���e)9�]:c]�aCP�Bs��F\���"'Q��<_,��īQVȟt�|�O"�fgi��ְ)�q��A�mVj�N���&���O*p	�c��5KhC�Ǝ�ߣ�j_��ծL�V�����[�O��$^Tz�rp�G�H��$�.��Y,�:M���d:Q�PdWSV~�]�ve�����������?}��Ge�lx�Ϟ=)�V�9T;�w>�?�.�3C�{8HXF��S6�k1�=�7�-�(�74��C���&kv��pm�K�E�ћ�U�2���y
yd��B���;�V��p��(��߄��\��U�tJ��
2k$G�*H?�(�,��Fu�Q�f��!ц�\���=���y�
�A_�:K���fw�:��*	����4JYL�a%3q}���uzx
>|k�8~��s���)�뎴~�Gd�B��W�3y��G����R�M�>�~׶�*���b�#�}�fm+0uP��Vd�z�K_�@���en���:n�@���O"��|���*�:k}&3À����7I�Qix8��l���a��;Rp������	��u�z4�σ(�5�z��ԯlgqF���K%
??2@�JB�(!�ap���u��p%��~��Z�Q��[�/���k��Va�:B�<�Nxe�VBs�}��o]o��T]��JZ��%:V6�EYh��b�%D� K�PXㅢ�asÚ	�+��q�^�*G�:�mCF���=�m��Q8����(o���S)!��jY:*>� o����1I*'"O��p�%A���*_�	mWT;���Ū~�R(�"T�l#�s�kK��d����E��������Ϟ������><�T3���jV�/67�� �*�� 橣"��10M�> ڭ�(�I�����/�%w]�]ha�2�������	�IS�᧕&X&�(\��Վ��JR.q�u^E��G�p�N&u�����h�RX��ر;y4�C(���e��ۻ{���Ф捍S����.��Z�<�����>ï~72 �Yr5���M�8�pR��T�4�OB)�H�'�#רǱ,a/��;�76���O�cH�l�Z^M'��C�PX
Q�4�%�4��Od®�G}������H�q9+�����̆����3�n�N����S�]+�����%KV*B�����_4Aw�psw���1AK��8�H�$�`%�5�䄘R�U����_DY��Fuo8pv�����刍RY�%8�4[�	��CQ�љ�vo�S}�dK��n�ؙ�⃿u׮J��t�<>:Y-�,#?q�E��3�NB%�"�p �q����7����.N�,C\�4�Uj���pz��/��*�����bR[K�^��8�렟J�t"$CU��BQU.�_���6������[z�f2�\U/O��vU,�$�����x�l���HZ�ܟ�^����ָ?�r��h��`ɇ_]��@.$g��<�Z��(���k�K�8�C��5���C��h;<<"׫	,ahm���D��ؗ�jlh��j6�I$ϓ�tA�a���S$X�9&��*�8�]ʼ��^~uy����z�$3
e�������gF��1ɷn~�k_{������H�����o�����ݟ|(�5�ww����$��c_��|�{���o���BN~��_���}u���eXzt��1r�Y��6�%o��Vl�.��� �t�(���N��ak�%kD140H�S��
����o��z��*��&��م�Xk�.`�������^�h ��K������]a�����՗����-�/TQo똃~��%ì�#�橷���=Q#�Y����_Ă�̸(i�3���ڳ���L\�s��;��U�^��$�/T`)!�.��B�|-	�Dz�".V�n^+=<��Lm��9m������%��R#׉<�z�Vٶ��lh��>�E��5��rS0��v�z���f�|K������Qf�����`�ƺ3+�7i���$&1�#^����_�O7o���Nn�D����4bY�J*����!���;͗l+�1QV���ǟ���Ca���m��H��l9�ؘN�GG'���0�:9����[_�D�D�׉�������g?;�A^/�~���o�(Bd��<{���C�KK{c���k5�y�����g>󳟽�Ǆ��������69�Lc$�D�R�pV�Q�8�VR	VyC��n�9(iU�fKg̅�?z�t�ƾ	AQ�vW��lYL�e�'��R�?����i��л������;F�a2�B��.��f���-��P�`x-C�������(����Vz:��|2ZW�54���� �(yw��&�X�_R���q-��;�o.W��${I�����҃q�����H
\��Ƈ�~����
��w��TbI+�w����V�l�8��$��{Z$+ˁ��ʒi�:�#����A��C:c�e-'kckS��ܲ#�e�p#�P���ڐ2.�A2L�0�w�h/u@���!v����W<a�v���`���spp����������h`t�a�cu�J���J��@�b�}d��lb�h
��~k$��ӤM�]��Y�>k^�2���+Qz��\c��=ĬH�E�O��g?s�� 7lo/.��Ӎ���J�{�M���	\��ӓ�Z��)A"󅄪�����T�K�D2�q�GK1�\�\�,J����qc�)+��bΚ��a�M�p��m�Y��� z��P��"��.lZ���S��1O]�i `ۚ�z���C���l9�$���)��/���g?L����7Q�Y+�
C�pG�˕>��|���N�'V+N��ڀtrAa؅j�Ssݥ )�>Q���Ƅ�!��Ҷ���E�q�׋�B�̵�
�Z�7`��a$���>�8�n�!���s*����"%�|Їi}b��\_l5��5�
��,�A�)��wdXB^��}�L��R`���c^�EӃ��y�+�Ss7k�]Z���*!�O�
 ~�8����.>�̳��z��v����gTlA����R�R�f��)�&fP�Ecu	�{�0"�C����v�E��u���z���V΁�Bs�L���d���+o��}6;z��qh�ݭ��p�)I�����\m�Z���Z�� Xi�ei�F:˕C�R/�ʛ��֤�����	q}�����Z��eNOҧ�[K��:@2Nо�S�yD{q��a�f=1Ñ�s�8�����;9��j�Ud�tӎ��'�+�D�`����G����lr�P����Ϲ�`%����1��א�����R�j@�=U��퀸a�b� 7�R��%�ŭI1�~x�5r�ڪ�q|9ե�)���ٙ4v����
NOa��4v.�a���Z-�sg�b�'�Ƴ���D��Xm��G�>��̜'��$�I0ࠟî���p��LM3��� �D��x}��i݁I�p��\�����gމO!�+��0�wwwc8�g}�Sf��=^��՝������X���:����2�ʉ���Iu0�~ٽ�Wu��<�t�mkUH����Yq)�I܂��:b!�Ƶ����qG�qp�ӴV��@�.<tt�4L��G���b��hd�:�y�q/Y+>�`z�7��y��$)�:,��b%��-}���
q���Œ��<c p>�����@[��|}1>ryuJ������YƲt���'QE���	�g����(�{�mw*���g�� �Bn�G�4�[�Q����Y����ƞ������ҩ�1�l������j0�J��&34�U����U�7���l��W��o�gOh4�`'\M%*GL(.�)���x������PP�d���
͵�hJv��1&�R�M����<�M|��
\�m�QC-ej+v�m���aw�{��1��p^�F-�,��a�n4c]d~�6��_얀y8U�a@l���ޡ�-�4��CQrw���(r�H��|�<����s�)3��w�u%�^�=L�@~֘�H��m׾��{�� o���?��o|�?�ỻ��������BӕFٓZs�����q�����"Q���"/~�1c�&�.B`��+#
�,��c�Z��~b=�pe]����%v#>���Y���|I3�C�$�����88�> @���1R���H���YtT��
����é�2�YE�9A+�2E�UZ�xo����߁���ʜ�bMvjsQ�L��1V�r`��+ETy���5M��Z{[��u�>�vb�J��U�m�4����P'��ۍޒ֚�5V3�m?
[�X�Z�)�^���vm//��g �����}�K_��>88���K���մ1�;F���7Əhr��Whs����N�I1!�(*������DV�us��ZG&�&�ec��2)�]su)	`,�V��lQ��R|<����j%<}��`l���D[3O�Y�*�pA�����P%[۸�/�@�+�$e�|��|���X��ظ���T3�"�2E�iD�:������3Z�����c�\�C����ĉ����03�O��Vs���h}U�5Cu�*�#�a��5�-�*i���]<��B�ş(��K< �B�d��ٙ��Q>�:���-v67hl_��b�i�S(q�xe���1W�ymԀ�|(xc+b�ٔ�Jksm�}�f���3)��K��"#g���O�N������ʚ���g������~iD�<��Jō?AAE���+��r�}�F�έxX=a�$�"c�ڵ�]�q��>��[SV�sze�iƗ��Wn�����n��w�rN�q��n�ә��^��s`f�����쌆;4�|�F��ڑ�ʍ��#�֥��T8l����Ϟ=;<<��JDY�y�
#������޸s����dC�n~~>(ᜩb��J$�& ��,��8d�|ꎙioІ?�v,�H�M_�@/i3xW�Q��Dذj6���+�*Pŧ�^N18���M�\�e���r�Wו�^��ϣ�|� T�K/����_l�� l}�d�����`���@���sV��P网����-����I]��Ԋ���ȨW"=BJ?ʐ�ǡkN���9���<O"΋P�+�6�"���H\�0��r��#@��2����K����<������mb�ᣆk�b�'k�U�Z�+����a�á%�]Y��7OX�C����6l��?~^a��2���U=X��F��j]�ׯ(�K� �:x�h����rkJa�"�Tǃ�Y�bcŪ�Q�vV�^Ye��h��1�2
������Yްcie�����������"���#3�E�����Y�,�S��QiD�r}�7A�=}&�y��t�� �/],̂q�?�\Q���,QIp��QW-��r��{�.�0u��+Xx��r9_,����+mKɸOk�kޑ�>��19_	fI�mM��B�	�0���ׇ�,v��"-C\,N����|�����*�`�e�i$*�|��T�@II��RSJ>?���L�!�6�In����U���� f1���WW�ؑ�W*
�X$���t�h>_���O�˲;����M�N�ʪ�چ���YU�ew�J��E!��2��AH�沜�W�Ӷ=]�4kOzYo�����|ڟ����l� o^@�L]������s	e�yӼgy�U�T\�b�ĉv����2�ū��n1�@��[��#���j��N�	����]]�v�yޯ�f���2I�eYJ��#C���@�&/,:Ij��_�mP�PpqWc�@$F
���jI񝂮X-���՜RyԍÍzv�Nh7ZR�U��,�IO�����s���`����6���&I1Z���,�
`�Gw"��_�D!Li҇��\M(��d^�B���,�"��F�z*lc��w���H���W���rqq&D�Aʊf1e���E�{[�;��!Q	0�b�3���P"8�	e�^^��?|���>|����h5��m<�p�3[Y�,u�9������FA�9�*��P0?N3�,W���:�l�΢�!�.�&#A�j���l�.g�Ǐ��"Y6��4̗tJ�#��pj�BUz`s6$5�A�Q����Wq�,V��UlmIti�1�G��&g�,�Ĩ
�EQ.�{�<���K)WV�R��,Ty����������|l\]IL�&{U��`{{3��A/��u�d�_���}~~.�Z�MC�<�C����K�����P����Ψ�RV�P����k��vz,�:ΙH��7E0�Z*cc�K���8�%L%���	�_5v�dm�^�zy|ģ-{U�Đ9�1�w-�G��Syv���7ݢ@� �¨�w�m\^\Dq��g��jvUL.f��*��>�w��gzy_�_��:����@�RcX��5�t$��e�j���#�I���!�����?���ח^z�O��O�#�ǋ
G��a��� ��z 2�}U�"��C���M&�֖��FHe��WY��th�8��!������a�}oGѴ���~ºEZ-2m%�e
�a�䉰�ONONO�q� W麬�$˃����M�SVb�*?���5�a������mZ�[�+��(�a�H�C'�.C�M�kަ��
�Y�p�c!�E/*k��h��Hj��,��Ly���?1_���Q��R)����ؒП��'�XK�`���t����4�N{�����^
�R�5r�J�H�D҅<�&�\w��w�|1Ƕ��/>{���'�T�\ڱ�C�Qy-I�p�ֆ���-Pjd�d�:�e`љʊ���}�t4?���`����;�@@����
B~=1���ŕz:��+�>Ӹ��FyևX�5&�ZU����r:��#�"�����ˍZ.��M��)aY՟r�����Z.��tG���3����|
Y:���l�(�.���}Z�8Q�G��?~)!	��`0ހ��~�ӟ�?����l�$�_]1Í�!��"[�Z���������E��~4�99���:��4zLkV"2�����Bk�Wޔ���S0� l�o���l.l����_N��6^YI���g'��WO/&8_ �J�Z���ʹ������^{c#��ڥB�m��$���2Kg6�8P���pۄ
$d���h=��b-���|*#����7���B���E�Bf���K�G�so���&ގ��4{0c��P0K�
����.SZ��U�O��(MR���!]?�\bR[�����Cn��j����T�0���g9��p,8�UY��#P������X<�\��9UP0�,�IMlm���@��\�hu�󥅐�fG,
q�5ֳ�q�r�`� �T���2i]\]����˜LN��ٯA|jZ��Ό-��I{�û��׸����Yr��b�1bJ��Z�ʫ
�򎶚,��_!�ⳳ���hb:��/.N��Q?��L�s9n��4�e��j���|F3��E{�T���W�?{�H����`���q��hC�xu�I՚H`�I��K�k��2�r����м+U�I��n��RG!Nt�i�L��ڳV�̵��9|[��>�s��s�]���+�)O#S���P��@B0q �V�I:Zqֆ>�SQg[�h��B���Ze�������,d��\=��^J�u��(FAL%X�펩I]͢p�����^�ֽ�:TvE	ՙj,�[*�/`\5�AR�L'օs$�6�lM&8d�J��0�D��bRo�0��)��!c�i�Fa�������:��:�T��c��'��W��`v����3,+
����5^�� {�����)�����|č�1�����	.=g�mo�J/�]vD#v�����khqf	NiM{�$����]P��CWU�A�S�8'D��Ů�s�����k��64 ����2Q7{���h��g=�WY�X��(jk=�����p4�^ђ`*�/7S�+krr9�+]��q7���|���ڕ'�����ȝ�pq��ςn�.�CkÙ�P�$�4�>a���aP�G���X�5�a�*�̟�P�d���\S��[W?N����@f�5>T��% V	f�j�U�}pY\I�� �Y)��$��`ؔ�VO����ʅ6w���T���.�	�����~�4<Z=|�X���@Y
kM�ժ:���!f�U��	h�ݓj��_{��<��w��q�H'k*Q�*6��{�3�Æ�7^��k�+o�e�ŵ�v��d�V`��Aދ��(����2����-m:���r��ck�/璯��bs��Z�|gH�k�bZ������*���r�\���[ŉ�]�D��R⤇�P��b>����F��3n]f_CcY��~���&�ݞT�o�J��*�A��r))���ָ_[��g18\�u�U�{؆~����M�V�|�-���ۻ���$Ѡ,+�K�r�{��Y������$������/O��n�D�3�&��Ѿ�=�*�W�>��9Jjòٖ�n��XC�P��O�<y����	֠����Lx��5Zg�W��GLS9Z09Z�vu��AS#�+�je$e�5�y��6��A�cNaNӹ�v�^Ϛ�,�b�T�ͭ�k��9ᰍ��{_�?\�'0\<���j#t�Iz��Rɢ�X��[�]E)�V����|[[�o�������e�(�����İo�y>zDg���LV5� �f�����$��Pn��NK�MR�f�2H�Y�ZFX�pU���v2Ţ`J1����cc�0bu��.GT5��t�Ej�$2�7�
F�1(	jv��R�~��7���뇇�����}�	F�gw]��v�p3���n�9˙��'�\|���%��^��^���H�c�)f��	��V:��Zx�W���j)��Ƙc�'�={F�P$�Ja �������w��}㋯cK/�y��K�$�^�{-��s��a��z!�ϯ�&B�F��K�A��4�6���(i�J[�V[����Kk�㤺z��*�k�B[|����U��
�|�kg�'�E��0��Q9	�TeW��,��X����^�|w���=R��	��2k�I!YM�,�
.��0�A2���=cTq=F�2g{�V��!��?�T�֗K����quQt{&;+(���=��������o��- ��@:]����Rd�M���+���n�����߼�/���|f���#�����fj_����<���?}����.����E|��DhaSh0�L�5**���ꫂ�k$;�� ��|s��b�+��;7áa��5?ћ�M���o�������E³���=u��������/V�9��@�;��������g.Mr��V�`�3k���ۄ���	��dR�)
R�7���(�Z�&w��Ôr��y�㹆+%�rw^�K>V��А#�Z��,`�0��v�ί?Q�Z�n��3���j�O'���*m��Gf^���'����� �c���K�q�����'�L.�W�[h�)U'�dꌁ]���	�q��WM����
l��r��Mf������BO�G��Pf-�K·2�W�֘:����ۿ}�so0qȕJ�kۃ+�h�Ļw�?.<=��������B_k��ַN}tF���[�ަ�ɢ�#O��V"I�]���Gq������������I;>>ƿ8M����c9<��櫋�J�-6�������A�Űy��V�L	�h�Dތ�#��U�&Q������K��G�{謷������4`��K3p���q��O�u�B�(��"̜�am|h�8D��rA�7B��E���/�l��}��[ס��It��r�Ι�>:�
T���J�X;�+��+�! ��	��Iȱȳd�8i���r|���W���+P�g�@G|�IN���Fo�hѻ��Z�/�;�G`�9|׾Z����h����1D{&�ڨ���ظ��҆t�i�u�5�``E��ZG��@[�=�]���C ���z��+G^��z�N�#2|a�|� 5*Y��p��J簽��>H�W�²��5,h8��6c�bב󺜙(���~]��4֫�֕�:�ǈ�qܖk�o#���{ڼ����Zl��^�'��!���1XYd�qif/��p�nݼ	��?���};c.�N�%��N��4���Wl @@�T��hL�KG[{	�Z����6���*ɭ&�6=D�k�t
ZD����d�u�gZ�LS�Zd��+�;��Ғ�Q��t�H�;<��Ue��'�Nȳ���A%���t�����I�b-���H�{VTG�����3�Q�n`�%a�����Y�m�U&8W��ӟ{���v`'��RY��!�<de	���3H<��d����!�N;p4���sO����7�7��+l'U�V�Ĺ���\��7��d�4FI.j�O����8p]G�_��[�L�*�ݢ���\hs��i,4���4�_Y^^��<}���㋋�M��M��DhS0߅v��J-Ԧ�@n�V���H�v�����ǟ�]�,+(~�(Q�w�PUl�T-�8lֳ�r+�;?����¼��IS���=�5���B�	Ñnc�*�9zGm�&�
$��S����b�	ՠ�岥�j�k��Q<��9�u�hwgGH�
�_���ポ������;j��ҋS��BXKT�3f�����������)N�/����f猈J�qM˫��_�%OG��O�g7L�b��F�ۆ�>��ĸ��N����y9���lv5_�$V Cݩ�U3ʠ�%c�Cc7�?88Tm�鬓��~�j��X;����ڀ�j��yow����n�M�G�x8Hc\yyuu�ZH�K�� �ͳ�m���k��8)�o�蟰�p�=��� b��ǹ���ey�O�S���d�e�\��niMVg�V��Mvc� Đ����L%��XX��>��勋_|�����+8	�d�jV���l����
[,ˤPt<YoJ!~�;�v���N�p�X*���HHgo���O��d����f S��H�0E*���SH����Q,U$�x<ܙ���
�~쪶�Ƀ�C�JB���t����{z4���Q�3(DB�*{}�&��%�pu=�Ɩؐ�2�ȱ^�ih;�V0��E���pk�������Xh{�'�#��u����␓�<��Ph(��RF2NB.#Eʐ�Zw,�0�0MM�Y���xbn:T�S+,NT�zr�$O�b?�9�+2�4]^/N__J���4�����6��>ȳѭ{C��j�qL��h��)������Q�x��\�ESJnW����|����?���I��/������d���τ��7�X�]7Q/�bw ����o����.���?���>�E�]�R� JzT�4Zj�{��J��WM�`�D���֨lZw�<Jw,o p�Ƈ�J#�p9������>���S�\��X����V6C�$�+�;��Y�V�G�Ct�2�yg&7z����Ԉ�$52�I+*��[��ݻ)�G�� ����D{�Æ�G��
�CE1��j�	d(�C�-QZ�#��ۮ��`�(t=�ܭ.��op���H�oƦg����s\���J�d�����l���������~��>��ۚ�̗��E�,�9�bK������5��|g��`�vV2�M��4���'�)��Td���?��W�Ō/E����:?������w�}p����~�q0�!{O٢i�:�u|���N����?+X>��r|ڮ����ק�����������Aee���\�6���`�:�Τ"-p�˼>=��ZvS��p���C��_�������,�4����k���Z�i��p*=$�����b�`��Ǿ46ZpNNk��j���GCc >(�߼��s�������Ƿ����{��Z�	���S�$� 뀑����>�i�rXK����*� D���ϟ����@�2��9::��9�8��V$���ĥd@��,�Q��	Q!J���h�����5	�����"Z�LNЋԸ9�p҈�0쏍�~u�2
��/N��d�\8�w�V�H�ۗU�X�u<��oE�%�p���;��	��T��fY�!��b�æ�ق9w��̈3��8����f�x�դB��i�1n��|W�ߨ�S��M�I�+)�1L��n�Fv�ɔ �^~���U�baGc}5�u��,��N_���sR��(m�\\[����ST�A��Q�ʰ5�R0Թ�yp��נ56��
h+�W�%q�g��V�Q���|����O�%���?����d:�?;�(�����/�����>��3%�y�����o�>:ك�O�hwwG��$�wŐRB[��.^j�'O���>�Ta�2-Z�yG[�蝢���Q�s_*���gk4�;6��Β_,���������bL�o-�%)�^��O��p�T�=S��#9�/A�v����k+j�b_�!m�;�J%��֙�u�A�7ˠ߰*q\�������X�<���3-Zw�]%B��+v3_4*���FUA��IQ�[L��k�NܦA�U=X��A=K�[ܳ:2n8.c�L3��<>%Xr!��J���!cy�0ǽA�`8�qFV��ph55��;�~IG]QT��!*4��YK5�JN�\0�NO��m��X�+%�XV�u��T+�yI7n^��1�بL�m��$j�k"ЉV7��I,�"a{8#�gF�"��q���X0�fg�c�~ц������-X p��կ��_�5%���S��*/4�ZW��@y�{HDS�q�&e�>�SR�v���]�X�
�=dB����ʸD�f�6fHH��v-�d�6�OY�F>v�;�%�k{��V�c���˵,���,q^3�BUS.u�k��MŦo}J4��{bl��R�{��/��� HR�lЀ���Xh�X���_<y��)T���+�NӀU���T�g*��6�zjkiZ��P�������77Z�ݙrK�[��4Q̑L��m���gX2o�Q2s#�d��	p������#��~�EL�L��z�����i��D�5����M1���q$<��wTZp�XJ9�[����N��q3S���f�W���#ǭ�t�O"6�/�n�����uuu�����P��I���->fC��Ι�&�/=�.�bì�s�0�H�g;����o:��+�Ctƍ�ܸ��v�����ۘ�$W���!bH
4��6N��.���{��5����q#�b=�V��9<<$��Fgl�Fn>��Lɶi25���U_Ӹ�~�"_0"b���4���l�+�n�]-4�Q`2[���-�e փ�4M[�Cܨ�!��жσ�r9��b\�]�-�Ӯ��\
w?�;Z�!3�;w�i�ӈ]a�_]!�J�1��R��s-��!��f5����>!��H&.��d����J��b�k���VE�<8�� Y�p��޽{����RP>%j�i O��'''D�FFOU2P˒��6͸�T�sX\vqq�Z�O��4��4�i�5	�$�27����n<s��?�X��);Ͼ|��l�Ǐ���>hB$.7m)���~'׼4T�f���D��ck�s5�/?��|������T����_��_A&ϧfޑ�������X�'��?�(wv��F�A���"2&��@yb�zΒ�<���'-�f;��z-b��I)�Z��Z-� Q%��9�n?���C��Z&St�ħ�ϒBT�Ϛ�� <�|G� N�,�E6��X]��Q��c�`>C���kc����>(O���DgDNAq�ꌒ���;�	���WyK������b�!N.����u����{{{w�����J�-p��b@�J����h �	UgXq��e�Q�QQ31I~�п5� ��u�.�_!T�޽yc����AG!O-�:�H�c!�-��Mu��ѣ��S���Ј`�?y�W8���I��b�xF��[���P"�*��?�_�w~g2�vD�=��o犱��˾���!K��F<�z_���9l�v�0Y���-wv=�Q�%�Zr#������Ç���?&&W�a�e���q�9LA.\�����-s���~���{����b�+DƵ�J��k%��×7� f�c�UĲ޿{kR�F쎾0K�WW�1o�`�[�/uk�5:��%���/�����S^р)҄N=
�r|l{0Zz��)ckb^l��,.�����]�5,�
�Hit���Z��@�1��<\r�R�d��Xy��B�3�Wc��TvL9��Ʌ>�N��ÿ�q?T�ًz��3��F�ӥ���N���k#�������`e�#gDX��.4#y�%J�2�9�&FM�M�(��b�Y����(�㢇�c�'�U��4L'�4Ź��=��j-���vjm�k�8>&=N���H��+8�B�r#���O]%§\	��0/�>�x޼�ViB`z~�_~��/�������W,���{X�������P��`Ġ9�~*k�y�"�O�`�^��+�)װ��ӧ�g򰾚QcD���Y����AY�y��Y����S&����$�\�s���v��,c�P>PKR^�x�#�\b7hs���Y'�<��F�^�w(��[�k�Ƿ��)��+�EX�	5��k)�3-!V'D� �|Y�34��IRϒ`�V�T�z�֋POڮ���wi`�nFU��b|o��X'�B%f $���9�`�7C����5�,�	!���Z��f��⃮[Tы��v_B��X��k�>je&�ȃ��[���p��x���iЈ�E2P�����i�Ѩ�����V:ߚXmuc�=U!-W-,�`��/�\�׻������p=ta��C]O��q����$~ 47y:-��E�-�����N��kYb�6�"+[ev���F1
R(��D���/����!��f�:�\W/�?4X+krO;���і��U���Ԛl��ʌ�1"tY�#I�RkR`��oڪl�M\/��]HDqM�2�1����0:|�v�M�.7��Y���գRv\����R�#S$83����r��#P�i�
��x4�Z����0u����vR�EY����O>�����J|x�J�T@��h2?9���C�UN��G��4�/����	W����ZZo0g�e�=[;�C�T���R�B��S�a
���f�������4��p\�W��*j�E��ۯ�z>��{�!������_���ELWm��ǣ���r�A�m�
/�x�o�b���{�e�aX0���V:�6�P��WUQ=�	���2�y�f��ٳgB&�3��L��7�s�bUM�H�='�㳗/_}��)�t�˔M�W�e��u�Q2��D�)
l]m��isD�mۗZM�?��T/��,zB�mbl!�@��Dl֕��8>�� r�U�����ܾw����!&>�t�$Έ�8:8��w*�O��'T)�˛7o._�|�F)��j�T7�'�1���z�L��U/h�\���}�W{�w��J��k�-sJg�4��b'>I��19�Z�Z�(�EW7B�y	����gU%+��P-W�Ujwo��<�4�ȅr~�U��,�!����zI�˯j��/F�J��JUIX���SK��(�VWg�U�]�i$n�"Z��ǭ���5�`M�TI:��N͂ ��;�,x�&qI*-���S%�/+���ݩt�іD��D�ˍ�7G�B�Q�z[e2�]5�-��u�ヮa႖�\��>i�ﺳLa0fT��h�:C�'���F�H	Q����;��$��q��/yppt��1�O�����f
%��U�t��1"�̿�>ף�V�"Z;��xuz�/��ׯ����G�q�qN�uus5{��\�VH���X`A��`��ٳ��
��p {�ֺ�[�:G��x2��|��Gâ��?��;�o���������[H��)�#<R�ۆ�j@�ާO����/��I^���zyhZ��:|�]�m�&�j+Ď�� �lq��Kq�$�d$a+-+V6���(��~2�����H�����+װ���ث��R��i}}�
���<p�!���^���T��jk�N�p#�O���%�#W�E��P�S�JD�}�l��DFۦ:Y�=�b�X�ޔi#cbmF�,NG�G�s1������z��r�*�:�f����/�$p��y7m0W*������gk5:���B}i9��h�-k#���g��2s[��s��}�j�i�����֥}��/�>F�~�m~�N�K-�,� �ů��Յ�����L:'(��*_&���^�~��a�[��՚u�~����;��"-C@i�m�5&��׬[zI��77� ����j���_�nƚqâ���Ҙ`̖L�Y�|!�H�&&���\�@�-���?"Kɦ���u��5�i �Q�p�`�1���G8t��C_�����f&5��R�b�+)e��[��|L��������j#8X�W�0V����lgD�VP$1}�f�xQ�]A��N������,4{p�z��'#Jl	�/���(�k6��Ʈ�l�fA0��V#ᄎ�_É���t��a�.�̭!�x`�w�����	X�m���y`�{؞�n���G)��>� ��Gnl}�Z��>Q��ߢ��c@J&��>fbp����W�?1�+!�m�Z�؊ӎ/2�Ës�$d�@Z���;��\N���1̆m��2�(���Vd�pV���bh������T������������w�_̍��^��k�q�!3�  ��IDATQ��	Q4���������>��c|e��g�7����jB��\��I��x
��̯��=����o�K�zK����t��1W��CX}��֔$���k��ѭ#�d��s�x��#�Ar�q�ImSe�G�0\��/F�W�Se�q,RF����=�#E��}j����p>o[26DN�qY\��t��n���4jD�kd	C̍-�������"��[�"��s��K ��`��W=w�l�ɄA��j�}Ԩ��@+S�U�m7tB|�47���5`<TSDe
�e��icݸxB�Ų��2���@�����
��������ު`�?<�}�	W������(hg���hkc�#	k�{!��,2UM^�I��`�S&6=�mle��>�UVa�������EftT!cF���*��.�=�m��������Ȱ��_�$��Z��`�0%�@E}i,NdU�m//�3^���G��Á�$L`k��>f�cit��뮳<@j�2��d7F�ˀ���~
A�o��qxxM)��,�s�ƆK͵��2�oz�եU�0�Ln��m��au�o���J��=��M^��+jt����#aͷ���O��Bu&���¬�>?f %_z�i��ݛxF����s]e� �W`��ݕzBu�a>i���\C���7��댉��g��$h�ޱ�b�̽��
�j�Ն6blX��ue���-V��:�k��o�:דK��h��&}��	M��t�3���O?�ȃ�n}_#,��N)8�Zx����\�3J���� LJce�hˊ\xG���;�{�g��("��g\5�%K9�J���̷�������#��i��r̡&���bZ���j#(���Q���3��\I�6���ڲ�%�/�U�h,o#������`�95���=v�� ��<؎yJ����l|���0)4�<��<�1·b�{�|l����t�hIh2�ҳFPd�J0d}#o|ssra�a��7�ܹs��ݩB$���Q'�;ִEԔ�������O�>��JIb�ONN�='��jY��P"�Q8I'r#<���
=�al~,7V`/U��i��a��l�T��9��֠�����kU=�^�~H���β�(`��-�s1�ʮN�\R�@_Gx��J�0~*����u�//)�e���ܿ'�$]:��t=z
:<�6���i;q���6;ŷ���r��e�p�������z�S�ɳ4^�RP��yb�P�]��d<�"j��� �1�aќ �:�i�qMT�r�"ϴ�؛L�>��3E�,g�I��%�i�..I�HVp:�żaM���/9k��@uQ�c�a��@n	�NUpE���ٳg|�!�h]��F
6�H��o�7o��_>>��Q���?������KQp�0Ɍ�8/4���,SN�`h1Zq~~�_��o��o�������~��`?��E!�d$EC
bC0������:10��z��r5C����3�N��
&G0Z��P:�;MG=��R�P˝5t��4���b�Ѫpz(�q,���FN��gY=��굧�;�yqZ� ���3Y��T{�s>iEP ��+^���4:Nޅ'���vZ����Ͱ��G�Z�0��M�!鵶��B�#����Pz�瓧����bپ~���Ç"�ce�/�eu̅�=
g�����V�ΑJ5���FB�K�j%��9��ﱚ��;v�5��"#��Ҵ�B��
"�N����JoS!<լ��(�u���Y"��z�/�����v|f�3��6y�)��ΕI0������Ƃ�����J1��~bn�+����<;�zx��G"�|�ݨA�4 [�^�"����+��d��7�b��>x�����d#U�wΗbtV�V[�5��'%���B���h?˞��3�ê ��R`�`�D�j_ e<�S�8Ġ ����^����5�}��ixZ&�!�[�%�wL76Dfá�S~���3��&����ԗ�̤<i�*?	 $u]g|m��X��H�5�tF����
*��@O�>#�Z'=l����'6�4����Ā�4xX�ËFMӔ���ə�R1��
�uj���R�����S�ۑ���� E�|sd��A���(Y�@�0IzU�]�I�=�܇P�x��D���E���6���Krð�%�q�Wn~
�.����`��Nw�� �A�-�Ǉp�@�j�炚���/�ވ�^KO�4�)���0&�,<8�n�Rl�|�$�@r�Kaok�"BZC�㟬��w��b`,Ə���5F>�+$u[�9�"�$�C�؃"�(�V�,�:����0�H?�a�4�?�P��D����aP�]J���dkL��Bg�3m��ǈ����u��A'[:�Xm�0H\ޤ�������꾄	;az�F�k፻�P8t"M�U%���D���|Oj�W�5�9`+���Z;�(㕷ݓTB]��c�ߘҕO��k�4��\�Q<�d�U0u"bA�GV���aAˆ'	/DR#G��X���W�Y@�� b���Q2���U�9�(�6>��҄�Ex�o��
_�����6	z�Ƅs��CeNVML!)j�Q���4�v��526�~Oh�����ثE	#Nx�
������|��j�;�ڄF�kx^�j+�M��ںGM&,����b�N�CB��_�-���?�)
�M�������X��j��/Օ� �&p��ք� "�#?��
ᵎ��o'B�� �tv<ό.1wD��X��[q�w�PTn��a�CV_��0m�2O��h���0/z��)*�/A�$ھP|�V���w��&+R��j3�]�iw��jJ���a��n�X�k& �ۇIԀ(
_XJK=�^��T�B
����j,H����;~�l�7��O?{�����w�G^��1�L$~���N�1��+��{�}����=� �̺aBlD'�!ߓ4(Fպ��H8'a��Iմ��0��'�L��y�9��R�Y�h
�D��$V��׫e����<����bܝj-v�X���tt��	V3/d
m(,��1K�d�i�0�D�� �3�gY-t��o7��{���LT����v�����S���͞�X4�Ԡ��(��m��%ͻX��gڍ�TښD?J� ��Xo�1��uO��ﭦ�	u�c}rr��Ě��������s�j���>޽1�{
H�S�1`1˺ �^�H
\rƭ.Ep���8uup)�0�o����[W>�'�;��1�ϓb��O�<���r��G�F�`?W/N�Q�4R�V�Y�c�ƺZ�v
��ȍ&cwq~vq�)��J!Sת��Ӯ�˧"o��d�W�
�����i`��T���X�����*�(���3�*�"�%��J\�%��s��b_
<ctRQ�����t3tm,yh.G�=:E����=�?*w�}\�oC`>��@	J���zX2l]L�--���R��´5�)���V�x�/�j9� 6�%����{��ճUŖ�?���[�����8S�`(x�]5�!��Y�����ݹ����ttC�J�f�D�c��� �TK�Z!�����ŮX?{�zS�~1��y8d�J(��b���{'wpz15�������ˋ��(�R�f�vć#�E8��TV���2y�h!��$ ����������_��WBЁ�k�
'�^_�����sP��V)���G4���8����&[|0 �^�Ř�I�p������	���k���g��)	��MDt`b�N�)$���<\31�*3:���u������(����Ǡ���Р�G���x���{]�BH���*�_�b3<�m|}sI��(BUWe�NZ�ݬz����饑/%Qm�N��ZG�y�z��bG8��Ó8==~����3�����W��E۴z�.�A�E���8 ��/�����i�":r��
��2��	[�;Ȋ�oy<~eR>;;�}(f���I�_����Z4u)��4],g�_>Sp�Dr�&�I&��������=!�J{�Px����j�,�q���Ը	HcZ��wjN�W�: y�Y��';;��C�+B\�/r��O�<��F&� ���X \���/2))��8	��q�¸L��\qY�cf9���1tx^l�AQ���,W�U5��u#O-�!ee{ik�c��:R�P�dڛV�F(\�&�����+�.���s�#L�ׁ<O�޼��7�� b�֑��p�X�J�����	�VP�^�-��S�9�˙�O��R����u�z\~dE �:2�޺�hh&�#���ջ�4�%�����Ŕbl����.���81kE�U�/r�8B�z�Kv�M��=��dܣ/�tņ��[ݐ9�r�=N�3�ì�������;3i�j N�ϯ7>4[Ɲ��#h+2c�hz\OT7X ��M�p�N��q�w�	���v�55-��O]	8�5۬��N�Խ|��ٳg8wu�~���?��?\^_��6�h�\d���օ�~}zzu]Ca��?:<>������ġ�w��ׯε#_�,װ+V����R�=�L�+&���I�d8����"ߔ#6.�l��W����usY�Z4��i�Ū,FC���`JC[]5<�/��R�"ܾ��;Pvx�FZ�����NK��ŧ��$g�G0<D�B4���[ɭ<(h+5�[��@?���'���_LM�X.�N��2�cgw���"�	�Q�$y<��R�e2-�R�`�7M�	�{�i"6�M	����u~��D���m֘,�H����Gg����b
����gu�Ӎ�<��z����B;Bc��O��],=.��pi�W��U;�) $##��@U��x�O���aֺ/��V�,�َQ��ϾI�N�n�D�^���,)B���d�ms��YB[{;hEU[�i�0U$f�8����Y��e�v���k<�Ym��ֳz���8G�n�Z4R܇8:O-W2yqA#rr��*�5"z�T�j��":�J�L��I���g��q�`U��/iEXl,����^�
jMf�V�{� ����{����QX+����q#hI@A�~���'�Ks�B�V8Ǿ{Nw]i��$��6���>I��DVm�1�Hv&����m��&���É��JR|R:*��Km���J�L��4n������1x:F�T&��:��΍�&���^<�\����t'�@�5���P G���G��߅N�o�9�	z�����U�}%BB�'-�RұLpg痯���;�Q&�����DUH @�}"�7F�v��Ra�������ޮ��$LE:~L��Tr��?
~s�3/V���5I��&�.UTz�Ӻ���������իP��)Ð�ε7CrR�&�Ms3����Xa�K�T��������&9����9�]�3�h�1��\� �W�褰�(�,S�77�1'�H�F��zj��Ј#��nx>a�3���*��t�kq��`9�1#�����4~��H5�A��L<�b!�Sês�q
��a��=��R��r����U�8�3_(XO�I�߉
	o��KݺԦ���Z>�e��N�aw�6��q��.��q;�!d�W	��<�N���P$� �����J�<��	��қK	�,��rG =��gB�zuu	k{�`��rT���R�iFB��H��5��X|�o����p�.��'�&R�Ga�H@G��|.r Lv�x��k	��I̡
���4C�&��L��%�Q��W<�B2�� �}:�ΧF���B`"���V���vN�,d�4 _�j��Ӡ{��%YC����j��/�x� ���0ҧŢƺ3)F @�X��?}���ܥ�2�$ϴ^CG7��\�"ʋ�(
����קw���G?Թ|���x�~��rg5Q��aF����!b-��x���.��4]��A$�mⱨ�ޥ�M�٦n�"a3J
��rӵbZ7Z1�#�� �D�I�U�����0�Ę"P"�hzz��ڠ��eIul�4~F��tN�-jP+[Y���\f	;Vp��������� ���?�SM#�5D�/I^�mc�8$q���"zpQ�(�e��:��k����1쇫��B�%��u0]�U��ǡ3VkN׷�e��p��wA���p�#�#\
6�IÍ�I�7�����I�aPx:��}y�p9�k̙֣�����th��ij���o��D_�P`���\�<��Il���3�NLwB���zcfej��N�w2Q�$%�h�n�bk�"K5Ɨ��,�ͫW�0��&��f��P��(v]�N��\��W���kD�a&�L��m�;V�\_��6/�P0���[�.���/ʺ)�[[<�۔+/zϗfToǄ���� ��O��"@�Z�Y�w7	��\���}�_��J�d�Aƶq>�}L[.�bL�	|��Dm=��{B���Ǆ"���F�P֑u��]ʳ&�`8"Y�*�	��I|4��/&��}(�ˀ�\���·�ܧ�N=ʸs�r%X3�䃔E��j�PsүL�+Y��A#�34�;�!�n�1�Uȑt`6��!�Ǉq����LT��;�Ҽ~�+���ŏG��W0�2cta
g!��Z�Q��,�l�n����8ͪH�p���ӟ��g��������?��e��Ŝ⢮+�X?~��!����?d�Ę��C&�0���14�{�AZk�
�3W~�X��!}�(b�+����ח��^��A�`���[�N�\�Gb*�$Wb���O���!l�	��ҋ}�C$�6F,T��s#�� ^^�%u�т���'OI��*%W֯G�&��T��wq�,r�,��6�)�ť��1s�cN=���t^�b��UzjQ&��m��u[!F
�autE,�[�j�C��M��ΌF!�u�*�H�(syܰ���RJ2]�D��VqS���>m�����㓱�7��1m'�I����g�H���JoV�?�1C����s%���2	C�8��5
l��ުʹ�2��(ɇ
���Gr&��^��w�娏�u6�����v��A�}*�9�Y��@Yl�b�\]���O���^�o��Fu[�]�r~j�����Zf��($��ƙ��V��r�^�,��/ز6�	��J7���ĉ�2TYk��\�L�d�5�k{�Ɨ�%Q
�[�M���5 $��]1�N�tZ���w�I�THTY-�=�?��n�V��Y"��=3��k�]d��g��e�`RI�E>�:�[�/��ͣG��jٖ�A�Ϟ�4٩�3i�u��f皲�S3H3aX�3��&��*I��/+�z�j`B��5�V֭v4n�KV��S��^��z�Y��˅D�E�����j�'_�4&LG�r��L`�$�-��7��x8��aҟ=������T�k1���(gPp�M[{����j\-�%���'�j�!U��/������b�pp||�<z54D$��+�|��,�M6U��٩�G�O�ղ����f���QS qG���"͓4׌}T�֋<��]KVsZj1��ngo|5[���}���WLU�A�A���<[ΆC�@���a|<g��N�2��`Q3��?���c�����z0��F]�i]��,��˟�5�E�J�f�)��j�a�;�4�rĞ!���yQ���Fo�/�c���2K�45
�X��F$�+P����%7�L��/�����5��'U�Π��3�H�ϝ =/�Η��r>Ǒ���xzxP(���`�U�R4� �֭��B�sG�d:=�)�+»�PMFcbD�dBM(M&�v�S�l�7g���t�h6�z���2�5��ZțH�ۀ.璣�����6�L�=n��'<��fۓ:�쇕�3�t��]�V�7˕���x�Y.�u:,�;c8!-�U�i��g��*n��ex(�S�)�ء{���]ݮRل�u� j�&�v��C:BD���z�t�l��P����o��c��w��I֫&���	�ϖ�F�9��¦�;>��y���1�"���=�5ef�n$�����A1�i'��%�R�R)p���I�B`�p���ܹ7p��,�k(�b8���٤���u'���T�s)��c>�k.ܮ��W48B������IF��Օ�(���GW7b+/��:���.�Iݵ���+�p�r>��Y#9��x���q�8��`��&�� w�����ܻ��xN%x;ሺ`U��,��(��A�
	fL�;i�=R��Ce���� x8Ί���e�YC嗔>Q�O��uבѾ�\��C�P�f�H9x3-Vj����H	s��Y����n�:���rM
���f7"��\��o�U���M�$� o��D��Fr�\�2����}��ד��G�Z�a�=z����,�v�(�wtxx8��[�t�u�]F�f�o���v]���c�L1�w�+6.����e�b?1Q�8�S�;i��m�""w��+��`4�x��Q���cd�Q���=::�R��b��6��*cO�Dr�ZH�)�v7�Yh����l�P��	L�-cX��1�F��bk�7����
Y�k�)/���6�dʶ��z���ԄN��8A\��c��]�����������<ٴU��d<����Av���.7-�	pc�r��Cx��X#�J�ꅾ�p𵎌a�hw�\)K�8���w��;�'|&�j�9�����z.4d��T��n&Z��f`K?�&�;�iS՗�N���$9::�?�g�D]�Nhݮ$�� ���5�~҉��I\aqsys��a5���u �1��|�9��{�{���*	�����X�Z̮"r&ԊT����/n��w&�ԛM.���z�j-�KYMX����S��%�2�e~��� � }wv%����*X���C��b��fP$����"R�at�p#�/�pe%,Ts����9�y�Y&3p����fnB�[Ǔ���W��P�Lt��Yl�d��X⸩�����>{q����}�{X܃�C�F���>�Gd������x�*�n��b�I����҈b��KLh��Ya�/���Po�|���������RV�Xy�����}�Ӽ��a��U�`�UaY��LH(���������CtMF�i�U^�E���ؖP�𘰵+'ӛ����\۬3�|����a�:�{]-Vq�@!��{���Ĺ�6�6��'�=�Jpy߻)$JE'��gw�n�N�P��k�0��sg���T/$q��T�l���T��H4�p��K<��X�D�1T2��]A� �]��<�D��n��=|�%���7�/��RAE3��x*i	���e��թ{%n�l6W��Y�:�^eS�bdZ���/�1��N�E��]3Ɨ��A(���w���j�������a%��]+g���fq�͏����0"_:ꈠ���MzO��@҆Hmf���"sY1,�>�/�p���U{���xL���D/m`E^�lq�YU����YY��2�%�;#���'�JAU�ɦ���d��j��;�X6���Q�Z[��؄�V3^Ϙ	��:=��p@��V\�������G��x���m"Ȁ	�ϣ�����x���q�pp��.�Dg�	� Vǧ���vO��i����ڳ���L"JW����{��xw�;�=� I6��V��T�x��{�.�ä�L���ȒRK`7�ש�M��S�+�z�d��'�:
�e5@�&���j(�GIG�ɐ:��\�"#k���B�-�6"�b�pH�����x���N���y5�����^�Q.�~ ��3��� Ǌj�(<��ц:�
s�t#�V��F]1��N$�̺���!�]��$
f�k�m4a�d!b��X@cޏ�����=��*vU��!V:�&Z�E�z	�&�q�{�U��.��}���6��q��½��~]9#�k�f����P)����>�'{4�X���Ji�}����[Ĉ��>
���$�
�V<�ܵ~�HI��]�	g�m���!�w�Ty��YҠ���!W�Z1���\���Cbm�B�",=�c�r�m��d��e,���$�y�Ws u��5����E.}�>c0�QA�⇒6��@�D�>t�(������	��8��G���O��GF~o���V ���F��85JDn�R��jO�B,�8*�j2Ճ�����P�	��v��j��ܩlH��M�����ڞO�u �
�|�2]���[
񾝖!�nk1�Ћ����艣�|�G��O:C��y�p�T*�j�z����-��S�\=��=���I0�%Q~By�饢8"�	6�V�X���-�eiLR���R�8(�T o�h�%�7S��n@���� (-h�u
鷐u��`i�fN1LK��f�M�(�c����?��O�:��u$րY� ^��p�v$`yl�u�LT��kCXaSX�������"C��>F��3����QN�	�-�x��m�]��Z����B�H�$w}-�$ε�y��%K-��	!�
���
��PL��=�]�8Ovw#��'�>D�5�*c�2�ȸSY�Z'尩4�pE��U��~D_κ2aN��U�h{va=��>H8������x��z��Yz*U�5ؐu�8��1�c��#CD�8غ+��V�\�F��'�&ߵ�Z4������%�|y5W̚�Y�˵���`f+�')��ey�S�x�k+��}vrr�+�9{���"�g�/c8`|GZZ�>���O�v�� P�P4�qf���?::��o���� ؁9H�7Y�R(Ɩ+���|���5�43�|
O��0��&������"��4�x��p�3��K�OMۤ<5�9#���MXխ�AZv(�L�!ׄ�?�qֱK�o0*2Mu������hGi�c�%Ԫ�t�'j�-�����D��l+y;�����썥����ۡ4sa�������ה��K}b_YMp8 �!�F��'�̓�d�IS��Uc����'��W��6^,&�7ؠ�֭[,dY�k}�����u$x�3s||�)^�� w$��)3)���u��x��L���=IF���{�\.�O�<��]i�Y��@���L�&������'�1��=|�O���z��N����FlKc<ԑ6U`�$]�ȶ<���=aވ�N��֨�(E�W"X#��S�1k=&Ζ�0�)[@�a����[����*�W�\�z�8�|b��dI��vU�]�XM��J�����?���|�'�׃zH=��?���^�F��;w0��/�PX��G�da$�f�Y��i3b�qK�~;Ɖ����׻��{�� ��D8��Pk2��4����<6r4C�5� ^~8�A����-����S�qKS��c��"�tSH��fS��?��׾����zw�P1���\���?8��hE��M��J�1�zDS��ȣ�L��������U���%_���Ò�co*��ߜ�����ϓdb#���o~�$��2=����y�$KkE�ƞG^J��=���D����21h:":�4=��_k���
��-1�;wn�v"����d�tT�$%��z����~n�RK{&�C*,����.�)����Q�$���	⍰,6��N��:<�����L�X�2���	VY��-��=�N(w*ʙ ��e	 �.b.��J���@<Ί�o�b�F��+��J5�D_!�ǩA�`�q`�ы��C̍����43b+�O��FP�����H�j��'�R�:�B�'�l�U�l��4��m����/8��H<�e�F����jaGq5���&���Hx(��Jd�t$9�t�H����5�NtJ�Y��c���M�Ҁ�z4�ÆvM�N�Y� �>�K�aeCWp'�$&���ѡ4㎆C��*�aS�I`k��M�ã���E��,w�����ً�3�? }|ګ��羄����+�"!`E���r���]`�FC��_�!�6���2�s��/=��5�	ѽ0!��a\z}�گ_�K���;����SU����}A� ��6�J�X�y���X�,l�c�m��mWzЙ���,n��MTBХ�j��c�����}V�Ӹ�i�p�R�ەz?��P��`�_�Ue{X�#�"	_�q��)-h�B2A	R��`GK��ՊX��re�QNR4L�#�MMh~FEpŒuF���h��6ly9�b�Q���Q�h�M~���+�c4hB`4H��f��&x��B��Ƒ<���<u�3��kG"� :;k��b+j�.���!B���Q��Gi]B
^���7!`5t��5���8ن���9�Z9�& ��D��B
C;+ ��Z���d�ƍ��^� ��I"��jT��A�R�n�$t�|���3�ʬ�|^"�D��i%,*�b��co�8�%˔@=����ݽ��K	����s�Z @p�bI�ɦ�Ҧ�?�;��dh��}M�/�B��XIn6�*`<���嫝�᰸u�(��=b#�YZ�WtD�on�c�J]x:�H�M�x�f�����77���W�����s g ڶ��c��&���I�kv#&N]i����4�Ӭ�%�,��%�\��Բh*S���}��V�|�?�e;M�oz )g++](���z���*G<��hy��LYa��s=�,gv��e�5L�w���J�i�� ���쌼cr�%-������\�y3�"HL�E�ū�ף��47�'���C��C�Ja�Y�0����??��!ښ<j����z������+�Dk1Zu��i�v�_��$�`>�������I��՗e���'}~Sc�+[2T�|ϸ'�����O�b��!!F&G��]��N���z�;��� ƨvw�Mݼ~}��ga���`o� ��p~)lܳ�r-uZI�F��׃bȃP�m-��r� lK}5]���Ne��V��0��ʌ��D��r&�6�8�[*�8�hl��[�K�����|��_XH�J���ؠy�5���5M��״�[b��P��qc�f��h�bcA�/��x隫��}]ٿRO��x�D[�w1ĵ{�uQ���h��i�PHFj��Q�L��i��vƒ
�J�~��+��z-�/�s�!�ֽ�)uY�⃨t�}-�07Sg�ZD��o�!�N��P������h��>ڔ���X_Ȗ�=��/�<�t0��t�ZO��}�J�����Z��@��x#�����z*�\���~||���o�N��/��Q'D���Ҥʂc$$��DD#�p��<�\'�3�u]6�(G(�x4�������'wy������{�F}����!��o�ˁ���?����w�~�m�M��ÇXk|���~��'?�	&�������������{��р���={��g�bQ��+,�+�i1n�A~>}�������X��E$�<��uR���\7�^]�M�xs��ګ�Q*���6�5�6j�J���Z�K)�j����LR=�����(��&c�C�'1��`a�|��(��H��jii۳�� /���Bj�)jeP������#q����'b����Q�@�b���R�ʸ-O�V
���^���ß�b?\c�q��}��o�������d<��ip+ƃ��L��ܻ���~��t�qX�a�>6��Ǐq2���/_�ĳܺukww����������9.��������������f���o޼x�v�6-w��p��e�#52)�Q���}�{�.c��遠����?ݺ}4c���"`6��N�ܹ��(k�F����ˇ����&FU7�^���T��޾}G�r�0H�+o���9�?H��
�\�9�J�Z7U1�%���ZFc2��%�b��,Vs���W+E��X ��8G�W����t�x���WC!6��j)�X��O���w8��J�� p[5�y�U�u�)�Y?I��#�X�T��-�}/�ט�|/�(���z���E�����$UR�B�S%ރ�0�Ku�\�86�3��z�CZ��$����Ebs���T��;�J�i�J����0�Ɣ�U#�6�XG��*�S�N15EWn��"X�aCR�mE���u���I����#i}m���j}�����xd�ēR@�sD�OA�^ A�Q	Ү6��S�E0bF��fS�Y���]��6��3�R�=L}OԄa�Ȳ�<PUݚ(�Z�z��|Ƭ�P��à3�F��|�m���q�MM?�ϰr0�0a�c�<�Q'��>�~L�l����j֩�	�A�6J��x�^u8A�h6�-�ݺ��F説����bXk�_����8��ʎ�1?���r9y�~4�L���L��}��B�pZ���A,h���X?�wv����6��hX$����?��nJ�4߯�~��b�8�@��C�:?�u��Χ�e#���f�G"�궡�~��K�}nC�0�~MP���r�xS�0�È,j1A}��	�~Bxa'��v��V��7�2�s���[��Tw���m&�E�fV_O��m?="��5!z[%yd��aق���$2k�ߡ�3^L��%�j@7���#�m�S'���9��ԹxÊ�(��I."��y������E�NV�m�	r&�8*���ỘXn>�����:W^22���ü=ì���X�J6ϊ�Yۚp�ֺ�8k&����Ejm�9H���1�D����"���<WZdEM�e4bl|�:*��'Ԛx�c��,e�-퀦O&��\�1���.���#ԣ�՚v���hZ�c�{-t�..l�Fxlk�7se���?�<U�i�F�<�w��h<�T�R�K)i����P�s*	��F�s�3���$����(�O���)7,c�L����>�DΒ��:ٝ���k�;I�uЯ����1|0f���5~�"��wQ�lv�����l��ƀ�喨S)p*傻�N�K�NC���X�101c�[��暇.�֍�q��;�/��cga�h�i�4r��蔔��%ڣ��W/eoOR���9w�6ˣpF���W�������P�v���؋�.7�z���O?�r0��6��܉v9�iչJH|�&$:izh_ޅn3�'A\�O�EίR�}�Z͔߰��JRt9Wz�X>�]#`:-��F�6k�R[�n� ��܃��pb��"n�=�V��D�X��q��V�pG�$Ӡt�z��nD��A������4��ܧ��%�5�>\��Y�w�L�㌳�ʆ����M"Û��2�ʬnl�ni��Y4֏��E�rH8{,g���v�=Pn����	l���7� �H��7���V	v�z=e���!�L�E��9�T�s��@��\ҹ%��;�g-D"�d����FEN;�V,�h����B�^U"�=�z瓔 ��!\:���L�P2��g�t������X��E[5��,)��� �;�!���|^k�䔓t�Y3�F\g��N4.$��R��i�Ӓ!-�L��F�ys�/R��#{NP�;c�&�QI ��<Z��_��2y�5
��\�������'1{3�,���9�.W�o"�^6�R���xZYs��Sy@[��п��o~�;������ã]5'��ps#w|��w���o��{1���o}��4�\�`�$��9�Vp�o|��/�l�&>��o�ʂ.:K��ի�~�������o�փ����V�zh#���}�sD���8��w���\H�1��"[mĽĐM�@?&�Í6͚.�1�����w�"FC������5�����6�l}aG.S��/�"��$�4�5͠Ňe�9oPa~0xl<u��/�l&�Ȃ�9 V�}^�C@��L:�h�~p2��zhJ:����F������Ν;X����w���LI�*�༳+��eS�&a>�uGw��LG��W�`<���[(PSP��P���;~���=��19<�w����ϟC�����i��:�L�';�������ϙ�"I&��@5������ӧ!��ﾋ��NƳ��(]����E�<z�ca))��?�>}��#@B�zkm�h8�Η�L|d�5ڵ�Ȭ���{*�2��qYm0-�3�CÕ�� ���R�xF]YS�M�����[o�i�x�<T�0[?���"�7ym��TXY9K���*)D�x�4�bY((�;`��JjE�_��	����p�j��24��8bF�h��q`��U�������x��p�&Z�K�+ueޣ|�5�!h:ZJ�O����'����[SMsJ���i`��!Nޗ���%�!�=<�U�4r�qw�nNrr��������O�W7����ԫc���r�hz��!	Y���:E�fg�h��ߍ{����XG������~g���48^iV,MR����h �xb����r���g֍����[�7z���1��T�2T�C )�d�N`M[�����5.�ҟ|��hg�[�v�
f��9*�/��w�����R*�EǍ���?9�ޓNkڭEѶ$�n仇�O�>c�E��ө@��8�+�y�z�����}(��/��[ߩB	�B /��>�ܿ��wt_����9�-ſ~�����/]�K����{���W����-jWO�@�,Z$ �,O�8�o;nbX��7�2z�!�N�cau��N�"a��S)���J�w�\&�n���Yհ���c��$�wYGY-g��,zq�p���71���u�D���5�ayR�Ҍ��6
�p�Y�^���4tڱAz%D����c$����M�OgXAp�/+W'�+t쇸��u�I�@QP\J�XNo�q`��aO�4C2�������Z'�[{�)@y�Zr�/R:sK��6���R��U+��">?H�8�!b4"�cft��Kz75I�~�T�\*�Wl����z)�=��<ى%-gX${�n�ze~2����O��1�
k ���j����5m�v�n?	��5��Ȼ��9��4��V����j3��Z\�B�n9(����׿��0('y�F��K�'Ϥ�ź�X�(���g~�!~J�"+ �%q?�#=J��*�D�V�nƨ6+���͆�Z��r����1���;˕4�P��'W�]젌j�~g�5H��,�ٜ��Z�7B�b���H;�.}���Ϟ,7���iS�]	�D���pJ�`��L��uO�oH�U����G�)65��X7��h �0+W�,�*Z�f�U�e�)Z��-���N����ݾ}z��~����n0���w0�5@��C��$��q{�S���2ԉ<ٔ�1�,��+�3��6jwqqM��C;�#m�,��۝�د���EF^jl��j�Z}}c�f<飼��h5I!�1�EnPx9�k6��nC�w(� �]�Q�ɎVvGGG�|�/il�.{}Z�Zț�����5VdCԳ�6�Ɛ	[̜t4b���7�I��T������U�����шMj�����X�

V���#�S\/��9�%�3,��h�ua�r�y���������Pˢ��b��@%=��>��}����gO$��]ų���b�
���̒*>M|7mխX�Y���7a�bA�Rj�*ɋ�t�]�Ϭ֊���U�)U��kW8I��z��G���H\K����y ��i���ܦ���rb1���g`R��	�I->�rBeu�.A%^�Ɠ��d6[\^^O$^G�*�*�7�P����]�����DҜ� �=x-�k�,�<˧��)Я&]ՇS�^1�f���qmlf���ɞr�K��-�^���t��	<Żh�L;�9_���VҩcJ+�6��k2Q*h2����>�M%[+�;�T�.ofB���xS�p����0o�痬�b�M.R�>�B��H',�-�q\J�s-M�&���Nipqqvrr"����F0��z�^֍oo+���a(3�V��Ȥ�8S[�w���zm^�����w��n}�߽�I�m��=������!L�
�>��;���pK� q�)�&�c�}�WN�
?������ �r��KFu'�����Nޝ��o���G��xK�/O��l� \a�Yn���
o!j0�p+!�/�/����f���9�qN��¢����dϧ[������N���ǹPJƠ�^H�hC̶��=�p:��3��<=KF(a��Ό��/-|�����=@9�J�{���M��S^:!4����9E���/���� v�^?y�L����Fw����W��)�{���NYtV�5-CJ�V�3b}���o�&#��T�d�u`��q���y�QJ��]!_ο��nU�M�c�t�O
Ţe}Ҫ���J+�=xp�J�����p_��[����	����P0��O���?��1?�^��xy��)1��/i�_�5�D2�����`\\_^��x������+��}���O����-�	o0Ε4Z��\\�FH׬7�E6���R�N7�j,���b�0f��4~ٝ�ܹ}����ԸFuP�Ӊ���\^=y��O>o�&�F�`���Xf� mNN������We�0c1x��'ZM�.ɳ���,�C����eC�Y���F��>�$4�8g���S,��XR��9��GF�L՘JHr����Z)^>pLUJ#�,�.�r��qbU��/��ؓ���B�`Q���S��?�O�,v�~Vi��6j���D<t�(��΅�n]	JF e��4�l��dg�[U�;��t^�L@�ft�X�Kµk�?	Lk�Qk<��\K��=�MP�j~�j뻆z�"����d�p�1U?fJ#r���)}�=�&B����Y�$=
^V�\��D�-V.�i"�s��Y�b8h�fmEx!�T�Y��4$,��r�~�>$Ga
�&��u��nZ��RX�\��˅�����0�k1d꺴+)]��b0ʅl|��~�/���I��n���ӧ9ln8c���<P��焏\W��͕����.nӊE��F%qch"�6��:=j�@�]X{���Q7���(֦?zn>���\��򧚈�r���k�#D�]��ձm���m8��(V�����+�E1X��N6�A��_�[�1�(���<b�n�ZD�������vb/�«[�I��`{i�.���F�qo)7%:��bj�D���m�y�K��N�a�T͙��k����rܚu���O��
�(�+e�<�V�A�8a�1t4V�D��1���Z�ԛ8	"h\ɲa$�R�avBHN���O�Sxk5������)���05��!�nGY����kn������-���pG�\��Z��O��~'E�ߎi����ᎌm0��r�<?�&H���7U�	^��:�ږs���g�	�5<�3y�Y90-���!��7�um���h�E]����MU��_���k�ȇ������@MH*v�.���Ұh_w�2)��~��L�m����V`I! �!R�`���r���f�C:rTR)�{A"����J�����ˀ��w_��={�����z['�k���0La�ê���cV��ө^!V4M3�㣏>�:;�)��H�^��4�;��Ɋ��V��6�n�����֘[H��@���װ¯��G�+�&K}�	a�Uj=����Q1��������0�A�`8��(�8ɸ��^�x�,wzz���[�ɟ�:�7�����࿬DG����f�3O�X��
���r�f͑ٙ��]cŖ@�L����Ue�ƤI5����ӫf��q��#=��XuK%kI��E2�Db	 �v�;�|��G$�5֚0�D��ח�~�;���Q�L�u7��+���[ښ�����+�Clf�*d�6
'��u�!�����U��4EA�����Qf������a �>{��ݻwi��C����
�����;c�T	��]&f���j;@��{��L
:��)��q�" ���vh��#�em[�D{�^X�qD�c��F�]]�ɜ��CT�Ԅ	<|��?�)�"k��Q��h��G��S�fp���I�>�N>�zw�o�CGB�(v~0
7!�oy:ؕ���d$��R��%��� _�ztd��D!�� ���Ё4-JT�U�u�ke��c�ȳ9PLԀ7PE}�����e(����A!ƾ�*Հ�F�	b/E�_)P���},�}���&/��rqX�J�8ģ����ы�-�bA�-�6uo�a�C����������.Lx�mI۩�Lv9	a;���W��� 3��S�(���nv���8�JZ����x�E���4B��l�������f-W8>9�o]ߩ�������QzJ��E�6�|]m��"��&Gt8���T{)����y��X�7(��z�kL��}r�ېSTd�*��Z�i���XƁ�+�r��٬#"RO�@�r�>�J���c�Q�$��j�vF)M����U� ��#`�7�<y�Ho�X	�u��]ܔҕ�kZ:K�/q}uC��-�F݁�ր�!�*ܚ*��a��#���k�k�R�QvŞ�,p������{��'O��J�2�_�4��;�9���bi�t�N��4��|�שve��{
�P��)�d9wwoP�������0�&#�1�����>�*�_�_z�I�j�����ѣ��G_~���J���zF#��Fajݑ�m�*e�F���Dcq�@��a8f�n�;�u4�{������r�O>������{29r���_��?�WV�ɉ#��ؔ�Hw�����W�),�Rl<���C�]'z�� uwy1�L;d���%�Q��;�4>m��Zձ�/�����w��(e�@@�^LnM�(P�h��:�	����B�у�:�����:���mǞ\�)�ԺО�Օ�NWk�U�M��׮[`=\�vE�5wQ>k���V��-���1^O��w��f��T�h���7�ǔI�fD�ѪA��S�\J���4�^����|����3ߤ]�Ƙs"��5��l�R���uUy��2������iv��vo�8Z_���A,3:���Ic'��W��Gӽ�!c���)�n�H��]��>Kh̝h����'i��aA\���W�';�~mü-�`U�i^�IL)��V���1�.��S�n�$� gQ�Y\ŋ��äϘ��a kT���JL�ȍ��y�����_����Ί�9F��#��0���i�Xd9FD��ϙ�L9������g�Ϲ� ����*l]�ȗj�)JM�o!{������d�m'W������/�4ɷc#�5D�>p�Cp#�L_�
��g���P�ܻ�h�SDf���E��
c�&޹������ �	w�A)׌{�b"�x���|I>$'�������XRA|��ɶ	l= ��2P�:bHһ���tQ:�֑�'q�7�|�,i��Iޖut�< �IҾ:a�%���4HK��bl�?#���$?�[ܪ�y���iiT�o�D��sm���i�遟�7P�!�QΌb+��
݁�!��~��q
�����Hj;-��Q�q\�?�.�ő#�K���e�;��`w�n_j� ��q�7g�b=�<y!�.�q���v��_
r-TAR���Ӭo`B�:��0[�W�|&�G�N����~_�k��L��Q���?X>�[k����i#�]�v�
��%z��������]������W�k��REogE�����1T��/G�%�5����!����TI���"gW��t�E��w�Ŧh��s�T"��E)���&χ� a���1?�[&S�H>Q���rszv�!���D��퉷#>�o��������Z7w���W�ݷ�z��Y�=�npn3kBFB[b�b4���Mߝ��~7�/�MQ�����l����D�]�.U���P���x��3��\�ǎ���p���e�:{h[[�D��2�}5�<�ļ�����c���?eQ�^�CR�E��4N��C,�Zö������'�I�O�m�F�M�0.�VZR��6f�d�y��X�mV�j�������B.�%�/m��j���SG[T�E[os �����Il�|a5���j5���I����u�Y�]�/������~^�6''�9�(V�uqo0]Tk�mi���#Ϧ�>N�u�"U�^��FU�_L�5�}�B�\���:q(
+Y��j���J��1���v2�t�th����bF��+��P	.˝�eg���������-��2�M{���jE�4���T�&K(k;�L��h���	�����ԉ�8�_��F0�e�ܢT�A5�E����6#�FE�#�F�W���]ή�:q,�z::���q�+:?�� �@�E2r�ـ�.���k�x��U�K�,��5b=�Z��h��u4�2}'�6 �r$m�僁�ҫ$�Vc4�ڃb�u�4_9�b�Cu���%��-*��3�͚zT�۹��`ߺ���$����ND:��������b�{c�1�F��Ft�����7����@L�CT��t���ɫ6 O�v�I�
2�oԗ�E�bX�������;����M���Y�W��AtՂ8̡ጝ(�igJ��gf(g<�mF�\���Looo�����7k���\%g�hzxt���'xK`/w 70�ly-2�_7�p��E�^�]��v"����zӛ�njȀ������W��Eou�k�)��Џb�&B�.k�o5�>����T�s[� �%?QUnꪸ���o��$�.5���?y��ѯ����7)?�Ne��Ґe=����ku�'S������r�ׯ_����ʄȾF�qkbim��ڷ�#X�Z�zS��0���i��n�lV@��`��j��4x������+����4���)kK�1���n��Y�j�F5�^m�ko�b.rm F�Fm#�g���d0�+l6��q�E���]>�� ��tPk_�x���˟��/�f� wMY�����Q{�@�[�]=�+��JWm'�lW��+
�S��צ.7�3��v�"5�X}D��P�B�5��s��gO$���-�&�<_��,��̡h�H��D���]^�W�Ϯ�6����f,���G��ٟ�����ޱ����?�M~��ߗm�������2*����^��T�Y�uQLe�Mq2�4����Ϯ.4߆��˻�zyW����SX�ic�H�,�x$��삕��N���1�k����>�����H�����������,��U�]ס���6ݨ�5�c��D �BU��N�5�SY;��г�z�f�WJ�^���.����k٘�m�4�.�D�QO�k\���r|{P����
$*hz+�A'��	KCܪ��oL�v�6C��ٌe�ޢ."�1t�`-��7�u(,5;��~�DO���bX�]G���-:���8���z��η?����;*�1�2`{;6�� ;�{ĩy@C�F��;W3�af¬����!S�x���WK0�<R�_R�)Z�.��u��H�$C���Wc�n'E2��a�C�W����SpW��\�@���[�;���_p����w����Ԝz� .:E=-X�t��Ҟj��$ɮ�����l��G�?Z�_�&�hR��e�F̂�H6k�%��w�����Y(�]n�8�4�{#�W;d�|L�U��6�7��z3O����լ��=;�j4���r����5�)0�(�ҧfU�Ѵ���@cY�>��VA��G߷��N�[;�|h�������@B5
�?#עDm��!���ta%�mq��>߁^�2g�a��I�[�Rhm9Krzm��.��s��D	-8=z1�,9r�#�	�w �I��3�sGX��3��G�aGn�9k��rԝQ2%����фX8�b2�;�Ѹ���������_!vN�L��0 ]؋���E)���Z��.�`��2� �<�|E�\f����N%I�x�C\L�Ĭ��(a�cC�t�������GH�-�Ζ��*�	h����|�����	�\���R߫�Z����.�%�ZM�8����Wv��Y�|�c��5[-r�vR��@���t+I��f�9�4W@�7�m����W���f`����1|�)�a��w�~���7Pf%��8M���VȺ�Qj����:2s1�ۏz�l!@��d�<n���b?��X���N����C9����L4��� �h���~|�6n{��=�;Jq����[dt�Aj}�1���j:L�#e�%y�y6�[��0��0:G���N�.��[��jC�&�-��H�M��,����#u9Ľ����g 562����������hC�ׇS%��:�|.K�����v8��*���c.w'�>��UϢ��wS@
�
�h�m��F��vu�my+��;�����#pl�.�=[��]X�|	�=��b�t�B��}?\��=�p�ha����[�_a���^���p��j�'��ӊ����F;ĩ4��/3	[1��|'�u�'c5q�M͝�U�����F�#FW�[�ͽ{����w���$��� �� �N����oUI�$p��'3}��}�kjZ_�L�߀��m{��O<�u��@�w��V��FP���&�E�@�#Y�/������mL��UDKZ6��������[7�we��Q����`�O>d�)<{�l�\��*�ܯ��j�/g�uǍF�edW� ��eX�Wy6�on�:'����M�7�,B�fH���|��iL3�B����p]d��X�JrB/�=�O��]��m}o
�!C�xE[�>O(#A��5�=I��%6��4u�x�X�I���"��w�/���X�ފ[%�%u;ID�J�LX4���?>>��I��xu����|H]�(�r�z��E��\G&P�(F�g�t���u��:�9jޱb�WL4(,+��@\F!���v�Ϯ��L<w)29���+M{�#�Bƥ�,�"]�^Ct��)K�@ͥ�/��#��D{��.N'K O-;��d���T�oy>�ZfP��S��E�l"�"/�Tđ\D���&�5���ϧ�&�I���Q�H�!��/����%�����[����B`N~��]�O?�Tr�^�h���g��;U�ݣ�)T�K|���!�&ퟐ@�Ѡo�7�;<<����������+�k>o$3�ˇ���"/�7���t�}H�a� �4}��KR�%[����c����Ɨ�ȣɮn��B�^�5�{��V�J��\s��>�w'>���r�i�d����e�rψ�i���7፴[q=�{ʋb�GP
�˴<��-�?��d�I�qG�-d~D�kp��H�����u���i��␒xRgQ3I _��t�X�an�`����7�_�m�%�>"������v�7�7���Ϟ=���'ϟ���p�h��tnn�7R�s-U�A��y�F>���SA(�M\u��喝9�"ltKh�8e�o�'I��Z��d�/q�\ �/��!�D]Ƀ�9��a���[� ���)͘���nH�Hb�œӪ�7�0��f
���0�}�����F�막>W�Yq9��YC�: �ʷ.N<3���D���5��,��Y�J��_�Ag.J��|=h�1�E\�W�;0�x���^�\��[��ܜt���<�����^����Tm�H�ul[�]�	�����]�$&��76��f8Ɨd�v���	��J_6y�AO�y�UZV��0�L�t�g��t�+SS� ǥA����cJZ��wj'�f:B��w��B�����x{����k!R��_�0�;�a�,(�CD����;�)�E�Cӹ�:���s�3�­F8 ��+�������\ �o߾����-���5�ӛ�$J�:�2E"�i�V��Q�˩h���4}�m*`�l��t룁*.���t�ьG�(j�܆��!��c��!�%���5'��ى&�&>��y0fp������{5,���`�^4��{��Uv��<�z�̷�?�(���q �֡?&�����5�)i�_ �/�56�H�hsQm�+��-�ͮ� ʦ�\�lM�S�q��ڄ�_�;��ZS�O#V�7P�6<�m�V����]ޙ& PNhF���8H�[M˞*�@=�6��J�*�Ov@LB��g�Iؐ��a-4ӎ�����,	�']#2]S��E��>�D-rn�(3��b��G�n�"�_�SO�B%zz]u��ڎ��{��ؑA�����3�*�-���F��ƍ�Jy�dT���Z�s�y�dCm�]�]|�"
�ߥ�!]�CS��`�a��?@����3�S��a�c����ƣ;W0������ ��N�����أa!|��iq�o�q�}�� wP�˶ePƢ\��[���*�X$�r����*�;�#�#�+&��ȵ�r�M�{t�4��(FE�������j�(��o_+j-q�p�\�r�5�l���d�L4�˕���� ����w2�q��E��o�1����W��cm�,��G��ˡ��V�k���	��U����<'�h�%��{C}�,�gW�W��j�'i��h����4SpӦP�$��YЛJ��؂<�͌(���-��{&�\x���8��9]V��w�6n`�7�,)�f�ǅ����cXe�x�:,��Х��Х�O�!R:ݝ���{$0B����q�4K2���F�LgrBLcg�������ˋ�;92�(I�$�	��#��|~'��GÉFm<zDu.~�JI0�k�=�%���k���vG�R;I����:φu}�L:�҃�Jo�`}�jkA������ُ~�����8q"�&s.vD�	���i
K��:j�m��l)0�r��Xv�U�?b�(�h��z�Z!�g�(퇲��i��QC�h�x:O�\�e�G:���bU���'�/�Q��� 5���bA��T�Fmf�*6�o�r����X��)ʪ�Nd�\_ϵahz�d���x�2�4��´n4��L*T���Z7-b�#�T�_��Ҳ���D`�P(�������y�A�d����F���&e���A�_,7�7�NmT��q��o��&t-��p
�q���`I�Z0��+j#�S׽�K��w73�B���P�ȗ�k�f����7���T�Q��eUk�4�-�$��q�$�m�R[�%�����{��M[1Eg���;$(^e�.��tt8��F�]VX���G�ۄ����Z��(5d�c��F��a�)������q~~.{������ӧZ�
�[|��76a���V�Z~q�$V��(G��wš��#��f�ǝ�����WV����bq+�����C�m��˦M���ڷsE�0���]����+��Bv}���J#���F{J��*~�f��Bڛ���Z�_�|��ŋ���k��+��F�|��4�{�&�4�钛^�nh��.r)�����ŏ�bƈ�x� �G��;�$ {D�d0�م<�h-9.����f)S$�s�7&.L���^MR�4�������ȓ�d:Oȷ
U��'X�|<��!��6��3�<�a/��2�p��.�q�J)��+�Ҙ��p�E)���k̥1y&rg6Nrb�d��јӨ��h(S�����!�>��SK��C�h��� 㿺�תH+Y��y#��x��7��ʩ��>}w&�)͇��f��&��T��~-�7���]ܝ���H���{=~�D-�I��M��(�O�U6;���)�}kݦe����̄������A��}��izň�!�����M�#�2~�ӟ>��ŋoD���g�}����P�Gyų@�x�.t��5�q��D@%b�iv�����p0:8<�?�����/���˯��O���6"������}��7o�p?ˎ@
G�biiB$F�����e��އ��c7f�\����Lgsy�@Y�Aɋ��.�1�_3@P�xX#n"��$E)������y�Tr���G����.����#�,���39t4'��'*�֥v��v$���mP[<#���vj.���("�{,�l�8��\������.m�i{GH�B�m{t�S�#����c�t���\��	�-�C���c��e�ha�r�������]5�+4�1M��M8�j�[�G�g��^CwCNM�_�;s�;c���!�g�Z��[��!i�=&2L撋#���ڌʩ��j\�2*$WX:�G��j�,����8O"�д��� M7!�bj��>}��Fs��i�,�b|��z���d���`Q��T�첨>P~�d����Tob#�h��'V�X[k̠���j'�8�(x�i25�z+�@�~��F�2�#֒��P
M���Y+e�x����櫔��7ˆmR�[��]]tcK�;����ʇ�c1��B�R��q��)Q��.�l~+�<Oһ�&T��A�Z�LE�Ѫl�@���tF�=�%e_��W����涝�M�FhN+�h*����tw��k@�@�<E�[0��c^}k��M�V͌|e���~]����u�ba|-|8R{F�v�~4�;�1+߃�X�|D%r�����l�]o
�JP�i�I/M{`�a0�=�����\*c{���*���bU��#"=�:�b�`^R �L�S�WQN�r"���q�xM�= ��CcF=ι��O��F-��YF���"�T��+t�f!Z����3?<Le�%S����W�� O���+��{��	C�v�n֣�d�������z�����.=�
�󺔰i�E������ޞ��� .E ���k7�.�&�+9d�Z���h�� �����ѧ�ȩ�/'�����f��9�J<��hf},��bK7ɑoF�ƽ�]C�)��(�̡�N����pJR�6}����ŭT�������_�ӈ��í�a6�9�!���G�5]p��o%<T ;��5�5�U$�F�����)�c�G�*v�d22��˷�F�D99z;bCf�g��uVc�K�=�{r�k�U���\iT�w0���������b:"ڢ���
L�2��ԨG�PቖM�������l{¦]�"�:���i�'�nQ��v� N�w,EM�%�d&��5\b�H8E����̳��l���+˵����%�\��g�����x��ź�Lb�9�� �6�<�(=Xb���4�OA���s0~�{��+S�M�=�*ĥ�J6qRj�B�m�͋�o߾��%���N������E�T��l�΅ \����္^�3w5�,�D&\VV�(�iS��ʜsdԠL�@?�i!�BGW+��)^�tZ���栓�4vS4�,MzWF��T�Zs�Y��ԗZ���'I��'�1'_RdM�S.��~��W_������@���d Z+.��Th�|:V�G��y
eک=��u(Q��C����� 6	:��8c]�(uĝ�cBt�Ql��X���Ǩ�+��Ƨp���1��'�@�4A}���
���Gˋ�j���W;�"���:HoX�.p�q�Eu��52v�N�b�|)=����r��'��f�4I�U���m4$B@b[�[�<��������O<��q$tb���/���JR�L� Wa��X���B����(�¯r��IHQ�Ɗ�Beh닭 Q"�K&��x��NW�@O�gcCT�Y����lf��h�gϞ�Q��ɓ�O���_����(L�עAZ���B�̅#��9XT��5�#wyM�S)B�F��/�����7<����r��J%���X&-+�	��b�@~�|�2�2�@�R��Y���H:��|��5��r��ޭ��XA�s���R���7�u*����"��o��M��STak�7��Ψ�\8��Rb$(���o�s$��P�Ӵ��ZICF�:�!�j=����~�����aR���L..(ϕd��)�,��.%�ɈB�A����f�����`��>��K�!����#�e��4�����u�M�[��Us� H\~�D���ZT��Q��P�&7 ������8�o�MӜ�=���PS�aC��Ƀ��|��}{?~,��/~O � �k�H�#d��K l�3�Ξv,�!Z�L�|�>ۍ��3(�������_����ʨd���{p�'K���+�o�x���O��e�kz��`e�BC�#��d�K4�\/�|�*���'ݓ�G��UaɼR#p*��Ƭu��_�.׊�\,�T��4*仲Ĳ�P<�a���q2�;M>*���2�q=�e�%�I,��L�9(����G��)_���=֢�ʤ��ZO�9F�3��.�7h�z@&f����\�փ�+��t��EI[�j�`�|S�ֱڱ�ӥ�z�	��!Ғ҆����c=�{���?O�e�(֣�i� )W)Q�a�#����n|&Nh	���b�Тk}+s�+{T�c���U�ɺC��*�C�x83�Y{�������"Ɵ�n*�[�*Vΰ܇1PNl�@5��˴)Q�d���3�	Ez��+�a3(�R�kl|
P.{9��z�8�  ���p�מQ-�x�G�a7��	g�$��n�����4�R����\!�%��6@t��m��9��PQ���r/9�"�>�����qU��gʺ�u!�����!�FT�EG|�P��ξo�aP�뙂,*[ۮ��`c�]x!��n��J�}y��c&.���W�v��7�|�*�A��^�[7
#	n���z�&��[����"��L�g|���=�淮`�0�W���QB\�9�޾z�;ٙ2!Z!���|sn:D����gXBߴ����-�;��/d�ճԐ��Ҩj�E��-�/��&N��&�LU���Ц�b�$C%f���D}(��7�6l^�)	�N�N�#0Kݘ�d���4�,h>͖��t�c���"c�.i�Y�#�IGTy�<[�)����p�!�q��#���1��ڬ��qd�1�`��[��[�N�N��8^�M�1l���z�!��y  �Nqm"��خ�.���lR[��F�y�^��j<܊���v�)Fa��X:���(\.I3�gv���s�DpgXNL�)v�i����W"��2DШ����Pu�h	)z�>��z(E�#���\��hv��@�����m�����S�R/N�!k���Q��z],9����xr�|Z\7˪��L���x�ZT+Zp���]Q77�y�Zy�R�O6���j��ފ��[�름y�e�!�e�(�i �{f���NT��7��j�ɚI���-�� ��G(��y���w_�MOU݈;U���=`j�ǵ��u8Y�"��d�aw �끷�j� pYj
��n�vQQ��魬w�1���ؠ{&�������^�d���jԅ�PK�Ȍ)
�6�o�#����G<�u_F�?!��U�Ĺ�c����lv9�[������׿׸Tu���Rc�U�M&�Z�n�\�o�u�X�D�Gɽ{'WWF<��w��f���d�ֳMY_;�	�̒
J�sS���аq'G�13)�L�Nx�*�Y~px��ny��\�L)Zq4����*s��S�8�}��� H@2�0��(j^'�;���|�,�Ӗ�)��sp�	�H@�B�)����<�5���$	hc�!�x{w��5W��o~���߼T8OkG���2==y\:��p �)��p1M��bd�x�m�Xs��DeZ�>:8::�m�X�.��jS�j���\��!�
K��Q׈�0_�]���^/�-l�M0��Alf�*��y�j<�8Ab ŮF�e���s$Ҧ���������yR�>�Lū��\��Ϧ�Y,�2�@��N��u���not3_��_�{��$z2]_'2��{�&�{y�!�����Z���Y���8�u�Dq��:~R�>�Y��LP��&IZ�0J&��!����/g�*�Z����f��u'+vD�B��k��S�?��/����ڡ���r8�a0�*�:����1K�O�K�}���O�?��?�_�#,�n����\V�H�:VP&Y;E]cZ-��5�W����k���'׷�<T])��N[��v}{SP?b;ȭ��v�2K��������,Z a�Sf��#-�Р���#��,��]�Y""��Ffl3i󀒐kȖ�կ�嫯����gf���$�r�`@y���E����u�����y�H���7�Ŀo��)���W���i��7g��T��q�j����z!���g����&�<�7B�)�����]&[�[�8�;�)f���X�%f�����' g�NI������ ��>/
Rfn�'��L5c����b4P����oz0�I|'�ߙ.cªpy>����9�ڵ����H�5�j��#�~��?����0b�������#f�����۳�K�=E�1v������?�T"Y%�I�)b6Q&�MݸX!8�m�g����/�oW��у,���ɱ\��>��D�$[I6s�r5��߼y�t��Hr3sA�
�Ǵ�>����|�^O�<���|@�Mt|O���7o�����\�����߿��:ڼ�W�M~ʴhk;r�Ѡ��F���Es��f&��5�р����G��z����ЇW����-|�Xޖ��j��]��N��h�-���	j��e�<��1/E��V���U�uq~~)Z	��J#v2$e��#Gխ�wȥ��tT}��9<< !�H��/��B�A&�N��;M&�G��TM�LS��,�?$�\⊓p�t@��蓋�q=
:��'����vb�F1��zVFG�@�{�_E�B�8S�.����I�=Eu���a��8b��=������]���Lփ����eǲb��:��v��"��-���M�=k?
�DO�X5<�a�ֈl��u;E5�|��^Hl�Yh�r�h�����A�[����eVP��zF*���@d3��g�
���{.K�8U��̘]�y�]��
Pdy$����9�)M�������q�%�Y�D��Ƞ#��?�Z�E����8���FW��dn�����ǩYT�D�l�8.��&y6�ה�X%�ș^�|���:Q��T}k[;ݟ�|y����8��t�X�>11mјۍ�"p�؈����<�W�:��D)�x��E|2+ɔ ������z�>
��!�K"�'b�eQ�� �������-ÀA&X�Yk�+u�I�.3�0�oE�m��f����C��1MAYぁ,n�_�N4�[]Ov#�:}1�1��E��%7���-h�a�|B�?}����Hc^f'L�Оq�Z?Y�r�w�\��Y3n|a���.��!��}��u���;�`���}J�Ṣ��25��1�<�E�<u`�����hYd�K�#��r�F�Q�K�	g�Ò�8�X�> n�-2���D6�L8�� ,8êG�#pT���,�=��tF��:����]�_BH�i+��ޝ��M<��I����t�!�c|z��HF��r8s�Cd��{�n=�W�4��?v����,������v~M��ԁ�Cl��C�ٹ�l����(�Q�xR^�q�p
F##6�'��!TU90��?��;j����S+����b��?�U�͗x��Qȕ�'�F��
�H�cȵ�tQ��,�ł��b��l�\hm?��ʣ�5:-�\����ԯ��
o=�	���gLF%>	��\�ǟV�Dt�ZGP��0"�Yb��ۖ�IH�v>9��Sf�u��14��W��e�\�N�" ,�,�����z�2v`\u����p��8l�.fWO���c��"�5̗�\�������ū���>]�]�"l�d�����F�$�r%G�ޱ"��AR�y�*�(BC� ������i7�l6[.Jn�u�q"�=�*�]q~���x�������菪zE% ����m�m������t5�<M�6ye��2��Y�U��i{��T`&&;���hj7��ʷ��JC�o^��	d���
�l������C���uY�����:�/���d��A�T��b>��_o��mW��z�LMS���cXA�Q�y��.�=�����z��y]j��b_^�r�Ɠ�g���8FoP�S��m�� |X��z��Ӣi�N�V���@�#t��SP�)웺�F��sSr:)�Ǟ
��I ���g�3qܚ���Z��!��s�.��kSݰ��sN�ɀlU6��S��j�e��RL&"�kה&��Uo�-k]A��(�TΠL��ޔ��0ĳg�>��c�����~����I�|�o��7NM�	��U��^g 
�=AF|%���o8�"�A4\hm
-�@X�}���؋u��\��[Nq%�c�Z 0K_�F[;���3M�~���o~�o��F[��U]/S߮��u�%�as�i���Z_�qho-/��Ņ|^�>��������|%l)%O�iel�[7�7�'�沲������J�$�L7���5$���F�&�J�R2|�C�G�=Z�1_�W�딇�:�*$�y4���V��o���Ʒ�q-�0{�=��I��xTe<���4b�]�{��|K���r�p�]��=#żD%���nUw\]�h�����jW�Ն:H��8�\Z�� �"b��������	�I��v9{��Z�������Y�$À�n��r8v�@մ�xs;G�TgL�(L��'����N�y).�e����Yb~��I����Ѫ1\��e\X�FM��{�eٳ����.-��VD[�p�e�t= P�mkw*4�\a_r�����n��i�Q�ju٢,F��(J%������+$-d+ƴ<�Ⱥ��J�f'�c�+El�E�T�߀�6�i��:���W��CjI���xu\n��q�zC�M��7��7��N۪lY�C$n�=�SC�ߠaw�2`��N�!�-���<�xR�46Au���A��|jJH�"�8���S\�>a��S�-"2��6�<����1�������zErd`܇|"�=�I��P/Std��b����h�sb�Գ��Xpz���<����8E/�����=A|��g���sU�o���=���\��$�:�-�����9��u���ɉ(2���M�<��\^d��G(���Uj<�%�%tA�8���-�T�k9�n{h�{G:T�����z�*�Ün��I	.��z���f)�d�Մ&��P��=&�("c�ؤ��?��^X��.R_cg|�����h@9�P���G�C-}@����^
����c۩�vm�w$d�Z/,x��!�`w^���}����\k����m[&�?�n���t6w���0��<��1���F���3�<6R&E�5/B�ˇ�5��Dp_�m+X�+L��&{mK���+d%��M�-�(o��S{Q��v�QJhR,�4I��o���;;T����w��2-9�+�B�V|K�oH�H�{r!��q�<��*2�v��5Qꐀ��	���E��hsE5��j�N�#�����mT�r>]#���8�Z7��g�eV)ƾW��r\L�c��w����a����#�B|��>�3\Y�Ͱ��keZ�m��]^��$ǝ���M���`2>�H?�����k��F�y��n&�;|�J�L%a7�0�l�↉YU��ΩM���@ڗ}���c6��<L�{{Α��Y'���ӿ"m�p�f}	��Y�a���S�,cC�S̔զq���[����EId�q!�0Ͳ���"�����f��=��MS�.�`�J���u���g,A�5.`ۆ 7\�����~J�Z��0/*�#��5�T��9'꼕������M���'���h��y� +NL�MD��
������N�]�o
绷��ҴM�b��R�5 ��%�x
dl4+�Vi��X��:��FًG+.�ww����,�b��4��C�#�+�`񝘾t��,Ocp��RzF�02�|��T<������IY�)���4~��̊��0�G�� �GI�>�����W_}����w
����v�UC|�ޔ�����Io��(����|��7
8���|�w8M�޿��YlJM$EM��e��-m\����Z� W�f���APl��_�ţ�[�ڎ&�MU��0hbY���&��@����bspe�h<��
mުuC0�j�1�T��~��ޑ��*�3�ɞs����e-��F�ӈ�`���vh�,���%r\m�>-�v�dzH�����̯o߾;�����7oސ�B�N�&�rrTi���4��$-כ.G\Ҋ�T�x���,����rnz-TԥjK9y>�N\x��&����,�ti��LU*�b��?>!�:�JC$"3=z�������f3y��uw4�I6���<��	$��ˋdP0���u���´۹y�YxYڜp�����1,Z������k���@�!��L�6����F�6)7�|���s�GC}�zP�L��^�e$�IL�t��u�+�*��XAǢ�5��j�U�*œ�(0j�ñ���uM�=�'#�,��o(]�j�7��IΩ��]�k�eȥ�V��+�&KU��X�8�.�9T��A.�&'	�##_��9�qr������G�˞?n}�L����0JWY�x�^���n!���z����~�����)(�I�l2-W���Z�F����g�?8�q���_��S���@A��$�.�OK�ʖ�9a�]/�r�RR�ּx�MU��"���������wg�c�����dh�:H]�g:�M���u��F�ߡW����rc���ZE�lC8F��c$p��;�?��_�`�y�X�ِF|SwI�L��_?��D�����Ha��ء����K���Ǌ�����"F�`�kE���y��7E/#�)�������,����.{�V�Y��f�,{���K�E������-Fɦ��bɭ�^�в�N���)
������@ԕ�GQ�, �+s!֎(��\�2RY��̘f$�V�m��W�����2��T�D�bS�"�ʂn91�,�~qm���V��Qz�)%��@��laT���=!m�&wz�
QX�r�ȜY�
.:�C�W�!B.ݔŋ/D\<x�@����iWW��S�z�:�2x�rF;7�'���,W����JO����������?d�&%�.9�����ӷ쨆�ѳ��J�n8�7��x9�S�$ަlHL�9:ڿ��O-�Ƅ�u�4M�L�̨�V������'OP.�Xf�?�TOV��u����ˋ�1�j--W������L�Q/��m2!��U�0��o=c`�ݧP�<��h����Pt�jU��E��]T�g�������i}�U]!�$h��O�~*�f����-Rڵ��eHZ�i�6[��fG%���⦣AV%��	�~d<!��~�&�E���Ġ� �dm��y(�cF�v!��v;�� 8G���X�.�n���b���sY#�Jkσ��X�K,����b�����A���vGQ���d�۲>w(�ԇɔi��hܱa��l���A��������M1x��&�1..��a ����r6����%0>)��M�4N��I�VBⴼx��z4�th9�Ȕ@�ZB�=�u(�R�&�h�0��~HV��qP���0�M���Imz��D;z� ��*�PT�h(�b��UE���Y�G�UD�蓡���'��ꊤ�I��(���;������>�&i2��ؤ���	EY�Eq��^��U<��e��!5zYE������6�-l^}^�LVaNz"�z�
Sc}(����Kc1mb��x�8���(nAkje�t��TKv����4� m��{Tg� ��wXBcvgY���٢}��.�6���!�վ�����w܍��������Tn����LOB���*���2_�l��C����݄��l�1��"���¦<*JY���D��=F;s2��8���
��`�2�ِ�� !ձ���EU^�\}%q���cX�m����q��f��=[G��#;�����Pi{Fs\^�G`�T ����v��j�������5밾�h��B�E��
���#hKp��BmO�(�FC��,*�3օp�q��^����x�E�z1�������~��~�ǈqY>���ۃ)����T��e�,cg�C1)MO.Xt/ґ����u;W�7�����+M]����!��us�T�r�Rhݐx�۞y'1�T.k�܀y!�9hČù�=ôJ|a�%�n�P���)���F��������ͻ;�jW��2�Xlʊݸ�`=�鴹r�iB�α����f��NT�=��N[=L�3��k��x4&��)0z��Ѳ��E�R�zj����>i�A�)�KL�O$R�a�T�t�͎�t�T�\��d|���0�-(�IFY�s���9A�B�!������-(Ye��_�.6�����Zi䑶�'��}u@�d	5M� �|m�A�	փ�bM��sqK����}�A(3!}��J|<����t�9�z5D��@m�ɈIoyU�O�F������S�L�{���]'�̳�9a��ep��S�����|jĬ� �ݻwh��������jST:7����!a������%�9�O-�w�={���}E3��_���p�d)"�9,��X4ⴰ���ח�f���\L�#K��@�aM6Om��'�A4%�k�������p�굊�N�1���o��E��D<8Q-w�u���ɒ����G}4�N�D&'Q�1�P-x<G!�N�A\Gͬ�G�
������Sr<i��.���+�Y�W�J��!�J��1�X�{)���&R�Y��b-{�=�j���b�;WE͓�R%��w[���V�=uZ��k!f[H	�8::
�"`I���p$c��Ty	̕��ȵ �8��@%H'�K��gA�0B�x.Tgb(�J�.��0�����<v1 ғ��W���豬��l�0������U�Г�(��r����I��۷o?��s�_��_�����
�m�]>��c����i�|��a�I��:0����t"��QH���ЊL��k�Ԭ�E����A��q���J!�j<m(%9O=a_����7��&Dϑ��̌��Nއ�Y�Bt]k�(T9r/��Х�J���"��J�(�s�+l��T���ز���,W�(ݝMH���|��3���$�������:/��t+�7��V?`�(+��k�+2ߠ��h82۬��d�#��4a�̬�$�3P1K����٢y5;2IT�?FC,2���tQ�j!�G���+ԃ ����f���1�k C���qB(Q�/:���wW�p}��k�����Q ��W��9:���j}o�'O>�֥�@��b���;�u�sB��|`�X�f���V9<<E��O~,�O7y�l���_~�;���,g��l`
�\kp���Q�>OL���fbE��c��[�����/[���#�吻$�}��]�A!v�����<8Pj��dL�9���.dBx�(ue��:���1�n�o��3UC~�+É���X���R��7Զ��D�Q�����E��M��H���F �4ԕ����2_*��|~�v�E���q
Mhi�QAw����+�����l��"IK��p�-����rnY�^�ě��g�&�l��G�3y�ȈJ���8�rz�c�g5�D	8;����F�!{t\^���b���Rt���=O��%^.7Q̴��B�]��7g���H"ׂ�bI��` �ƨ�eHT> 'H6!��"$��?�m����1��\�ҌÖ���3Ǉ�a�7_|ɑS|��;�PYB!�0t_�����"�g�4>D|�η�N}g?�a �p�ku�	�#
R�\�mʤ�(��d�����g	NNol)�ĩ�\Qԭ��iF���ŅlK��f�s]Xb���A��S�`���d|��~l�GB��ۍ��zT����g����+�ⰳXj[�<tn�0��
��;?��J�ݿ���;��v�R����-�S;���
���5�Å�,~�.��P� OwHd\�jw�}����)�,ۚ ӝ+z&<r�#ēq��8��2�a����U�,�����ĪOАZ{���Zȋ��b\3�x���С�.ă�����
�t;wʃ����h]KbC��Z"�[��rY*���v�%�q`}��{��w��6D�2������!�v

3Qn7n;�t;��9-��`	��x���Q8�Lr`��p����ą�(t:����{)p9$ل+�;t­�<;ޗ_8�ǱS�0W��M��51;�Щd�^x�M6�1d��ԑ�6�ʊg�v��?D$H �NM��"��XO�^TWH���'�c�NƿxD��Uv�	������_N�(�;<�&�;�C�����߈IG*���6�{�����5/`�Mm���ݐl�0���p<��;��ZW�
�u�J��a5K����Z��N55/���Ǐ<<�a�V*�G�=z G\&)Meg�e�@;9Xp"u���������߿z����fU��t�5fAdCy��Y����;Q28�rX� �$L6
N�+���vS�]]��=3`"��X!�<,-<�8�i�D�~��E]=X,�{{S��U���H���H���-^�Q�ߌ`L/T]�����y��Qb�x�Y�B��<}w&V�����lֵ��y:�T�nź��&��Į�����y��xzz&˽�<�n8R{�*�y4��'�If������p�6v�(���Nͣ��s�@ Dc�yp�X?�f|X�����˵ڲb��}{z}=�o�<:Ѹ�J{J��'#��^mYŃ|]��OB*bTv ݊"��l&�WS����8t�O�&���'�*|����Z}ַ��D�Ri�i�ięy��T�+�o\�X�H.������џMu7� ���>��tv2O�#�ORtU*��z�C�W��D����Ll�1�S�]ʪ�O����G��ng:ȋY��mzy��R��2-���2-�ޘҌ������Q����r� f+nۛ��/.fb�ӊ��95���bXJ=O�����-blBLCYV��-�t�6�zS��-�,V�Z�����"�h��&�W��#CÝ�٠�d���vj���UG�@���ϝL"���3W��ã���CV3����l!��J��2�4�,�L%��Lrwƚk_͝��Ҥ����~.k�mצ<e�D���@cq]ޠ���w�_~�e������u(�m@�0Y_��Y��l�ͮ.����~��?���~RV���n�w���{�i@P� m?��˄�U��ԖUmz��d�q'>g�V�i��#�6gf��G�0YP���b�����w�߿|�N�<ۆ�ԲK%+�K/���S&���Rh3�ց��q(��,.�_ڙ��J�-E
uq ��P*�y�䉬�xq�^����;$��ij}7�e](�o~��V�j�h�8�j+�ӊ�RQic�2㐲\�	�FA�rl#�[��TƸV�==�B�o"�T�Һ�5�ן�\b��#��M�Z�X��o�E$�H���j��w�ИF+a�����\��lv-Ӓ:��	v~�pw+�#�!1���H9 �f���*�3ZS�ޠ���8�d�{o|���K�|�!X	{I�j/.@c��>M�L�=��+L�7%(�iَG=�m�]G����5��N�����6S�%H���
bNiZ�	���'''�� �S�8׎�.�zu���P�r}�fQ�;{���G����}����?{��Zq�F;�D��LB���;d7m��\D�! �,��Ԣ�u�˪)�h�H�'rX^�zI\!�\�b��c������5+��Q4�׳+�s"t�`��A�a����X���rM�:�>z�oo��޽���|��H$�0%�'\�40�����$dBy�"�~�&���{��1�k���J�O�˷@��g�90�H�}�LV3��ݫ[���~��8q�5M(�1�?�����+f�Ў5"颦�:%g}۴rr]�@-\�57�5�y���z����Ⴡ|X0k�`��N�|Z�c�͚iZF$kO�G$w/�g�N�]���A㓾<�4�(�������D6�z��=�*p�\o->�����^�'�b_y�����Xn�Q� �BL,6�̅E��`�#y�����G��=PѠtZ�@�����B �`V#�K"_�F�C������f1f۩�;��*���-j�hBȩ���.'E�x�U��"ߒ�ba�f<8&�=�T�D���v��0��k�4N:�.<�DM�@����VE�p=b_}�0�������`�NQ |yq���;hD�s���Z�Ԫ98����7�{�h�6�V�Z1���Ùk٪=�X�ڃÓ�M+r�w.�.^���g�b�tP.�C�z��m�,�a��n��l��I�-�?}��k]3��i��]4��fq1��Y$����ؔ4
�<76�h?�M��}��l�7�m���M|�)+�g4&DQ�n3�-�M��5a�-0�+t�A��]���E���E���%�ZK����"ji���I!'g��k@�q��~�����$a�ދm:7��@H�K9E���.�!�b=*�m[�\���`���R� "���١��̖�Σ����mOc�b����ݼ�̵�ᅚ�{c�|�|-o!�b���v�u�y:��"]%��j]ϙ*�5��ƾ�d�;�c��nl)$Bx+X��N��$��>*��ց4����m�T*bj���n�lנ�)g�
R�߭��,Sj�g���g�)4Tֿ��/�^��JXnT�'� 3��	"�?\&̘ך���~�x�Ƴ�-��;�ҐfI)��%�Ð%swr����E�7��3���+-�[En��7�0dWӡw5^�%�z��_��%�f��v���c��k!�_�z0��Qr���� �岗 �9����'vm��Y���j��#�@���k����z����ْ,w�Y]>�G̰.	�pd���
�a4.��V�p�-�L̾��v�U��;:�H��O��냉��?�ݤ`V!�X� &g��F]E��4&	�P��m�/�gҵ�.�؝��Ln���;�.F�;�\f���F�/"��mj1��@o}~qzvv��h��M��%;����E�I�w�x����ViQ(I�9���JQ����7�\s�7�x''��D9Ol�����[����"w�'7͜I��K1Zd�̍]�D�i���NT12*�%��{qq������bő��T��L(��x��ŧ��)q��}ƞd?�S΀`~{G�+�kvW�,�s�k���3
n�L2W��db�:j�)� h�5 ��ɃL��t�T!4k�m�,͙af�<M��m�s��;��E�A҅��^�>"��{Ǿ�w�R��(e W�[r~)cV&���p�� �e�!2N�vqGxӍ�RgI�jy����p�Fa#Ϟ>Aĳ`�G�"րn���-A���-=�H��0B䅳3Bh���Qة���IqD�/q�eZ�|�R_���Z��.��r���%�Y����=ȷB+'~��&5-�4K�kDE���6.D�T�E?pV�Y� �l�oj)7�&�6wz*Q�t���%�s����zp����?����������_��_����g�¶璱FL��f��!�##U\׷w+C��G��̓w>9�H�:vW����� ���oN_�|�\n~��_����6�6�M���Qbم0m$�@���#�|s���Ek|�?X4��o�!�����枹�A�LN�[�)w�裏2�c�击�$7Q��ŭ��Vݼk2�ԅ��&����]2�D�GL�";�D��t�D�	�׵��f��%�Mr�v�������D��0`v*I<C%���?DOMH��xѠ��:B=�
6'kN�6�8T�],m�/�Z�`#ԩh#��F�j���@�<2�J4(W�A�2��7^�[G~���łۀv�gX��}��m����|
>�܅����c�̯E%�� ;�^B����`^I�e�(	 ���#���.U��1<eT���������/�R>�zd�{��t�K	�\=z􈴡���T�#K è4nٹXF�=y�Dv�"�`!�����?���B�L�\�|�駣�4�?ĝ��
��b�Gn$iy��G�	�&�0�@D(�����)���\��{�O�8W��'�v�M��B(	N^�ިv˲Or߄7ea)b@L�+&�L{�-+�������bw&�1�)�d!D��̓��OQr�x�θ((T������*��e\	��
���d!x�ڙ���v܊z@p�MN���#ՠA�)�Z�%�.ĂЍ�ҽ�0S+Y��#U��53�4�]l��2{�uYtE�44\e8��|琂�̀]�\���r��3�����-k��LQ�A�r�{��\�ؗgq_�;��4���ܟ�YDXWڞp̜�)�y$�����5�$�!�(�/Ŭ�3ʎ���hEX�M���&f�����F*��t�bw:ύf#,"�x>HC��p�c�fX),S�R�Y�6��A���^�V��j����j}��rMy8-��9n�F��h��[ Ș���:e͗�� ��E!
�/���;��AU�u�#�{��cD��?�ӝ�]��x(b����T��f�	b*�Q���+d�B8�r�Xֆ����:��N�s�.��;�YО2R}��XS����k�ղap�nJq#-#7����<���J�$ۦ�}ۗ�d�����G�={�Z}�j�6�h_��*eɲ����L��̥o�I�p�D���%/3X���N�Q�V�6=���ZS�Z�����f2�����(_m��T@вol��#������ �1�8�8;9��S�z"�i|*`��H�Zm�Z�E�6�E��)cl�4�5��}�Ѵ^�u�Z[�p�t��9͟���.蕧���b_�k�P��(���r�r���� �h}����~�)m}�����O�+!���{�/jW�[#@���w���Zq]�zo 3���D��Q*س�1�qUD�įD%W����Ь��L���?��իWbZ�w�J1��(_��H�]>i��l������~ǁ%��>�B�}���cŉB������j`�"���2�X���cL��x��<L��{�k�E�*^�N�X��[7]�.�df8���լ΃�Q�]u`-���nn��iKE��VN-��-���lT�3�����C�S�����d-*���-�R��2�h�E�&��_�r���w������A�X/'�S��..�⤳Qc��`�ڸT��
`�޶Mg
.�ޣ0qu\_�~��ݻ5�p�~�r��LF=�=�6�I*[Q��6��I�\)�N6Ң�H�\���v$&�����P�b!�6�����Ng��X!0�}�-a��`nP�Wօ:�
b��\��#���.��_��lzqys9��F����6e��" �#M��~aȜ�t*�l7�Q6����{)�* ��b�پX}���~�R����F��6�}�E&QzB�S�'�h�`$�wS���PƙB� E�,nOoo�O>��'?V�f]^�s�~RtD�"�4 L�4A�#���]^_����ë���ō
�t<���+]���v��V[b�O')z�Vb$M����o�^���Q+����#�j�Į�Y��6r���ͮ�~c�Vx�f�W
U�c�<��\�ީ�?�0���v�x��}՘�D+t��.޾}+_����}_ܡ<�i/��<;���7����@�q����TN��ⶪ+�F�Ǉ����`�r~��U�kf����4�@Iw��eƢYE4eӚ���L�4�ˢy����խq�lK�����^U���QcF����N+mv1���Ɋ!u>�v��{]Y9�Z�{���|}z���}4�}{6w�Rk��ի7��[�ev뻾ݔMD~Bd���Kڛ6I��bwͽ��^гb P�Brh"M(�I����3��d|$(�0��޻���r��y�䃉T�XOuu��{#<|=~|ϝ��;�����I�;��:\��������6������O��6�w/߼��gD�&avx��w�C��(�г���G��N����{i�'CZ$eZ&��{�7�3ps�E��%(>�����yˮR?�1��e�I���u�d.��5��5��m�Ռ�=m���P�P�E���l.w��jvmwb�����lR,V��b>[.ggg����{r��:;="	����rV,W�ugI���d�Y�%}V���S�vU�e��Ú��e����tmX�Ǻ-�u��lr��ɧO����N�����woޜ�=��$$i�0��](�i[��ȷd��R :�B�\�H��%�����ɞ O�pc�b�k��(��_��������ݻ7~����|����=�"�k4�����V�Ɂ�v�Q����>�!x�l��T�t�� �(�/�*=#s�f��̰^+�� �Y�B�ӳ8�7h�3�=puQ�b��|���X�Ξ$����5�Nd؛�`G'��{)#xr��f^�� <{[���)���L��KI(�(�YE�B�1@&U��L'� k�0�z2�1��#�Iu ]�Y�n��{�")`!+�b�.~��������+�l�vʴEn�&� (�%?��],cp�Vx��T�䄵�L�Vq.
�3d��D����>�!ul����֭Z��?/E;���;��F�s�������|�>S>��������fO�<��{!�� f��d��PzAEH�2ǰAI��?Ҵ��;�׷o�����=��B����ۘ����q��u������㏎��T����}�H��$�	)�&j3%R�ً�s����IIH>+L&3�aA Y��B����0�X�(I��+H��+��ߓQx����s:���6��Ii�%bZ5r=��	-H�qB��S%�^�)	�����:?>��״�e��������f�	*=��J������[��-�����󎼽�il�4��P���G
W��4��u�se&����^���\KS�]-�[L$�A��8�y�;@��̕de ��6=��ِ
�
y�8&����./��w�\#)�����,J�(�"j����%È�
	5���Q�2i����6�y<������L�P��J�axq_JxH�P^ڛn
	R����lԜ���"�i¸�ɟ���O�PT��z�VCWBNd�\�����q���	a>}פ�X?܂�֒~Im^�T+}*�~T¶�k:�R=�0=�%�{�Ҷ��1��ȏ�<�}���=�� ��X?njr�S�Z�&�:���� I�v
���͵:oĂqhiC��r���L�\�18�3�<�ᡛ��l���ĸ�!�g'̴�2Vȓ��W<��B�N������͎���K1���c��0+J6qL�>$��7}̍s�p6+�C��ٮj�"�ֻ���8����$����-1d��ЩƂ[��Q��y+I�%*��@�״ ��(V�,����-��KQGy�r�^Z^z`I�"V��#:��<�E6&)�xR�(_��d'H������A�r/�I,�4GZIg���=3�p�u
�	Z��u ��q.¬u{���O&!??�
�\�0K��H�d4n#o��X��G�l#�p���BDd-��A;=4����W�gr�j�ȕ��!������Q�L�u��S&�(��X�q	���b^;�t�7��sZ�E�0U@/��$b�\Іu���;�WT�6�;eh��a���ԉf^�������s��:��&�+��+�L�S���t/��þ*�.��b�i��<2�C���x�}b`��px���>4�'J�wb�ce����ɨ��jAx'��j�K������0�:bU�p�ۑGq#��@o&��pp)�c�@�B��g��@L�)*�?
$�/�����V��*�hK~Y�����6�R���5m�=�@���)Q��kX�9O�EB��];!�#w
�!�p���j�hؚDg�����+��N�[�����k�QO�����)�}�^�}�(�)�W[u ���!3s���� ����,�T���i��e�8����f���_�����g*qH �:�a��x��dU����T:l�{>(Q�-�hʘ�S�hC`t����H�����mOoI��l��b ']�xuD'0��U��*P���'��~����~���|�ɀ��2!�������e�?9W��02^�¼��J��r��?�H:C��\��^.��$�OB�A5M���u\���}�c��L��2P�d��V�A�	b��`�yt�,#��~sq��s������ŉx��nL� �;Χ�Ǯ�r�O\�9{�����׿M�Jl�N�vly��B	�,W�I�(Тk� ���3
� 3'������씊�^�.�����b*(K�Is�x`,���x� �2�O N}'���l�`���@�P��G�)L�d��+��ַ�@O���'���8��^B� K����=�J��=J�;�P�����a��L�M�_��)^�7B؎P�����a�1�]��u��ڋg<űbG��Pq8eҶ��\yͼ2���hWN9aS��n#m����.��u����QH�*ޑ�ҀYQԫ��p��(<-̶ڦ0���^��f���?�"-�OF��xa�]��rb��0�u<�l0PwRˠ黊��xt��"��t�%K澎�8y�:Ȼ��dv4q�gDK�ɑtsKXH�H��t�=����-�泣�����홻
�:;�d�{OOϡ��w��j�'+�����0��5��X �!�`3�Xyp7m�N^tR�[�OQ�S�����%��S�?
��y�~-{�2$v�3�C�`�:!�@&ݦ=��<G䗅L f��n[ȕ�V{1��W�MM�X@u#��^db���rj�NT�{v��C	"�-a�k�����R�r^&�c��J� ��F	ʙ'e8'��@�7�u:�D���""��ıI5�#�f�,�S���vcO)�B�˼b�{�쀞��r�Sp�H=@?�:	�J(�,t����4�z-���"�;h'#P<6U3�A���yk����Nt�l���p�,�@�U�?��?p=g�A�5F	�X��+�F�F��-���dp�A�M�rqdL�pV��B&�Iuݡ��|1�&}����t:�0��f�y�l���[����\&
��-��}_�T����~sv��&v�=>
�)7t��\���o�"�g��>I1�P} ���RZ�nO�:|/�OA+�b�T*��
��Z@ ��B��X���!�^�V�D1�N�����kۗ�F�N�~>���ׯI ����>�"ì�>љ�f8�0(Ы��'�@��Nڻ�|f'�����\��dV�:��)�z��Yke�L"+6	ɡ������J���0�-i���4�����v+z�46g��K�ʱk#�&JꐼAa��$��5�0���8��H�Si6�wy|"�W.^�+�����,-}�cP� ܪݳ����(4�Ğ��wR��t��'!���u����3�F��� ��Pn����a)R�a��������񸁓Tg�Ϟ=��� _�\����^*��hH�q:��L$�J��{�k	#
�0zy�����4&��昿זZ�L�����.��(��/A�YwJ:q*����j/�#��n��Q0�)�h3�9O��xH�8��b�=�N&����	2YPJ�s�fE�E�2�e�TU'9s��|* �C�0�
��T���3���^��>}����β��}���$"��*����<�S�^K{�8F=��
<m���Lv�y#kZf�p��s�����Z)��x�M��O�*��^[r
g���G�^���a���M�k��#)�S�.�zi��p��J}��}�ŸJ��j�s��"c�C�>L��c��6�-I��G�a��y�q"����)��8h^F��e��AȈ)��\ ��8�hjh�y�1k+f�ene��un�2p�M��.1�0�!�yX~�X��'j� �'����(N����M:�c$o���g�O�#n�?�
ĩ4E�;�eY,2�I�cFA����g� `���i%+Y�ش΋�ݔ�+�L�Z���GO�<���5�m�iF�M�t";v�wfn��zm�)d6����d.P�t��gA|�R����Չ�c��z�~�a�,Ï~��[rM�En��i�L�A>�rI(��k�$�žr��o����-����=l�(���W�j�wu����������]�|�n6��lNt���>	��#� �-��<N��:|A�G; yج�uC7IC�����%+��j�C��V�j��R�sl���y������l��?���ۻ��v�T<��ܵw��T����;����B�t���DV: a%��S,��pe��w�H��s2�d�͕yj\SUu���┥���o$��;���_����	�"��t���;�ߖ�|u����_��;V/)��r���l��{��k6]���?>0���`����Vl �"r�Ta?l������i��b���mE��{���d�����|�7�р�E+w�U��]/Uw�J��+A�d�;�7r����	)J��cͶ�=y-����|Z1
��A�����k��y��O��-�t??��s$�b!����RzU�k-%'��eJ���W�D���#6O����X�	���P_���m�f \(+��ż���������;�?L��bY�Ǉ9�8��ims���0C�-z�-"���{��c9О���0�=zZ�<� r�$A�a1g>�"k�H_C����J�����"�$_�Ǆ�~?�VJ�%'����2s"qҤx=���#&�8Ū�M�I�����Q��Q�&�'�D[C}�$w����JTbu5Z����j/��A�����5�sz[ú�ѯ�Œ���A7[t<���1?�gC9t3�"�^��M����vSU޽�C��=K��ճ�?��?��}����v�P5L�2�?	��͂�|���߽~-��q��!R�l�y4�b,F[�fIpL����G"��w�_�����'�:8;��qB�S�`Ȑϊ�%��Az�1���������y>��a}�f`�
һpbmiG�s��z�J/唿/p]pj9&�"�F���R�,�5Y�!�i`I[= 0�$�}�|A��R4
�*��r�$<������}N�αKƆL�&��[��9��څWNf���/�;��t��tƈׁZX7<)p�H��j�G�1]�s�1��N��A���k�c�&�Z.R��9�ƌl����
��~�C���h �h��d���m�t|�NV��yHJBJ�CF�X<�i{f'S��P}'w�o���+Z��O_��g�~����Ls�Lq��# :��֎]wl%���D�����)j�#��b���6��dc�r�E��0��sUK���A؝F�9x咳8Vu|cN�FY�h��2�Vg�d�rz���rѿ� ��M��ڮ�����y�W6����~2e�Eҹf8<?P�4�ld�5<�>���£���V*�љ!����y<rn���w!�� O�'˳��4S�-�"`{�D�tϖ�\��+}-n�֡"�b]
��^���t��;jڸW���6:`��^ɸ-��Z�}��S�$vTq3f�-YyNt�%Is�ȇL.����2.(��(��:���koG��iJ���;p��.�__;,���1KncE�ѱEI���1�i��,N�G-�(�w1v����v
�h�N39����]Ҋ��@�n]�n8���{�a�`R���#�ZSpud19�1��jI1p��#o��j�K �,V���qGAV:�y�A(�s����ۆ��m���08�[��lH�-˔���ܧF�>P�B��hw-�2*(/���7�v���i]V������=ȍ���H���*^@�YK��	m���-�:��+���:�Q�R1F����<��GXd,�,����L�۠#��o+�������W؄�b�폏2s�uѣ��.D�<���IqEq>I/)��c��΅Q>��f͓��j�8(E�c�a��b�%;�����4�1͗Jt����T�Oâ��f���}�l!�89���/��E��ˀ�E��U�zEÙ\M |�0r���IA�<|���1t(�.�潍�P�BK�M��Ł�
J$���[M�B��ǲX+U�0ja���τ+�:����4�]����u+,�7�?�X�F��vN�nT1L���k���E����-so���5���T?��������O*)W�pu���-'�m��)���$"��e��l+�Ŏv��?�1�:�H�`�L�P�hǺ4L`Y�B����p�<-���T��A�a�@����
��Z�Q��`j^��w�޽z�����˔�oj�	��/��[�54�QZ�A�Ut����|K���{�9����ܑE1���n�e@XҀ���<@��h�b�x��,��3�5M{q�Dd:�sV2�E���X=/���i	�-����-��̔�[���@�R`l��w%��WŐ�a ���'2��؋��x��v=sNǢ_�6B�?K��.I"�}��D��iTV�ȹ�C���wXc\�*�z��YUL�$�T:���r�?���o�R�ߜ����.�,�}KP9��Ҿ�ӧ;�٬ǡ{�/��;�]�\Um. v3�;Hb�B4�f�T���8�ڎ%vZ�YèLH�A��	w���B/����۷t).lN���~ɸ9����Nry�g�Y9�'9�� �:d)Qj*l��N(B�g�(��1^'F�bp�S� �oK#��A�݂�́"A�I�xqq��{0V͞UPІQ�l��~�={v|��%t�1�X�%z�*H�x�0E�$Ǘ6��%e	|�*1Z�DZ/�7[,q{��Aj�xR�XF��-eB�D�Y�1�B��c�*w����r��9� �Ne���i��s&W�Dفy���(�Zz�Qk��:�- ��::@_���#�  W>,|�)0�����݇렐:� �[.紭���t����L���vYt`���a�q>I�v�ؐr�>m����o�Rl3[�藂��]�������Ӣ���J�J�i��X��\�y\�Cj���(�0<y�z���;�S��T�p�Iq�x��,��*f�������A�T��dT�M�����6�3+-]41?�+��)k�yx�8˙2�X~PR<1��4�;!�oZ䖌��%��G3��Y$��U &���0K �rF�'.�F@?� r���4`:�Q�Mbc�{#Ւ*f�P�{�2�0a�pH�E�72�U��-_�
+ޏ�������$�m���X[��p9+<��0�ۦ�Y�����b;_q)��˗Pȉ$|P2���`"C����� ��K ֑�FBE��ʓ3�_6{�n�Yt��t<?��SҐ��ʥ����s�t�dO*�)d��]MA�a�=�AXmz���@a�v"�e��GPÑ
K���5Y�_��W��\
��=/�z��:6����p��d�|䰑�F�༐l����I�[���/����%�!p���n ���O���(����&cO�V�f�9YC�7y�Y&�����٬���|q���F�B ߗ)�z,��,EPFP`Tl.`�tq�I�El̅�\��aDo�DQ�N�A��]�tiA�
x o��A^9N�:��r�N���v�WZj��M⌏U(Dy�T����������r�W�F 73W�@ �a�AN�:�M�0�l �$�����E�o�y�Z�͚s�c�����e�=�B���W��ɂ�L)M��4�_S�53Ť@2��8a]7��0��e�#��E=Ϗ���!hfz���P�݁4?b����b>�P?
�y�d�G��6QR��èw3(�"B��Ǽ�ƭ�icX��_���M��,"�#*�.�؜�x��_P=Z�����2�Ͻ"��zz��u2����Mcjl���C]�=�55I�S����hM>�I����єJm.QC-33��aћ��,��3�l��^$O"oe~`�G-.�ٻ�31�����Ο����:�ݶ�]蒋S
��V���
G�6���A�D-F@"������M#H^ٙy������;�Q��L��]b�
��`f�W�s�Ԗ+)�T��=��l�5Rŷ�M��=�\ ��r*jKf�}S�\^(ec��׮�*/r�	�=��|"�&H��xx�t��1�*-r�\��Mù�<(�ϴ?D��ر����.6����:gq�`��*P��,A��vrۑ�H�]��K_���_g�-d��.Xi���i�Q��T���@�U�@�"�rv$���̲���2!Otq#���}0�#�D����ΐ���}��ݛ7o��|yH�ru"�K�*�ɜg��؉��l�Tњ_����m
@��(��ǟ�kw�Z�A�O�LS������|V-�N��V�,!-�#���W0�,��f����W��~y���{h�y!���|W�P��_Z��cg�U�л�bRL8�~s�A�G�G��uE����ș�<k���K�`�T�n�^]�;��_�e9��� �BAk2��G�4$�Ⱥ���h�w��}๭n I�$i���_owi^�n6)��r�[K�s`N�/O:%��޴ '����-�fsF�Ai�}Ӻ}\�M�&�1�d%�,�Z[�\���Ӭ��.����,-H�z���&"L3GAʾ��!�h*�7��d:�-EԙOp6e�LH�g2�ww���lv$I�yע���t�r���#�ɴ���O�������X]Ug��WO���'%W��5��;aE�3Nz��	=�kWd���\��gi�qܻ*Y��j�ڳW�Z�΅��n��!�no'}8-�f����ry��2[%R�iz���5�!r�n��M����lJ����J�J6'F�ҜH�������������D��~�;:p�ɀ�R�z�,���e�3�U��~*
S�nh��x��t���]B���8V�$�e0���K%!ޑȠ�=�~i2�n�Խ�0EC���y/����C@�IU`6Ź�w^=}�T�e:�3�����>`��e:�گ�y�<Z��<���x^N������N���!p�����.��D���a���I�H"���[	���Ȍ�5r �H�%g+al����Q���P��Ƕ��5���Zz.����%>p��I6U������B��d���``��Д@y4q}/�3arh�ر���]^�������h��F�N:���M>����?ZS�68��Gco��כ]�6$����:��<9����wפ���Α���`Z�������>y��������׿��< O�e��s�Ihp���3�)K�J���Ơ?���	�٦�S��H�����I��uC�JʮN4��Nء�8/	�U����h��n'��.x;
�Q0q�)t_f��G %����'���>�ȣ� �?�s�嶥�����B����Q7���],GI�2��zRC]E�A���^|����~�&����5�e�j?$�4ۚ�m��@���f�[	�>�����I��k-���0�&�*7��tj�(.�g�����@2�y�B;���Y0��u��T��t�M'M��O^q�EwS|��c[{���a��k��p��>&2� �X��"{2^��C�Q�����dyiq��p~	�ޣt��M�+F�6�_Ȱ$b��0(>S�s�+
y�iҚ�s��N"Frx��s���k���on_�|I�|��L��0�a`
�B�K^��B,�0�s(�Q�I�~!�L����Nګ��o�� X7�Z>�;�d���HW~��Yҫ��L�eC6{�4�n�*�;�"(���m��#&3 E�e��U��BA.jy��f�R��x�4 Sh����s���"C�9�,LV�xU�I����(ɪq(�̧%`�d�H�H��kK��t�{��˝/��%L��Q	A�dP�´;5Q�"r�!�v� 1�@[�S��p��v��~�F�-��
�/�'����IZ��Ǩ�N�{s��$p�t�I�P ��TzE �J8�ƙl%v��B�~����=���T�y ��谯2/bZ�g0��hO��D��	錓����:�������dOج�/�D���I�=|/�~)�����T@GC���Y?߬X�,�ֻ���%�v�q�$�1!����\&ƨ֕���c���Z��o�yļd�8Z �$��&���p@��4u����[�;r����ye��-�M�{ܬ=���,��eX��aH3�>|'9�tR&����D��6��P�-u�L\'��!xޘ3A1�?D�X[��\�B��O�Y=�z&��g� ڪ�x���,�6h2�X��<���҇�0�97'�,M?%����b���L��n�$�w.�K#�;���,�����T�K���*����:'<�W���\��ߓ��}��4��5�d�,#o m��
�z%��ZH.�����+g$��T}'y
�S��A�»(.d*�����ǒ��6�fZK�yB��S�VWD�i&HV+��:�i����|GӉWܐy���q�TK�)�d����C�3���2Kw�F�vʊ�K�gPљ�v1��H��ǂ�&� I,YI#�g�J1���+-��]dܫk�*!;]f�,C����������[�-$y�x{\�A=�W�&�w_��&f �u�*7"{qI��Rx��-�5�'x��7�r���9���l�e!�-i�@O3(?�¹���hٓ�f�cA�+�EA�B����d���F�dH09��:�E;*3؝I��mM>�4�j�"9�A��5��u1ڎ'r	��ES}2|���sف�O~��F.�߾���9��Q��xA#[�k�Z͇���f�fr��Z�jH��y��X�qW�p$C&�)G񼓎�\�W�����h ��ђ��6�[��Km�]�pJra`X��}���g�����$@J�a�?.�e�'�|r$<�R�Sc����Q� [�{:[���a}�=��cU���F�8�
js:+��4�8=��vP���8�fx��!�l$���Ap�77���,��˙�?��?&�ip1Jg��9;1yIan��L��m%�ݘ���Ȯ�~�t��8c#p{HFc���g''?�я���7<%y� �*����@�H]��A(�
�G�4�Y,Y�a�� ���  ��΄,2���e
0ژ�W'���b���Dbpuu��s�R���8�6k�\~
�O%�Y�Hel.�(F��)�� 4Ӎ�Oʆ@Rr��É�?�9��F/,��'\�BY���?�73A���p{�.���};f����x��<¶ғ�[ũD�\�`~��j%,{KVYd�@)��k)�����7(��'�Z�gE @�>],�Nc�ka�����[v����9� �w�d "4h�(��ƈ�u�n9:�NV��/Nܼ�i0`z���Dr����[cz2��XG%�q�m��V���Nj�EZȄ����.-l{��m��_ɵ�;̤��������޾������[^����{�3�|<�|��pŀ�`Mia{��5�L�\�WBdD����5y�� x�̠R��Q�zP��6Zf���A���r�{Đ�"��,��<ځ�*B'��C��Cfq5n�Ơ�"q0�ɛ�' t��&(�%�N3i���e�k���@2�IBAAh-��2�o�7�lNu ��|�9w��qb�#�bp�f�օ�G���?B'8�O�ČN�޽ �Z��g9�0��i#k^�@�NG��_��B�N�P�Ct����o8W��[r�B@�G#��zء��N����;�3>N*��������A��q$������w�ٹ��emP�V|�����3��C�R�׃Љ��(�.�kP@E�a�/%�W�]c�J;�2}��r��4 }[��w�h����f8��Yg/[yK�Q�ࠀ_�Q4z��F�I@�2��t2�?��$Q�_�t� Oڋo� ��9�Jr��F��X�}�4%�$�b�rr�nQ�9��I.��&��Ȝ�f�D�����u����;a��;m�t�)37*�ɔE�s�އ:�
�'�^]h�^�m��8(���t��+98�8��?U�M�5PM�F�g+��pз$��P:o�I�X���D��oh�"'N�D��U7� ��B�%I~����T�zx6�	y�����{��\�6v����g����"A@��Bh�˴e�m�a���$�kA�����9}�J^a��ꁍ�T����06��oDj��"6M�2Cw��%��F�A: ���G��qv4'�����4�Y҉�T�:M1�FY��C�Y 3^��	�5�������u�w&�i`��ر�)87��`qSe�r���]��p`��>#��U����^|�v�Ds[F�o����d��Z�ѯ�z�K��[�ˍzR�M���h�MŜ����&MK�W�|0��В��{���<6l�Q����r�-Q�t�sfi�]�+y��	Uߤ;����̞���U��	ͮ�j�j�<�76��6h�z�X��ف|҈K\��鵩-�5�E��E&9k����"�[l&��)��Sf���J���ua��F,�}��?���瘭�-`'8�ǣ�(��lk84�{�m���0Hi���1��gk�x �̳H!�bT�v��z�إ��<N�p(5�p^����ܑ����"���Vy�M7e	�1����j�r^��k9%#���v'���@tʌ��श��{��i]eU҉8 ���s�j�s���N��n�L���<;HR���%�[�X���5���X���	A�=��P��_���+<bX��N�D�Xv�o扦���$�v�%d,Ro[�G�^�Mm�Y  ~R�1��kg��	I�D �����v�Ys�������4g�d�-E��]˔RE�����X�U7��Y��f_/�N�]-_�
�$;Z!Z@x����zWL�0�����Ƴ �^&�y:q�r�C�K��,IڦeJ7���鳧�9h��o���ǟ=�xc���|��r����a�pSm�̲�s�	����Mij�8��u�Y�����{E��g_0ab)G����Izzz^� ��tB�c�ti�n׷t�>���`"��$�=�G� ��C�ŧl�R;풐?�da@��C�
��p5�=�r�����J ��7�Q�<�J�L/�K$'y���̏�\L���b5����e�'��b{��ɧ�}D�:��;Ჭ��|>#Ol2!���޾���~h�d��0CW\�S��J$�۠xf����q*�^K����]\-hK�=W��NLi8�����Z�c��)Oj~@���B+��p���o~�����"��A��!s�M�d����a��0�G��e=O���4}+]$8��I�'��H����O�yy~quu��Y�����ޑyfn�U2�p���u�O��M��	Wzx2vo�w���v6� cH~����n|�3p�:i��kZF�Lz�t�ͦ�I�=7
j�^�`1���M�g��{&Gs*�]�a;�"�'O�n��)(E8-cT��I�^u��>�y�W��rI�@'��L�O/aY�j��w"m:@%P��bv<&��r��Vi1�暑a�$�@��ҡ��^�a�2�O�hǓ�+e���G�J���H�t1�n�+���m��G��
��3-��f�!����S �=Ɍ�g�Z8�3��Q���H�2Y�Ip���$c�2@����2�r �\R8镛�񌗊�']_5�zM���� �v�����3/]�?d�t󸾹�V�]-�������g�t���Öӂi�ُ�����]�3�cb 8eF2�,X&�Bɭ4�#�#�Z�����R�@�Z����J��R�I�N���al�,~g��^�j��9u&���@�m#�:�+��*m�-�S�'�6=�����)0�Ѐ�i��T�8��0������_C�!1� �lbO���)Zvnj���CB�H�ׂ��G�'"��{�#uD���$C0����sdZ#�W#�!)��$W����K�|驤'���ʸI�����c��= U�����UI�����ng��Eq���INO�XVB��ߎ��f�0�{Kjc� �����Yd���#Í���k������ҫ�GU ���Khτke]���Ƕx��~F^�&N�E��׮�LLv:]j���I��lv2t�<D�l�{�h>$ˏ�%<b~n^���r�b�4ڢ���m�׽z�@:jI����O��'��g���x��:�gP���X��x������n!Ҧwww��\�*0nq��a/��]<g�I�8�c>
S�}')�k��T�s�X��^��VpI2���ղ@�����i���eZ]�
�45�Nj�9��T
�1��kEF�#SE�e�E�<�f,���2'�i7ᥠ�j�D���N��H��R`g�y�6J,n|��&����f���	9e�`�����g�j� ʟS�'S�ʌM���妭R����#H+>���z��j��'���!f��FI��Zr�a�ɳ}��Œ'��g^ow{rw�|.�3,�<Ǥ�x�|9�=�b6�v�Z� +�h��n�٢eʰE��M���3��u���8A16{���^"�����)�h�ܛt
�oe%1��	�>��JM�����U�?��?�[
檓S�z3K]��JLDk5�fLgH&�JA�J�ɾ+�#�?��S{ht˄@C�z��X@Kx�1��x�gK!|+r�9�a&~�B0� 7t:�p:M]\�~s%c:2g��X}��$��f��!��y��� ޕ$�>n8������4}&,����0�]���Z"4�Q�C�<Yl����HC�m5�M��'��"e.�aCZ����<y�	ߺ���Cŕ�7_�:��\[j9�}����J`Ӓ������=~I'��^��]�	}�Ì�=���ʒE=�O��@"�@�i#��b.I0�Љ(�AF�$&��6���N!�A�}P�v����`À%�������Y�d(�2([5���!�1�{R�q��\�螚br���!U�k���)=�4՛YE<�f���p�q��nYs|?461\�q"�.�Z���9-�[Z�>A&h�nD�u�TkA���V�-/],3��`���JڳD �iP�Vt2t2?��r(�lk�f��h��l`'8c"p�R����(� l�2�#"��t�"!���������?��(�_9��.�>�X�R��
k^��"�⼳)���iy��4�<��螠����9��?1�hC��̖ݰs}�\�<Cv7�222����E��X�\:�a\y��c�g
A����$��|z~���(�����m����� �9�E-8����>�(�@�S�0�|b2������?$�x�}�P:�{�U�@���#N���������ϟ��0�i�d��� 0��_������q
^��)�Wu��2��������{��z&�+�Tg��P:jI����'��Չ�q)RlH�%r�ҽΖ��3ȉ��~F+
}9�F�dϞ=���~Bn�ry�.���D �L��P��]f��v�:�E��4����<}���<-Ni��O������Kr�IKH[�1�-J���%��;���S�w7�gR�'���3��w߽B�&��J}��u�ld�,�@f)@J�����Jl6- �2�����F��6�'��Z�@�c>E&�݁�*:=8t�����^��<�����@�����O~*m;lg�so^��C̨�E
-���}��4������'(�Y���-X5��&h�U����üR���_��!hu�s�Y��O��M�5�[s}��\��t-�qug2-��6�#oI�Pb�"�C ��*K��Ce��a�|�UP�b`�+��Л��>����o5���<���Ɵ�ɗ������_�����aE#L�:
J"�.Ԩ;I"@� �H�X�t�� #����jdr�و�Ú��"2�f��F����^�(z��r�D�9��0t�w����~��ǫ�)cj����C�{S�/T���Kوw�\�n�����6�^ưЧ��Ѫb�g��x��)8�n�\XΨf2�nƞ�����U��gA��FؽT\��:İH�f-�F�I�y�Emg�v0�@̚!�R��@��cGK�\�;q �����E"�hxW�_Z�1�� ��`μy�zvR?��"�) 9Q����q"��|Y�'-�0h'׿r�q�����`�z���0ф������>����*-mF.l<W���Z�N^�����2e6}��'��a|QfVǜ�lD\�����$����ɑu��0B3e�����.�E��$�'E^X��2���2���7�L#�7?���62|��?�}t�N�Q��c��yTC���/�<y��$e�������lY�n�EHx᱃�Z%K�_m���K!H@+3S��9�2d��3��m6q*���5�xl�������nw�#�W�nȳ�ھTN�g�EA�fzF�T2��!6�y����I&��a4�}`�.��r���o��p��ؔ[``m�G�C&	���y��^�W��U�����`����I&̴�q:�u6���
�e�08hVE@��F��5:>�J�� @�y�'�/2�|��"��G�����`�͠���{�i8U�9n�աj�VƢ�x����.�F�=�d�y�3���5y%/r�|b���w��_��p#�1S�cc�Gs�FYt�Lmײ�\�T���p_�ث���p@����i9�ĸ#&@����L!a��o�[,hkc��B=���̒��9�U��6��r:�fPL+~��ĵ�5�C{S�����<�d4���Ӻ���w{�GcA��*po�<5֎�*��FXE;�A��h�q�o߾�jf~�N�ԷSiL���8���|F�.6?��}O��˖�#z&���0�5�G�ď���;�;�H4W��Dٜ|`���<�t|�.�L����-�o7۾��4��[r⇎��t�����������^�J��/@��3Nf�/���r������ɜ�0Ho|�N�4'���@��Z��t�=��oZ�.�uȎ�[V"}]W�$W �=>��R����WS$����.K#� 2 �:&�g)Ls��N����>v����+�@�:����7�NE��ZLpІ��\�ZsƧ%�"bzEz"=���wP$�~�p2]��a4t��u�Ò�!��\��zezv�^��S? O�t��Ar|�x�8��E���X)�W�!�rOVS�mr����C��i3Qo̔D�)��J��U�}�5#��!����*�O-�My3h
2T�0��������TY��zsve�&v�� �P��#mi��������ު(GI��%�+�(I(M����n��霻-��bQ,��?��gW�t<C���]Ɂ��'��Q%��Qb���?��/��5�g�$���c��
�����lp<�������F� ��m ��&q����z���'�O������>�SQ�ݏ]1�x<nxlB2t������}!���svѪ�&��M�|1�><ܒ}���^<�޽y������/�V��ܹ������C��4�v�*���w�Cǋ�����;���d�,�Ŭ%�I|�� ��Y�IUrɭʳ9�m��~��gOI��Z��e���2�DY�8b��w���L/�Ξ?{zyu��2!v"�r�V���>P�F������0HRi�����˓O?{�ӟ|B�a��CY�4�)����\NAG�,�NN�%�����޽��o�T�t&�&�gOΏ��#��驘��j�O��ò����" �8�)³��7��I%m_����g1�vt��/�N1wo�:&��'o���:Z�)�[��2���!���-�s�� bF�ٹ����y\�j9]��N?��O����tuuy��GO&y!�2ONZ�T�G�"�֪v�ߔL֓����#��'S2��pZ�ǮN\vr�^OO(��;ڸ��1K\�����,�M'7����r_l��(���M�I&����o�tZ;��b�p���Á�f+��y��o1#��d�f�t"� �g3sy[�]ߥ��d�9^�..N)
b�|�ft��������(�����o8������ram6���z�QK@3,�rf!m������ϒf3x?L���$u���y������Wo蝛=���?�ǟd\Y%-(�3�SB'���>���Oy0�d�0ݞt/��6����T#��B/i��*�ސ�'	bZ�r�.W�e�l���ؠ5��@LdF|K�d�}�I�%!�t>��۴b�]�YW3�2瑱{��9�;��-YQu��EՄ��r>���mɥ�����۶����VcW푊�����eN�ͮi�ӓSz��-�{i:DVt|�p+��;6�6��������:��k.�pY�3j�0�!e[���,�X�<X��[_�h��ť���D�H�A���h<(p�B�\�f$>�=tjq��a�"^����PI��^� t��5D%�r�5�FD�E�:#��3+1=L�u��;
�������r�I���1�/f	�_��;2(]N��dZ9��T�MԱ|άN2,m'>e�0��1u���t�?V{�G�Qa^��ۼT)��SPZ<S`��Y����#���k�0�HlP0�>̱@����H�1Pw��a����r�N$(m�%��}��7H�!e�@�ɲF�E��ޚ�#8�S�L35� n�%�]�)��d.�i���)!��{v.L��8�N�x�h{L��	y8�H��"�#ૹ����_�䋟���?'�#�K���n�(˼X���[f�E|":{����^t�G=�~�2���T��q*��Fǿ�޹S rr��;�wnGN8�m��3�+���-��is�ix���s����	l$/�y��Z�����V�B-��)$3I��<fꇶ#s�;Yռ,��C�l��Y"X.d���H����s#N�a�� %4��ya1,Z��S8W�C�0�+�EB,��^c��B�Jw�Z9�l  ��IDAT-�ꠋ#�b��|~#. ��%���8n�F渐P�����XJ܆g�)�ɑs����������Ҫ#���aI�[�qHQ���x��L�>C��oѼr~z�`�#z����Xg �[��:�!'5��3�6-3h�0(�0��Qm�,��z��5�f\�����4	���r��dZ��S�Ѯ�C0<�x�F`�,�]f���n����m7��3�9T4i�$��q�\KN�w�M�*�E̦�$��ݞ=(?"���%��3��h[�ӔB��̇ ||Ǝ�P�MYN�쾹��0��BkP�>��Lwq�)��I;�[���-���8E�Ή�W_��!6��׎{Z�Ar,��d�g�(��`o�$�;��s/��c*�Yƭ4y��E�TM˘�4;>=e�_���jE����_]:-Qk�����g)a�,�:��ջäd��Y�K-含�샶*���#@̒�i�x���1�dB@�`P�V���
���)l�AiHt+~OaM�4�0�9@q�	�>_��|L�b�,�6�p<��@��tH
ߤǏ(�\d�)w�9�f�Qu�����i��3�� �k<K���s���euk%p֞�	=.$�����Se��堸�0���_�]΅x��bzX��Җ~B$�ꔚ�ԢSz�0��C��\%���h��l�C�)�=�6�" "˒lL[��ô�(*���Wt�<3`�YX�E�
ag@�"�Du�	��,��˼�1���A�2`4�
}�W^�C�4���+Яr�Nh��'"U���Ӌ������yd<��Ԣg+T���β����nH��Q���6}��D���|q�??|�@�*Pf\�fg+��X�A����S�N!�����^˨�Hٛ*�	-)��_����b�M��c�}��$��3�ڳ�Wtͫ'gt?Ϟ^Z��N^#�pL���k�pc��[�ƛ�R�)ʅ����F�Y��v#�~�f o7����@w���h�h�=�%Y�̏�_����s
�'��~����A�干�p�,�>��>�⣧��3ac�E��J���'��{h���̳��M������>��t%1��-�t`�?��*���w<��:PDA���T��7Pkp��utq����w��Y�NkBO�9��v��1A����zR�2r����4IPA���)s<�) I��O��ŋ�fn�N�A =%�i���@�syy	�Al4�l�	
T�|�1������X>\;�>�)�8�h���{n����x����p��Ȁ=`�[8@/_�̳�իW�;�]�J8����1���@V�$��� F'�d=y6�%i42�3��n1�1;���4?g������d@VN@����E#�^$���	w��&��D|��0��k�B¼X�ۅ;�m����_��_B�Ъ"����� Z� ա5��cmiAr���np}}Mq	��At�|� 3�h)h� ӛΎ�#\8���a�����K�=�CJ���^s�z�����ރi��G抖�r��$��O$�P���+�������/9�����'�*��<�#X�^Ȍ����Kic���_��t"0�:Qz8޻0$^�lh2B�G-d��e%��+��(���k�>��+�s�%;��Ւ�a�%�`�f�=�\�V�Iz�ZAiG�4�����D/;,c�՜"d�̠�G�yPXM�G�k�1�ۏ����D{|�������A�6�Z���إ�ݎ]>ՠ��q�%.�H�K{�#}��^ycsr8����Zv�<C˸�:>�a,i�o�(�;���Sj�
͡b-�)�
�� 4�JM�B3�L�*�ڎ�PMG�H�<�e�"�2���������"�9�<��mߠCu�E ���NF׭5�� -ב�N��,2��7��ق?��?z��� Lj�
�:�C���"-�LYsU���S<�j
��9�v'�vPZ�\U�#�mm��D�$}�l©ǱT��_a��p��c��Ɓ]e!�^�A�f�"N�
��0:��"�ʄ#B���88kH�ua��j�G%u<�q�^��뇃
�<�p�����W�f@�\U��I;��*�#�M�XN*hZ��G%�D�谆ң�a�	�u�X�����N�n��BB\�
\�v���$&Ed���9b���i�2K# ��7�ɷȝ�~r����w��d�p�Q~�� =
3Gvˈ����DZ[;V�jS�M[�*3D��N�h�R��A�P��JP���d�톢���5��R~�)R��E+͡�`���wNo$Zb&��y�XҺ~�����#r���=;<�$����g�n">6gА�M-�t�J2=i���&2}eШ��:l��p�- �	6ЅC���q�^;��#��d�|��tS�x�9�����Nz� �ŷ/����,NdzR���v���@��͜�¼����єc���YD�9��Od@�vFF/0ѝg?�ݛ���h5/��[w���j>+g�S�O�e.��^�q@^�>���\��ո��O�AX�z�9�M|����%t������2=�29eB�#d�m�@g�d����p��L�Kd�1"�h	La!����.�֥��Ch�\e��IB~�qbV]�d��Y3��!a���tu�h5�Q�|K.�e���g�y�P?�
	��c�Ҿ+hQ1Q�+΃�9/��� bs���5�֍�lۙ��(K��Ou�ۧLF��D���RƢ�b�~�<��N���xxu�C�CH���r�dv}���*ɴ8�` ���ʷ�:L��cơ���IZ#�]�I?ne���ɘ�0x:vDl��pV�8��^J��~����M��� ��w�V�dt	X<"D%G���ߚ�̀�"�u6�D22Ӊ�8JA���t�y����BV�c"�Ǥp'��\:���Zm-�xy~�sʶ��b�k
�R
�5�m�>�Ϻ��7�ӓ�����ׯ�����m"�>���.��j��uC?��!�Q�.u�jJ�!Eѓj}W�ɳ˳�_�<;�-��o7E:��J�}��sCE���g���byyyY�8���煉�v1��f�8;?���3C�����]�d��nnxvĴ�g�"HK���<�v�w]����3WW�'y�U�Iω���y�p�(u�$���s�4'��De:��0��a�&�t��X�����tyqq������d��'�$�/J:4�O��c����)�ɔUi��0%�ݎ~S7�]]^��������͖�krf9'�VwmWd�ޯ�N/8����ړ��~��n��C���������Y&-$]�d��Ȟ����HuRLsZ�L��2�Mr���?�ܙf|�U]q���h�N��Ew�z��������C9�N��jQo珷iMaUʭ�$ק�'��mggt�iO����)��l�֪�}>�4%cp�on"�#R��@N>���������)���MNO�����>Mzɤ� �e��Wih��[���������duG��~1Y
�|������\�?�Qn��LV��6�5�O�l��糳��)-�۷o߼������	^,,�\�㣥u�g��ݫW�����nΏ׏��L<��c�m�yb�&��P#r�<�ٴ�8?��<�(VO�֠"��Oo���	�^R�-�gd	���ԋ[���d��tF��PbJ�cI_�0dibU�i����~8�+���v��[����܁"'y!��NH�����t�d�<�a&��2]����W�W�L�'�X.�U�VĨ�^�'�5[ԥ��-��A� 3�#��W$�нۖ�j�a��CD�-3?�M�� ���BB8z>換E1�g|z���}^p�q�%y�y�K��Ւ'�_=]6�{��-�''���
�kr�fYf��l�Б�|���~���V-����;���������韹���˜M0�(���Z���9���&]�^o���t3,�<T�����F��yhL�+�t���}�k��sZ F:	�Չa��ʍ�E8M�5:+#�$�b�D�J6��	�jخ��h5���Q�Э<F�q����|p�$��<�����1ѫK��i�TzH3f�,|SS8زԱ�'��g	�N�9*a�B���0��k��ݥ����%��h��Sin����1*/��R��F�D��� �k*A2��l���ܣCw�����4�('[�n�Df����wYjo�q�Ԃ�tD��^E����h��@�%>�l4=�x����m��:��r���%��9H`�/��/>�P��/Oķ�oZe��_2��J�f�p8ۃ�ˤZ��D�����;��G:�i����2��y��|�k�ԋ/>��s��W_}e�p)$�P/���b$�Z�ҭ`[X��jL���!��A��w7����Ng��P@3��BZ���ͽ!�!�J|l�q)v�$񐻎\y���h:�c����G�tl�Dyu��PrP��ux���)%���˒���k��e���ǐ4�[/E�� zH5�PI�L/&��I�P��)B��$�CjXD�j�Z�!�F�(��9��A��H��t{h�^w1q��SM���Ŕ�w���`щj���'P |���j�"��V^ڳ�.m�t@�:s��o4)�)��ȳ46o�"�<6���w^ӂ��x�q�38�aH��%�`���%^�B>?�w��r��M ��U���U��vL(l�R�Z�*Q��\�4IX�H�r�'Y�{t{{���U�4#8��̬�X���s�ݷ�f��%VJ������`��G�FDX��+��cZpΨ�0{��'�΅�n� ��G�ƴK��v�3n��<����E��e1g�3�ubS,��5=�G�F��	Ku*u���I�̃���S`f,f�tBeI�6?x�K:�O_1-(	���� "y�1�Oƞ�^@�$9R.����vW�|���8}h���� 	'%��gui���)S*�-����^�������2@Βڤ#Eg��}S~��+��WL��R$�0��Xf�A���p��t�� ��i"0TPB�]�[J��n2����t��8U$e�ղh�1�M�������^3��4AJ��M�~X�0/Ў�#~���r����D�n�������Kp[��VH�c�����"���C�������� $r�6�t���E�h�ck	8��qY�J��/�z�{Z��r�Z�2VҚm�?N��z�h�i����l2(g��G�X�T	-do�� gۛ����J�@�lPN
�����m����>�@䋹T(5�X�����`/2p"�[��s�L�i��#[�e���@�Dm�$�5r���p�#3�:��D��2w�	�@�׉�
8����d���
3�"���tB�����mg��h;�k��)�l �UPT6v�;CW+I��W4�s�q�u��8ͤ�΃�x�(I\a4��3)0�
w�������X�x�4�_�vk~��o��m���qO���d�$��Td�O��9�Z��ϟ���
y��	�ֿ��)����Zry�� F�﹄Kj��1�x�g�I���ܾ�Cqb%-�d�p@���Im��G���$ʍ��s]��a�2C���\.�<���
ׁ�5I�/�z����I�n����h���M�q>��� {r�ytvF� +�
�|�x��方��E�ը��	]��jt�k2d�n�W�"�2�	}���ԆE���>̠�j�ˎ�|�1�|ܦ6R
��ն�t¸W	�,8�3����v
sqtL�x1ک����*��i'c�G�F<����B�h���N��9GG>�Զ�nZWG�Hpla�&鳍\j���t�_|����Bď������=�|��%�6��٧}!�o����X�Ldh�yQ�ⲭ��ճ$#L��U��M��?>�0 t��e<���7ӿ��|��f��=y�c��
ur��t>�J�������U"�DS�Q��"�-/��F �.�I?|��F,(���Uт�~�z6c�6���t�'��q�-��+?h}�>��͛}��1�N���k[	���q$I����+H"��<l8JiZ��Vh���I+���+n�_,R�l�E�(���f��<%f�y��в3����d��D���~��?��?�����P�C|PL^��l�����t��D
�$�bĭ/�����6��]�Ʈ5�x��G���q���8,毺Q\��)�x�v��#�vc@�5�!��?�(���$�M��+�������$���)sr:5�*�ʜ^�!{eJG8A���FǾ��0-�}�Т����:M-���`=����f;�0ӵN��}���$�V]ӗ$�&c�iv�!s\a�7^�,q�d��<ۗ��'��!�L��镬a[��aqG�C|$
�ʫ�FnJ7*OdT.�v$�B�V�s���B3��x�����V?�ltv3^��8�8�1I.� ��_��������.//��_�|9�x@d'{E'@K�c��� ,H�`=��B>�:��KZ�N�����g-�ҧ	��y����P{z�v�!���1PM�R�g��H;��� ���ǖw`�h��5+�A�4Zl�#�^�}� l�SN�h�{L���кO�QClt�� ����������!����qf��)Z!�	�NU�.,#�N<���\*�^K�X�����EyN"����!}۔�����b��v4(����Z��W�54d+Nt�AA��DH k96�.^Wq�)�?[.���ڹYJBV�
���j=�d�T�E��W7(�q�����яZ;�P�F4��0������o?�����Kۛ6I��b7�\k�ަ{�3  M�Q&}���N��H3Ap��^�k�5�+?~�{��i1BTZ�QS�q�__����m(3D�r����;l��K7z �Qȇ�ۀ5ԉKHc]�\����
s����I4z�tf'SgO��+�yj�[0�+�Fk��z�����,_m�s��(�����1Q�!�@[�,w��W������g�`���u�pǶ	�+7{��d�$*�4�L�_Nj��|)����_~�x���`�v�)]-��<C�XO���es�$�!���� 7'�W�S�r(�G�h|��>9�(��B��:��8)7�vt>���{B��,Q�����:�Kш��2�Ng��+-��2�0�p��q³�U2A���U�L�3����1v�k�.j#�wg�7C�G�R?Ka��s�1�]�ա)C5>�FX:��y��2��URby�^�	��r@�����.Nѕ��d)y7PX�P}�V#�+YWӽ�h2�̣�K6J�Sm�t�3���v��V�U)$���4�{�<��Rs�幹���``��b�dc�f}P��9�Q��H��ď���d6�F��n�驲ȡ�CD}��q����1����lD�ȴ)�ir�1�k��2Q�˷�[��P�آ�Χ�j����n�]�8.Ehբ%��� P��$ɍpw(nl�}p|��v�J�u!.��-1��S��mb;E9t��h��}=[,s� 4�:�0�z�;�"�Bﻐ�����o�b�PM�!�V��*'E6�;d:��ph��*��(��lz|4[̧3��`,k�B+cӪf������7�}l�f���d	�h�����s>�^��Uy�f��g��I����%ϟ>}�?���x����g�X��L�a�UZ̪���:_���Zɖ����%�c��w���d���T\�i���[]tL� �x����Z��g�&u�"�u��?Ҫ�av��<]N���.����i�I�)�j>	''Ӌ������Ȳ�!6���:hUZ���� (	9�NlNNg���K����>��Ϻ�v�XN=ztzv���'����Ͷk@oۈ�)DN�,y���=�s�NW�+�/^�,��D��J��B,�Ј1X߯��I�n��k�w��	Fb�ê���:.��w��ҩh?���9�c��GG��*�N\���a8EL�Rwç�:�`����}�3�3UhMe��D\�؜M�?6:9�%��ݛ7�&�mU��G~�?Y�eY5�����W/�>}��~��O��ǲw�me��%�����ٳ�g�G]���k�GS9[r֚��T��C�f��Ȇ?<ȕ_�x)rs�TN��W���Щsl�ա=7;�$+k%��������b������3�)9>b���Ta9�3Qp=��}#��J�u��ľ*��, �0n�9�G��b:YΦݾQ�����2�񼿹����
0�\�꽞Mg˅|��Ǘ'�Xl�r�y�]��I���L4 ��s��a��MUE���ĹƔ7�;e���6EYM{�����|�;����v��_�~��GZ�#����0fR
� �@�p���ۛ{p}4����&�_�z5�D���z#�<[�Ԗ�S�;%�>��	M^�����l�����~����eqt|Tl���j�V>�޼[}���?��o�~����woQ���)¡���~��0I�����_����U���˰ކ�	P[�w�rٳӋ��ۿ���o��ߋ���N\�=@�ɘ*�{�����z�������_D�'r�k%�Qi4�Ln}D6�d' ��h3|3c��ԏ/O��G鈤�+ȷ1Y@Yʭ�fZ+p�Iă��ix�˽F<�O��=0��ne�R?�����vM�����L����S%�9u�4�bo�𤘇�>��,������!b��B���&Yӧ �����I=K�C(QK?�VǑ������ �䉋<l؋ޛ��k%��M/ÙZ�ʟ�ϩ��P<�����O��F�WZ�Y6jOc=��^?B�Px|%��vز�iD~J�U�h<�*d{p��(� 6�@�1��;�����n[�*+=�D�췺��������`J-�)�$i<����)�hj|�RS��#�����H�
�	�Q�=p�QHX��ݭ�����կ~���K��o������h*h�ξT*N�}�Z���6���3s=�͂�j�#D���01X�h(F��`<������ ���g��ݴ1t�f�d�DǕ���I=��u�����EBj߱=�F�Se������|v�˅��!j@���CUeq@S\�5Y��vN#/0��^G�|a��U%~�*<{��ˣT�&y�����)�|3�T]W��R\M붖a��g}���L�cC����R$�;(�������\ٺ���C�D�8	�	OfC�N��?�I�K�s�D4H��N�"M���ҕ)�y���`n���K�&�/�Nw���U76��yU�g�
լ��������'Jc���H����7�?f�G5��]]I�}�y60�҂���	y����'&ono1���D"��O����:�����lZ*��^N���f�x��M��D�E�l������z�!�|\v�}+|w�=��Sϩ��b1H��)0(hRl^�Ph�i�&oh��(���'����،h���;��wo?����Ǐ�����Ǭ�dφ~yr\�w��O��ӓ4��ı�F���~��J�-��/�=i1��|�l>�Ҵ(P�ݬ�w=������d�@--��M�����
���yլ��N�y�ڄ;�v����(rxd��2�8F��4����^��x��@k�f^ӓk���V<�_��c�Yei����
���}���Үn&��`��/>���3�Y�.M6�W4G$3�������O�&?2/<F�'�ĭ�2����|���LԊ��`� (��KA4q���%�ܴ{-�$�av��d�:_�R��oˬ/Ǝ�AM3��5
�_��*ts��ew[��o�`�Y,ͳ4Mlo3d4ן�a�:D��S�]K���ノbc�*�?��|��ѣ ��L����E�*p4;"��)$8>�x@��z��ɔ�׬2��1RN���������C-+d%"%�'/�[0��zjZ�R����K����og�,���炣�Da#&�'O��y-��1]b�
�.�lVѪ��*X�r��8E(uf����,�m�˥��S�y��iaG�>}*���J������N���e��r%�G$R�G���]�B���l��Ã��v�e��Ϙq;���� �#$i���X���Y�,u���ry���z����(Y�b����m�u	Z�žȥ�aaT޽{X�Q��8uA�
����O?�$���53���RFF�>�2NS��>�=�z>{�L�VUnD����/"#חey��9��r���c�]C>�RF6JWH�������#�B��55�:cSf��F}o�F�j*�7�u;א�aٴ
]i?�f�ur=��5�zYY�vدZ�����^_�$|�ꫯ���%C)�?������$��t��-KG�E	����s���x��3ˡ����	l"b���{1�Ls�FČ�܃��yg�tr� �8�X1i(���������-ׄC�?��sy���GR�f�O��Y��{AT'�bٿN,�Q���p.ao�<��Z��d��䩏*P�{���k��`�C̑�tN4����3�E�V��z�;l���PdS ����H(') /Xvy����s�K4��h=6��@�a�Zh��aGB�0�#V�RMUx2��f���VB�r�}��1P�ך�	�;�<S_�u� k)�*��^���_��꽀�ޯ��Kk��ѓ�����v�����b !w���[�5EE(���R�4�7���S��������ﾓ�-ft�(�N\KT �!��_�X�2z��4ҟl�m�3Pb.��j�`$��5-�6f��_��K��̉J��7P������v�_1E������*;��k���d�᎖S���=�T��<���0{A,��񴦛*_�a4�āv�6�1�k�\�1��~>��:��A�V���G�q���L^<n�q�6F����`!��T#�����#�E�ǚ�)�`+�@�L;	��h��_�1��묓)�5 OtL�Tk�g�=�׻��U=��(��2�fww�aR�ZQp7�3:���T��D3X�
�Y�ԍ�<�kf�ͼH�(/�')+��@��]��"?|��7�P���o�I�Ky�/����[����ڔ�g��06.�(����釼��e��xw�* t����w���9�h�L����Р�z�0S�}$�O��@�_e�9 =�i� �wt&���ȪRg�UՈ�2Z���P�X�HG���Ꙣ�(�b壥��=�Eq�{��t�bL�$��'�I�1q���)�b|G*mFbE��
���8�":&�kus)��1��k��uZ�,��k*@xTu)jW�~R⨅ȓ��.d���	mde_��h;�)C�CHO�0����-�"W4���.�Z�a���g�'��I*k\c@���\O�I�d�<�5�^�N�6j����>g�a$C�l����Sz�kĀeI���8��cP�?�UbZ�3"8rf�L	g&�:�)[�e�;R�e��<>��"Xr�H��Di��t�SHk�Q�O�5��-�-�ϗ�`�<��g��ro�S|�
��lTT��5_n\��)J�����aD�$@���ȜNJ�J«��:�3�)����իW��9���kg�E>_^��IO�o�S����9�l؆���Z��]R`^q3�)K5.qbE�j-4����rm�-SH�@}�^<Ԁ�V��t�h.̀Z�#�E���JH� �ՒJ.Hɤ����Y�s�Az�x`<�AJX�<�ƑbV*�>fʗ���-f���9�\��QWǷN�V��9�m���c���QG��)��(�w�b�� �i,���J�7�1[M/�9�m�L�j�Z���~�6�v?�3U{ݳQ���#2Aw�h-�u�6����[i��	seX!�o:EeN�d��z�F	C�� �ĥp��m���\�T&��E����y�����g�&���OZ��"
І=@�wD���|��@1��.�d-���*�m"��E��ݦ]��mK���y��NC��؝�2����h]�44m��&]g�ڥ�`�f�]�R���ʴ� a>�dZ&�]��ˋ���'G�����#	��<�VB��&�*�Er:9PU�zY�y�����V3�*2(��W9 ���ZōM+���<��8����O����c^O��������M��wa��T��'�#L�6H��&5�ھ��,�Zt�t�d��U�����t�z8=Yy�V��C�G�s�a)�Y@$��ɫWO��x��Y���Y��t�3���~�M,&���eV�'gg�l��ə�-FE���>�a?�.�=9��sf|dq�//�392������/Ύ�K����J2��ʊ�q��n;�T}��T��K���/IwVSH�x���q�w�w]��,դ����a�ې
 ���3�L�$��a�Ub���M��7Q~ߢ��b�i�,v�KdI@�y2g=&��p�7���� �� b�݁R���V>5]�@�r��4�x�����-����.�(O�T��DDev��>}|!ZE�-q�e_��O��I���^�T~�_~����R���hZ�r?�j����N	]Ef�J�C�P�hH}���񣳫�Bs�:0������1�\,��>N���'�B��gO�ʣ�9��S���B]L�Z$X�D���`����|&�;�YT���ً�,8��'��`^G�]|@�S$J=+y@��8�O���湒 ��Z���Q/���>���\,��l�]:==������諸��8��X�ijD�i�v����.e�\tK��MěK�V0{He��զa�@�vf Eg�\V`mJ9���o>@��{���G�wB!�9|���O6�;+��YZ��g-���h�Xab9�Z�M���� ��«���Qݲ����a�4��5�ŢA��{o�6�~�]5����"��󗿺��ܯ�X@����[qmb�l���i>��Y���jV��fZ�?�aP�li�NN�~�_0-B��%^�lJy:��7�#~uu�i��<�nd�+d������3V{��V��I/�R��3��e Jk�{x�?'�+l샷��h�����^�۾K�a�8�7�[���e(J�<|7�b{�+�`ђ@O���)��!˛��u�ߠu�L!���n{EC%�5��p�4e�1P���0�;-'�-T�^��ƨH��^lw������U��^.�k�G�+R%��@�ƊR�c��C
H�2��K+%{�R����z�/?�o�����Z#�A�<��p����yVα�9e{��-�Ȍ�n��VOoFh�Q�N��.N�2#�F���<����6���~v�B	��� C���^�c��	����̦L��#�"�r�)cN�����v>l:�<��'NDOs�	:��8�����>%,�HB�;�d8�귿��\M>�!�<�!9��pO��#:������#YX�}H�A�-�>}���c���6qׂ��и�GU>���pJN�e]�m���0�®�3��vhM�O&C�H!� �#�gG��F�s���M���I����M�N5|�4M�s�Y�����O��a��zFs@	k�!-j6.9��� 7�U;��DC��E�&]�`�d�������P3��E����u��������]��j=��Ûy�X��@�o��?��o�
�x�z�`��0J�e����{g���h��A�\=ֳ�`e���/��bI����|-f � ����e���o،�Ț�R��#�<��>䇂�?v�d6au���h=�L4�1�	�$�0���
m��� g�?�Y��$iW��~c?�LC�T({5`4�I�o������c {�6��6�!��؋�@��ϛ�f��,Cj�R�`����	ܘ��[�h�@�Nm���F�aQ�H�sTǅ{�*�):�*�X�����U��+f����@.f�U��}1/Ŷ�f����O��
K	ptj�<����=�4� ��H���1���'gk�Ww�/^�c3��C[��6J��|�j� �8�ONu��MI�B� 1=�j�]���
g���Z� HKq)Tⱎ�}���UJ�gi�!�2tzL�@�Βy1�;s���g.�Yá�(��ߝ?�#��-��{C��jd?��^٠+le�h]��6n��q4�I��֐w��r�ȍ���h�cO�gV)�Te�����Cr.�$������������EC��90��!=�"O�&1/k�ښ�|
?��#g�Q��P�T4q��V9��9�ü6_@�#46�h�wn��b��A3��g�A�9�:�<u*�9D|b���A�oO��$zc�U/p�o7��.�?#!H�d�Q�C���V���az���]<�7o���ܫ����X$��O�>zt�� �W�[�d�D=ܯ�ef	�*KsB�4�!�i½�ʱBƔu4'`"�ne��9b���-;�f3�SDU�Tq"�$3R�"��:��
	�5�覅'�w[��#]^z��G���pO�Ġ���>�z��Σ�cz������e�4W����ިċ�;��:���j)����?�\���)�����bp�rAU@
|������tu�I~O��/�1���q/�b��0
`f�͛����sNe�w��Z�1�T�z`��� ê��܃���d���,�&@Y��b��}x��1�s��Ӊ�
c+�^�#R��ٳ҈��e~��_������>g�	?���%(�HόVM
�A�pC�&�S�p������vy��n}}}=�'��2�÷�aO�N�P��G�bl�V�3�1�@��.�:O��@P3��dwR�M�/�)��^��,�{�1y0lQ|��7�n*P��ܳ|D�R�^3X�咩I
�k�5���`���n��<����S�"FJ��&�- "P Z��`�J��L�L�B)0�,Q�rቈʃ���y�Z�Y ==��y�������}\&+%x�6�%}��&G�E�ʲM���L�L9r��Vjr;ⶃ�J4�c�)�n4F�ot �\?�6��@Q�ǟ+����v<����7 �Wб�6��������|%Z�5 ���-�E/�î3�丫��<��ꁵ9M{�T��v0P�V!!b��u��� 7�g�l�|�~X���������o������x�WR��vX�}�W:��ɣn�rr�\�Z�fM����NL��=P'��B�u$}�VR�e�M,$�y�q8ZR��:�W�7�\�ǧ��8��Y�؍��\jZR��D��u6e2Z�0�����`�v�JdfEMh���#�h���M�*�����.̴��t������-���|i������p���Y���>����N�ºw�4˫�p�6� 
�0v0�?�t�,|ah�bľ�c�AaM��HH3��Ϝ�Xhؓ�FNü����н�8ɧS�d�vs0d%����$#{2���ݟ�!4�~�l��/���E�Y�bՐ:�B6~fVۈ�E�����Z�x����*�������g�������_����l�C��ڞhJzU�Ƒ�v͖"!e5D��& /�~C��A	+W�op~~)��)�N9������_�U����I���_.�E�����ٿ��c�����H��f?�֠MKD��)�����a��Eo����g�5sW��E^��w��#L~�����u��ɳ���7�~����� ECD����zi�6�>p�}N5�)'����kM�+���|Pe1���t3�>�.hHU�W�E =L�kI��?�0kZ�Hu ;�V~p~FVjy`y'G�Z3P�X$z�[��,z��Iq�h�P���π��4D$�k鎓��;�5]�����1�%+�^݉����g�%>#w�vV�R�x���'�q��m:W�E4��L=���6�@�������'�S�h���A��S�%��8��:�o�n�g֨�u�/%g�����' :W�ۢ�O�G�����/N��炏&�.:Ah�(���@?_���{��Jc�(�� 䴪̻��b�Z���#yp��1
LY&.�l�!��ˬ�~P���]���`Iy���
_�~D������
.%jP|-+�6��7�!u�3�8�I�&�?u5�$2���2�_S���PQD2W��d#�G'��JN$Ѹ-��C��v�bV�ճ�Ϯo�ե��u�|��=��:�L�6�y��/g˪� }r)�}�J���v ��x�9ўd1�`�H�SI�D��I=����=�v�$��b����Jy
MLk¦�6�b�y�0WR��ZT {	���j`����h��v��MD
tdT�^�)�=3�"rUݨ}b ��H����eU�Q��%��)��mz�_�}<��j��i-�W��,�~�b��pW4���d��iq�6�ai6�4f� �B�&��:�m��P�y�1����Q^EBt~4��k$��NS�͕�O� �t����)U߉�����^�>����O���x2W�l�3>($�Z2-K?�&�l��ݭ7(,�p,ኆ������"�ۭ��f _��������r�YS�r�
�GR�7�6��r���PV���@,Ĥ���k��׳�jNO�ճ���Q��{�8��m0s����+i=��q��*	ZZ7��@���D�z�A� Aӂ��k�,9�jZ%Ϻ�W(�٢�~�>�@����d1��8�2�
/��G�m8�L��2��+�x��l��Q�)���uj�M%��кV'�f��J��]��f�F*So^M�8{���|Y&:X���‴H$Hb���t6��*��W���
e�g��4I$i�J9���g�*_��ibY�HL޿��bE	�'���XL����b���"�전��6(�ǐ��K�x7iL�q�j?�ʜ�c^G��@�(�You��B��1�:>�D���>�/��J�Ǐ�xxefUy2���L�wzx�?<���ȓn��۳	臷�{Q��C�!��d6-���n��l��E���Y���f!̋R�c��g��SQ�C�w{��s�S�I��+�yح��e}�~�~hz�^��Q��yh=:^Lgb8ڡ_L�}��m���D��yq$=�G�v7�}����ˣ�b��D���?�@%���AQ|߀�gO�'Y��o�jR� ��o(�0k��۽�٬o�v���t9�E�=�<�M�g3�%�#������K��.�6�e4	�.//�v}s{͸`ӘM'�RV����a_T<�ȕN�J��6"�bϢV,��s��j�6{m��˹��Z�&�q����C�/BWf��=�O	�*Ȍ���˗����Щ-2�mr�@��qNed��I	����v��b�~�ϖg'�P�m7��4ĦRVE������z{���FeH��ڡ>=��V���I�u��2 M$ֳzy��j��H�PM�brc��D}h�I��O�߀�N9!a�� HS�`xXa��n(m�~��/w����۵��"�5^6�z�
�вK�c0�)�^5j�|�ܹr�EY:1"A:(Xlr-�C.^�$L�E�X\h�U�I���@9e�t��'������!�U�0�����w�G����7[��hNY|�("��\��m?%���߽����w����Ѿi�Z�R���c�8�Ϸʽ�+h�F&��Hr��qh�+po�v���̇�W�N�]Y �N+�٬i��E�)���KۮEX5���"U0e�k�>qrW�g�0^�����C��-Q�ȗ�3�qHC�)�\g�:_zǱץ<і�EL�r	&���aDb�,f��U�Fp��2��(5]�����#�=u�Go�8?��+/�XZ%�!�O���0�w*~y��۞����;D���J	Y^Og�-�#��~�-A
xž�{�+e�AL��(�;�k�3�Du�R��\B�9�B5�^��!+49��ԩ=��NT+�ۧ,�z�]Cp�sL�o����&�STr���������{f�!�<��DE�kH� ňY# ��J��Y]��{��f;(+w]��!K�pz��jH���g��j��f���z���������(%M���믮��~rt���w�����󗟉�(�+ޅ|D��ŋ��b@~)�̚���Cb���5�����K5��fXE�n�)�V�j}nXŜ��`TJ��w��[�W�L����{�G��� ��t��ԁ�%=ֆ��n�'e=F~�����������o���\�������]f,u��X�6m�b�aG�b�
h�|�JH�]�"��x}4?:>.�s8Z,/�/^~�B,]�ET2�cFĶiAqqQΪ���'��}���6���X�bʛ����]c<좑u�h��T��Ɍ"_�N���v��}�c��Ê#ݘ�S&�G��yV�D)�[�b�D�F6�hF��X;��r�8��b!���~�n�(d��T�I�+�Hx��VC��S��"��T��|7��O��#���- = ���3�0�iW�J?��LQS��*Ҝ��(5'�L]�����-"��ݺS"<Y��3��o��o2��0P�ڒ�P��V�m�ʁ"ᓐS����(���n��#�Y�<\��2�rtyN��\��u�<���ysy;⒲XL�7!{3��Y�!�`��p ��V:0%�ʂ⥠��p=;��₧|�C4�DL3#���04�E��nUr��m��"�-�O�g�+':*t-�@��/>��0(��w8����^�&�G��d8(�D��0��%?�&ܶ����~�~�l?|�~��ՋgO�ДOFL�q��Y�0j��y���n֔�J�f��-T�Km(��U� �/v���x�|Ye/�,�'���u�����IXY���L�Q[��F���P0D]�0��S(�?d����ִ��فX]V+k+�"]V9# X��j �`�(.b��z'����6��0�|�Xㇻ�����O�>�RLנ�ο�����2>��ئ�!A�Ps4+��V4�����v���/�s�����r"-�O$K�P�i���Rƃ�U��݃I25��Wq��X��ĴE����pJ}Ϗ3�Q���%���Ts������Y>��R0�Un��C���������3�6Ǎm۪F�D�ΰʞ�ό���Ɓܸ�7{h�㣣�Mabr&��xg��
;��B�I�l��q���"/[���O�?.��o��o����w�P,}�1s�+���g���Pqtd����F��պ���W1��G��1YŽ�M"m������#=K��	0D�$��8:�rB��YU�!���T���K�U=2qо>{���n�O����N0悡6g>�ɒz�ȵӓ�AzN� #��.e�Ӕ"��|uv}�G@������|����D�s��,K�I��v���#a�����
݊�B.�S�P���}t
��S}9֕N�U�(?7���Ì���+^1�߻˫"���a!޾���I4&1x*c�7?�|9��4�_�:$k��aCtAzw�(K\����Ĭ����|�]�'^ �dE4����V�\Ύ8�m>�<�1�5��$���SA5A/>���O�>E,�s��Mug:c���̗w\]���t�=�.�;ʭ�LÛ�����+z �8gH���舛�"L�o�7�����p	?}��K���izJTc=!W���7���)9�n)���Y/�w25�QK�Do�!H�
��J�Dv�w6 .h��.���6ŵ����Sɉ���w����.az����/�6���A#\:7��sS8�z��f�>�\����g����y������[Z�|��"���w��W+fi�ny3,��b��=��V�#�lJ�F��S6^e�:WV��M�xs��9SBȵS���䪈�l{@AOT ����D�By~���-����!e��SM n(n��Ϊ�z)72?Dz��g�*4i�����e�;���+S���^Dӑ>|`�	O
�#yE[M��0v[��(�1�
B;}ٹ�LnR��pe	����ؚ������"���3L�J��� ?��r�fG`�|��Ų7r�/�Q�?X=?�7��(ģsX�8sUF-{n�o������d�!3��L���X�����-�n��γK�&�E��]7��8y~ʍ;M*�Z�y�j�����|�f������+�mn�G���l��q��2�䤸��Oޏ�
�,�h�ko�_w]�[�
6��Dږ�� M[o�e�L��,l�ƟX=�o��Lj�"��4J�F47;i����2�d.�~�&v�����0..��1�뗗����o������/..O�<y�2~�{�����ANvj'@p�����IE�;�D�ypw��{EU���ыQq��*)��GJ�O�:yR��t�W5�y�IʼZm�k�/��]�f��?~�蘛�?�c�0�Й�X�M?j'Ry�XW�J!��_��a4�~�mD�}x���5z��)��B�0#4�|���Jd�;>Zr���KtC1���5�#M�����N�G|X�	@Ό�*3<�[�����PiM1��a��v&�?o9�8��à��!}a�Y<I�{ (�5�J������pk[��g�-�(���!�1�̋Z93�Q/����6��r�Lu��"�2�4O4��|]m�|v�g�fz��M{M�F�+@o�Q�[��t0��z�@�C� ��)�����!���o�*�����U�s�in����g�N�n�xd�Z_���8�@�Zi�M�HU��@K��S��M�5��:�6�q��6feƿ'��v�2B��m�s����σjd	�<�8�D:��Í�&/^���ӈ$�!"M��j�	�M��Yłf���+��J�v��L+͓��՟��WM�� c��I�`�ln��;W���S<<��_��~EoŊ�����f���46|���aR�ˢf��,���Q���6�csf�,�2~Eˀ �(�"^��30����Bj�@��W�4"�MۂŮ��$n*r7��oP|Ӡ�� �D=
���H4#qhz@ �˦�E�Š�N=u~�7���r��K+&����\�����0����ϳ6/c�J� Hf:s���d|�|#�M��T��(V�[����n誏EKd��
nQ����|�m���D�P�9�{��v�L&I��F�����t��Ȑm���ɮC��z������)��~U�sr� �H"A%m��TD!2T��(W�Q =�2�s���c��r�����]w�f���}�^���ȍ�q0�w�Q���^Mg�ܮ1��N� /gs��	E
D㍎�*%a�i5/��$��u)��N���@xi{�L3��/*��:Ycz��c2Q�2Z<�@蝛����&�FC���6(�Le!kC���D�#
BT|�E:gz���W��t�6ϴ��	��w�A�#�O���g�.ʆ{`dm�o�L���	�7��~��Y���\?f����qM֊�Wi��E9)�ߋ���j�t"���&r{����ۮX�W�)���F�1/0���p�8�{K��k�<�ZX���u��q�!��>XWWo�O���6:QT(����w,J��h�q��t�6Bf�V�>چ^�Z��-��L��&���8!���2m��s��@���?q�����ן7���œg0N��D���E�+|�Y�\�wʭ1�T�������v�q��9a)�`T�	,�1ţ�vdtvJ��ˣWHE�j�"Af��OQ֪�����Rp	T�^�$�T�߷�5��6�^!e�
C&&	pT	z&e����e�Mj�Jk���y���@�V�n�$N�T*�7�4��hQ�p ��r��EeNi����({9h��b�n7�U���&��]ȃ7{6 �H���b�Z67�σS�P�
�z8�7w�j>P�����5��R�Z�wj3a4����1
Ý�x{'7����N��8����f�f��G�)�WԙR�`���gO'��_��_��'��/Ć�t���^\������P��]7b43��Վ@���,���,K���};�D&��W|H�D$뙄1+�\f:��F�a���C�8�M[<�r[|���\D<rN'��#��
k�dw�����'^�N��֔�[(r;k|L��fI=�t�N"�&�G{۾}��͛7�}~�^��{�<q�"��#wys���!�/��w��y�n���)/k2+C?��s4_Lrc��S>�0W�8�	:��+��݊4嶧��NO1��9�δ�y�W/>u֚,:�+����������8����g���:q
�jl��q��[��*C���
2���E�~8\p�v�����#�j����c��#dZc1Xg�t[m����� �6#GF}�h¦�SeM͎6ʍ^��A��(u�K�q�Kq�u�5F��P#u��S��#��͹;�9g�8�x�
��Zb�]Lhdʓ+�;�>�d��Rh��e���ܧ��X�z��i�̨!��=z�7�7��ū�O����ϗ�D�{q21�|<_��8yb�Iv(�*>)����Da����b�LY�҉�2�wI��6=5�b��SXV�	�T�ԥsevQ�������]�mU332x�}�� ?��׿��ֽ��G�b���iO�+͛�yP�}7��D�م���}��?�����O��+�3n�E}K�YZP��{��nK�6�R�?�\���:D�w쌦�ô�Hi��� 1,�xz,��
��|��m�r}�5`���a�i�E�O����ŵ�)v�Û�g�HL��J���pd���-���T�c>Y+�L`4(�Ȣ���0�>aY�3�t*���R�z�b��~v�&L��ȭO����*�yOz��#v���>%ǭ�8�k��%��%�O��������W��2��G{��͚��^+�׌%��Q��r��u)��37!���Jn)�_Wnvi,�$ �>A�o���dZؘ��8P+��c�+)�Yf���8,�`y�Z�0�}�%��<�{�݈��ف!Q��{��߿�����w�|����TxL/3"��́�Ѧ�������H�2G����V��NN�g?=��Ƣ4�
_���x$yмD�`-���-����<�&�`s�p����~����b�R����6xb�@���2(5pD�KH��@�J�0 y�U�O��C-��j��4ѻ�l �iO��Ų�Z��5ؙ�n�� -��;�ާO��h�����nv]`�Br]{� n�Y�?:�+�Ѯ�l3SZ����3�1GK%�-P�����I�O[�/�y~)���6Z?H�z��Ǳ��V�a�����0l࠳A�SdL��i�蒳å��MÂ5Ee��<)l�]���n�i�	2M�dW�5[�e����"n4t�̵%Zq�6����u��>��sQm-����4�yj=IWRD��5l�Uf|������B'WicԵ2F꺪�/sg�`�	���٭^�wmN��#�Ol�����y	#���;�.�%	V�=R�e�o����G_,��r8����޽��3jN����.	�+����:�KJZ�i�2�9�fL�7c�y�" �Q���/u���ga�/36��'�����dW���/1A�P����[ �LyT�&M��'�j��o���-����w�b��� oأ���|�����#O3�A�W��%�����u<>�;I(m5<������&��s�4E7�3���FP�w����C=��ƀ��C&O�� u8�ȥ./��5҃T��ۋ�We�r�+&b���Ѵ�����6DT��j�����Ex��]k���`�M�f�9�6�NEC
�"U"<9�ܗl�KSt�~	�'!$�s(���٬�XT�D��L�N;�T
nl���n�="�P�0HHg��M]��i�U���k3�����O��R��Z��9�x��Z��}sOAݫ���&r��Q}C�f�<��G��VL�sAh8� �H?��D�p�8��9�׌��0^��<�؛�LI���@Hl�m��.�zK��Dwp�B[�g���w�F:4����9 iŔ,*ZÛ�DI���d�n�������j������2�_�I�����ڻF� !�7�����ɥ6(��e.rfl,�QøR��5�dZ�7� �1s�ܚܪ#:@�@�[�U�%���:4+��R���ݾ�W9���=�Cn e�K�]�ɾi��Lמ�-� Ģ��G����'�ȟ��\�e�aD���ӽ2��z[	�A�<��\C������E�=���@�"J/��Ϛ��sfȔ!1P��ea�
s��>ŏ�`��Ƙ����V�ˍ���@}^7�+�`���\j���ܞ����`�0"��G�;�F� �C�!�|d	�.ANzcLv�<@�/JcId�=�p������w6P��`Y�B[S a��c�\>�g�O�k���X2M���cY��5�X����`@B߾�p�T��P��F&ŗ��Pl���ɣ�O�<Th4�{��J]&�_���=y�}��!����
�nM�_�ܮ�7�7������d��)�aQ�r������t%�Q��23���v*��B��[r�w������~�u:.�W��9����&W �1�$Z��1�w���!7W�8���;	e�Z���P�����g�˂�}�V������+3����V��`:����UI[ Z��:��P�۫��6G"I^xO��W�į����)f��Y"89�*{5�EeD���R(�퐿�ƈ�Ѯ��p��9�#5+�x���,��X�
)k#T��!60�Q'4�m�XV�v��9���Rߑ���'Vz�!�!)�1�E�,f�_��%���fLF �h�i���0K�ϯ��J�99I���MP*���d��oDFS�&ɒ��n��Y��t򉻎nhp�L��(*�{wVZ��N���=�HS+���u�_�$]i۱{C�L��B��S�e\�6�3��K f?�NY?��iםpLHu�HP7�uu�n���cUu��Q��7����h��}}���˷?��4���Q>�õ���LqЄѓˋ�ϟ�={����7��a���q�(ߞY�����{�c���Ƚ��C燺��4X|A�'(>�a���!�w!����"���iqG���)��M����֓Z����yO�z�&�T<��pbtꛨҥ]���[�$���x�^�Ѽ��`�E� �ͤ�S���bח��/��,�Ta���"�Y�� �lE�\�Q����-M����>�R�Ņ����'fG�M+��ZZ�)�@��߮�2)�Wc��j�f���w���U��ov�Ό���۫�1��A���Y�n��H��n��"`5C�GM����߯�S�ue�V�V�-�����JI'�'T����Z�m��~%�^]�v��f߯������^���r�N(zԛ��*�lbh��c,X�f�t�m�m��(�.fXV)-ud]�z�� 2�M���l/��~nc��a�-�V�rSG_$��}f��fT�Zi}=t}��U)��������߃OA�*9�O���uRO����*o�����[qXW `�S;��N
�$y�X�J�w�`��*�᜺qH��7�Ι��uY2ң���uksl�#;2i��=�.KU&��	�-c�l@�b,6��w� ��g@�U�}ꇲ�g��S�����E�L�H	x�m�_i�e�t2�L��<��p��xH��oums(����ׯ�P~�={2��n׍xp�̸�o����߾�}�'j5�:���7��E� :��D�*��ܺ�<.��أ�0>�W7w�Wןn�o)~դ���iB�y.�P�![#��:�B8wG��S�uP~�L�"�V��lD��7JX��w2��Y���(+�9&��}�Z0_�����𶬎�Op�nn� �tڔ�A|Y�<���G��#����P"9����;��@�g����I��D�,I	�m�=�sz{���ׯ_O&3��T/U�eʩ���ޕO��#�Ъ��'��A)m9�q,��Lۻ���r�A<c�Vc~*H�����ڡ�ʕ��3^���Ug�\.�ٮE�2�'*�2B�Y�&���Nk������M[gI��W��[ֶ� @��b!7@+�'sB{"���g�lzt�\m���� w�"�_V��_m7�,�ۥ\��S!'N�������v�k�}�ψj���z���y�č�i�xd65�O10T����	����'+�ا?h�X\&eп�p����;?/<�"F�a�7�5�,s��D@�������T������8;��:`�Ӛy N������W'�����h�T��岨&q�`ҟ(���w����o���n3`^PT� MW��x�v�6X��J���lb �L/
0v��6�5N�Y*v�������v��$A�yf Y���Z�ғLv�Qe�EcZ��%^%�|ތ;	x%.�@I�P��e3g(�*�	�����o��%D�3�r�"��`���lT��-5�I<8ݔ֯0�y.KB���3��Փ���[T���'O:f
����ֳ���W����[Zg�gv|O�aU�D[f�3$��d�9�������b�,xb�)�0JZ��x��n�wN����NsS��'�l���~e������?�u��gp�7ƃ��Vg������AW��|���E��r�J����-�L�W@s��NBg |��~�Qccgh��@�|?�aT.��-UJ�|���
O��O"�.�$��U�0�nnn�"��x��i�URE9��&Ů�{��[Hڠ�G���6{�99��pb0J�g=��Q�ˌ�µ���5fP����O�V:=vh5P�E���Q
Z8B}�eoN��m��!��6�),�Vq���|7��(��Ϟ?y����ř,����
`m��F����E�g�<F��hX`Y%Y��S�xT�n�(q��^!e)a��zl�@
�������~˫E��o��mV�TX4r���q-��]��
�7^�����?�1:*z�U>j9�Ѡ�7����[&��D��$�˜�������Z9��c�F�ĄK�h���bmw��HW��0���$�Uu�*j�c�ݦ�$?�E����,q��j*�-�A�ǤK�-�e/)c�e�xrZ��!�x:��?��XR�>K��4L�ã�Q�(RI[Q������bm�.�q���޾}���#>��oū�n�D<��+��7��1��=�M|�Uhc�An�@r1E���n�m���*d{�`y��Z�F��A|�N�Xю����NPBo�O�3#��T���0mR����']�|�9��r�_~������F<���[��Ԑ!}�����z�Z��)�P-�����,W��_~%�Dλ\��nuq!�c�ܽ�r���ʍ��+�u�x��;�}w
�B�Y�F�LtAR���EL���t�&"��m���y3�AI��R���r��*�U�?�}����-JM�z�a$�a�3��#��S5�`_�h\i��˃�#�eG>|��s7���s��aC����eEXah�p�l4���8�iO�R�B�g�+���K��
��x�򛝦3����S~�Cb����t�|6�w�Y�T�www�&���>GjF�Of�򌓺de�D�)X�d��Dt�p��Y�7H��W��$6����_Θg�6#��<W\�`�j�*�ɛ (E�������%�\�<���������Kg��@�Đ �4~wg�AI-*���'Pу���/�e��:��/��>��TC�[���(�}�G�D��`�q�V?�Dv��7�ުX����2m�����R�4�r�S�e;���g>�yƋJ�P�	u1��5AC�4j�F�@�D�c��Cr��6�%5�>�A�6�~\mp� ޘ��f�{���!NǤ3^���+�l���};��!�ZM�R_����Ϥ��Nj:���f0 `���}����q��(uŒ�b
��ߺ��3���7�-#����O� ˽��׿!���7��O�$
�&Iw;L�/3ά����F/�����h�k�1v]�����^�R;Y�~����Z~���� ~]e;��\�F_�xM<�NG��[�D�7}���ey\ҢϘ�8و��bV;=��[�M�{	��޺&�ѵp/�s���zd�{FG�!_:K�Q�����Ç�f��F�r�����S�G}E�u�F�/�֛�j\�p��Fг�~�lafV�g������3-K:z1��]�z����e��q&��3�9Д�B�ޜ��s�,�(�<+�)�(�OO\L�]��...滩3���T`R��:1Hp4��	��E����.�St�Ȭ^�hm�G`�x��\���p�Ć� O���W�4�9�:�S�	�zB�	ڈ�X�)�]�S1F�x�����o��߿����[-�g�{x,�6;���0�A� �.�G���F�"n���9K��Q����f�7���Ϡ7�6�6R���|Di^��A!}�ๆ�Cb��,���5��3~{w���kRD-�s ����G�GO�� X�u�Aw�����C�L��|J�-Ҧ�H2Uߦ!Q��!�Be�� ����r  !wM�&_Oxy�(l��ke���t܎�~q�/Ii�9��ӨT���@��
��5Op�Z#U�`�{cK�{v���̍���
W��7�d��C���W�چ3���C�t��3�Jo�������AY;������I>��p�՗�)���(̬T�s��:��ˋ��Ѣ~�i�䨣��e`,�H=(荡�V�mGH9�d�|�q�	���Xi>�(:�; ��ޘ���K��#E�a�HB��"��S>.gA,�9��o"���3�����L]*�P�'�*zk44�	�ʟ�7���l���Vn��t�L��z�!j��[�%�F��.
��zFY��y��<���2aaIf���+��@6;�+=����I隔,�R
����*f�h�ִ4�N�ʕ�Vn��4���W����i���5���s����M���?3�j}uu%K�H��\}QE��S�3+�P���5��CiO�gg����H�!�A-{����x�
�z��x�������=u��7H8�ٺMC�
Ҡj?�t^�H�`9\3Knh�:��TF/���h浹�� �I�YB0F��~[���2Ѡ��2��yX�(w���5�<܉��Ɖ�����_ŉ#-2c*�"�9̪��>ev�$�Z�?ѽk�����p,6�2P��{0������x���6��=r�,͗Y�'�Z�M��0~β4G"3Cl��TE�+P3?H����㯾�J���9���!���9�����xd�>��$�G���u��2������e[����O�����^�&��w1�`�[%���U�{��g�Y�lX���-�R>���H�oǅ(n.K��y�l�Z&ʹhB�U�E�?���9�vԤ��!	#�-�@�Y���a��M3z��'��^Q��n�ͦ�gg�Y��"湛��������w.�2*�&�C��@9��޿b�>l%Z����O�g�OD�������v�'.��*�B�lQ��Y�q}���w��13VZ����X��5�S��k2��NdT�ܒ��V�邏X��:�P�G`^�~x��?���x�U�O*q¢\�'�O\=�����x���ܭ�� MLK�D��F�a�~�٧�_�������n(�>�M�L��M��l��P=$����Z�0k�u�,j"@���0��7W��)^�I� �U���\�lͬ�#����H�\�ڍ�g��=�;�*�ĺݽ�n�O�#\__���F쨢/O��<�c1�#V�!��^E�\ѹ) �J-Q��kf��^@Q("3u+��f�\�i,��[��CGI�����)�heV��m����w�v��F�-�37�2���J��!K�]Қ^�_�!nG1�:���8�����q�mכ��~��&���yYWu��jGŔ��&0��/��~'f Wd١�y Ƿ��$���Ǐ��n�n����E<t_���L�*q�Bę,t�������<�3�*)��������;��(Au!�������������Z��ɷo���f�m:m�h��ݶ�^?�gUS	WKoqŴ��@��5����R��t������T����8��L����FY�v�����5����a(�|}g&�`h��[A9���W�Q០=ͪ֨�1�Q6N9O�ՏJ�<zLj�b���6��h����DD��@JԫI����v'�#��0��2 �:\�C^G�Ȕ�<kyy��Z�:Y��İĀe��3Y�I]����W�<��!�lD����i��!$�$�Z��L�� ��Ti>�,�9A�� ��&�E�WWF�.*]@��֭��tS&�2k��S2X� �p��e$̎�kw4y"D1^����/f���㓣�lRm׽�ۨNR��DV���*�j�B�����|�d��P�FS~:ۧ$�`UO7ww���5͛]�����g�� ���}x�����!^\���u�m��~�IV���]�;U����b��Ц;��y�ڨ4c}HX��7�����|/v�������䊲�;  v���=�UXő��S�	9��1�a��C�B<�1���t�Z���4�P������_��t�g%8i����2ϳLp;��j���QY�fp�<:W���ǫ���Ƴ��#1��V�d(�%ۤ��c�\�n 4~�Ɯ*Q��`��tnCs�^�i01y�%U7�pe�z�t��b���{|�2�A�'�|�t��!�q`+� =��b��p���Z;6��q����G�ňsyl|��T���@��C�8��>ͬ��+ɛ�@o����0���������.ɤ�$�0���2�ѐ�0�׋F��j�d�o��2�>���#��7�K��8���f�f����(GajƸ��.xv�V���x6�b���t��gnc+:�<旖�D%!����"d���At�Dݗ8/�lu�a,ZQ�&S��1'J��믿�˿�K�[ �2Zd�Q{p5�����o5�����c&�i��'�e�)&5 �<y���3�P�`��Yߋe� ?6ʞ����� ?P���I�]���� ��ʩ��_~��f-~��({��\���h��䒀Q3&U�k��.�{]G���'�B<v�N� çR�D�EΦu�e?z��X!每<� �k6���-�
>[�6@�#*�G[(k�e�#ncY�'O��+0(l�j zq%Oq�/�2w��EK�"xn�R��[�>�0/��X.�5-R�@������`D4�;g�`E�l����h��y����g�N�f��a�!���T;�	\5�J~"�v�� �٥�SR�bq$� 9Šk��Ʉ-�������ū]Χ��U��^^x�#��W�S������%����iZ�yIG, 5S3E�;�[���̿��3����7W?��Ӈw�[9@Jy�Dd�
����q�v̢������R8���Ҩ��$�<�/���f���&>l�<q���� �Dl���J���R<ꐐ����6�����J�bH(�Q�ܵb)�\l�2M᝝��|�*C����ӧ�߿e�X�py|}�@�Cb�M\+O�R�0��C�^��\y���՗G��u�����i\�Zl�a���*��)�m�d�t�+�6ا��=���0��A�����>��C�	e�����ݻw��Nq�r�4C����Rڛ��]�؉J��lZ�в�<�ŉ���|2$�p�R��C�k�"��˵�C��:�)����.�Sm+=�7�(�t-c����m��kmј�ظpN�	��t�΂�Nq�}���J9r�ʬѵb�>}�$��I�-�nV~�y��ut��cӑ��o����_�e+%���ϩ|�%='Kq�W��by��ا����/����ļ�x2i*(1>|����(�8�I
�j/�����V:@�O���S�#/s�����cpo��]*������0}�(�=�Fߧ�O4F�uZO*Q#TƦ'���?2���n)�G�g�o�`g�>��60r�%־Q����uK�o%�H/H����k�l���*��(:)�h���[R%[Ǚ�'�'���ӛ���J�r��ß�j�:ȍ�]`E^���߈u����$�fB+6�3��|���A�.��ɯe���e�)	���h��`t��;4�̡s��Dҕ��]��@d#����
	���/I�A5 ��o��9�@�z�̔Al}"뿘�<3)_^���%;����؏�-9X�%�^�>��~����+�����?|+���7��*�S�������Κ����b���|K�2vZl�����]}�aM�WS����/��@��c�&�����F�����Nm���?o��4q�����R��so�Tܻ����$�ܚ�Ʒì�rMl2�`�"u/R�*Kq����S�%ʘ,U�f�%�$��j��Տ?���Ig���oid���xA>#V�� H\X��|��DEۍ[�����`����J�X���B���`�\��F��E�&�z�;�:�
tH)��[P�iVi1�9B�Aم����~+)�H�Q.d�hF�#D ;T2L���$�Gʌ]��T���x�_\\�6���΁�p�� ����o1����3� �l� ����g3�X�� �����������������b���7C�K�'��`�Q�����FS�(�p�C���rj�,��h̽�(6ʤ5�+�'��}d��:��i	ϡ����A�Q�qjʽ&[�vs�I�jh#�5�'�hx�|RS!Q�lw@2B-�v�!�!�m��������D�Z &%�*i�hJ\����}�qL�8�4j0E�"�������I�8thJ]Y�J�%�Ȍ!�S�b6��F$�5`���[�z�!��w���m�|��{c�<�F�Eg�J�|��i)�<yZ5~o��֦ak����W��ef�ϱ�88x�(�끘���w���)��(ő���N���ܩO�Qm��t;(��)e9Z�c�� �!��%�8�5�0���7�M�|���8��
�z�u�]�[C�[J���ٛ5I��bq�\*k��m�@I��d|�3d��d2��..��fz��5��E�ݿp�Ӄk�$��ՙ'ω�����M�������������8V�Fe�0�f�R�#�����h���)�{ql�|��cM�t���o!�%�^��
�:�]���EpL�(��O~�%����/���c�'p��e�rw�� 
�^�������G���+:��pK���Fz�_~�s��Q�'��Ύ#J��05CaV�2d�^�zuss����Wx�i/�Х0�2,ǽ迆$ ���Y�8��yZ��h�0g�F;�=ݣ�A�F�nI�9
i�ha�U�%��H�-�[����R�s�8�r[?vKD`�9롱�겦g �R���m�0�r�$B�,-���_�M����x��-o�L�e�!dҼy�ѱ�0c?�K�7���԰<]^��Rx�R�>,�S���0�8���P��:��r�8htI���	���k�)�������d��P�
����x�|ޠ�����Ѿ`ר�`���z�]�N���M7#e*�(=��P�P;�O�-��93@��=%qS�B�gQ�jX~nt
�Tȶ�����g��S��@F4�����/K�@�NӇ���|�M��h�l�0���B��p�1�&��%�9�Ov[�-�P��0���UU�/�*d�Ό��Ҷz�����0�vЊFf����8�*���]�֊���`���
� �	�F�b�x��eO9�$_���s��~�j�鄫��C"�kJ
1&Ea�N��O�('�qh/�S�xL��z�m���D�R"U'l @!BȄi��C������w�>>�g垞���ؖǡH���=���1H���K�o�-�?-Z����oQ�^��w���!���q��o�v#l���^:N�[t0ue^��(��lo�����I�����ͻ�O�����ze5g�PӴ]���Ezܶ��E�8�� �u�!�W/��6l
O��?l8{������������W�gt.ga�nw����l� h� �m�HE=��KMf�@!�P@��
�������9�9@��"fƒBc¤y
�bt��eC7��:��MZH��f��<���-�,O�������͙cG�3k�	~��������΃4�,�¢��x.� �r�������ANj���rL4T@�P�87aΦ����+�,�	=)AI��`n.*��6t�H@��x g-U�<�L�d�����iw�28Hrp/�ZH�Zd��Tt�.�a�o������_����}� ���^d2�+��dYg���;�"ɵ�R�R��i���J�{�'}��;r�x�Ap���zG�U1��ŜG�
�-�`�Hʣ/9�a2e�+ȁ�w�+�tmeM���6�k��؏�b有�V3��Y��;v���e�݋Oɝ ��Ka1?;.��6žF�����:3g�wΚyt0:h�D�i@���n#Z����=���
{)�S����!�J���U���2q��-_P����߬�8ԉ�J
X0�A���;t��O�<�!���d&cY���S�&��	�%�򊳂T�|y^���z;tطBi��p�V��Ĩ��₿���?_�[��3�4:�#p�}WO�����ɥ :#�Iw�m���
����	�#��C��0ώ��<�t�ՅX���~�������F�ii��`&�z)�5LQ
B����O�<�^�\��<ʾ�Z�l�$sl�͌8<�K��@��ƈ�.ELǶ�n�;���~��N������3�v��^���sj��/�W<�e����圔���ש�d�]�`��AV�eS��H'�c�q�q��6̈*L���O���A�9���r6�i�dV��Z�f���q�ɰ�C\.V����nߵ��?R��s*�8r�I�ooo��{<;[��R��!�$��
�D���K%��E��,���U�����19[u(�?�^�zt%�E�C3=C�ZK�V'@$��
�EV�4)7 ���:�����D�񀣝,���F<
?�>.uJvh��]�1ޙ6ݸ�zE��!�TXkxDlt�\ݴ�]+�=;^G��a�C��/�JVu\�+e��c��a����HW
�с޹Pp��d|�>O�0�W^�#���j>m��d -��q����)���a�� Y�Ts��6�U2��Mȿ-i��kԖ��HgK*���b<I+���,>�š�t�#�&��^���*�C4N�1b�΅F$�B�a%ǝ�sN9���;o�Is��|D�2�W��+�ݛsy/`�-p��u�4�b-s�|�)q��W����]�7��[�c�|�E��C�*�Qf(/�Ga�+8����nK�c"�ƴup�H�	Ͷ�3Ȋѿ�9KL�ĸ��G����82�Y�i+��þ�3���A#2D^jH�Q;3
���/(�muP��pbIK���"�Hg��*��sNa�tM��^xEi-YA�+ s98J���=���/~�����g�9O4�eR;�]�>}�n��5��z؟1��Wr��ݚ܁���W���C��2I���vM�t�r� ��ksl�؎2o�xI��Т�:�}��}Q�C�+H�3�-hw��l�����.��"OD�E5}u�J�xX����V0�ۻ;��q/+�ݬA�DeAo#6F冶���Gk�)w#��b&k>`��hKZg-\G�
����栀#��iT��Na\��l�	!�P��[�t2�
�A�=��Ӷ�	��5���ę��Ȅ�sLC��m�- 1���|;@k26���I���y���*5�R3�e� �pКѷo�{:FB��yqdL��Ƨ��E1s�C�R4��R��^�%H)�i��]JH	3��ބ�{�|xg����ᩮn�`��$�F�y�x�v�����9}/�Y��8(j�O��ȳ��Uӝ��#)��gб��N���LP���fsr*CY�#M��#�q��C
��L��������Ҕ��9y{�v�L�cnF
	��d�HN\���Z���>˜	uu����8���ճKK�V�3��ryБep8�<�H���=�2ߡ����a�%������\J��8�� � '��@�Ӎp�ȳ��}d�8&��t�i�� ܀Q�1���u{mD�#��$'d�����fu�(+O~�������P�WK��Q_~�zu�P0iD��ن�-�b��
u]j(x���wn�[1&�$z���2�O^p��I$��2�m��6�I��D� ;�<�/!"�[��/�q�6�+�:C1M��Vq��劷�I��=r�L��r���bu���i�ڊ������sQҞQ�d������'�p�_�-�XPc���f9���><>�S%�rE�i�,����H8iAP���o�0�s ?�MP�^��q�t�W����#��~h�kiAo`�!E��p1��$R��̧�mKs��LB���*����f���]@|����MvM���W���z�G�=M�sm�Ŗ�t��I��ѱ�:�Ì�e��ʠQ
Wg�Y.	�!��9�%Sj;�ܣR����m�� �d`9�isB�"	r��?�N�A�N������NY��/b����rH%�w�Տ/�/���M*3�YJ)�D`�a���+`20h�#�4ݤ��N�{�@,V0k��x�(G���25����8I{���4�=E�Ep�?q���e��EئO4X9]�\��^HA!�{V&�٪�|�����=7�J�A��hg�,re�#�p�r�+p� ŀM	��%��*�EN��%�A��Y�t䴋��9w�(� � �y�����dGa����QC��c?Q�Wj�U6�5�B�������Y@������f,)
��a @���hV��F�0$d-���]0op.�hR���0����7'�j2=d,9FuP|ʔz�)Soo}�y�qp8�I�C�t9�F��&@f�W�
��3̈́������"��p�v���p@L�<'=�|C��=�C����S��g_
�h�L�I��D�y<���!���ĩ��r���8��a+�5�����C�W�;.��DHr�Xj����Lra��;�i�Ʌ�����[�%b<Q�A4�d��3c� ��y�5g�H`�:�wk��88�r�E�Q�+0|�NȾ qo��h����R#�)g�xtY� ��¼^ǣ�2<�0[Y��A'���Q��:��RIa��#��yID�17��Z
�,��kS��|qV
ԗ��ln?�ktl=��=vV_.VN�`�阶�lf�E���(b�zl=��ϗA/R�M��eX�BP�0myآL��P5��s���N8�h)�rPb����r�	�.�z�AD6z'��©�"jJ���xA�m��d�
2nǨ�Ե��`1-�YKDjD1���B).�<��4�5|BdNK��i)9ي����3֜��m�^��lG�2H���)��]�^,	��i{GP�N�S^�^Y&-�g�p�0���Is|+?W�/x��ÄK!i�����Ni���q��ЏAi��(���bQ[�-��똗>NF�@lJ�b[�������k�2Y+�Q�d�����
�}�:aús^�|������_�my��ht}�����{hf�,�/�.]��7*-�����7���s҅�>�߽{��q��Ջ�|� ���MD� �a��̟�����?�p~��2;d��|�L�6f�ӊ3�&���-�'F�����1������5��v��(�5>�w,on�q��36+S4��i�.͊eށ��$���?�i�]�K1p��~�;�1_�A2=u�	z�?�o� r��ʨFL}*�ۡ^�!De���F�i���B�^�x�n�<K�]�v�ab℡����#.9t.|�5�|�,�dP�����p�I���N.b�,�:0��"-RV�)Y� �a��p��z����Z�	�g.w(��%�V>*a@f7����֔�N^@H�ڡ5����2����l��22�i�B�Z'C�/�qe,2Ȭ�D�g��1H�C:k��ЦL��������%�O�[�/��h鎋&����$4/	�A��jVXey�+�\�ڴD�;Q:��~����f�7A��<�k<8�9�[<�}V�x`~:L|�t�[���ΐ֚��ְh�T�L���1���K�b7��,��v��Ns���p���e�v����U�
L6�B�J��c����!�б*�l4ө˛VZ�zٍA���$e ~���u61�8B�D�b
�� 5?�R�?�q�S��D�d���ʆo�|@&�_"̨W�nM���LZ�1h�����bu����v�1�0Ƣ=�C��`��n#�����B�Kk�R(�cHC=2 7�������nf -�^�K-s�x�yW�I�}dK �ucGF�B�Fw28��藒�֛`8������䚶c���*E|�]��C�s�I�u���$���x�6�ޕ����&�(D/�����<~�hj'����(�0J�'O�'�(s�_(3r�6mO����oA��Y�k��Μ�Ԩ���$�a���aΜHsa���s��e%��=r8�8�	*IQ���9!�I�Z���P����J�ߒ�O�H��4�^N��@'�5�L�`f��`�N����|�8��L����ݤ(���[�����&S-�H�#;?H=`I-��+gQǠ̃О0cՐ��7zPS3���X�o*�M#I�8�z��Na��7n�.V��ց������п�T�T���oT2D��؏ÞO��%�ѭVd�I����e!���$�(h���@��٬�n��>mWTu��j
�S3t�ʪ�+|zP2���|�pN���[$f�"�`A��k� �.HT%}F��<#抒�,3�J�hf��R����uE� ��r�?����ぼGN�-���P�.&S��Ǣ$g5t��R�K��.;�3/�ι���a�F�C���:��_7�B�;r�y�@�0�����z3��(g>T;/��ɑXe����q���q}w�ǰ�/糳�� ������~M���hyy�z�v<�����.���=%S�x
*�%����vU����~�����]�F�����#�����4��n�jB�*9J�^'�R��@��_��P|D'B�q���GVnw�����91v�������<m�1n�[��?�}�9��,����@�=���a�������@�F�<��O���P@>�W�5R��[&
�$t-O�%��l����.�>����S�Xȅ�Ȱ�ˊ:;_]U塮?9����ryA� ��'zD���%��ӂ\���]Ə�>p-M8����	Nz�.��§�[�0.�-�l>n�ݲ
*�$HʭߨK2X�gxMG;0�d|�X�/�jHO�����H�WҾ;8�},*�\����+�}(h�<�[c�,$�G����:Z� U�z�9�H#R���1m��e��r^^]�I2�)Z�$_���-�c���T���^��1d0I�iB��
���97k�d���m���'V?�?���l`�;@�Z�`.KiF��������0�!%:
�(GD[iP@���]�777U�a���ق����sҪ����N<�
�F��:�k��D�h1�n�NrdWAg�Ȧ�B�橈	%��$l4�RG�.;��`�h-3�n��~0��<���BG��jɣ���^r�X2��Q?�ƵԒײh��lN`�pe�Q+ޏ����sp���Jg������������Gs?�<ح�"a��k5KR����$��4�5Ԇ�d�9�A��ނ/�)����X(36Xv5j90L�3��ZROʴ�X��A��ZRW~��3��L�A��p@!���0�;#H�'+���wf�,�j/4��Gz�o~��b6��k>GOLd����p�鸽��4.�(Y��*9A�̎J0�������:&t'L�����EX�3@�NDF�.9�W��-�������!͹���g�u9+� �!�`N_�M�p�'�%̆�����p5�����HW^�ξ��W��\�C\I��?nכ�������Ǐ�)�����w�wH�ҝ|���4�`w��ge�\�_ض�T�ȳ�g��
<so�T'#zJ�~򓟠FBw���'��X�Ȍ���q.��z�}�a�Zi�nw!YAz)l�8�:k8ImrT�7�)8����^;u&9���e+	��!�dg�u��>?�"d�ȼ����u�K"'�K�k�+�>�wǮP��ϖO���$�.|.#s�*{��~S\A��^{�$�w�Z��%a��I��jd�:��)�m:�akJeM!�C@��e&%���QB�R�r�:x���:��+Qr8ȁd�xW�-��Mf9��/����;j͛���+��U�98��`�E�'���֊�cB������܈�	����΅Cp|�*��;�
��J&�����s�J����#~@M�|F#;��ɬ�E��Q|�j2�iˣV2���������.�P}�pC�Dnw�t�N�`�����~^ov��LΞ-
e�6�
�K��J���ET>���X)1iN�^���%@�s�3�1]����5��*�"'}e�3��rˍ��ڗ���B�@���~�d�ر��p+�̞�b����oK�������4�(D��g����<ω������b�mU�m���qn�2ү(yGL��������%��a�Yx�;�9RmBg �O�'$�&:M��\��!��lb��r���)$��X<�r���X� <J��8���͚����5+O#W��,�y����1��Z��8>'�B{�&�O�� W�sau�-%��~!�o�m�Ŭ�ɷj���;qp������h�)���I�����M�c��YI�K͹�� �8
�����Bˆ#�#�8��Bz1*�����#w�e��p��Ä(�ݙ�_g�\�υ�ցVR]�<�Zv<���������M�X:|�S�H<�����b���bQx�"���HO�s��ɞ��/� ��!X�C������j���JQzG��X�	�.��$�Q:.���9y_j�}�'zp �-�'����Ȝ�. {pA`�B��9�.�:��`09�	�F�vj"2^0��d����x� :a,'�Q�pUDFm�H�B1��xH��6�̸���|e{�/})��9J�X=<�:���И�/���q�ub�s�����<8j�X{r�i�(�3Te��=��w�k{I�,�K�+z�BɳH�<�>�_-�
nz�[�Vk�N�SN�;����N�H�C	YU:&�a�&s~�D���5ܖW6NJ�t��\#.�"h,8��2�V��r%�����_*�ȴHCD혣kb���\C�s;���A�jV97��þ���9�����T��b�x�gB�����ѷ_]_�;D*�K %�d�l�� ��g�� p�hY����f��R�9��KuK�B�ʔ
i�+���k����P�iqn"8��=���Z\��Ĝf욥ED���𘑑'1�����Di�@8JO
i���,iY�\���)��Ŝ�:&=��n�4jI����w]b+���(��QG*xK�p�G��	)H�ʹ;v�P����f�^
J��f��]뙏f�")�g�(2��R��j��TZ0�c/���LK�ڂ���8N�R��E�b�1��6����	g0�-��q����6t�=�K7e�'xC��h���P�F^f��(��(L(+",h"X�i�3�2W�GF�Ԙ=��#A�Qp����G�,��ښ�*�Y	$&��C��~I���*����x��35�?`Uho���,k�&�9\#j��4��E����[��]0����͵[J�G&5h�$c���0f�~�;M��>�ω9^Ð�����&a^P�M7�N��b2ȥԡ�v|은o��1]�!�u�温��MCzei���^a��|60:�(d����-�c�I�&m�OQ �H�W�`�i�l��,�#����/��o��o�^�^;I�D d�5�r@�9����w�޽�"$�!ל˸�"+)�BY�� x�����<�jŽ�d}x2{Ɇ��%#�����"�,��D �1q� ���{��<{py�/��/���Bj���n�?��_�}���ݽ���&@��~�M�^M��4����)$$���\�*�T7 ��cK�|�ju�����W_�Wk>�T�+���{v-���L�`�P�-8�����='F��)���	��q�tzuF�s&����+�Jg\�/�5iuV��L��@��#��OTG�\xc���굅��V�0���� D{z,3b$ݘQ�4����?���5p�IA���q`o�3�	�$H;�9E!C@��aҧ"�M�g���UlZwLd�������K��p��I�u@'l6��ċNi��M,��LG4�c�7�i��ͭ�鈧�K��%ie�$d�T�s� �yk  S�k[2;�� �ڍ�%�p�&
oh5����{��9l�8b^�TB�4���%�νk�e�,��$��2f���yѵI�QÉ�}y��?�]Y�wPZW����3�]�r�(������@�����A�?��uʁ>5)E7Ihz��9���@`�s�H�u*��6�4L�AP�q���������_|An�7�|�����ֽ�x��bf�k�Xh;COCϓ��ѭ$�]�Ro����+�2~�xBr�dCX1=O���j/Q��K�� ��𭫲0�
=8R�̡`�\��#c�x�T�k��^a$}#��U=�8��Y
L;82 �=�C�e2��aGo��J��c6%��eHSS T�-7�2t�Es�ZNy��*%&ޞ�F5�S⎇��<8�6�E�U����'א���m����+0�o�>��C��=��K'=���ep#�$˚du/��*���)~[8��'u;�L� 51NG����ѣU��H[ZH����Ӷ����d��%m�� ��������Ե��������f��F���;;$й9��R@19Z�9Gk�՘�F>���3kΑ�:�o}	�OA��cb+#��h ��=Ud�D���Y7J�U�hR`EL'xs�F��A>y]p8N1a���}4�dЗm1<�"�=>�J��6vZT��n�Cq�@�iX�b!L��ئ0�9�>y�x^������vN��مtV]<�� �;(�t~>��z���~�����h��� �H1p:;[nv�>f��Ud���H��b�N^/���!�қ��ٹ�?>�ϗ�i��N<+G�$ M���y_�Z��l�U�����e��/�g�����s�^v�[6
��j|ݞ'It<\���ˊ��N���q��B(�1Rx���q�Ƈ�`Н���n 7��ϙ~����o޲�)IC��!�=�2x��'�/΋�QiC*��;zX����= ]��1����},���>R�Ys�+=ɩ�$�3����6H�'9|�_=-XM;;���V��z�c�[G;�tC��4����B%�%7��)��r�q���������B�|y����/��V����z���j��[���>=/2:����?>l�a��nn)׮ls�{I�PS��O�r1�𓢃��XV3�sG*:��xw�}��x4�=[]�苎�h�E"���䑉eߡ�f6[R� ����������Zrbk<v푤���n����!7�Y���Q�3ҕ�ggu�`;V�5�T�۠�EMw����8Z�z��(�;2I}�����3��6k{�H],�yn@��l����L���h�Y����Cє՜��ٮ�B-~<%�-6��n����#�F>��\p�<��wB!���:ՑIlҡ�8�!��*O���?��D����C"YB�<�����ࠢ�I¶�#�<:Mp� ��	]?MZ���f�=��EBI~I�����3��{Z��.d.���{�"3g�C=�^1"����b�N'-�쁟%&�J��&��R~��jy�S�E�"&Iڝ�e�"ڛ��CF���3���2��$2�@%ޗt� �s8�a��3���
ʟ�����]dH��>s5��as�N��eaQr�f�� �#���Q�#���H��a�}�Е���eQ�2�C	�ikFĜL�4�MS�i!W��^�K� ��u��0a)���-�6s��nR�D^���PK�:[))�~��ܕ�Z/���u�u�Z��,4!Z�t��i���7��ț��Ǐ��}6�#��>;�7
�E�,X�dD?It�t�6�R�: ��d�ffa�8)/��-���Qy[�
E-����*akPA��gO�i]�Ҕ��m����~i�۳�pN��tq�2���0����w�7�{�~�4t�)R��OJ���y����*I.�E��`So��ЏOO���N��݀��U5Ph��--�G;�E��h2���|1����� �[�=R������뎂f`��Jf��~^IϲW��R���#�5M��G�ȗ�������|�|��x���2�7�R2H�',�8�A���"�L��2���ڊ.���S��Zfu\Ҕr�l2'�f�| B�v)X0P���&��s �IVZȐ�O�)�i�r�ܬ�ygt������l�g@�m�n�<�3�L�#� ب�∡�h>���ٌ�bR5`�=�#
��:C��d����C�����+T0�t�qR�w ��`��_(�d��"�� ?�V�ny����W	��в$N�uy��5��r�8P�*�{�#9?����Lb�R"H1ļ`�8�l7g�Lo���.c��f�$ђ��{-T��Q��Ut0uǠ�QƝz�HBp^X�-�e�����P�7�l�h��NiaX�����Q�.�R�ڙ5�у�d��I�_��@l��$s���m��ۚw���y�����b?�I�I߬�D�p��#��J��ɦv��LvW?�L_�]D��ɨ,�(8]�ϛ	�|@H��T������F?/oeװ� ��A�M�|>�*8y�̃�Q���3�ƃ�#3y�܂m�<s)T
�MZu�Fx�A���fä|�%u(�'nI�QJ&N��$������ٜܢ�����/���N(���oi�/�bDI:���J�&�p�ΖnV��)�;G��8g s*0J��(�U^s�r]��r\ӭ��\E������4�Ķ��B\���k��3�G�3��0³a����r�jg�Ə��1�J��B���س8�� �X��B��(�����8Q����Bf$e¾�>iA�?�N�s�m�A+��T�O��bWr�W(x�aG��`$;:���F�)�st((r
��S�?e�a!�� \���ʾ�Rtv��D�qhs�U �UW<������X|4��}la�9@?���Rd��h��/1����q��u�f����טr�/�s��7\+�e] �kxxL>��iAn���P!o���M�G͋��s�2��| ̉�C��uN��d��KIN���\�~2O'3�M���ɒ C�$qNgGBZ��+6*�"و��NO�M���E��g�y�L��0$.��1����R���u�o�\�����>����ʨ}F����t�Iґ>��Y>()2J&v���u�a������c5U�r�2�O�*��	�\�o�'�]=g�gA�7Ζ���`���ۄe�R�r&�n������hU�#�C^� F�c;ؓ(x�///�`�f�^)]ԙ'��G���(���e�������'pL8F�s�!�s8��۷@��A�`����?e�M.��������}��~���/I�"�\��3�/yҫ�Yd�YA��@�8e*������~���b�w����p�SȤ�����h���?U�,K������X+e~=@d+yY
�V��NH���ִt�_|�-;�E�s�kI���xR��Q�� �`ν�g�)�p��U&�͠J���ˇ�[�d�J���	�*	���-����b�W�^��BR��dzϬY��N�#����x�fmQ�g�[����Oz!�S�g��m��Y~�%"� ��iM��PKW ��jj@>� ���B+xaM�AP9`�.��V�h����4������y�PGб�/+��6܄��!c=y�"�2PK�1�B<A�0��kkeI����1�
�];n�vyℜD�W���Yn�� ��`a�[ha�S냙()ٯ����ʊ崩�~���8)ګ�N��dfD��10�Q(z �LB���3>�tC+�l��9zI1�^Y8'61��0g�)�vh�x���Q=��[j��9�`���.��4�m�	3kp���Js�+eU�lY��r��̊y�����.}9���$��~�����p�=3��	����Ȝ�4�w�ɔlA�(g�]Z^�N��fmy��5�������t[;�zV�Q�lb�k�`OTNF1�߅�R���?�3��N�b��A鞱����bo�<�t�7o���׿&���gjk����i��� aq"�f��ͤ�a�隢��f��߳~���$&P�0j���/�hq�Z�x���������m�hȢ��_��1�hI�$Q"��8X��򉿏����>�+�M�6ݹ̴}#Y�<&=�)O�*�d��������Ͷ�q
Q����������a+ih=�ϴ�,���;���*���EW�Ŧ�m��3�H��ϟ?�K�:�&鲏���y����ѲТ֗ ȋ`��0��p�\�Ag��s��c2�5p��ۗ�QQQ'�h��q7=�77��<]$Lf�O¬I�D�<YN�tA:��Z�jP`�mk��XŴ��=��� �GB�9�߲�T����d1�n!~ʓXN��Ӫ��M�@8����i�3(��ļ�]0��$���qC�F��6c&cPX�؏p��S.�$1'j��F8)Gr�P�0�kJϛ&�������F�	��}������s��r�u�Î�����5Q�
�G�?kN�<���s���@(���E]p�'�/�Xy�`h�r���m{���wG2?Q� ��i>a���͖�t��e��0�wp�ٶ�ϧ����c:(�&D�GN2?D
fV��B���"tu�׽|����~/L�S:��t(:xp}�	�s��d1���d�N�V�6�(�+\ũ����`X ���ʭ��]c��<����"��!�QF�&h���2*J�.�A:�y3
9��d�K2�<c'��zyR���~p���p7����>�~~k�t����x)قV5�^a�qv�A��p��N��I�p)?]e���.ڐy.<��I����R����B�3� ��j�QkO�Ɵ]\]p�W���4ܡ���l���atLjS1����eA���G9�oM"C����9��u�frtk����.K9G�e(�>L��������s�j˲�N�<����S��L�<7i�\O�+��qI��~[����c�N��r2Q�ٱ�і�������!�Ҟ�Y����7�HgR�����sj���O�AcK׼�\��L�M��Q����A:��4+�����l��#@E�*�,�3��8�_B;B{G������\��9N�
�L�. ��e�2�حF)��� ���_f����㯖^%Trv�=\|Vm�W��^>��7����_�ׅ8kI��Xz]���=���۷����$��]l�r�Ն��H�dܷQ��ӣQly8�.g�[&P-J��*�:�!3*F>ˏ�"TϮ�<e���Y%g����n�<t��vR���/�y#���~��Fı<�O���wH�={v)�i-�$�^�&��,Y��=,�$����=��~��LOX�̲3l�������>}��U}xx����z�Q6�^�%E?��!��8��3���[IasW��vK�����`���s�$�*t�w{�M�SLŻ���6��PG��x���ao����s�HeI�2�6�t��{��+�(�����v�Z�&J��3�P��结�RR� �t��='C)�e�S���*Ys�������'��s�qN�o��H��o�?��l����ڞ�na�܈)�#G�<�z���t��=�Դ������t�����rOC���|��݇��h5�??=\s���gz �|uq"�ux$t�o�������{�+r)$��v��2�9���?������i�'.�2?�w�ϯ�8���c����g�?��&��Җ�]*�L��YV2Ud����|~�"�v^���3{�͌� d���k�G%��x�qw�y=_6���ӆ��~-�,p��0/*�j�4+0Q2򾞷Rg�y�6wⰉ�(�3���㧶�(bG�N�g��Z���w��	Љ��k��F�Pp�rnI6Gί���ՐM�]M�wP�jx���RB��X�>S]J�["���c����^��gJhX��S:,�c:0��&A�U�0F�-�-Í�9�%F�CB�-��� ff���j���u�8�aIs/ ���6��d��H�g0G���>#�&�K���B,��˼�;ň�f�͊iE����4�@k<O��M�U䯱T�B��Bs��J�Y�S8K�d�hg ��E&�RdUP �"'�� ^1n3��FmNώ_̑0��Ix賵R�[HSL��>*� �P���7 Co�7�gQ��}�`_n|v"BK�yeA��m�t��zm�2��"x��x
��2�d����$�D�?��9x�,�۞w�mɵ�d�	��-��kpE$ΐҕ�[�\9���!k��C.�ܑ��	������p�J��΀c�'��������bu6�t��_��/A����d$�쒿S
�ń^��1ׅ�"��{���g�U2�F�.\S���c��n�E�t�
��G���L �>�N��� ��N���%�|���	�N�#����+u�) Z�[������ l��&2g�L ��C;]�K{�l��jX�р��% s�md��Q�RĬ^����ej H0�C�2G��������`��Y@�B�b�ﲑ���%���+(��S^Q+z��C�YE�EG��&�R��,!�1��v�$�H�b}����T���>"��#��&G.h��9�/t;�e�0#�����'(�
�p���f �Z�Q	ʱtQ1������s��M�6z���L�1���4��R��N�y��Y&v��aهTܨ
K)�Z<d �]ʀ��$9��!U'�ƽt�9���������s�mh'��ʍ��sF��p}�Ϙ"�Y0��D&e[�u���PK���c!ac��ϰ�|j"�(R4��E�����Tw��h�鴼�f��g^_�>|��O�������"ɒ6�Bԝ��-G�*=�)���% ?�xC`7�2�^9g �8 ��ɸB�㗜� ��䶰bq�p��><�?�Vuh����/6����c�1�(��5�˫g+	�����e�gu3k|����$���u�}r��!�m`w���g��R
����;v�<7��$b<�6��b��8b@�þ�]��g�$9�FO���8Y�N��>�L*1j_��<��� �p�y��":L�
ۣiR��jb��c�O���̲A& i9_�s�r�����U���9���D63��c·XE�Ҝ#�������FŦ%��D��{��O�%%E^/��<8�U[�G�R��ʹ�0�m���tJT�t��2�Pb��-"O��u0p�1}$��h8�6��A��Yl =
v|��t�@�/�:[���7x`�k�s��ye��Y�k�f�≧�d]�RD����/�/Xh���x:��@���W_�w��7��nwb�y>��Hc֡Q�epdm��]���x��J�t�b�._ˋ~c�RX�)(՜c;˵� ���E{�0�&��z-R�C��i��#����C�nQ�D���M>����$���F?�~�]�)l���\uJ��|m<��d���hzw�0�7ggs�QaH�ɴ��N=!��-�lx��#��L��.��K���>��>52C�B�#lz�/��Odi�v���(c��)�գ���{FV�������9iϾ�C1��z}q�=�p�A�i[�홼��*�{y55PH�^���/8�(ot�(]�O����x��aK:�;�` �w��xǍ��G�n
Z��b�*����*����L�y߾}KZ:�>�
X�O7��{ʍ�(���F@�SI[К���cRT����>��U8�y��a���B�+,�2�@0�k�T�+�W�LT/OŽ ܥ���Q�}`������P�ʒI��M�
�:���Z
��?f����߀�D�H����!�8!&���o�E����DWK�|������[yg��ZGG!B"�?%���Vf`�A�ظ�Lfy��C����S������>uqqAצo���o�?%�)�t'�@��2��0�����#�Y���u��ze�#��� O_�GV��OS���Y���uW<*���ԫ�$��\�	�U�ʀ&F�z����LD�G�X9�i����|G�bN4�>�9�4N���q2D�x�%��!�G�g�/Eh�c�Z+��:�z������5�g�V$-]���,+d��S��>���%ő-�.ˌ#�\d�G�()���"�G$��2x�IZ7��%��bҎW3�\�u�e,(�E���g�ޜ2(���)d8#���3Q��*�)su$���.Y|��G�WKbڛm�������Ť�����vB-D��8%�r��ݜ;��2�!7
����8�D�o� �_�;�5z-˹��KēTj��u�Z�h���|gi�"�\�A�aa�"�6��v	hB��ۑ�Lh��ii�	eCkzm�2�A�.l�\(C�44�oK�hsz?^[y�m�9���ņ�
����>�{C���O�(5aq ;�������ׯ�D2�|^8�$�/_������	�,V�	�q�[ �I���R�_��z�џ���W��y��?���v�5�w��F�&�4��8_���rcV]��;�q<����^���O^ =��Da�B�MKQ���^�m��xII��|��T��l��F\�Q�
�ū��y�VY�����L��/�D���`�i_@���(���}�.�x[R�@���ft�vY�����I����x���EfIF���)H`��@3 ���ĥ`�,U�(�9А@�.�"�h2��@>���PښIĨq�䯔%\��m`�-;� m��NŅ�x�G� �����z�$��1*S�8nf� ��<�[B�yI`#���B�����j�4�����r��=��k`���:o��@��_\��ҕa�Ĳ�
	��r�I�ֶG$����V\ϵ�X2/~��*d0��[� ��)I+O<䆤�4��n]�6�G�A���$�!ṋ"��_���S��f��X���^��x�W�9�� �s�ݏ</�4�:^�~���1����Q�2�'z��<ԑ�.�CZV��z'�/�s�la�}\��W��I�p݅4F7�={FR��L��S+�w7�)��'	���{6(e���^�g���;Б�&+��]5Kfc�1r��s^h�9�py�s��f/V�f���,y<SYs���l���a)����Gλ�U�t�ْ~�v��<���/�4����"i#�5=�u�]�H"��-�%E�7�ŋ�����=�S��(���~+���aps�]�|C[��&u0�!�%��Y���Q��y(����ŵ/��ЭA&X��H_�-���J���eRP�uɶ���pi*d}y���V�b|b��etE�u:/Xu>��HmV75Ӟ�cC�2����|Q��!XE��+��x����F���A�Mݘ�	��1]��<���i%�\�P{н����뻑,jU�p�zn��$��gC�FmT1km��G/��U��ԃ��E���������F��HJѽ?H�FdO�4;fSX��1w��W� �)��4g�%)��(J�ﺽ�;쾃�x/�4 �Sƃ$�KH��蠆�RX��|� ���A��I.��o�Af�zC��B��0� ����tB(X-�BJ����<��lHuT>���cۂ��0�����Tmfv�S���u�p��馗Zь�49
<�2B��r�2��%�5d�$���O��Hn�+@N�u{!��>u5��i�+���_͉�4Bq�;��:�Y�y\���,�q`'��Eˆ۷�>������j��<Bz��~�'1VUf��Ҭd1I{���q/]������8i+�U}`,�A�}6;�%�ޑa�<�)���4�ry�ٱ�eCƂ�|�]�o������V�ϊy������ϟ������؂Zx|�#=]p6��|zz�摌�s�M��߽�~�)	���0�),bN��<�	NN�gM��{�8޾��t�8��%#Ƶ������淿���*?�NSx���:{��9�?��[頬y�bU�ߙv�'?�	����+��G�譺a�����LjS��w�0�����������~�(iwk�f]f�J��[�M��w�r���������H�[A��0������+����{H�i�v��=�jO�ex+n<����o�3�e_K���������-�h�F�s�x||j�}l���=�'�8�NƐj9��j��T��C)���v�������-kΏ�ǻ��q����;�����~0w�]�ꚽ|�7�;����\�~��l���G���J�V s')̔�I�V� &�a�x83�	[+�����Pp��F���c+N7�PhK�͚峫�/_����x�]�x(�ɶ;~a�٢�Tp�$�*2�w�P�U��Է-�kQ�-�#[�+���#������cA{-�ٺ{��4�Z�{�c���Ԏ�X�ʟ�􋫳�W������%3�~����/���v]��_�.�-IѺlHaqi��9������7�<�?ԥo};R;�H���a�H�8�I�e��ydA�%S^}+��J��:�Ư�����J�ixc"<���t��Y��H�d4� �a���o��Y6E1��@ixR�Nج�V2F�<�NR;�׬�y����A�a���e�Α<9ߔBG�J6��]ٕ� 	��+8˟H�叼6�:m����
n),1N��&%+ <}�BB4=	}R2�B~���~�1'�9�C����0�Ԟ�(�"}5�ڷ�̪�Ղ6��	�@ȽnN@��s(2raL� IY��P#W��M6�ƍuSFmײ̣�h�-d$���;g�\�o[ט�[�@��^;���-xD�5�cy-aj^M�3���cM����pMd�	-'�%�$Y��4�k�#���Eu�&,<�a)���C������r{޼yC�/WIRQ���A���(�[I�pj���bq&<�'��''�<?�XpTU2:�	�����p�������3p8]�P��͍�����������d�jF��hfg��x\��\�TT d�(=�����1�0���;����#z�p���?�~��nڎ���C����q#}�������R�@)_��8̤ߪ�9מS�l	i�HV�ϙ礬��-�J��H>[��xvB�cUWt�+��"����lY����7�޽��|X�_�X9�ٜQ(�BM���s��S�G�@�V8�)K��<O��f��8�[2�uIb?��-����kuU@F���B8v,G���=�]�q�l���5&��&�R�oH��8"����ǔ{2"�ɖbF�����K���f��ZrGvNOPP_HkGⴚ�����Fv���j�Y�7\�g���.u�mI�hvu	b����[=����%�9�j1�r�f ?'�T�W�>.�u��-�<d�KfؤU?{� %��^�����~���~��kV�ȑ����"����<�jBmCÄ��Dě�������h�9a&�j:r<����b����I�v7|�!�]po��l�so���������<��=y�׾�'��wH�$����K���`�H�ۖ$�s7��Ŭ_\q1���e�r�lrdMI:��?n.R8_-�� MD�]7�_J/��U�� �ΊK�����a�&������� Q�撓�x����>���W_,g_�����9gHg#�aϜω4�s:�g��a�D�3E�%O
�t¾��C��J��?n�����"��$�46��Up�K��(%#y!!Cp�DH&���<�̖(9�싐��I�ؘjC=s��6
.4p͡�������^�)v<�"��٬��:��z,^��Q�^ېH4�ۃq���=�����8�:2g���������@��U�'��N�v��v������Zf>xf�����.�WQ������F��3�K�2���D舳J�2���k)yk��!fx��'I�%eMFE'����������*�� Xc1�7bZ������C��L����D����W��]b�)��]yZ%�
�O:J,i��h/Y�LR�y�?�  ���e�q��X���|9���A�d����!2�8������rnu0�U �#��,�6:�*j �y4���P#�Wԅ�s��̕��X�:0+�GkNismq�[ٳg�W#���Z�9��9]�1}d�����F�B���1�ң��'�5��:M���f�@X����Z�K���T{%���Ӎ����ݩF�ym��3kA�z���I!�ӳ ��J2�|�:f��XvS�2TKT憩\u�.푡�B�K;)J�G�[��
!�w��}��F�)��d��1��?r�HkH�4�.�AN�Ҫ�{"���d�yv*�6�;��ڃ��ŗB>���'�ᡑJ�\�P�-^�L��P]1�dS�$�v�p��l ��?q�+�]�cbV�o���[H;f�����>}�6t�GI
v�j9��Ç��C�)T�?5d$/�@��:�
�.�,#v�u.�� �0_H�+����fH �YJ��<Ft4H~;#��~%��U7�U��l��:H�2��qbk�3�;%����\��	JR���|�Pqp�i�p��0���,0]p�XM�U�C|�G�5z�0T6ԫ����!g�`�l&*t@� @�$��<q$���#�����
����CJ`ݼ���B�D��U����A�D	����C�2�=�z��
M$�״ܨ���;~d�_��X��w>��L�(��<h~�]g��J�o���b���h�:[�..//!��o>�}G\}>a�) ���{0�
(J2�^�� ��s�J2�� �_XC�n؃�3�<
��a�=��C������5`_����NǓ6跿��7�|�ß�onn���� R~۾݊�sq�}|�)'N�Յ�'�Ѝ�det ��I<�s>�\L��l�|����g/_��|���X�����m�㵥�Of�R����-����l���܀?殷 �D��x��`�k+l䤬�A�����&1�%�pKri4�<๐R7�n���i�RF'��Fj�mRpG����q�^����L����~����HZ��i�rTH��|���>~>�X}�����Z�+�W���lQ�[�&�vcޅ��H@_�cl��ǘ���#���Ӧf�N��7c}�z����b�k��	�T*�d����	Q���"��b�p�l�w�B�;��&
��ƀ��.p.^�Lx�^�`���uZ���M��V<�Q���+F��<�7��V��F%�	@c�Yc�����+�\��ˇӘ�j2���tH;��py���� �V�k�yx��>�	v!)��~C���B��X���)��3�z�t�q�P����}h����Cf���_~�ybS�xǭQ��9]� t.x��n��*��`#���\e��U]�1B�\����wE�*��p$@����֐�gOdQ��݈����2z�g@i�*�Gr��.c�!!I��ͩ�B,nb�}�`��<����p��k����,�8��G�-(>QN�h�뵄��Ϲ�3rY���NY�4j��ަ7#�Z#���������DZ�Y	�}i,��bjѓVoH���}��JCޑn���1/��7L^�<�G�0���N@<u� �$�I��H��+���2�(n�$��4Jrr��uF��31������)�������1��������
�w�� �8��M�l���iì�\�#H=QEVA�<D!��[I�g��RA�&!x�ڷ�_�;a?�.Xff��@�`�9岰\��r�9TqB�_H�n��@s�G|�x�=&]5��3LP�N����z-;�ܵO���Z��=����0-���~�������믿�;f(�J�_�[`�U�e	���ۉ����҉+/ֈ!K\B�'���b2^���~xn�S��*M��x%@U?�DA�&>A�Vͧ�ɒ\�� �Y0Oe)�.�Y��(<�p��E=�/����Q3ew쥷1�2r+ߧ���f9�N����6`B����q�Da6Tc|���::�N�ܤ8���1̳�tt��AI%,��'�+�������3��.U�3�S��]�8vv�C�'�)�����m�u`���55�Bl�%;ܘ��c����A�s�2��g�ox�L2�i32\��`?�eb� ����4��,��W��謘�R�%pkW�<I�� ���r�f�8:s�+Q�:���H��nJ�1�~��Zџ����y�9�W �q�A�@�C�G(�)s-�R�ح7!<EΒ�@��&�Z&��^���1k��#�>L�Q�I+n׺�Е������af�ES��[Z_��a�I\�6�%��U�_���)@�k�ق�B�	����[ˏ�%X:Ԓ�G�.ZxGV+F��^g��yӍ���޳�f�=�n�g��������޼���0�Y��bK|�Ʊ~@/g[�LY�o�n�;l�{����!��'+kR~����u7����-��!P���W�-�n�ʻC��Grj�P�|���F�賏{�lG�
�u_�NڝBMI�MY/���ise��n]h���Ǟ<���UM�����9r�dj��>�!�)z�G3,h���4AiT͂��C�o�jVֱ�SIW��- ���8V�؉5�tI��1M�;(�rͣ,�ef�m���v�'K�Te����4�� �`�7�=�g�� s���Ok�Vƺ���*���l�@����K�Ȭ�}G��a�XҊ��s�pnWw;���!�t��'���p4H� B���&1i�SO�=�a>�2����톢d-�^!H�2+2��>���Goo�y#X=1�<�X4U%�C7��ʻ�����j��B%�)�<���ºU ��f��yrz私��Cz&7<��9ʌ����"Jhtaæ`�K�g��B8�g��bf!\ж�~���������[��vؾ~���l��������t'�^p��������_={���S{F'g�4�xK�
.������_}��7����I��&L�Hz/���#�H>�i��Db~X�t.��V�8�Cz~q�T��jy���<����W6�*�@ꢔ��1'�ݪtJ� �V�(%w���K��|��D�p?,�'M=��^{bKe�3�'�pk��5����v��c��\|Q�;iRd5?�
��N
��Z��j�R��턂 ��4Ұ|��h�W9�%u��V�:����E<��l���'H
���D ��~I�l�GR9x�N�U�����4U}y~A �L~8�LL�u�$fA�����Ȣ���\���{߀-f=�jh4W�GqA�|�V��ϴP*@{Ծ��l�ddvg�L72���g�	���URW'����/���2��)�Q�n	^���<NP�+j�>-�|����E�N��s������>���~�(�b���L�r�l9L�����/~������:ÕrN�ڡ�]Ϟ*	}���ٕ^[\�iB.�<#�[�ݝ(���<��j�)����F��_��(��ǻ=ס#{��h&#B�&N�Y�k`�Ò<z��(KW�B�Rf�W�+��%7���R���Żw�d ��e�m4��p�L^i�GF�;��N$	��G�G�
��L��{4���P�EB
�WȭE=�$����vT chv(�E�4D����QG:?�¼�s_syd���@�V��_ۨ�E$h��_�)�΋l�P���J	XH:�,��}��}�l�WDӻ�ۧ�㳫k��ȥN�� �T斝�ԛYS�V��~��dg�e���M�'NFǢb����s��>N�������Q�Bz�קn5N�a��f��\��8t��R��6�Y��R��z<�=gG�Ā�4�\��y`o�Is�����������-#����fO&�j������W���E���i���'Lƈ�T�c�z�B�ZH��gE�0��:l��ʻb�v����$�R�x���N�����eSowOM�^^?��Dr���9�J���	,��[��%������n2O�D��?h�L�y�磮,���T�JOh�{Βa/|�����-e�N9%�N��X�"}�+�{�v�#�įJzh�n)��V����\|�J�a�%��JK9�iy ��7������-K������P�̼(� �	E9-П�@�~��sm�M�h���`�IqO�12E��5s���j���(WN�ɧ��T�S��o�u<\Sr�,��Ǡ�.j��>1�w��$>��&F$Z���)�u�	ip��*9��"�#u�090��eT����^�tʢ��u�G;^�D�d�M�d8\J�%W��9{ۨ���.��MER�k�O��/I�b�cB�5���}e�'m�Q�J�bv�HXL꼸�4q"���xss����9+�}�4 	
#-0dF�����?qk0��YY��(e�P�	*j,>/�� +�d`���VtE�0��X= y0�+O�a����0�GF� A~�� &���4w�Rب���{<�cUy\$*&u�,���������Z.S�)�j�g�$�:�ж OD�ό�IVҩ��\��[ʹ�i��ER���+��c�����V�х=
��!Ԏ'*T\�Dq}�dhF/�O0?���^	zd%ч�q	�#�]s�����PG$���C����S`ye�� j�sh�~xx�ʂ#HW #�!��:y2רxg,���*���eo�dYr��E�Y�KUVem]U��F7 0�� ц3��L�|ӯ��!�h���M�0���F��^k˪��z����'��m�̛�'_?�ܹLt`��!��������6!�
�P�(߂�H�S,6}V�mW�^X��O���/*�F'/q�2��lԩ5�+�P�c+�cAr�5耎cH�^��K�]�W�mc2���	G�ZX{�f���F$�9��q!]��cb$t(�3�x�(G�^K�ĶL�!V	���G�U'θH|�)L��6��D��"��a�#�>��~�H<���S�4��t��Ƃ�I�-u8�XtS�t�O.��6:�'�خ�~��w�>}J���oT\�|d kS(	�9I�`��UVǫ�YaT�N
rf4iBssH_��^ݽ{���駟�w4���?����`ǧ;��8:�O.G$����m�瑥Đ�H+�������i�ɲ��Ė=>>�g��eY�h_I'Wm�2`\�ycP#u���4E��:ش�镒���|�HE@�|��g��7�\L�9�B�4u_�u��a�!)�����̠wEs3�D�Q�춘�4LK*������o&�+Qx����D.,%����� ����J	[#dIt4f�GΐX�����uQ	�A�3�Ө�wAJ16��B�k�z�y��;w��ۄ`�
���@O�AbPs�cr��B�k�j��I�wk-�+��6�Q{��P�g�n��DC�I�̚���s�3o!<S��0С����f����:)�8�F�a�V�}�R`R=�`�H��F���j�i��	�HeT�C�d�Y�Wy��1@"2��i���EG1�#9�9~&�hO�
k
����:I#��������uQ�xt�<x����m�����/�\q�v�}�I��6�O΄<µ�f��}[��#=�z��~��]ơ�چBx�Y���� !B[ �^n�,�=�
�-IP|�pt�*�r�	�v�V]>�#�����F�W����kX���G�s�W���8f�H��W���|���?X|�l�zܧ"Nd�:(���!ۇ"P䊦v=H���.��(��"Ɓ��PD��S��S#��B�yd��r�3 ynf*f�ѨT�P��ز�T�sp��|�Mw�w�.�-�"�?�#�2��E1S���&��Qf=��l@9�"䙗q�����Ң��Ȭn.&�9^��� [hC����p�߲Rj�V�����M���z��'�m;�5<�4䰼��!���~@L֩����)������~Ӿ�*�&ޣ�_�H����id��Blʺ�Q����~�[7$���~6Ql�f��E���J� ���`����pC��=y"��Q�8����&�Ҭ�����xs�'a�w�Md}5�|��!�]2xʍ��w�B�\0�g�۾[/j������� CT���Tm��l�P(���Nts4!���G4��B6dZh;��9I����v,�k*~,�d!;lR��D!�9�XK��� ��ܴ�6#��\֠}�,�յ�g�(Hc�������ٟ�5Ϋ'��+�^S���.c�����VZ��
L�.+7C��ݠD��&�'Ұce�WP�?C��*�mFp�����C6�:s|�'�8���5�`�V��30�=���Nv��n�8Y������v�
�xVH�pղd�}C��T��P�,y-���Ѯ�����������Y2�1;'"����Pf�/���OOO��Dt�������4�� �s������4RX����8s63vZ���h"6�k�����0��^�X�S�7G���Z�L�GXbҾ�MlA1�(`���f`v�2^�1i]��i�|��/F@T�nb�S�-Q����C�2|��]��|����sqM{�����s��If'���"��	��[��K�]�� Pܰ��vGJ.�)tѓ����z��b5J%�|A&N3�~t������P����qw6�Y{&S�p`���N氓.�La���;�3�=f��t/�;2�%C�s��;J�Cm�?nH�Ͷigf8�������0�����)����%���%IH&�bA��k	�0hT�׹�2��Y3�N�=�͕o|�{�]4�j�EY������>{��<�Z[�)��q.���>��V�>7���P���L9Y�z�V�=�u���zCo{����l>�h@�e�8 ���^��|���H�],�ֆ�~�`{��2�ϵx_A:0{�b��.�1۸QZ�d�px.��iK���`��QK˛ >9m�Y,��#7dK�|��$�͌�w-U��*g/h3	7��xց	p�\R'd�EbN�j�^���|v�r�7�:��>��K�{.�Cm�1�e{���7��c�5�_�1-�Q����+Iod����iC��M�7�X��ۚ�b��$�����|3��n�	��Av�������*dM�Ӷ�}�
��ܪG�(S���[�B![<�Q!��ì�!w9D\ڲW����{���o~�?��Ǒ�ݾ;�/���K:?o�Oo?!'���ͮ|��||蛹D��d����P=-�d�z��O߽������Do�^;�Ӭ�sݾ��.����`���'�}���W��Y�j����_3��V"�6ܤR��GC�"p�2���?ܽ{��<���*�zK�TnbV�Z#�x��Ӌ;b�eP�
�4���Z��:ا��Vl�@>����/�t�x��Y.��]�2"L�YV
����Gh�܅|�A���a�T�P� �`}�`�A�c����Z�曇�0���3ĖMf����^�|���}�g18�9�3��\�����
̀t�3OL�+Z��,�3N#�N�
�6��Z/\�ILH�M~����Uk�&�Е��D�'A��a�XP�|H|5����?Jb�ik�N�s����^�\� �_�u*B�����9w��`��v��g�F8��Z��>�v!]��&{��Jm�ƅY�2�V��*��RYy��g�߬]p�-�.ʏ��#�Ux4J�g>���͑�}�_-f���#!G_w��.gb�B�~������w�5��O>��	��3G��~�۬ֈ��E �s�ҙ*��U�%��K���d���%��؀�͙�����{$�oﺭ�C;:9^&��&-����R
Ei�<Z����t=Ea� ��^+G�[�-�fw�*��:�����9��J�B�ꅙ��ێ������i.�rV��U�Q3kd�;vR�31����mP�6=}��e���(7�����vf������d��0��1'�P�I��vm	]ģ���@�MD�p�DKog�!iL
��=+�5��vCp�p����~�C� ���8]T�%i��n���P,���^+��*1�yyv�C#@�vL���q�����"'o��hĳ�Ͼ}iB�I+��yB;�@U��7_
�m����@Ps����=�p������G�2�|���Ҙ3���]b�Hp�;8X�-4�������M=���|���6�H��BO��7�G�$y���QH�3W�A3�^a��Z��>���c7�l1�g�[����n��=��!�
�Jzu�j�fFH�_A��|'��2���FDxme�Q���BN� �3��	X�@������\�@I^�$��o���ɱ�>L-OZi�؋�a���L+��hW�ǥW �{���x�V6���̤Zo'�)"�$)f�Fh��Ģ���IE�ز@f��1�_�sT�T��7�z����sK�0Nf�׊W�&,�-�M�ɤ�՝6ʄ����|S��-3��:�%��`lӗka�ب����(m��qp�km~��VZX�G��s��y�,���4�R.��#��o%/����v{[82v�~��r�NNN��ãe��1w��&R!�9%��5���j�+CM:�h}Qa�s��u0��3����:��r1k}��,�tldYb�E���q��c��O?��Xs��Aȳu�;r��ޱ�IⓅ��S�9A��Hj��A	���`Jp��\����3n��;�:`�!ζ88Ե��mW�ѳü,��~�<T�li��&���xӐ��3P�8�9�a(� �'��'��G`+��*SW!k-S�t�;mS!�E�wܞ��V�@Bb[;���9m�5(z��/���b�����,�@s�2��\ʫ�E�&WbYm�a�,U
N�Sst���j�V��5������L�}���#�5���k�;��^��I$k"�D�3�,rʥ��Bf??~��޽{t=/f	��|�j�^��,�0j���	0�p*��Ǘ�N�:%����F��µ�{p��{8����Q��d�1� /�-1��tȅ7�BWB~&��Y����)P1��=i�'�G%���>�>pr�Sd>�	�b��8�W���� v�� 	VjI{Ơ5A��:��ke>ŉ��A?��q������.�mEz�Ν	D+]��7�ԏ�N�U��sZ��GT$�yh��h�BD��WW\�=[2�ݻ��##�;Bϟ?���/^D�Nifz�]�Z�`����{�Ǟ��=n6#���С�yl�fB�A��k���)���L���4H�®jܱ#���m�n�C-�I�&�|����y�����ϐ���u�۵0�A�4��c�z��������a U �:m���!��;��<I�0q��z[����4TT��L�Y� �?X;�R���iQ�Ӷ�["%�>Fm�N<==�u��$�W��$"��A�u#B՛�{��x����;�(��1�t�o'��k��Ak���f���f�j�]��'w��A=�|<�(�͉	�`�+\�T���
5}d��`L�<�v���9�w��v���0��� �F����֖)���z[�4�ޤ52��9�I���yu
WOZ��y/�든�S��4-L2f��H�s@����Tx�f_��m�냻�n�NAR����IN��;
��3C�@��)�+...��&��ѣG��1���&��{�|�������0@�6\{x��#p��zNw���m#gǣ�6�}F9p� ���S�9�k���,09"��*٠4l3�C߁.�R�����&+ I#������+	�e�l2y���H�� �+�nn�� ��W�Û��}ǝ���W���b`Q�>�
���7�f�(/i2�LP����v�>�y*G�F^�m �R�GƎ�G�>O&�-\��*��Q`(>(}u�<LZ 
WByu~A�;*n��L�Y�l2:�R,��h���:7��-����b�,�����GZ�x���tn+f"�Z����Tp���T�yG�^�������{��yA��M#[R�Q
�}�;;�Λ*qu9����fN�Q�t�Fn��Jg� ��X����i��~+$���/c�Ub2��� p
��6(o���l;������x�6*5a�N�S#��@{�������
����k��V�|)��nn�����8jI�X���ǔ��i'�<W(��}�����k#���Wk02Ş��E�6��[Q#�Ӓ1��6�:D�ǐs.Y#aF�-�:Ћ0��|���Q{�UZ;l��n�tn}嫤�4&���A�lN�^K�̯�ڐ�/[x��J��'d���Z��i�ث�h6�8iGERΊ�0c��Kn,��4��JĢA���t�m�Ny�K[���j��SK-��¬Y|�y��"0K���4J>5�4�
,4��捔�h��m`�-t�\|��t�O����Z���wz�dfy��w��ɿ�E�ȩ���G���n�90eo<Xd��h=m�=Y��m�ٚ\߼�  ��IDAT�'_}-�Ƞƥ3^�A�qP�a,B���+�7N�����L.7��ɪ���~��R��p`�BfI3-Xz�U��]�ܤS+�p�г����M\��`���ڊ��Vd;��MyB�����P`��]��4�Ik���>�+�n y(�k-�R��m�5w��X��j��Hі<���_96qpx�����&�H��cG��6����/�4��a��k�r2�(�P.I��z���G��BhꖓcCL�æw��U����z��]\m�{��l;�5|���˗o���ɝCތ#�&�$UG�f�vp�֕��CJW0��-5䳉�
��A�.��*F���^ai��3An�ԣVe�&2��eT?�r�r&���d�|s��Ez��;$�lq��/*�]p}��n49C�D8�v��v߾�p0v���l��vþ�¯�C��u��ԍ��TI���j�õ���+�P�6y�zVJu�������Q���^K�&�Oh�tqv��jl���U��=%C<g��_�����	��v��95�T.lv�f��"M�#3HX���ܧ�m���qP�׮���~؃,�j�b|���K�^�����I%�$�\�!��Va?H�A�W'i���q�l�B�F�z��6�Q@~�~���J���CZn�G_AODK���c�4<���/~A\�gZ3������!b�F�!;��m��Y��=Yb'ԝ��1�>q��=8X�
b���K��I��///� !�an�&�h'/_ԊBZ����K+!$'�C���Y���"g3i誚�	q��KO������7_�k���n./���j}�8\̖g����y�Fܡ��av��5���1��,Q�ywM;�\��j-(����:��w���NONqn6D�w��h��w����M�9'�\%+�����r���H�A)��Ƣ|�h?�N�>ۢ�]�B{��,�t��U0f��84��.���l.�' J���auFVSZqN�Ҕ�G3�������� ��H�+E���0��&�L�\~���о@�����>iS��9x�Z��9a�Z��C�eN:�u�N ��hD�
�	���0$��������ޜ�n���Y�f��
d]o�-���P>_4�KZ�����E�������裦^�NZ�S��")N��fQ #�d��'�/rfO�J��?�[����D#�c���B�������U��efm3������(�crdH�j�|����J���5b��_R$�j�4�B���v�����x��W��H?��$�| y�A���#w�"��<��2�;,�;z��Y%��㰽�:��!������������{(��ɣ�����Կ8{�碝/آ���l�Y�3tI�x�KP�o���T���_̍E�	��#H�bQ$��,�L�o����b��Ę�7�wHZX>�c�vs���Bq�J�G��Ih���Si�6/5@�pF%K�G2uK��I�G�th.�`�D/�?&��XR����l+7��0i1qa<hu]7�I�*�o�i�.Y`��Zf��ר=IJ�?*o�� �v~O��6�� PeY;���m֎�}��AX���J���t۽�&�p��Wd�s1����u+�Mq(�Sa�	`��K�6��0�^i�[%p7��$��%i�v���I�%�\vB�����0�T"�>f:��':�1b�\��]x`Y,|�n���ّ�k*"%왚�}�����+:J��r��R��F�z�e�<w�����#]H�־9�[�$�v�հ'}�����!G��MX����BVM���"���d ��A�E�	>�P�ݲv5�YLK2����1A��ު�ޥ���(�jQ��86q�wN��kd�����/-�Id��1��? ���wN����k������wVs|��3��/�h?_�湼��V��mm]`�K��/`�O�Z����0$&+�:���ð�Þ��|�Ҷ��,
���H$��é6�,*P(hR��̡�WL|�qV��Vb�r��6��aj�����O�w��r�0f�Xc�l�X3�qք�J]�u�L0��'2	���)��eB���)x�#���%�yȠ(2���]͑P7�L�	��ǃ`�$�
��X����T��g�-}	h>�����E\?�b�j��~1 �,�Aڗ��u��OH�ћG�%�|qy���k�L^���e �4d��\ �T�ҿ#9Dt��גx�@�s�9j��L�Z(�1S��n@�do0�ݨ���V�*��w2��c{cz|x�H���[fKG`ҋ/�����+�d���-�V�N{��Џ� ��	���Z)d�.���Wμ�J �fN�Ks���&�ւ���g|;<[�+i:���«��I_���&�J��$�n,�W+���GR�3���1�;��iz�����-k�[������5
�?;-q��
��n�����AbU��}����/�������V�.Ε��72�3��r��3:B�p����O�M�*-�����r3���oYx�����rSb�T�+g�+H|&����vK��K�sm�R��L\��N��s�;�]���t� �q��������N�Ms�4�߀D4��������;(軆ۡܲ�)Y�kdY������q�d��۷oӕt�iؘp�6v��N��9�"�.$�+H��HڪT�&���a<��$�9��[k�/p����:��1ot8P������R���Ɠ6U�ݥ��j�:�8}A"GN]�Pq-ɨ�IK 	v,��ʣȒ�p�0�vx��6�ë�������Aٻ�����KH]xb$4�
(�����;w����{���.xq��.��?�����qֶ�j��շgRl؋���8U���y����G�D�0��3>ŏ=�+i�I�-�d�{F���i��y����3�}��\|�h��{;�~��{����m�q*T�}�sg�^�bJ��t��VE�/��vZ�IΐE��d{Z_�q�
��&�,*,ńRi��b�+jJ,h��k/�^!��ʨ��4��L�').��4e��oT�kdҞ|� � �hHy�>h��I��Ȅ�
�Cs]BFg�J����C��&Т�<ɵ��V��շ��^.i�c�<��!Fo6����
� IT@��M��Ad`?-����
6�����X�T{%��9lET���UZ�b�2c&�Yb6KP��-v�}�����
��k�"� $Pm��e�g_ĦA�W����7�ذ3Ƿ��,�A�M0x\o���fǳ�ѵ�dջ��7!c���=*/�G'�����]�� o|�;�uGI3��l�������d+�<ͼ!�'?�	]���;dݹs���Ǜ=/+$�,g����aH^�DϞ=��<�w���BDo���}��ˁ�	J	�?&����xý��A������sG^ }���H]	3�2�AZBsY�쐬͋�h���bs M19��-<�>~��c�/
�+��DB�]�M��E�G޶$J6���L%����'���#8m_���O"\3+�U�����`_�'�Y���!h�g�����Օ�8_�����o��Czs�I��]__���k��v�E(��:��3�6\���͜�JÐ��5;�ND/�!���t4��U�wS;&�\Ei�xB��^d�,&X�	��|���U���45��ׁ�4��Z��$���>{����~��7o��½��nru��J0m�à��ح�@V[˱�B�o[�d�}� ~�����.-�u�����B�X���ǧ��]O�M:)��J��)�V>{,J'��69+ea(Kzߒ����0�b��i�\�Gy��٨�'��l?Ǣ1Z'X�F���|�d�X���{��g#6�	}���q"$�����(��n�˴�,�S��"尝�C 3A̵2n��X����f,�@"�V�=��9{01�PM����|7Z��Dn��v�k+F
��$2c� %�.h���ѫ�+�&d���a>������U��F*g��O9�+U�b�F_�����k"�e߶�ų��G�cޠ�'�6�vR�G�n �;�,en�Ϟ2��쪉��-C.��� ϼ�K��et��˙Ä����*[8w�ƹ-��m%���y�oRo:-7�*ϛւ����9��i�d%��ȫ�%��P��U���a�
��˅��xq����2��ɹ�^�.�}��z8����u�
h�ƕVI�Z7-�%A������س{e�Z�])�DT^KD ��ȉ����+~��&���˗/�?^eH�HBr����ϳ�f	s���z�Ĳ1�D��6V+�4ah'�)�%K���C06\�3���WF�A)�-�'�m�;��I��e��:�r�������Z���{�i�/J� %��E��Ο�����.��Lt(-����uEѵ�����xJL��@�$��?���`��]�;��F��F����i���!mw����nxqzz*%$B���б�_Idu `��"�2r>r�� 0IH
L�m�H8Яu�J�
��g�p������΃,�i��W�^��'����0�(�ꦦ�`�b�:��qf~���7�؛öڬo��{���7k�,h�3:��	��l1�ȴ)�S��]���Tj�"9#��Ҵp�e	���;���03ƅ�����]��}xkt��(*�V��m���c�F�GP�����/ts��[�سQ�ɸ�{��4l�f��
P����D.>n }V7���M�
:�_~�[��N�	�Ү!}.�����4�nu����~��Ctq:��\��	#������1��A�4��#�C��m�8�w;'�x)C��=ƼZ	dƻ���.g�i�an�{Dy����6�::�����PW*��l���ӆ��d�Y�gk􂯃����s��P�w��2+$�}��3� T��i�C�=�sG���O��P���,���i�ɧ}��Ქo~������1�O�w�:i�D"��̓{���n��:<>Z^����o��s��%	��|��{~`<fp}҃����O���xy~~�p�7,�>|�����[��ɀ�����˟����_���9:8x����z?o:"��\q�pLEM���y}�V�7/�߻w���Ũ=m�( ����ɼWcW<�c�f�օ������j3�Ŏ-�z��B`g��C���ip{��S)](j6��
�H����I*z�8���A�s%��5C�)�/����F()�O����&��|��V
�:��b�Eg�)��N��i!��-�Ҝ�I;:�n���+��6���w=�Y�˦�\�����M���M�b�d��>H��=|2h���<]�O�W�b�ð>�
��171#�2wW�W�
���MXX����%MI��������^{z��b�j�M7	�bj��r��!�b�����Z���nQ����bި�,=n�CW�1�@�A�Jt^SO��T��F�#*���&m�ZP������~W>��NiR�⨪���}�Tb���BSE�1Ym`��b�<����&�#�8��S*$��9�iK�6�8D���d9���7��d*�9qt诗�tk��0�L�jKʙ��%}4rY��%���KN4q�7v�8,�-�q����^}Ł���׷�n�P���>��pv�g*�uEri�<r���$�Z-nw$�[V񻵠(G)U�Κ��{���F@��v��'Ʃև� � � R�f��t�ؓm$/tQ$l�XS2˚#[9(q����z^�s~+i��L�C�B��� ��Z�ڵ�t�M�Z��Ͱ���-7�-*�(� �f�n��{�ؖ��ZY�5��I����2���4Ǿ��0���_T	AR��]dZ���!�G���iYU<rR�1���#h�4o3Udd!I���kь�46�CǠ��Mpq�q-a*L^���H�+ ��o>��!"���!2�zty9��A�����W#��?w�%u��ɩ$�7��~7����W��N���՘`SP�Y@ۚ�r/N6W�k����l�]v$�پ��'�..Nn�M{~����i�M��ۡc<�Gռy��������铣��ͧ��7���ӻO?i����K�1og�Sa;��}Q��c^�9S<$�%�%�݂uS�`�$f�݆Iz6�T��Lh�X;��tr�׌~�%���Q=� &7^Q�g|�А!O�����#g�Y��,�SZ;�	ۀ�����~��� �Q���K	cjK���?���^���J^rb��SkT/�z�'����,Eo��R�r)��r���QIL�\Z�l�dm�)o�3CQ�k����@��c$��X�kmd�}?����3������0�^�|ˀ����*z3�I.[��8G@�LW	����e�d�,��0MF�Dp�I��J5h~l��(�X�sF��:�T�1C��L��V��k�a{�
����
2�����&'I)8%�"����+@�E�n#R�ŋ����}�k� '�3��z��
S�A�A�J�L�Z�vl��-�%ʚ5�EO�f��
��y�x�t�e�rN	i7�&�{�Ĝ\��믿�ML������l�)�2�ZW$Fԇ�
`4�XN�>�h� �2�aɠ��C��t[^Ƞ�qcY>�IQX�ϰ���X<�T�7�`��օ�n�"蔡�CnU�3��y�$�a�#�ɘ)'�%:�a�̊�C&���L�).����d� n��T��^K��G�&�Ke<tC7��f�MʓC۾Q��ʴ�S�󉳉���RW�2���^��i>X�Q	�\�����&�Y�� *5��
\we#��v��`��v�t��o�H8*`Gg�A.�nm'μ5vp���lӖs��`� ��4p?(�У�6�L�
���hϜ�����'.�;��<�����7��@P��
6t�l'"(O��x�ÇC�?�C_0Xњc�Y��]�`*�g���C�6�6�vǜ8�_ݹs9��Kfb�wA���;-��)�^����p�ZT[�5e}�q\)R�e�N[���T���o���w&���D���h�r�KR�uq��C7�bL[5�gl6-}�B���c�7
[�v�s�>�������0{�w�y����l�%�sFF}�}�d��xA`�i�%E��rh�S����S���w���7�~!7c�ɽ���\�=�>y���G�����������O?��O^�_���h���ې�, �{�z���Rl�ҭ���y��_��Q&��u��l�P��RAJ��2J�W�-�i����M1�n(Zly�P��1��h[:H�7��ŭ�i-�	i�i#Nh:{��dE>K���],�\�<�*�E|�49!���਺-�����J4��Rbۊ8E.`���1��\9´pj���|jX3x��ax�����&��6x���Ύ�}'�d�@Ksb��@�1I�z%�O=+�/�J���,L\Z��L&�G������/ª��B�!�<`V1@�9�1�",
�~��ܴ�Si�ܰ�Fw�P �#�d+��E�ˍ�b�S�N1�.��k'7��6�d|�-5/ߋ0��z4^P�&!�QJZ��!@���7���`�éa���ё��,�lK:���ً9$�5)�IPD�*͎�R��wu�]�wk�E�q�Qp&e4�,��B�{xx u�i����Z��?�9�t+2ؐcX�˥\��p��(�����#[���F);�j��K�M�<��h���a��� h���a��S虏�
�N\] |��d���}&�m���j#���2(��ϴ �ԠL�3�qL a��-�8*��ww5>D��t���t�"�JZU)���'Α�h,�l0'q���A�&=�{xv�]nD�u���1�����@�m�Z�ӶQx" ���1���+)���9�&A^�w�v@d�<�Ng��F������M�[��aA{���������>h	�jES�X�������~�>����rؓ�		���!�����D�M,�2�^���9�o$;�	�g����=m�/�Ҥ�)�d��fP�B�+�7jUeoq&��vEj�$-P	*�B�v�Ө�N�J-����҆�X���b�ij!�X�ݙ����T�\nВ���x��E�.*�4��,�F ��n��C�����8��Q�0NFs���}��y~�,�:j}�[�-B��l!T2����K�|1��32�/c�x�u�$y\p����D�G%���zQ����pt9�.,!�)%Ke�b~� !0�ЍEJ9*�+��*vG�@�7M&�/�݌��NZ�4��d�1:EDÄ
.m��Y٠p3�*�T��3"Mc�؊��ke6)����Aoi�-?r�)�y$}N��q�F��6���W��՗_~����&���<C��r������C-����!��m�=�{�!���w�M�&I�X~�h@�x)��:���W�5�q0�Z����M���F�쥴X4!�
���5������x"�� �s����W)����ӂJ���~�6�Rv$�4&��!34�"�>�2U�3�����ƌ6�(G�J���<��,�Jʞ�3�}�k��u�[�G-���IG�Pp���j�D��̌�aW�r� ��u��C���Ӄ"m��ܠB_S>f�%uh�I��(Փ|�E�J���a�XG�����4�N:&[�� �EU�t�fD�jb�tj�X��0H��>��Ë/�_;��A��`��.Iڙ�v[)�`�
�&ۋl��ln"�L���bZb�b��ff��e1VC�����#| |��IC��Cn�pHs���#Z�O?��������|�;dĐ��/��/d��C�ѥlo��\<�[�_�����0-�4�ƻ�K�Z���I<H�W�]��M;}NУ�8!�Q�؀ʓ7V�x�-��mqf���^�v��w��}w�c4�cE�"y����շ߶�^���r�����(�xv}�vO`
C\����'E-;vf*�ю�^���r�8�k������'�q� /�<�-�({�Wʧn�kҾ�LS�E�!cvd1{�ѭ�f��Q1�r�ye^��L���(5�MA���N��w���o~�)��y�.���z��������{'�|'����s��zytz�a�m3[�{"�w7�䌒������������I����������囗c���.�zz��+qVE���ɓ'��c�T.���S��G�}����ISH�Q��_|������i�������)����ǌN:>"+�˯�����[������4i�,�6���E$NL�Q_�ߪjr�F�	�/�#Ƃ0i��C�\��������+�s�����/��=¨j�#O`�Πe^ِ���i�?��j�	��LM�`}k�Y����\��cy�Ĭ$���4[���jCz�{ÞJ%�>��Q�J�ꤸ$a��ӕt=ɴm��Z���
X�,Z�99}���溡o��Л||����̞Y���%h��ܪ!SG���f�PP\� |�u�f s�iq(\`oF�A��]��B<UQ����!j]���"4�(I(��m'�F�IQ�
`�a�Z�	!�Q[�	25}�Ҝ��{5fX%�*�Yn�f�b�o&O.�!I�
���M�!�m#{0��cQ���%ۜ$��#i3���Z톁ri��A�a����d�X�R���\�ns��z#=�"�ڑ������n���j�7���A#��juAO�������	����}���ׯP��f� ��[�#�=�-�$;ḡ�4�N<�3�~���H�?~̝��Y@�]�疵3�q��2�WI�.��/�]�8~�c�����N���j���;�t�
�v�F�V:�+����M^v+#�0�u���9��������]"	���G)'����瀤�"�)=++�� �H��/_b��:! FY{7!�|�D�;�h���������2EP�/E��������A��&���	!3�&i�y���S�=y�C2H �.�KP���v��d���6����
���4�d�V��#�B��!Q�4��g\���0t�߈ߡt���O��0��P6�k���� ĭ�lQIL�,�b��w
B6B��6���~��֫5���d����M  L}�>w�-��ܹM�a9d5ݿ}����&��`v�&~�ů���7�=��|<k�������.sAqU��x��,{]��f���`J�9��q*�os�:�Ԑ/�Kط��Ύ#\��T�����]G˦���ܣ��=C�9��8���L#�s�Cp���y;Z#�g�;[����s�>�Ϛ�KPkAA=�`�M%$Tp�~�q&R��Y t��?(B�e�S�mֹ��i&�&�]����|.�&��XЊ�*�}nrʸ:���F�?C�����B�Y�`�G��5��ej�;H�t�s9�4E����n��HB-4J!0�Ò�ז���*l޲4W�*2޲ǧũ�������bb��%�JL?�3�թ��Ý���;���b�� q�G�4�
Q�]]����2�<"��2IM�,��N��݄0��^0Y�	GrG��}��.��WqP�#T!�����0
���G�ܠl� �V��G�;<\ =@s�h�씱�v�}�5������?'��!�
}��� �E��?ă����|� ��EZ4���r�@�kHw�����Θ(��I ��g Z�^�<;g���F��vj�e�RG!�#Ruj(�b��D,��3e��(p�ک�.��lq9MY�k�>�WQ�)���d��
Z�'H�����) K*���.S��>�	^��t��m&�ǖK&�������Dt�*t��ڇ�B{�v��i���ƥQ�먴��˟&�?3�K�!���E�C*Dr���(փ�E�1hÇ�鵽r;�c\ũ�� C�5ʩ�L���̥�OO�>|���>@�e�P�.p�9(6+�������Ǫ}�\j�.{�����,�M����O4f�%�m�JH����s~~A���M���H)=�i>*X�Ֆ2�L��P�1u�u��㵤=|��@�I鵈�Z���d]��k��q@0i�����j(*X;��h'� ��!�J1x�ɒ�)����B�W�^a'C�?z�=�B]�E7*���p ����A=���+p%=��޽{O�<��m�.�q��>��.r;�߿��bA2;.����H�%�$�58�ҷ�\��Y�*3�g�֟���O�>}���Lu+� �6ʎb�O;�+��X�!�����O��O��]������I8�ߢ�z���������O>�{��\~�^�Ts.�E�D)>\�k�þ<�^�-��}��˗gY7qu� ,m{Ǭ,�%�q3�\��])-oiu�Zql6��z1W���V�孰� �G%�0�ߌ��P�ʡ<�$��E�Z	$lil����Л�ғ�Ʃ2�wB���l�DI��:��B�>b[�wP�9�`DN�k�	<�VZMn{-g�g��Y�Z��y���+Ai[��>�6��sgF����)���a3�m����yxh�ؼ���tu'��U���DD� ��<�E�U�L�
�����ut�@�H0˜l�_�yŒ��?�}$�[�K��U�6{v�Xr���5\U �w����O9�����g|/ip�45Q���n4>�J�"2�c")7O�t�nK�xvq���ˁ��~vt�0ꃥ�!�@�s�A�Q�\ݽ{B���_�<ĕ�51ݖf��x�&���DԫL�>Ґ)�f�_�>?���}�"A��� ������l7y�at�DM�0u���d0d�A1�0P1��,�� �7hDvZT�&@񃒋�6��!�L�e�wu�4;�2a�VY�yun��%�P3�<݁=����#���8���#��w��SIw���3��X�d:e��D%/�74A�Qev7K=h�k�0@KC��^ؐ�+�<.fsx�Q''���|�����~}�+FlI.����k�LtبFw���5�(�����%��ٌ�tf�r���=g�pY���ˢ�I�4E�^�͒k^������a2Jhx��<[/8z��K2����!�����,Ϟ=��![�f�?�A���ӻ��.���=�T\��M�7o�Ҵ����������w��.�J��¡4M�f�>d6��$�eQi�RQlV��2G6����&)����K$�^	ʋ��������V���*��讷�?�,�#�w�j�9�%�+^��;F���,ә�+CDY2��L/���O4��j���L0�e�/��eޗ���qW�1rN�7��iڎ!sg��l��ԧ�#�%Gʹ�1�\A�_!��ƦJ�L�\3X�j�r�1Kg�����M���X1�eoeQc�W�ȑ��Dr��)s��p�����֙M`�d8W�*��.-Q��T�:����r;3�S�v��qϰ��`���WD�9dWt?�=���'6��q��y�</=iz��]�7ڿ���G��ْr�<��U�"�'CX������{8����O
D�R4��h�� �Xժ]���u��9#iIl0�&��Z�C������?�%pv�Zb�<�(F8�����E�$)��2���"�t��S�'e`�_( ����������[Ⱥvњ� ��zA����}	�+*����E��g�U��.5ܾ�)�E��
�
��g^��kZ����!���ձ?���:-d��^gb�Ȝ��N���^s�B�2
"Yu�{�xŕ<a�`؟�'"`5���gc�I*����pJ�I����� w�d�/K��ͤ�ġ/�uj��O�_f\eqJ���w�����͊)�"-QK󍎥��zY5d��DFUB���Ͷg`B�Y��ȅ�T��D�x����@�$�*
�Ӟ|��\��D����XI ��O�d����W�)" �ኰ���|�
�v�(�a�ca�H�;�+��V;Qp�#4�����gt��R���Ɖc�4A�j��h��~�<t�2�&wݙq�����{�NN�AZm�C��L�9�f�似��ۘz�-�q�8�#ͥp�.�ʂ�O����ndY�Q�q`Z^��BM��㮓3���7�s�!�/�d>�i�Ѵ2ɦ�����v }��NR������{Ӣd�E����f�� ��m7KZ��P!;���{��Hix}vn^\��^���Qgy��}��������
ˇj�+��8��.h�Cv�Vz����_}F���I���6��}X,]�_|�՛����`|N�&�=�a�{ƚ�gm���?s �!0iz���>yz/�vOS��"_�=(�4�g�۷o/���\`������	��A��w�=yp�̝����������ç>��#]|yu��矏�I*���@6[J�J.�r�	9/R���Q�dHsB����JZ�#k�W"#9^\)�<��1�l�E�`fߏE^�B3N��X�Qk8����-)a�S��,r�R���EHT��IH3aS!��s2���Q�bI�`15�^���f�Z�CP�lK�J�Xʀ�l6��>�����1dȏإ����6�r�K.��=>��f$Ð3@�%jer��p�!l��4H��a3�����CIE��X�'�5V	��$!��0K�"�υ���,;�-�~%�B� h���8t̘�����}|����d8F.��wbL�&�4�zp�a��bӴ	#��nd���f6�7-�~ r$	�}��n�H�S�NP�$q���=N�6�|ͷ�r��,�޽�v\mwD�/j��,s�|��s�w+��d,H��-��6����w����t���_�H�<��w�Jnrݶ��+�~1�rˉ^i[V���xq����GϞ=b�ayyE��n�����"̮� a#��իW�1��3޾s����/�� :��ri�Z����8�mk+CG�A������,a�[�	�ᤨ����$�^oۖ�P��R�))[U\�t���/��a]˦ȫ�gU�>�������m�j�"�Cv�Ivo@�i�<䎡$�v�P�b�a�4B�..@J������"��q#����YK����#�sW6@�	!1�{��w�{IP��|��DA2A"��qaM���g��ѡ8�'�����O�[����U�j �X��Y}lH
!�E�&�w<��Ƕ������J@<���*&d�5A-�22̠��s@���rm�be%\̑t��������;�BG��S����>�#)Ӄ��G���o?'���'���h)<�K>_'Ǉ���I>�EZU��� W98�߹��.w�?�M�?|x��q�og�v~��*o0�8�3���Eb���`��E�)�u,��5��%*Ħd���B�:��B��b76�f�C(��<c=54ĥ��/�Ւ0���pN\n����Ĭ�[>`����k�G@�O��=yDbJ�1�K��:�X͔�(�y�e$"� 7ʙ֠�RuZ$��7�E�>x�dG��4*�kݧ�gR�^Q[�5vc�]�A���6t.���~�����%i�+�1��oPH�v镯��{�mY���"a�3"��nc����Z�ir�av��
8*NY-k@��p%V��4��os�B�4���J�W��+�*\�<�=�SXBi�G$�a����Ä��JK�]Ι���t��z�����D������2�)C�o)�^� vj�aZ���͙�}V�ڝ�WA��I3�AaMNjh����o���=x@{_e���7W0j���e-�l?���F�He�v�}��Б�A9�vM��>��N�4��w��%��HI<�Gh�e�B
�,���"{�]~EK��J�0<�Xq���u0x�B ��r�$�wJE�D�	V���v�_.��vx�ycˁ���=�����ٞ��X� �v��Aӯ�yC��h�d�r�Z6�$�����O8���X�!&&�}:BI~cH��%T��(.//U�`���3/U�����p8MbЗq�Q���d58���T2tT�"Q+=�
�v���}I�"�\�
d"�W���N�;�h�����aZP}�j�Ew�]�T^�i18�'���-��d��ռ� �S"�y�k�,��CK�on��$	/*��-�"g�?�v]�P�S��*Af+s����A�BӋ9��
������p�i���|��t��2�h9<-cq��<�sj	R��eh��%�^_ce�Io,��Ţ��o���S�k�e��eM�y�g�WY��(���d��S�F�O�=������?�Z�J��q@�YZL��}�ΝG�a�}����FYƉ�h��:;Y�<��^3��.��Pq�A9�4�?���|�t#]Ff.��e����72�j�y�JQZ8&�8!�h�hp�ji�(#�H��a�t�SX���2VhQ��&��}�{�N�^L\�6�:�p�������.����#C���0[�)WrAS����9��F��	��F�V�k�{��j���)%r-CA�4��=k�_S͸��Z��4;��y�Kok1f�=� 2��ߚS�V�����C����K����J��c�b
�e��H%4�]��ѨY��}��@<��86"���J��� 
���� m�z��8U���~�5��� ^3%�q�!-��:��V��S.���;�ݕ)�r�<���m��u�WD^��˗�̀M7� -����w�����MT�A� 	�$�����?������ᗿ�%�;a,��hB}�^��56�0�~�����h�úB��D��{)��	c.qݧ
� �����&��4����?�o���� �q��ṅ³��0�p�Z�
���W��+�m6�͛����?���!
������nly���CdMzt�կ���XC@�SX �̜Cߺ��l��Qt�Ӷ�}��M6��D.��=b�l�Փvlĩa�1Tk�����P����4l�ݎW��7��QiRP�6J����]��:��Y���Z�g�5*l��!̤&#��{o��ƞ��(�����k h�	�L�Ί*E̴CY4�hF)�pb�.�m�I�o�Z�Ě��Y)ïi
�A��^�n� �r��ȣ2�5(��k�2d�>ȋ2�[��rR����ه4F��]?U=Bl�m��'�޻nV7��U���!r�}���r�3�dTR�a�z�t!=�PQ)�U'<��{)�*�,���R>>��ר��m�XM1D�����8��>NSK#�dJў���o����;�v�����}Ž{w�<yB҆޿{�Xl6��*Y�ʈ�jhBS˞�7�ή�m��d}!�	�4��c���[�1W��,��4�O�L$x*�G7�'�����z��*�_�U5J�f5S�v�m-;#�qJ�n��o8�j>I�] =��\�˼E�*9���%!��L�����K[��,��y�Ⱦ��w0wm�$�����y�O�B�4�Q T%s$��Ґ*�q7��%L b�m"5�@_��0�u����k<�&t,�N�F}H6	k�+jp-5䣖�𐢷훵x�����z�i���
�ԫ�׾l��Z��S.�P-U&WJ؝�Lp�M!9���F�Z���Ҧ�l)��q�R�JpE}��a,ȘSQ��Ont��Yv��X�2,��x��*[���X[���k�Z=�D��^{��ŖG[e�S����	�3ҩ��g��z�-ر�
�E;9����w�"�,e#��Ϣ�v�17	n��I�l��k�D�enȼ�P����yE�	�	z�'q��K+��t�S>5�~�!�2��V8��/ބz�''S������O'Pb(*�
�(��gϞ�in� ���q��f�,D/��OcS����pN&�^��GZv��T!h��c�n��Ihy)��J��\�2��e)�JY����ˇ�@��J:��yƖ��f�T)�������
��*�!�yO�|U(��>��Z��ˣ���|"��H�l.͞�����|�Y�r�F64����."k1̃�-�c�a�$�s`�BPBކ���!�Jϵ�/�G��@Ԟ9�x���YX�����+�$xr^z鶋��4L����%X ό�u�u��º�u��fIjb�f�#=C�w�@z^�M�"��n�!N�Dt�\ړܫ�/��5�ds�n+�
�a���\���L���NH�����u/��"9z�W���Ur9o)�g\�3�����hO1���m'd+���t��/�K���B��c�K6�hI�r����;z�õ.���@$��az��&{u�LF�[#��ۍ$$ @��̤$%$���uct��VO:��ڜ�at-�υ�P>���@K+�W����{hJV�%y�h-{gM9�N���^�#�v��34n�b��h�Y���\H�txt5bv$�iɐeSA��V��FK.�i��q�-�}H�ӆ\��������o�����Պ�m���ln=}��T�~�y����o_|��7�_-ԖI6�z�fovKO��,d�OXd���e��"S�i8<Z��K��fuO"G���٬�f�������$v|/�M�*h�̅²��k;ly<�}�[�eC:KZp. (��3�~,(�n�D�)��X���!�,M4Q0�S�h��q�o�( ����fiT�83���ƕ�32�2�/x'�v�I�^�vP(��a�"A/�e�
}{d4{mF� �?��o��Zk;BQy�b� ��<�b��b��Y�m-e��C�����\��&���N�[�F���Q����)�kJ°S
W�}�(ٔ����lV-��U���e3ڝ��0�5Ď6o��4M�%�L�ٝG0r���m2	ڮ蔕�*��A�����g?�?��$	O"�N����'������<�A���e)h�pm�5Jz�f;��V�,Om=��Q%���`��Eɡ�!wZc�4l���s��H-\���I\&��Ҩ���K��̤�v6��Ii���m��������fLu�vG��-�m�d��|�=~L�)G?�f6��0����?���Ǐ�����~��U�H|m��F��'%�|J�7�c숄���J]
}`��8����&�[��\��l +��6�y��l!8ڈ���E��{H��t~G�m�3�
}��m��q�rՅ�T�V���lś���$7{O>E.@%���j%���v��9])��-q��5���Q)�!9�K��7u[R_P�$�+�)��	@�)A�;�X&��7��4cr1�����-f>)���X୰�fv~�w貃�R ����"<�24��8���!uRm���OW���M� ݍ�#t5�Z�'�hHtٛWg�L�e��Y��>V�JH� �я�7��K����ұfLh��V�>Z��"�(�_��K/OAbpilgq��C,���.�dY������h6�j2���޽����/D�ȭYNL��t��	ǆ�.#�|:^�Dv�~��h�VS�JUT)V�	9����)���Ԙ��Z����_˗+2LeZMK#Z���-����^��K��%&����(Y��!B�۾�'� 4lO�8N���8�u�(�,��XE�#��s�?�Ϣ�ww�������:ቄ=M�/��є.IW���v*l�Z�}��|�� >�LQn���(��<-���CG�N���J�O�n��ߋ����q�o��v�����#����*'����yj���)�E�i�]�J=�F8>S��^s�C�z3E���S��`Qj	Z�H���������!<����t�S�`!�W���ċ2���yfq��ID�:��Y`�9\���-�2]�y�4��6��	���|�]�֬2Y%u:���Q�?r��
Kl8��q�z#���l`�� w���dB5U���sd���'S{������<Q�9gvrFP<�$��go�й7��4�y��-)��������l6J���?�� Ѩ7�R��D��/_��A�=i5���z�\6P�Q�IVR�	����T���M��`�X��M��$�r�:'E�Ns;`<T������,N�W���	���@J~;d��lĖ���,}��p�w�C���٩�r@�&1�n����㡄8�"�L�k�={6J�;�ý����^R�5`���v A3����
.��l��<�Q ^-��z4��{=������*�}�X����W����@���~��E���ŋ0���
�q ?WW�*x�s�Q�DҎo��G���S��r`��a	���hu`u����''��+_	f�ĺ`V����;s�!�Pe��>��l>����G�
����N73��s�ڻw2u���O�l1jk2]Zm��	����LJ���H�.COC��
\E됎�~���:}X���[t����(7
H��� � H\�&���k%@�ӷ�1!�b�{YJ>y��JJgF����<��ĎH9�O�<�ϖ��>� ,�:�	|?.?�#������m!��߿OS�=����ŕ��0`MKpp�Zw�e�(����o��o��/��j�$�^�x��g���͜��6��r��js�nyE~�:�$��<���z�8�B�q�0%�h����oNn���㏇�H_��_��F�	�\)�0$oD��ZY� �Kc�r7iJ���1G��ޤ�V�I2OO�^Nt��s!xi;@�ab!4h�PKJ���м���e9Z�ۃ�*ƃC���C�E�YB�A5D%6I�5�k�4��E�fu�� p\%�lh���W裷��F��݆�>���%f{-������Ǩ�O��hA3���p0�	LY�L֣0W�r��i������+df�H�\�$�@3Ğ)�p���Q�iBռ��%A�t�N�U�'?,zǃQ�Tc����i��qOù׊C�2��� ��o������?��C��4Z:�|C��d!3
�F�B���ٵ����A�+�q�h��P׏��DXr]�̕����e	�!�l)F x`y�HDppj�2Z�n���{�ڙ�C{��1d�pN�vT���9??������w�~ӂ�2u��������?������/��}�����;4Z �;ƋKN��։�m�C��!U0��Oh�	�j�_2��d�/Z�/�3����`�Z��od4�u-�����Z�6�҃n�,þ,2���M�͆NZ+Uon����K�$(��q�Ǔ=@V�UJ=�iA�f��a�~6�Z���$a�Ao�$�� ���i�ݜͨ�}�>��~MA9 ñ�,ɞf<���$�A�>�!��'p\���Yk�O��@�ƑM�>f�"p��~�<�`{Dľ��� 6E�h��]�O.�x������R��=D��g��y��&,6�-�ΣU}��sq���2��=(*P)�;�р������_a,�U�����. ��;�^�=i��::��(u��1��$�C�3KTˋ	͓V�pd��0q�>C�-�fZ>i�Ѡ0�2�c�U�����
�,�+�ŝxY��M��2<B9�c�T��v������+O�/*/
fN�9#^0
�M���ja�
�8})�ꊤ�|�}�P�K�&�=]%����öY2��NT�ă�H��*YN&[Ñ������ש�^FK�R�.�yX����"y�e,�k|������$�2��0���}ަ^y
��\�8`��l˗a2���sm�^kUT��(ɠiG+�Uˈ��H(���m�|:��ݡ�߫N�9q��.:���<�� 	KW:-��2a3&��D�qvt���5YT=:��xW�4؇6a���7q�
R��VF�I��a("�t�9y�YֱL��槗��9-ѨDj����0U���cE#Z	���}�J"aY���bޠ�/0�|��g�1k�0���^�׈�bRhO��t�cT]�
��C�������n���v��:�Q���i��v$�č�,�#�ع�퐄�m�f2�8�9j��O-M9P�d��j��FS��ե�Zg흃E{N������ٴ�;&��-2��y������ٛ�H�%�b��K�wWw��pf8�(	|� ����_p�H�tI��LoU]Kfe���2�g�B ��ʊ�p?ǎ��}�Q�ۿ}�Is
�ݺl(rMr�Ei�>&Ra�Ni���D<�A�x��}��B��������۽� ���l�[�x.��Ɖ0z�k*�Kǟ>B9� ��h_�r����1�v�&���_SW���,�I���=�����d��Kb�~٬��g2�'Q<ۛJJbs���u�1E;-cy�2������\�6�(��&�؋-���le2
��F���ByKRqQ��Iu�ս�DBK�9�m�]�����Y�k�t57n�d���=ӓ�>=?��n׮���Ch�XT����h���H$G��ӌΦ���nn��/�2�)�c�]doM� g�S櫦ˋ|���pڷ���^��Z�HE�;d�aÊ4qm��1�iI�d�If{%�Y���oM�� k��@:���o��?'��dl�3��u��=j���H7����ݻ���>���U�x$Y�1Bq��ɘ'�%rN8�$�U�[y�M칠YW��'Xɣ-�%qe��N��x�y�'�łd��>yft��?���5qĎ��?��s��~���۷Pt��Ѡ��N ���5����8A�-��e2>8���z)~Ѻ��8O:neB/��4w�*ŞK�M�9�Aےvږ�ۋ;	*�P�� �K�7D�PF�VV̗C�]U�����l7�r�ɚ7�O�(s�N�x�$�J�E)����^@&�|�8�h�:w1�҉U��T���IL��Ȕ��#X���I��d}��9射���N��خ70L��f%)�ٓG�<×Q���}��r�f;/�d��,]a>�Yu�ԇ����q���G��`fe�H�4d�"Vn�J`F!V�H�s�U�|����ݒy���`����Ç�L�4-�u���kr�|���b<b�Z���MVL���~3��)x���t2�����z4^�)ٵ��`N�q}�����f���k#2�$
[2�Q��&��mWň���x2+F�%�ɪ��.I�t�w�ll%M�mtyy�㏯��4��I���ݧ�t�]��Cwҋ�+�v�iƣ�觓���䝔���J��$1�GhD������㧏��.e�m'�F�iD���r�#حΜ��(�X0c�A�� i�
2q;`���yY�@�]J��٥bԱZ�����é���v?�:ܪ����w�������{-E�!VǌN<~�?�ӟN�%�-�z��#�TU[(^ů�2���1b�@���6�H͂.��̥X�LҘ�*J��<tG���]�f%�C�`Jg��IZQ��5��ELlJ23�'ӛ�:FT��H�
�mS�PT�W�$8028��ܥJc5|��m������-��!$�6�d:�ܹF�*�a�#Ɉ�?K�[Ȓ���$�MV� �I�1h�CC;���=[|ن�$�K>.�����������[������;>km�n;$��٥�����/�NN�����wuu��d�~�f�?�u���G�K�z�,e�w�O��ٗN�Zz�)vX.?~8�ܽ=��0A�^�����qU������fI*�Y�Y0K���AkjR��R�.�M���lR���^����Pn�`�鸈�2��t��q�]�ݶ���/��l6�r�w�*�޽���k����r-��5�vېm߆ػ�(���8M˺����b� ��b,����k�dr��ֶ�U!��)��u��O���NH��C�NV!�_3,*���Wd7ʐ��#3��iU�=\��p�j��頻�Z�yh��}��J!%����Um��znMk�����eR�y��)D����<�z�%J��Jx~��Dk��q@�����. ������L'�L*���s�r'Hn#�Lȑ!���F�9�Ðq9G��F#
�H������B^˖�����`��rə��Ί��B��qɵ�Wח�\|~�^�=������G�o #�,5'��x�g�r�W4'bVH�q
A>Kk�T"��[�DJ���B��\���kQ� *�����B`�@��*�}Ė��
���=yLK˓:*��{Y
��l�X��N1�4�ũg
�t��l����SYG9�?v���5�����%���l>�(|4*ȩv`��=�r*]k�I��O>�����G\�fI����;�I���7In�	��P�/�;��DפxhF�|5���ցYNjՆ��okd�WN
N�^.Ny�G�w��ap��M%%��Z!3���1�Y�|�RXaaO�Ȝ�1�Nr��[��P��Faj��#ё{��:�Ff%u��&:J%V:�K�Uz��SO2����6�W2�d�X]�����)�8�tJ�E؉or1��X}��ǫ>E^g�r
̇"�l�� XCv�	�5V"�_)�s�C�}�)��2�$^���2�Z�WB=3�𫬯��d�+{-<���%�=d(�A`PNl���2����h�W���@m�'���d܎�D-nPжG���5���xLc�h�m�Z�2.��GJ��*��i�q�M1��D�B~*V&(��Ue}��Q���7�
D��Kg1\x�L��Z�=���Mݖ�C��j��սv:���L�i�o�W�0�~ط��)�P��žC���|Q��.�^BH �]ff��7���Y���?o(�L!^:I�BHP�$KI����ޑ(�c2��]�Do#�����{��8tR@��}R��J��!�L����w�>Hi+Υy-��p������s��ʚ�%�*PIL�l0E�dK�\�ԲE8ч���q�����$����$�6]*+��t'���`D��ҵ#b��-���H�x���q0-!�"�[�!J)�qaڒ�Z��o��0Е���BMglei�̛�Gw���A�ʾ���^���aRקv������>� ���N��X�ˬ��v6m�#�n@ֿ��m�T���N�P������!�J`�ҋr.z�M˹�<Aε�a�r�Lȶ����"�&�B_Q������b�_����Ln,�)>����������}TLD�<���y���sS�f>z-z�
�*R4��<��W�
��zޖ@�����N\��V�Ks�K�]][
ǣ�hȱVa����N#�u�Y�>��H�A�NN�0ȘT�w�YCf�T�{;�R)�����7������V��[�B�zr�!�ޘi"���;�ܮ5��C����L&A׀�!p�d,�+F}@�dDF��ᢽci˶Z2�di��0�0���טb�7�����舤����##4g{S�2�f �B�;��M~ �tWS�S8������L��R6.O9#O�>O�Lv���	G����0d+�C���] ��-��H�M�D��P���5g�R�G��縭�� Xbe��C��٩�"�Ny����M�Ny�#}ጸ��^��So�i�̗3'	qP����Y���C9%���H^Gl��Od�ìb7`��T� q�8J�"���bN)��<�&PO�"���"|s��]y�`���k���A��a���]~Rr�}�/��s��0/^	�Ec����#3EA�7@�q���N� �h[�N���9e�1O&�J p̶�����&Q��~�����2V�L��  3�3k�Ĵ���Em~!<��a�~��O�>�b�~��\ϧU�\����L���䃃>N�D�E6k�DpX�Q!T"�T��N��1F���Wl
׉I���o�$�8Z�%w����W��W�^�^���I�l�bBg6�%�#F4:������=�?	��w��n;I#��u���If�=h9�'YƟ~���w:� ?Ewr-�*�Om70a�%�eYϴ2��1^��T�P��xM�З��u[5�"Ե�% �%���7!����m"W���J�᳉�>�g�>�8�tBa"��Aa2�����<�������@�T�Ӷ�xX����YP��p3ҩZ�#N���B��d�J���5R�/�,�qCu��L!��N�򇊀R+N�
0 \�����ͦ�3��U�&������Y��S�ُ'O��{��!���oI߾?�v�TH|�	�:Z��@6%(��&�h$�1�%@rz������~�ۯBN�O_G:�M
vX�I�;�`mÝ�=�/�iy�8BM;��5=0$���wa�^�`������&�+���h�	�F\V^�"TS�E�u��3^7�7��ie�v�YC��4��ċ�
������� .FL���%L48��@��N�ԙ�݇������WXB���5������¥�.���q��#���q��t��K?|�^ƌXh&y�>�iu}�#��9��H��{H�*��|>���C���BJ��FVp#>�\>=�M���.�h~�iS���挕��LFXV{`{�N�6lՆ�X98�;Z�w��b?��3�`.�aqT'���Z;U�_E�H�*��س��0��*�쥄+����L�2����17�������f��#u�W���G��Qp�/�eƤ��\x���^K�f-L5��.oH{�x�^�r�	�*�5lD���J<t`DN;Sp�@,�/8i=�8� ��'��l�<���ɑOEN2n�Ɇ�Í�ZGy8�I2`*�Nٝ|H���p��1�i�$�O���0ާ�"��O�&���Z�<��dr3�%0N<b[FI�	��e��q�rϜs�DDW��HL��H�)� g�[ ��V%�mؕ[
�$�������r�'E^Px�M�uSm˫�l��b��Xǎ�!ꛞ�`�,�R���L4[@�)0�Jyr�d��s2	�� ¸�	r��ի/I3J�6z��-��D}d�U��9y�OIq,Y��q�8��[�M�q�����t*�{�dPZ�ÌvLG�p�Pnבg��%Bx'�e0#ׁDb�	8pN�$�?}ϣjG��~Ld���<�N8Z����^�f"�]�����]�i>��h�8����Ԧ�ַ�)���'��Hv�k��i���z���G�EIܢ� LLN�A�=�s������I�0#Z����c�>�BC(�u#CP�ť��NA���@b�|��y���ܡ�TV[&
(���F$aEޒ:#��K�
��F.u21�,���e13F�ϴ����=��1���ST� �AH~���	�w{1���n�79=>b�KΖn�7i�FvʈȤc��h>��sN�獒�n2�Ox/�;�ڄN�%��1I��=H!�{VeQ�IWڶ$o�V���V�&���3� ��^F��2�7�L��� ��d
t����퍤�4%ag�]W�G���AZ\c����jȜ�V988�_�'�~^��G�F GE�Q�2� V��ڊ�beQ&��U��ȼ��I����(]�d&��zWIi�,��-0G�+F��I1�LF��r��Y����U�|���g�=?>>���:??��f�{B:����%�{�QIqa!,�;�oR
Ɩ�:�F��S�X�����&F���D����M�l�$c���8V��g�/��g����^�q)(K�׹צl���L��\�I����El ���F-$	�� ۊ�#-%�G�aH�m������V�H'<I:�b�هs�H��=��E>����6���A@�Z�?C����l�rruE�a�Vw��� D@J9�(�c�$w:KA���&_�  ��6��~������cKa�
�	x��2暚�m��{�Z��e�����8k˒E�C�Ғ_^&�:�f�"�d������u�1�Ptd�,#����	#3�7�$��Ί�H��2�`dW�R`����h�k����Zh�(�$'r!�	��<hpE�xk-Ĺ뵂7`����}�NC9%o��J�ik� ���Ѡ�o�3?xYv�I'>���P;�RJ�m��C�����D��HW���^t��'���H�:1��X�K��������+^.�h9�ҝ_|����7�$�|��m6���o�PP䭔�P�������f��1p\�f��S�Ёô���M��KT�=���;1�^�"O����w�t: Ȁ��1��>e����2)���e�f�ƷL���w��ȟ�ǧ���0���ۨ��Ǐ����ba^���'��4y$}�mk9h�W�.ĲӁi�ۥ����t���#Z��:�ș�"C�ORf�8�g
�Q�H�(N���4!��RБ�'�g��5 �	$���Jp�d��zU�m�Lt�� �w$l�B�#�0�$��C!)㥀M?&�{x���u�m�l$�r*14��>;��N��h7~*�*F��2 (���-��>��������a�	ԅ�I�l��q	,a����A�Z�3I�hq�R��?F~�L*�*/K�<�2'&���+�b}kQ����L��H��?�@�M�2-��ć;M�7 
X:VP|L*�F�lA��d��D]m߃���*�[	�A�Z�A'K�G����.��puZ�cBj�D#xT��#q�nʎk�Y�+p�2�M@rC�Y��&���N���z���,)�o��ms�y&����h˒En7	-���3�ͼ����`�]R����ߚݰ��76����:̈́�_��^Mq��5v^BG�Q�O�q"�ClE.�T�ҝ�SٸF�D�{a��x����5[Ki��"$�YC�D�(e@��}7��g>�M�SYݿ�2��_+;H�%��8�`Ӊ��W�K}P�/~���g�7G�.�ٟN�|��c�ȩ�cB^N�h���QY(ݮ�ap��ϝ��~ٮY}��P�J�V�*$��Oh�oڢ�Oln+��z��ĉC�7���4Bz������ZY�՘,��Bb^ڦ����Zx']L��Vzt�7�p�Ua;-L^�i[7��N�H8�O�0^ "�E�	(�-�Br��L{�s��
t��ꊱ���d�.M� ,�|}�=�|"����@�#D�/�� ��)]m'���wn34�v�t2�}�L�L�1�,�4׷wN�	�������:ŉ����s�\p��g�@�4~$ ��)Q�)��C3P� J7�B�,c��P����:=)H�|�xl����Yz��zͬ�~;�H'��W�`�̋�;�,6΂k��zð�+�:h�<v9�g�$j�N ��ݒ���g��a����r$lk�V�V�|]�)�'���{Ӆt�ʼ�O�68 9X7����0�`q�.j���dXȋB.�i7�ׁE���7m��dH�[̋&�F����FwZ.�A�j7(? k�����Pk:E_�>%���4ʿ�B�������1������Aq�ŋo޼ 6MCks�c��:�w�M�$�}Le�:m=XW�A<�#���mS����ћHdyfb�4c�f��#�1�@���&%oM�Z��v:G|�K}�'����U@�!ϸ��\P�B6�T�TA���g�K2I�I/����R�W�� �B��c�HFA�Y 4�#/_�����^��~����^ z�d�$l�*�.x�A>�]%'��_���D����e���D��f!+$�|T��^�ɗҰ�E�9�?�f��V��j�O����Z:%�Ha����А�f�&K���R�a�|�
��7�T�� HN���ZS,G��r�LBx{�w�����$��^��!�Һ0�I(�����w����� �zW���-�A5������|!�#�C]��X7H8:�����kuvD���B�a��A�� ;LT�q��������
�R���$<LU) 
'L���E��D0`8?�b7��9��&��V��c� �;���|	[+�fZ;�7a���$j�&P�����t^��W�X��µ�uJ	������p����*i�R����'�X�9;Kqv�Ӭ���X�DYM! E�X`�,�6s��n��+IBn:V&�$vV5�}��%�H�4+S�t��x蹸ǂA��|S7������ݻwj4��z��s�������<L:
��#��68iRA�Y}����^.]��l��;��J��M��-��ad"�2���o�1ſD��*���ƚ܏4vzz:�������&�`��Ss'`��<��$�}o'v��֯ʈ�޳�W.xsZ%9n����^�mmrHϿi*`��-a���';z\�[����v��:���fZ���gi�C�G��ԁ�3չe��pV!bS&��/��v/U�;T[M�X�I��W�#���B9'���BආL�{F<�@&Nϵݔv ������
u�lX2��
�K�STr��	�^�-/��pܥ���^�Fx�D9Iq{�2�`+�S�C�7���U�b'�?
2hԅ�n��&s���v����jG����R�@�`Sq\B7hF�	w����bi�G$!�5l}��e�.+�-E.t��)���ъ��;���A3��>�y���	L�j��EN��n�dza�.�z��֕aH���B��������Dd�Ÿ�圕�r�����@�#��AN�)7��>�Y�\�������w�;�nP8�w�;�:~�~�ˍ���CT�=��o� ��f���AR�<"��n�Ro�� A�/�ٹݷ{��E�N����S4_Ƿ����B��n��)Ã�<'{-��w�������h�i����t��.��O��8����8������F--E����O��VK�AY�"ܪ���t:��/ f�j�q���G��P�� �g���~s&���D����*�Ie̡Ϯs�7U8�N��H'�z�u�*�M�:mӆj��1��vp�!ܶ�<�>��#���,�*}�3�i��;�9.��dq�vo�j�Dt��~���;\PmZv��8uX]xʝ��#�e����.���'A��m[��ź2�7�!u�JI���F�@���v��5�����d@�k����nӘ�o��P��L4rM���t@d���dJ3��W2zu���۷o�]QX�8�q����˄�R�����\^_BEOK��c|���f27�t�rV�����E$'
Ϙ���(Dq��ܘyzz�������˻�ˆ���<�^rW������Ǽ��������ٮ���m�U9}`��wR��=�'��m9���A�p��`n9��z���ܸ,�ۮ���$��#�I ���1-�4�w<�G�;�+���X�p�Ϫy���������F�0N✣�,&�<RZE�����U�q�jW�˜�{$n�&Wŕ�8��ʊ%Eב�&y�v�,+��˞N�ۦ�qvv���[F��T&�5���y$�%���'�IdT�f{�<� ��5��dZO'���1"!�s_��4�H������L��J�"@���jj����j|<�|��'����_�n�c���z�s6l-T��,s���$�up�"u��u#� ��c��g8��`-�/J?���0c�h���L���mGb����t:e1)��������М��[�o6�7��zx�7rO�gV�ĵ�P�%�+I�P`g#:�I%�Or����m#Ƀ��Ƃ�y,�it���6	��o�K
�*�A�Ş���(L�{�����1�J�&��㣃˫�=�j�#FI���;{T����!k��0�Qb���qJ���rrt���I*���-V�%��sPI9[O[_�a��M��,ߐ����ù�K�S<:�"&�]/�ZV���Gj���	5)�m���I��$}|:�ӽ�d�HV��6��pAwH�N��8���J
�>��3��8اEhM]��\1޼~��ey�1�TPn��0e���?�*̗@`C*m���'#����$ ��+����+���/o�z��py�I-A�|�$΀gq�J�dq-u�Т�*q�jF#ʘ&`i]�,n�7mDq�(:�|�)
Y-��>K'���I�Ѵ���uI�S�/��O�5�u�޿��/�{��~�<�sZ\o�����4���R�,��A0̉��۲��������^�q%�Â���b�"�ߙ[e>��Z�RK ��2��oQ%��Le:3kS2��
�� ��잹�p_���@q�ݘ)7(.dX�A9r�%��Z��=��eȐ�9鵻*֩Y}��rJ��6��e��$�>�ۥk��u�#F��B��Y�����p���q������XItYb/�xچz�~&:�˜d�y���M���B,���u�	�@nI�H��I0�ӊ�I��h��3��ф�FS�!	-�*��ޱ�%�4����{�oʄ�@��؍%s�$!9�Y�w�6��./���K�{��<w�}D�U8P�9!��2�^�d��<Ͼu��r��,!�9�1��z�����tyź���eU�&$������|,�n|֒lC.:�on׍�dŹ4!,G���ŋ�W��6�����Ů���;9�'�e�b,����˻���G�$E�m��r�o{��DpO	)<�9A/9P���0$Zd;���i�"�z��H�����-c�hwȾ`|
������Q&�:�Q�ng��s���ÇI���ԏ�4?)=k��i���-i�s�3�6(���*�l�w��%�X8��C��"MJ��ȑL%"؋`
��o8G����@ȡ����ZPKCZYn�V`$C��u�0 @g�w�e������-�1�M�`�!�v�r,�"{;�V9�t�^\_��J� _���)��W�G�P�'�N�*-���Ʌ(<��'�+����I.���\F.��V��6q-�䈷H�C��j�d5X�6��qA���6t|�I$CK\+Q]{�?'�)�lnx�s��4�ĉiW�r�������Ue�<�8LǪ��}O�E[=��e
�8��-�)�N�R�s9_;%L��,�`��(��#�ף�*�a�hM�;M�·|1�ɒ�nP��@������.<�Y��!�ã�t��W�#��C�^��B�B�o,���tvOL[�&�Bj��!��W���
�*O$M{���+
yY��ct[8_�z��@_6�0g��DΞ�h*ؖ��6蝺G�s��gr�C}X�O�Ԅ#�`I�x����'68x�`�0�e&Fp%qC�[;2̨��N��҈������^���:���St���w�I󄌘e����Ų[�҅�d����	�#J�Nꦵl�0�C�(J�פ2N�V{���r
�h�NԜWT�z���m�0;�(��Y�VN፰I�dS�Þ���$@�_�f��i����_Vy��B�v����aC�*�t'`�-M�
*�-�6_OL�z�K���S���Ӯp�|��ka��X'%P�U;0�\0���n�瘥�Tu���9-?5~)@U��X,�mh���s���rs����ժ���B�����,�#poIL�yҰ�G{T�0�
�0 �B,d�A�#>���Y�Qq%�RKq���O�p����-%��6�$��h�믿~����O?����G�E�+ٟ##�r/��+�T�c$�N�fjg>M%v
D���msS� %�Tn�$��<%"�����R��hU�U᥷�)�|�I���8��F�����A9'�y<.�i����AN�����bZ��JI|�e|"�TY�ٳ��&p�6J�M{Gߘ����'��sZR�Az��5��ZA<k$�2���p�[�ޢ����v{;)�r��є�M��D#p���$�pY�@�)y~h���贈��	-�X,�̻�]�:�����O��H�Dλ)i��T��~��g?�����OȘm�v�4��
W	J����˗�
9x�+�a'��J�2>��O�zY�#��W�^�f����?����x��0%�ψ�"̛nA�E/:��A����()���=s�[�H����H%�R��r�`��@ ��w}���=����?����d/�#�K�3�F�6i�݁�x^y�h��{�N��`I+%���ӷӂ��C;A'���F���.HG����~Ǣ"z��@�(��@qM�2��~�CѶJ+�� ��m���Α�]�1 %���+�q�q=����$�Ppf1�J<{�R�!4[U��`�G�k�f~�v��ϼ�^��Q
}�d=��~Yx���S��H�t�C0�����isφ���R%��/���kԜ{� ?�'.�kk���C���A����e��tr,��NR��2`b�®[|	m���H+�&���0�*�W,�9�HJ����P���Br�q5��X4�6�SZ�y�,˚�y^���KZ�-Í�N�ӄ�.�Wܟ�x��b�����N&E�a_�_2�^"X.KC�L!��-n�/�/Vذ�B/�r� 8�W@�+�%M�H�$���:��<y�7�7_|������?�����ϸZ��r}{�l�W���%doi�^�'\1�ӟ!�?�]y��Ņ^��.��Ž�W&N�������H�V����fGGG��?�<E�#�8�{|pH+ �����t ��R��٨`.w�F�[�T|��W���'O�������������oJ��-������]������ A"C|_�����`���r��f��u�����[ �'��Z�l����E&0t�b�)�$�b��	�,�$�%6e! �0�'���#��b�^�����٬c�Чdƚ�@��aEd�MA���y�1иQy��vr݀p�,�h���ׁ�p,m�2�#O�Ľ�Lȓ�G�T�J�5���V__	��Δ�Wn�=�Ncn�Wf�Xኖ�1m?̞@�2��t�2?�M<h�����F����y^p��v�c%L���D1cn ����=Ҹ��PKL$}�
*�uy@� j����Ɏ�o�<�Ų���-QQ#Cm�-���=F�ڬ�����<��$�G>bd��YR�s�[�}�Ӣ�t%�! }rf��Hu�&��O)E��w8�r@�����)әQ�D�L���
a�� �n�u�D�E3� 3�*�b�v�WA��A(�C��o��ڞ-�ח�68����ݠd���/^f�܀�.�s� �o���\a�f";�Dne���O�F�>I��	�wAsj?�䋶��˯�"h4#]O?�^;ҹ}����b����b�~o�S^䒕U( ����!��i.�P6B8 �I������cXs�*�_o ��~PR���~hR��M;d!ML��=�ґCk������ ���|�\�H�k�S~eY1,)'���zڕ��i� G�P�`g���~ࣛ�Iq�"xQ8'5;f��{�-*v��߰�t��e�O�x�l>ɴ�aȓT���_�;���ĩ�W҇�d�������Q�Y����;S=�t�j��4����⇀�@�$�2����Fr�N�������@ ��''^�.���h�Z��"����P����2�#ϫ�7-� v5ڲ]�mdk�h�� '''O�<"?���w�7UY������|���\㚻������+T�����2M�6��no�K�o��zI.i3�YG��wG1g-c�1�S��� ���ş~x�ffҶ�ڴ����s9_g:��dcSW�wW��|6�"��\~�D��gҶ����$�Uݐ�F��2�`ͦ��Q�#8IxV�6�,�`��eq$��pZ�$�gМ����<���-פi;��F�I�=�K&�F{��8�T�*Jjݒ�mԸ.���sTo�bgH�6���=-��)HJ��O1N9:KWu�J̀�jˮ��Vm�ϧ��wۮ�ԏ2���o��[z��!���p i$�f�E\N(@��i�-�9�kH�%d���'L�S6���ˊXN�Z�V����.#��4�g��	"w���s)��џ����C/IZl��[�T���PR��4�/&t��ٷ�O�hR�i��[�B<��v_Br���Ѝ�"cw#s���3C�(T x%�sz\�x��5�n�'G��=uGґ��`Az�5;~�b�G���ц��d�q�7���[v9����ܯ�]3#+@���c��������Gcζ���7��w��!e�)��3:���'��{e�sEj�A��"I��|���ܘ3"�<����<��А=�MS�B��T�8N�˪��?\K�<�=��E�˗���AQ���c������kƭdI~�8Bk-�$�֬�(�jz:�t<�����[�[:���C��9z�dˊ�F9�z�dqA�mID�u�n/�^�ٌ6��8�����'�ﵠ�#'�����C�������9IWh�&�Wo`�(�|&�[��m��P�T"�f�T��M�A�؟?}���v@BB0ϩ�}C�줂H��x�.xy�	P�������~�Y�H��	]1�V�cD,H��X��Jyti_�"����-n�uu�����t(*���h݂������#w���l>�9w�&y��Ev���x�	u��Ɂ1�vRn�2̶���8�~.X:��9ZC7�z�C�Rݤ^���ۜ����F�1�QH#���Gq�~Ρ}u��/�3�,�!QF��������V�c�E������yP�vK��{E$�	Q���q�1`�8�(]��Ǌ!M
4��5���Ӓ,�J�Fd׀��1d�,7V0��R ��8c�6(#@�V9)s���l�'��B乼4�������4�}�+x���]��)$Q=�j4��iL�����讼W�X�昙 ���*A��MZ���P�Au���}�9�MvdAG���!Y#���#��[Z����_���777��H��������3�ggg�~��w?�xuuEzFv�k�(<�`���zT{��%�H[�Q1��p��}9::�jAf�s�vI&���#t�S8svq&��pJ�d`y{w~~��U�@�xC;�z%a�'�oo�.>>~�x>�����o{��^~�K�e���=����Ŗ�P�h�y6�yO�������o����Kl�������ѝ��?;�$B�$z��][n��8)@bژt3xQ}��q[�l��h�)Z����6�+f/i2���cEl�ʹ�������b�V���{�r��T���&���n�c�>`�z'O˳�������p�ʟ݃�!�E�bm��,��L9#+�t��Vd{!�-����iY���
=:���7�F�����"������L�+�c�tR�֐�6���{�u�|at��,$�J�83Ok�1sR��獼�aØ��,Vq$��Iy@$U4��|�����!��o�y�_�aG�YѲ���Y���Q��jct�yF��&tO�i�YA�f$Pͬ˴e���a�-�b�c����
` �ho����0�*�g�n�ڎ���j�:�r�6R(�ƃ����F,r#9Nȍ��E
A�07�[��t�0D�c���_;��H r�+�w�9�$�{��$�)v�X7��S��rV�$� Hf}"`�w^����6� �����Np��G� \��y��i2���wHZ
���|�m�<i'2L�$�|��Dff�&2��OE k�vL�b%0��ˀ��|c�
I�P�� �)�ܻ^Y���;��n��z^I|�jp�FI"�3�/q��k����]�� � ��N�n�B��6��åw﵅�����P#R<~n�W��A6�1���_����u����F��:<����v�x��A#8�\���0V@b��\����9t@���iO�k��@�Xl���no�{-#3�X����/�s�������1����)F�ⷍ��D~X�Fb6�{-d��Q�-m7�|�N:�ζ�6�D����-j��uhZl��7b�[��t��H¡&c�1�"��3�@Y�,8s�K�"g��˿��2w.3�|�=ngh9���7���w���wX�,�<�<:yL�h-�$��: c�\L�4X}��&3��w�&�����"��Bw�{vJ�IO1�\H�����>�y�������W�(�痣-8\b��8���@@���W5Ӑu����"�b��4�lw)��|��B6qϻP�x �>��<HK8E�C98I��~�����IL�h	�J��![��/� �Fێ��f ˶u��+yIe�!��J|RnT�[���Δ	�v>l�h�FnrA�ևd�~��V�>���h�qJ,@O�FƦVh�0�BRi{HP�B"���S����G`!����*�y��AZA������Y���eo�ǣG��
pi��E�Ng��/��Y#^ 9y�g�Hz����W_}Ew{}})!���)�FN��)4����W�����?����l�[�͉�/��cn�'I�KI�7�n������F]_�|���%d2fNƋ�ˋ��>�(/�u|ttD��>�����(��##;��f-�n�^!�����˗/{�Wp�3�@R�'�[�Z�/k��H���&(���fi����O��!�D�es�W�_q��.(n���sW
w޵���\�<`�Ƌ�!��p��y!uN�Q�q<ac<�<��I�H�Q�����ށMR�G���Iu�7\0��0LH�kό)`�^TT1(�����/1Hm��>�uI�D�J�O�B"�D��D�	��@���LWW7�s0	��5z'm:2;����~��ܲ��:e��m���dF�)�)���
�u�{%��D��.�vn.�$���{M��Aߍ��Ze�����-9%�����61���JV�Ϳ��b��|/I=�w��@� A�)VC�\;�I���D0�4�^Zs����@I5�N�����Kᶑ�u�~�[+�c%c%u��/>E� ��?,f�ôa�e$L�
�e�F��-�I�f�S���郆ǃqJ����̢�v�Y�Nz�,��y�!��𑣇)`�+P@&
�ĕK�/�� D���c?Hp��5�p���p�3�3mj~�������7o޾��T�BK5���'��ae���<xa(�5SkX�ցN�S6$8���F��~D=�=)�����l
�HF���'r�{�+}{����ޒ�Z��
I��Ĝy��Ʒo��T��
�������t�(�~���Z8=|~v�l8ci�I�LL��� :������>��j���ge�*���Δ<y$zxj���1`hHl�̸6@Y��Q��h�
�7$D��A�`%-�O'ׁ��T�@�!ӡ9����c[&0^Ka����	3b�b&.nMģq��(V&;Z�j���JcSZ�S�w�{&�py��LZ-zOJo�N3�/+�N;�Ӓ�����рj���by�I:FMH&�J�t�q�H'�'}m��Y���_�J�7�>~�xu���˱�3���2�F���Gj�\��	|��o�;^[�Ty!pcd��L��{N���d����iO���Ї�PU�1�\`�	����:d�AO$�i7� K�Q}�u�)��_��.�u������a�(��x&�l׷Vր��;�:����X���`���	F��Ĺ"�aP��4vjjdj&���g�+U����e�%��o�g�����/�� vY��r�^�1
q� 4�n��q�����ͽ�5ɽ��ütX���
'd��T:��r;�1%�lA�c�f��7nW�SS���P@�ts�?�x�T^�@�O�4 4m�ԛܷ�km_��q4�a"�*�0tռ:����w��'G�`;-�.��aT9'�q���#/:�����o�(��*�u�c�h��B0;��4�/
��8k&j�Ͳ1�eI�����i�6(��ag�ӄi�2��L2�y���8ܭSg���q�xI՟���@�g2@�E ��^A��s_�]�_���V���j�w�p-���a<�]h�Q�����dd
4�^,`߯۞��$|Y�95��t��d�;S
�?N&%A�Ͱ��5�^z.�-��o$]z��r*��j���Q�L��Xn�k��Z3�����~Z.���\�Ez�?�i�������_�VkK|����|�Zn���ϟ���k��sf��W��_�::<|�MF�C�K�=?���鎂DrƖ�OE�چ��8=���p�j���I1"����G����?��zA. �Vߦ̒K��jɼ�d�hr�I��W_ѓ�!�z=��ů�x
>s�;ie=::����v������͟��]ې����-N���_/\Vn����}i��<[�<]ڋ�AcP���$���/�\&�<{zB�V$�"ZK���2���n_z^Z@Β�w1ho�S&���"ׁ�v�c0({4=�|�N��ģq�7���ً/��"��7�u�R�Ps�^s*�3�����n�-�<ws�MY��|��>����?�ʢ�{��<����=��IS�gS�u������:;�������}�ߔ3F��x�D���ȧ�pr������/_���Ƞ�W�>	S%�L\�)7w��@_�^/�����˿\�Ϡs��q�o#I#B��L�e��a�R��c�L�dX�j}{}�o&�;=yL�#	��.��#CG��`.=��Y��V��L�D�f>/����<9P�ѣG'Y%��NaDH��>9��_���{ZIs����Z1���!5�M$�ǓOH)�k��l����Y��0���g�������وs��f���ݜ�,��dD���tys˸$z,�^�OG��Ǐ(d���;9V�t��9tB��Eն���M���g�L^��Fwr��s�-w����x��'���jg��,��G�=�5���MF��>�	�t��ۛN�)�ӓ#�cI�>	|j�3ΡiגXҹ@���r�<{YBǮ�}Iv�k;�T���	��`��@�y:k��'@ �1L7f��^]�B8ustt�J�6�O�<!�G�����i�iB�C�C�FD
��3��F�\��''���+��E{	Ii���E���r���Q�Of�y�U�n7�<c�@�0S�l3MH��\�M�S��5��@e@?0�=Q�!�C��q��$�=�l}���ͅĖ1���q���R�G��hT�$�O��v�%�`'�kE�;�5+g����6�x��YiY��YÄ��5
�S�g�G��l�.����V�����!rK��jN�f�d{��N��(Ԯ�A>*N���5�(]H�7v]]ݐ����k����𝅈���`��g�2�N{��n�ޅ�[��i¨���8E:�5R�C���"υ�'|BC b��ձN౪^��j�|�u��0jH�����$,	���N����G����pB֟4$-�Ic(�'��;B�Q�)I[�Ϧ�b�)�xB�Q�I�#�!�N���	�	��Wӟ07<�Elz��S��ݔ��	�y]p9,1�d#YR	;Ǘ�ȏ�H[�SǮ�<]���%��7��~�)��#|s�{R5y��M�����3:!���v�?%���vy�'���no��	ww�kZM ]�zy���9~\0&s�"�:�\ǇG]��}"��d2��)RHPo�#�@��'TP�-!��8��#H�&� ��ac�7۪��G���n.P��?TklL�FIoP�����y�{�ؑ������a	cd~#eV���k;�@;��B�j�t|0J�_5�FD�+�L���F���x�/��Ʉ�_1��C{�eN{����4�z���kap�r���	���n$�B��:y]!RJ+���a��2l�9�b_�@�C�\���܏�Ek��ˣ�C��(���S�����#1�{N�R��p���Iz�t�p2�L�!W�i!��C���������ɴ�'��li��8���Z�)N�$�k��m%��
P���aj wu#�qba�m�k'���3�;��#u��tVP��u4"��3ɲ�j�,�4A���a��Q��5�G��������&���J 0QS�a���\�g��m4A2	��E:pØ�+����Ss��$MaZ2���W��?q��b�%%�@��%3U*ề�v6E��Я�P�be�L���Ze6� *w�l ���3��%8Ғ��0����H����~qu+��M ��Z�������&C�7��V2h���hDaW4_RH�I"d�p�R'�h��H{�w�)�����m�z�=��I��S�:gۍx4Vey�z0�?L!�{DԌԏ��Ez�k���\�&�&|�wʺ"s����b[�g���mC���)�}�|G����ְcQ7��j�9�H '������05�2��W6O�����v� ���&r�eߑ���C/z\x3Mנ����i�k=�R<{Gf6u�D,⡎�N��W'����2$XyWb�@�$|)������#$!��+�u����@$F+r���ի��c
5�<:����c�����?��	i���c.#��g��Vpw�5�r�'yW�_���\�V�Rda������1;�����m��v�؝���E��Ն4�7���c��9V�jt?��;z��)��f"���'��*�l���8�AW;��ӟ���?�"�0�k��cy���゜㢐\�;`��������7oޟ����~|�}��~��/���O�����ϴ���J8�V[��ND�Ƀ���X[����5_�|I;r��&�
�t��YJ�0[(Iiҹ�=5�+Ɇ�o�]��yrr�y"B�plQ����7�|������}./Z?�{F�E�ʼt�Gے�?~�,��FIjH38k������O�����:gggg��克�/.H4u�,m��G��>����t����~��OW�8靴�t?o޼�E��Hutt��^O�	�[��A�I�SH@�~�H�.Q�e����o����f�?��}-3"]^p"A�OU�ȅ�|�2>}�����x��	0����LD��򔥅��K���tXq��h�hA��0R�PVzCf$?��}B�yyyI����YdS��,,�4�{ؓ�"�����K���'�=�ǂH&A�61+�B����%�-}�SҚ�~�Dnҥ��C���o6�*i>ڛ�8�|}WU
f�Ɠ��h���#o�L���aBn�q�F�^�E����̽6�̟����̢.4����̿#�v���G߻�n�'a�c�ܗ����0�R��(��q�0"[F2���VB$w]*a9��=B�L� �.��@���_I��9ww��4�&'^r��o�Pg�]a����!r�N�Ϟ=?�����g!�7��&���(��ȼ���zdj�@Q
Q��ڹqhXH�n�p�+����n?�����t!a�H�F�1h��9s?`Mc��0���ۆ��yCh�Ny����y��1t�/7L���CO	6�թ}���O�*��V�Y����\,<���N]���y��9�Qp��Rk�,�V���4�3���'n[��tZ��_�^�%IK%b�-��[��:H��S\0���]�V� �X��!�@��Q�8)�N��;M�i�,)���;�����m�Ʊ2�t�h[()R�b 4�Z�Zp����8Ŷ��G�� 4̈́u�*����@궵B,��1�\Z���p��f��������m�s�cm��nתe1�܆�_��p��9ޓf�+\��1�MHS���ڿb���ěɖyi*?<<;3���s�ku{%�P�w�ڶ�Qr�fq�0$ܤ������n�c[�u~!�	�U@=xg;I�D;��9qn�pI��S�) �<�d�<2D!ݬj��	���V�օ������8���y'Du':��b�H��P\xO/]̝6���{tiit�]��u�g�+g�F�:	#�A�4��g&՘�3�c���ГlC)�X.�Hjt�f��L�Rg1�a���+:E�vM���x��<�h���l7rH1)���q������ә�4�QN�
T+Dt $�R6i��,{#�A ��|r�M�$�.Ћ����F��	
�� ��*PE��0 ���+$��qpԪM�n��,~��ݻh��+�$j<��am���A\�3�\��Ńe�I��n�R7���e��%9���kGRI�k��H���:
�Rr^ag�rB��G���͠Y�|�~���JI�|��p?�^����1�������A�Ӝ��3���x2r;�.��ȫ�����Y�4�t[�.'�������7
8 ���d����eg����з�ڢ;m�u&4r>	���-��X8�X_s��A���_1c�m+�+Ar��X��?�[8������$��3�x�8L�����:9����!ybW�m�Mg����6�M\�����j*F�	Ȝ<?H�;�*ھo�i��əׄ`�Ӂ{�G�KBn h�HQ�NV1�*.���br �#����?Ip] ^
1���b|ܚgh-�0ۖ��\��h�������j�^ޛ���h0R��L
���}��@�R�H[v�`��-��w�Y���8��&�yv�ﲥ��z�)��})tl*�~6QL_AV������'�O�ǿ����~�H�u�B5����'�ųG���GO����|�{:"p?���޾}{{{��W��޼���]\�g��>{��/^}�ųg�F�ʁQri܄��|2NNO�X�4��g����������wM���������/髏Y�v�ݎi�W	KD:J��2��D$�?zqr|���	]���BSr��4:~r���x6�g�M(ޟN�?K��(�h��z	�r��M�˵����i�E����w<���#�/K��-��磏?�MI9g��$��,�7�qu�#�
�	��ے�1��_~���^>�$�;�Ұō0��U��t}>����z��z�B��GGG�ڴY�=�,�,��{WM&��}��:��G޿/���i�y1�ߟ.�'�����h 9��-kb���&Ƴ٘�����$��sVWk�$ ��ퟜ��}������ ���8��8���>���?�ok�����w�L��&ٯ��8d��k&5HZ�gn?���s�]_���뮝ϧ����իWP��?:9@�	9���1m=)�kˋ:AI��5�ū�����㴤d����>�����ؾ���H6h_f����!�CI �^��8�{�r�'��Bv�m��KMl_�U�xF-	E�:z�4�M[]�$�CU�W�{ځQэ
O�)�\�v}M��|�Y��]O�d��h���q��d���q�����������'��	��7�n����J�*��m��'���t�r����}v#[2�ٔ��=sZnW덀��EE����������h��`B:8���8k����m��^/�m�֭�I�$����������H�Y*d%�o�0Z�Q�ȗ�8�Z:��8>!��F�@�7o���ج�}��>AF,�b���Ѹ������}�<OR�}�胎=���1Ϯ��Q��0�kE��X�ům$rH$���m�4=�{����$N�9?D#���1̈́��-�?o*lD>| �E��O�=���Itĳ,�{*f�II=̦�� (
ě��K�*���	$�8Z�!��4.�\F�yk�X��O�G�c�_\��-��xJ'(/�����x������t���׆ZQ#Ί�#����5a
�����lr��Ղ��sM;Xc�.���[;h@�,W�26z���甪V�W [7��7-̷�G0g����B��m��X x@x�{���ԡ��R"[�4}�!�C;���֪S
��\�8�B^Ѻ4��r1[%ә�#��<#� S�'��d�����mq>�d�48+3�,3e��y�?�w�.@��5-��t��V��e¢��4֡Q�K ڶZ �iZ?zHi��X䭪��@�Ӗm@�E�� ���Rz��Yҏ=�=�J�8n�4�dƐ��ޔT�dT��Rc��s	�C��#��W�"�X��n��k�,�K'�	���DH0�T���� ]A�/db�{�[ґ�)\���"3*΄	g}ǾG[�do��6V�Gk�L�3Y��������rS5)2��}�߼�������i�d�eW9���U5ir��%h�����#ˏGZ<Z�=¥�-��KƬY��b!,J�k�[�g�j�ۍ!(����\��� �x@"�f�>,����3�\���OPC�@̪@7��E>b ^�����7̿n���L�����?��(�J ��doLw��j#d�Y�Y,�pe�-Y��D!A=_ ���~%ԥ)"�����@1"�â�<����M� �������X ŭen;Nb�ÆݛD��`1�7u�-�)���~E�#�4��#�%5�pП��V��~`kb�_���F�*�%��~��;�iɇl�����5G�{{L����V��B�,Ā�����]�!a�K�7;�8I��;�h��r�0�_$mr&��g�Ve��$L�2�e(Z�w�*n,�����J)����R�ӳ�� ��Rެ���"�jݑ���o8KD��.p�6ɀYbX�p�t��R��0�e���V� L�{Ehu�����.dBE����Z�r)��E�Z��4[�S<+�6�T��F}�;��[+��]®m�s@�9�m�}Z+;f��4V!���
�hk���!j�'��׸o��81��E̴kj̩EZ��A8Z�9w�^��onn� �`JǊ�n��r٤^����jQ:��ܳ�g����p��-�N�;�6$�QĜ9iz�0�w�On01ք�#�
[p��`���!�
�٩d�C��X'a9MڪZF�P���6Z�3U���l�^�2���3�>V����-�^���/��B��!Z���*�C0���p��)�-I��WQ�&H��oe$��'!iIh�����Gۊ-ӸY(B��ŋN�5��(�z�R���������$�ⴒ����dB��@���FL��������9-�O�G���=99���;ӂḓ ����S&�3��|��B�Cw+|4�w����b�AZ��b���_��_�O�=�썄+�-�2t�Z��eC�����e����ׯ%���Y=1'���¤[�Pa1g���3���������Ǐ�'�|���ܺS'�JZ�6F��|[��CJ_AK!�jLn4a"�c���m��pj0;��:%�qZڢ|��1f�%ҧ	�Aυ���0�wC��KRHR��$���V$_�碛Bb��L \]���`�e=І�E��TB�-j�P��D���'�ࡶ�ʿ�կ~��_?��NG$FB���$�X1�|���[@����+�G��@�XTdx�5�%gG���ie�f�<iE+I��~��g�ֆ���t�@YY����Ӗ��6������i%�XJOko�<�G��%Yz��P]p����� ��6`v �CS3�%b�H;�:�Q��X��7����//?b#��m�  ��})DrkB;�O�yv#�{�,	zޝ�?��qfp\6&�D����'�M��n��$0UT#�E7C� ��2�������ԚLJ	�3�-#X�'O���\O^������R��Pt�N��9݂d�����LU,���]�-1d�v�0���SQb��Tk,2�4[FU�|�Z�~F6�?h��u��ф! �G�
,F�U�#y/R5�߿��B1�P'Z�����2��d@��3̂ܽ �4��X�˞��۷�FE�k6e���[�,_��h�����Dwx}}=�t����BT�E{�����`�
�X��ZwX,9K�F�NR0�2�$�L�C�?�e���2���Ĝ{������
Sb�`ƅ�e�q�P/D>=��v^
��H�lzE��
B��C+zM/���53��h�^3��,�B�d�N{�w�P�ȘD���*>��2��P��Љb[�!β`�`�f��	�:o7��<X�F��ٿڟ���R�tN�Ob&�L�S7R���R{�, ��	�x���	7r�H�k��5�c�� R {�3��A���t�+UfI<#8X��t�"��O�s������{��tȖ��?��V���v{͝���	�?ϼ
n��}�瑅6�Rd�W��F1��0`�jy��
�\���V;~^`�cE�u��|(r���rB�1؉W��c��T�5c׀�ëQJ�^���+�����s{����m�m�#�)���/����k����抈t�Jf�B�c��@VI��
�9W�7��U���@��Y��ʲl��3������I�e�q.g�s�YY#��FMk��� ���q��$��̴�Ff\�<=���#E	F�@���5fVNw>�D�ݿp�����k�B��;������\i8�p�Y� `kx)DxZ�_�"(����!����8sMzsŦ���)��'��<���j�Ą�#݆�$z}�K�<Z�x�+��"�=���S߀+�,�`Pk�"i5P֔2��+���tx�^g�]h2�8 ����.���D� �� �>�xǊ�X�
KW����F�%3R�h�#]ļ�l��I����!ؔ�d
��/c=&
�k�N%3y�dę|y�2�r� Ӡ�H����ZQ:�iN� �p���]����l�����$�?�>B)���D�N&3�8�44�rKj~��_'���P��C o���]��G�\h�T�����t2���ک���4��<
�	3v�w%Y��2\�����%��<!1qM?�%�C�$gP�0��ʵ��tB���d���$<Hm�]��N����!EQ�+^0E*w��������)[�+9TM5�9����W~�������qWNSw��bSz�E�d4x�A\Sx����P<IrQ����\-�$n��N�mykJV��H��Ra�� GA�K�_�R���R�ڈg\!A�f8��*�%jy�3ݳǖWeL�Y�-N��3�i?zTIf=hG��`�۱��l���j�pd�r��g�Ǡ�����3X@��ea���nk���d�}THʹ���A�\L� F��xTb\Ѡ�駟~���(��׿~��P�!����F�Ԛ���/o%���w�H�t1;EK� t���65�;aF���ICB��A#���Wr�./�a��/�Fe@�J���Lq�L�h!�=��l���O�����pX�yUo��齃�vÁ4��K׷W��\�
���g�)jp�{������ɇ��߸.��غVr��xZ��MI6b����=<�7���v>�7�Nʊ��b��
�Jk1A�v�8�� wPu��7�듣=�����v�����?�M��7W�.ߟ��oW^�%�ք�O�"gy8:�������y��gV�U]�Ѡ˽�`����b�f��-��Ѭ�~���Ʒo��@���s�æۛM�߿�fk�+�x��膤F:><:��}�v��w�zB�h5I���}�����H�\t-d�f�l���2���x��୅��N=�R٣�J�"�k�����GO�s���x<���z��cfI�7ί}W��sk���I}��q߮_�~9���5������nq�Cp'�d�3 +�e�)���V춇��'�x��byMq½��'O���������f���ȆG������3R�t���v�`�����N�O��n}}���m5�j�t��"�3���v��˗��rqsM�r���������р����R��x+^;f<�����/���L�O�>���?�]c�A[�Z����M��xR�Y	=m�w�d�n�Ȇ���7p�y��<pI+�LH�������pz��sY��zA��,~��W��6<����pF����>�k�����.W�,�V�\��^�s�$������ݯ�����z�aC��1�L2��QŶ��5g���YMFc.;�:q����|6��_�~}~�t�zG|����9Q]��Xn6�{�����~��c��(ZZ�y@�x��|���lJ/��ʑ�wvv���ɽ�YYq\������������\��������|͌�2K�[�����lQɎ1�]��7G �)���b����E�gь�(F��,��6w9_0}�B�er���������
9��Qp50�W,b���CU�Hp,�]�� ����������I/���)W/�2�a�k�90��;I��ha9�)��5�!�֘t�p����1:r�Z���MG)EI��ZE��t���w���!��02��%��2 ��?�^y�U���0(���0p<բk/��fn��6V��(�]T��b8�kY�W�[P�<
���u��Y����,��Fe�����4RGKZh��Sf�Rǣ9��e�
4`OP�ʵ�kF�H4�̂֏���1gک�)x-(ܚ����Ĺ�\&z"�)xe��ּ�N�]�g��-,<"�vF�.n6uJ�uB��	���8f�J�x��ʤ�[���B^3���d�+eG8(���li��k>��`{o���̏��!�o�3C ���Y�rş�u#�%������P<������;=%EqsɎ�l�UCP�І>�v���:M�Z�T:N��m0��j��aܛ.�=�t�2s���R����>�S�m)9o��OON��Am2�I(&����9]�p�`Y���U�AF�ދ<N��Se���믿y{~!q� �w	��3&|E�CUVYLϒƠc��tJ�G�y g"ZVt#��o�p�|Z/��A{��Wed	
���**>�M���+��v�\d���@@�!̴�Vn7¥Z��#](~�ϓi �0BR���+$�`\N>p(ۗ:�/����&wi1�!B`�٬���9��4��`��6���؊�3f�����)i�K:Өr/��(a(1�^���L�g$ʽ	ea������drE�ׯ�7�a$�B�F"#�	�WNz&��kXz-eҢ�eUQ_��M�2h+�<��(��,Ͳ ��.��jݦ3�������-��!�h,>� �k�K�S�PSC�:��h1��\fH�ɭ�&,A���]��3d:@֞�e���{�`�cOq��շ�|h�5���"��hT4w[��=�V��m�J@��Cˬy&=��
&���d[��|�!.4���r\D��C���������$I��8���>�r|�rZ���R�%�p���\RN��@��f�`^��'2�"�H-K��3|Un7^�rYva����������iwv듷�IށDq�}��Ɯ"V��5�R���>M3Bq/͸m�7J�x!nC<i'}�N�Yd�)����Rc�N�VlkaF���&MHᲡ��:�!h�7���W�;���u��7���<�(Ac�yhs@k��f#!I6�J��)���5��+�=:%��u�r7��/Hw�RQ;R�8�Uz��G�S�s�t���ՔP$����Ȗ��>��S�
�*�Sz]\�����=O���`���`����2�?�0Ƈ`�;ÚHZ�v��e-��7-;�m�Vs ��^LNۻw� ����3޿�^�6�DvE$/Tg��K����+��� �h�ZF��CH3�� (��JH�Vb����k��X(�"�ӵ\]u2�r��Ւ��)u��X�G�}�駹xK]�%G�j�Yc��ݎ`e�~0}�ӧO�]&��<�G��X01���z��lhV�k�E��]����K���i�U��ސ��<]9bc�fn���P�!�A�� !���n����-"N��ˮ�9���_��V�1�2ݶ�2�CD��4��ܪ^!,��C��[8~�� ��T������|o��sp�`��b��Q��O{*�c ����$d<~�;�9==�����4!(�0'��h��W����k޼eV��t���Ԝ�e|���X�Q��~��=Zv��^ZB\�t�"'aľ4�Az=}��l�K�7ۧ�g��%�ʧP�il%��,r���x��#ڴ��2z=&�`�"T+s�L��yZއ��?�{!9�����?��U�#��� ʣ���Ey�]x�.��)�j)p�v�5�ˆ�R�M�Ck���e�^��l��f4��u�a�Jn�,�����w��ݣ�;kH�����y���E�������5��>�jGy�7�"����l+'��Gz^����'|��/���j�満�8���"��<���qL�}Q@N*��s.2� Ȏ[I��b�W��[Ak�F�����T��\Bڏ����.��8�5t�NE[Im6�:�����,K��D7�h�<����1��{{�Bv�Q�X���D�����KP����	ؠV�����Y�oe�9�\�+ڑ��,��&��&P\m���#w�|8��BE��8\�h�]<���=Z�&$� �A�A!A@�S���4��"��N����'�Bi�/��I���V7_*�J]$��uc�d���F+���eZU�x�60$��T:��VY��ۍ0,3TD%�S��m��X��\q��鳕���&�IE��*�v��,�Z�ߞ�,D�W�D��d���+e9��k޾mY������,aw�g���y�O��V�Q&��\��rBw�ؗ ����S��/��������K�6j9u}u	dM���-�פ霒~���<��a������֛�k���s�߀뚜����B-VK����%S/�t;T�{ƶ��q� C.Dsv�.//X���@�h��1�p ���e���]^��ꫯ�zEi�r��B$�FW��"S��l;�>g���Xn���d�Y6�� �븘��Rc5̈́���X���V�[7�|�r��?���;��J�X� �t:���b��cs&���`Q$t�ۛ�X���T�<��Zm�+��CY��Ǚ*c�\-d~]��w������$�@��]4�
��4,m����&s�AQ��F��Y7.vzƘ�S������tv����U��\	�#ti���V���-�P�9�����z�����;H����pU�fc����9�f�B&�z�Y������&�	7.���˗^TB���^`�����5X�O���~$0f�>�rj��6 .��2k�שǽ"�w@k�j�[Rh�pr^o��A��A��~o����%L�O�����UF�X��O��Sf�÷���r���4[�%Pz�F�d����%8�<�R�ۋ<28Z��i�VF�	���b�������a��H9	�����o*��0�
�K�X�6铚i`�ƭ�l^��%�3ʽ0Lm����R�R�Y,��`n�kˏ�H��]uI�0}Җ)�8h���
L�9"؞��1±WG��a�L�'�����!��h�c�HCQ8���6���,���M�s�o���,KvY����J�����Nw)��_gw��ma��(��ئ�*�s�<,�ڡ��d����C��{�������&����"X��L��@W�2gV����W)�-wԗ%7���}��c��_<�G�aϦ��T�� �9����%8�R�.J��k~�9-f�+��옴e��Y9d�-噹�Y�I��	�-�p�J*m�l���x��m�Wm�h�s����<!n�l7����f������]��'��+��:99z�ӥ�����u�������1�2�˺�7��/W�����7�Ų�VUV���`p�?�?����/�X=�UF���łL`U	34�Z�Ir~�ŭ�P[V�d:,�UY/[������� ߈#y�1��l��(y��F�'K s.�כ�v����̗�-��ݶE�1t�d��?��M�K� �UFg��[�d��2�R��������Z���S\����`>���1�Di�P�/���kZ�!��(����_���bJx�:$g��6�]��n�}[��,ڵ�4ź�o���v�Lh1no���n+9r@��dt�8fb(,�[O/vHR)I��r����q�J�PҙشP����uOF�:��?���Z���xȉwF��ݙ<�T���lP�#F����F���p���6x��*�g �0�VӇ|_�eur||tp���v=P��~p^��g�ů�,-��	�{�v������0B�II0֫�D��vP��1� ��ԯ�s�/��Z�<����(��`�Y�Zr����+��G��^"`�����ɫ���F����6<����n�+ϕ`J��uI���F<D��L\�e\hmH'�͠�����fД���fI2��&����\���?��~�{䭎&E�o(ॗ����t�}Φ�䅪�pTW#m����b�Y��B���Q��)��\)����y.y�@�W�8GI;�	�R\�ׯ_?y�$��?!�7}d��T�^�"бנ����$�]o�t�����1c����H���>;;CD�,�H�����у�/unC& ���HC\�}U��x���zLn�(�#���eP��6���B*dL`����<����<�S�;|G'�#��f�@T�T%���j�~}�=��L���Tf	����;n���8+��=�ippUK��ܺfOZz�`tn5�ⴠ�9�����p�S� �n�,�)?���ײ��$~K��4��� 	�D��T� QO˺�[�FH�����3|����1�%�RG�}��Y]5pq���iq1A{���A?���N'8wh�˴ ly�BYeQ��:|@FZU�]��!��)i5>γX��\g��CRwIVh���\Gc)�
��ZE_+$�{�5i�[�/h��+ܵO:�sl:|�o�ne��TǙ���(��h�^�_:�Bo����/_�o�S&�Xr��ɣ�I5�}K)%b�:�o�͗�q=��6J�Xd��	f$�������Q�it%�������2NA��j�-d���K�]od�j@j�K���������hF�����u�(_UY��t2=U1�0[�W�^�z��$�~L��m�f��\���V�2�e {q[�?z��֍�Z�c��$��|�Ю��XlE�%d�R	�B��v�B-��e��.�'J���EKmf�){��^<z�h:���ʁk&/�8��͐ҰT2G�&QĠ�%��w�.��5��%�����q)t���̧#��k0�y�� ��&Қ��ѭ��|��ه�@Α$\�7e�A����\k��0�X�(f�]�<@�whxӓhDeD��f�B����w@��	���V�켎�@�Av?�2�c�e�a3,�!�#V�uiA��IM�����8)!V �e�Z�C�m�H-��1x�r�e�d�N�������$ߍ�^�vy=��N]~7!x'5fɄ��x����΢e��΂�q��2�pY@�fK�g�l�"ٮ�7^^ ���I���"XD_�f�v�;���xp�@��F���rc����"��{�02� ���C�t'��bo�[:��}��l��]*Ss\5>[�w�5جI�6uIf�T |�(1��0�QB&�@�h�tǍ�S�w����}B
�t8�=j�5�rdR#-��usm,%BH�M^5>i�PL�3�Y��-�6��A���������R�LH����ْ�(��k�t�G�n���g�r��ԡ}x�7����`�1�u��ڹI��ۄ뺴1K���9�ER�ʹbo�G���vD-3h~q�xI�Z��2iF��F��TE��Ci��>��M��X��6�cK?�w��*Φ`�Z7/^���P\J_J�L�v6�D���Q�k��?����g����.���Ԋ���-�623�]u�[ PXi�`lZ-��0H�x���.���s�F�f莔��b���q��x�0��%�ǬK�*�ӿ�F�)�ѧ��Yx�h��(����M~��}f�z��������{'f	Hd
�tHVcL< wm���3r
a,i!�t/��c��VH��ʁ�_x��L%1]���'�R��N�g$p�D"�p�^��|�����{�.��F��9��.����$������D(\m!<ƣP�/���L�]�J�'��]��EkA�_�:���3|�o�6��ǧ���0�*��H�d%�\�𥂠!W�b:�ɚp���f�UE:�T�X�	��~�͆���ї�+G����ϟ?�aj���)�--)xj�- �L+]ƕ<x��XpC\*u���^�f��{�d:�2;���(����q!6�I�.�m�8X�ô��]��qD���p�AhA�Co�o�CDK�I����O�3�(��ъ�Bf�Hg�w���l�&�O&O&,�N���W|��@����z�Ȝ�d��Xq��(������;�)E��\g�C��;�'�AhCQ�e�0�Ι�A�V0�2����vB���������pvv$S�g���V����m&�4�����8�C��D��
oy�B�y��Z�h2L��Q����SG)�@��Jb�vM�̈���E�`�"��'�e᪲�D8�	vU���f���-G�ϼ�\��t����cQ��V�{&֜LG�{-uk�#3:�a�r�
	F��J�"-0�R�)iE��GK����9	�<7�W�rRz�Tš�z�X��y��۾8ŉ�\*yt��S�:�x�A�)�n\`�Bk��q��x�]1;NKp���mB�C�8�P������:�P�B������N:̷����c�pX��V��2����*�sP�x�4F�*��j�A�Z��u&�ja	��2���8n�x|�}D�I�9:À�B�f�Ǉ�4O�P�'��L�`�lѴe�\�L���B�M]Bv���[��rnv
Wk�#"#��<�,)�r"�j�Y��w�s�5���~��"c/�7_>����>�EQÜmĚoVK�4� � ��b�ՠ�����m�b�bSfHѵ=|�C��ypda]��>?˧��5�{wA/ ��A�2�߾���y�ݻ��Y;��9�y$zLuC^�~�HN�ө��r0@y�����Vi����8�G��Jz����[�M)$^�4V����P��4����Y_�R��ʑZ��R*���������f���1�&��Gv
Մ��"��7`���ߨpp�M��m�����΢|o��'L��^�J�0m��7���P��-?Π�� �"&f:,��q��Q$�Z�~
Ѡ��h��J$�l�>��.���A<���IW��q�.�GK��J.5Cww��b���(w +��J(F9nѳ2���z ߈r���I�y 8S���l���0U_|�!*CR���}�V�A~���y��lx�0 ��t6T:(����	'��;ʻ!�\�'���z$m��U| IМ�y�/�6![Z	l��HT�ܠ	�Vzb,K�+RL>,���Na�y�c���,GHX�2��i:�%9Đ<:�iΦ��LG	�)S�_KAn'��.�K�3ť9�`��� 9�M�t��R�54cM<�U3U�xHf� �hX��I��e���
ӻ�?3>�T#9��J���h2A���W.I�>�Vu��2�@������/� E��E�U�j�{G��P>�Ȫe��ɕ���o���גq��@����Z����ڐ3�R�jt��B¯lN��҄��s��
Ѵ��������h���Τ��`��%�Ό�@����Ax�&F���q�L��Z�2��n~��Ӊ��	Q��r�|�V�$������[�oM�Ŵ�Q�-
^_͊)<�`�a��!T�-H����gt����j7�Ձ��8��i�N��,�^�}������G�y���w\�^�6�^釬p=38
23W 1��)��pG+��S�����xn6���}�͛�����w������w����;^3!�%�?�g7������{���4חW������|SE(հ �b8���A�P���r�ޚj��|��T0����+��)���j�����e�vm��j��T���f�"ʰ�a3�/���k$�ǋ��J:.3pJ��f{��|�`����zq1hF���d�C�)���rE����� ,�-
�!�ő�G�t%�S�������d@�G֚�e�Sz��LR�9���*�U��ߓ���r�X�J���u�,����C^�t���n�ڠ�R����HW���{}�mi������l2�R^P��2�hD��do�We3�����D�b���ӎ��i�`)�eUz9���v���]��
���	�� <������2�Rz��|ssE"���1諸��:��p4�x���!,~2�.�m�XfA���u�v�-nuY��ӷ�����h�::��77�YY�d1�@H�s^V�p�}�][�<5��;�5c�
���Y�˂$���I�H��P�[RL~��u(��up,ruVȷ�����L���f}G��ʣf6Qh�v��,W�Q3�RG�5׹l���ٮrב�{���E�Z�iIi�XG9��d�XI��|�[�y�]�n�z�hE�yA��ey_7���7X!t#wE��1��*���P����܉d{����	���Mqx�wp0�뽽���8���R	���U$k���㽛G�����-�r4m�UYk�H�є��6�CD�g�Z:�+�+�&U2lh�!w�6���9���d�������͖���#�<�]��3߭��?��G�}��N6;���XG��W�`#ݸ���.��������3A�\��múi�����g��N��3��*��p�5�d������u���V�ǡ4� ���~4v�uV����c@
�����IX�����C��y	ÊKjjn��)��5��z�,�ރ�'��z�MU���@{��L�Ԯ%o�QPGg��?���lʰ*�H�o�-y�߼zA�OG��5b�v��U��3���:x��ӣnȍ{}�w�t\�)�u�ɋ��=�6��J�SaP垜�����m���tt}L��a��A���Dmd6=ݯ��'�T1!�D�նe�wH~�gjN
�i�H�<�������j���$���9
i�1�pk�6����p�ܾ���	ʆ)j򒶄���S:�Y��� [O�c���M�d��q���r��ޫ�Ƴ���5]���#�«�F���9��RG��0g=KFnt�m�L˘,F���x��P6#�F���[�Z����8Y���{2L���-��:8��xIpIE��2�P����{�e%�@& Yƿ��1LIt0y�H�1����߲�'�sף�7��b��R�hLz����ݶcp~ù�6"n�K�<�`���^�cXb�I̧Ӊ�0�S<.�Ó�m��y��̦��6��xBQ69��f��D+^j{����)�ݝL��J9-�Z���%)g�):%���)R��%��[��(��%O�J��-U�k����Ձ]�� ���͚��K�It�C#I`�1���_�v�X[���A�6f�u�Z��3/^~#�6݆���w/��1��|��b�H�7t�|{�� �&���V��<=�s0�iܽ{�W�ע"����M��Oz�����/��D��u���t�Z�F�ܨ�h���$5��d1yw�6H�9�8 O�~t||L���qP`Px�
�v�.4FS��5V��Md��������׿��>�g?��ׯ_���7Mg��G�{y��|qM�Ü��"�f8O'�^�+��9��r��y'���7��h��jQ���v:�G�j�->m]�dX.�X(�g�lk��Y,_����W#A&:�l7[��
��Z�U.?�;��+}�6Zኙ��Ȇ��D��a �>0z�0���Y:��+ �ԲQ"��~��{'?��)��+ɂmY{���<̂B3/������1X��.� ���H�p�+2�ۮ��Z�\L�gHՎc
F��e�(H˕�H ̥��m8�YY�x&Z���]����m�ge����l&G@�7\M��w`@&�4�p0m��l
��1��Ά�!#�	%m*�=��*8�]�0��6�uNγ��-'�{�$�M�.�G������7yt$��\�✔�#=߲�&���X�,2�H��Lw����b�zQ�t19��Zd8��N�⌣����i�_l�Y�-[Ą]Y�/���~��R�b5
fܖ�6]��|3��^J�֐��bh�ܰ�b�#�%þa��5#�0�H}`Y�R]{�칆�1���*+CR��$L�oWI,I���"'�WR`s����;�]T�}�^co$xZiw���bq��K�<2��`��tj6_Rl&ށd3�#�b_�ydt�� ����Y𦹎+@��_/#Z
�ߐB)$K"7�(/Ev��jp��BN�[�*o�K�&�Z��&�Y�R�w}��w����.6x
/Wb��V�إp�!2�n/��������JB��~6��d���"iض²}������m�a���	���~��Fo9%���H��X��ɥS�]p�$5}��ـ*^IP����`l�����3�@Tg"��Й�̣��������l�TJ���YU�S	
�8�z�s\�S��^��P'٬#���}��!���-���A�MV<��c<��B"ҟ���_|񅬞_lW��Iᣣ#���DXp�ȥ,a���4XRp�Hof��kwB�{`���7o7L%/+J�D/@�5s;�h�0( �3 T�~�C4��2Q��{�Mo0�Q�s0pv Φ�����9�}���xBo��:�pM8�C}��>� �5!ߑ����Tb@qe�xB�A�{�����
�~�m�I�6��>�\aS�hKa���!�l��L���,���K��2Iz�e-
7��;s� �+������-PX�Y��r�2| �� ~><<$�@��$��;H��^/�������#0�̆GV8��w{���w�|�� 	3=O�XTb �PB��r��B�Oak<���`�.��e㕈uZh�n�������<�:�{Z�M�c�Ӂ\Ç�2�^?��/��_iO��0p4��{�<'���X!���'�z�s.ٜ5ʹ��f���iyZ+�p��8��Gz�)x�I��gn���Ǉh���o��[������ �#�hɨI�pvr���u���Q0Έ�s�~
nDHz!��J�ܝ��r���-4���8��CJ��Mi��a+jò��������|6[n�#�X�=�w��x�~�v3���Y&�唨F�pU	�҉�IE��F�#7 �m�Ʉ���˅��hcͨ��)�+�����V�j�F""X�*;�tfI�<����8�~���;`9�*1D�C8� ����l2��3�E͐ioZ�i��L
���I���8o�A9�Y����ۋ9������@/I�B�W�R���I��V�>pnzӱ�Q�µ���$��`FE�ъո,����J)���;�y#(���Ĝ�>i8�$���1�*�pٓ��̋3`W��{��N�í���f<�EM|��*��I'����� �o$>���\|}�IZ.$�z��5[�Mk����0\I*��/���[�h@_�_������4�)|,�m�@KVH�`��Π_�&�!�r�����B�Cw\��Ah����ekG�k6��g&��H���!��rRff���Pz/�H���-�	V��ѱ.���������Df��c,}������bd\U:�8���ۭ؎Z�O'^��MX�)�\g��J_ˍ��2.V��߶[�B4(�����¤��C٩,�p)��@Ha�&�:�����W�ON����k���/���+��W��!�5��Б8P�(�qc�p�ҽ������?��_��K�O����/��/nn/�&!B$K`E����k�\��E�Ԏ+'�4P�����G�N��%�zC8�H#&�i�d�/��uJӄ#P(�5� `#c�����п7W� 9��l��Н�m*�8ѻ�uÑ�H����(U}Dm�.�D����J,UM��B~E3�C9 ���J��V��}���C�u�d[��}��4����>�p���YD��#$��p� nεJ��q�_U��$RZ�\�o�q��@�
��ꩮ�	�f���W�3 <�˄ {)�r�ʄ�V���Vu'�S�Դ�2A�h��g�_h���t��B��^'ܗ���+!yˈ���!���\�����[�a4y��#�����}�x� i�'��W�pK�������x�qό N�y�!iF��zm�L}�*醴���-܆�L� �ľx1�ɕ-WP���`��]�����I6����)�-��!�q�'n�)���'SN�r��ǌr���#�USQq|�H5���!/�lɛ�� �]�S�)!�t0��a7��>����>g��7l�r�G/?p6��zt���o���Pu@��:�J�_�%�^�ڝf���Nޠ��]��T��ۇcš\2�4���b�����e�>\�L��xb�KBE@�\��ED$�O���VY2��@vs�jڼ	��b2m`��)�ܒ�����jS�i�I˿�e椶;F�� `d֑����]c�G��-IסA	�� ^�������p Zγl��w�0����Fz�A��S3ވ�[���#���ε�v3�v�@r��Dް�ܺ�^y����pt\����I����9+8�����*h���GGG��)ͫ.��Yؗ{�3�><�G�(����B�N	��j�=wq�4Z&���unQW��xr޿������i�ϟ?oꑥ2;!���9�3�����1#[�e2�$�%�߀hܲ�r�W�<7��lK���W��o��e�zȅ�*��M7��������
���%�5�c*��Y�uL�p<-��ju�))Kr�oo\v�F�,�+�H�յ��z<�����V�\t/�!�;.�.97��z#�X9�%z.I!oEbCW{u}�����A�����#�����%Id�����Nh�d��Ȗ���˅o��l�U�[�����]�d�7��]ܻwo8��r���{�{���.4��XNDKD�V*w��9�����հ����:,߼aD 2S����̞#'�o�Խx�X`����J��R&�\��K<��f�+�Q��S�����n�|@tǘ^�J��N�˼�#�
��S`�������/߽~��+k�|莫rX�S�~FVy|�����������B�J�3Z�F�I� h	�i�/]���`j���1�����bM�3E���n:�#Y]-6�.k�b��d�������l��a^��(n-�a3����ۛ��ջl5_1��@x�%)���)7(TRv=�}+��yᐛ�\O�W}��N��Yq@"�ʰgH����L�{�j��!V�����b̋�}�50$轓ǥ���0/�@:�ѐ;�f�u��5�^��=�&yE;	O1���j��^PcNSf�����?����z�����?��?V�$�m�r�˪@~�>M �|�	ɋ�K�n����:�G�JI�����~3t#x]���m߿O��}�9=/���d��p�i��atͯ�W�'����/����[�2-Z��c(K
-�Vv;�����2�h2Y�tf�=�i[.,>=�_\p����g ���&���(�^K�qRjK>�ageQ��PV�^i�m\�_��y�4p���i��{��g�󛻂����� �G2�_��B8���ɹ�3�zN&cxh�㒧�j�!>m�u�D��;�0�`�i� �������ut��F��%j�=v�z�$2��ί�D,�
J��6����":�{��4Ո#)aZ\�N'�ү��-l��;q�8�NF�v��z+}3�o6N���g���Y.�w-�.���%mM��*������p���j����a)�gv��#BK��������-�A�a����H�@���9��ޝ��j��=H1��,�	9�=���[�
�o8b�wG2���3Z%R�� �x��g�}���O�����_��G?�").�����Z��W��G�-��,�Q�Ŧ��L�����d�܋�a	�w��N�կ���(5It�q�ᣲ�nUAJ����Q�z]�(�I��Zrm�;�r�u����?�iܠf���Թ=�RůA��Z����G��MjRugA�:��
��q����>�������л��$�~������nz-DΕ?��~�]m[&�.Ɔ.������ґ��SJ��d���r;oW��dnܽA�EH;��q����Mo\d[o�$��_sus�{�zyu+��@>w�)�\�=]���	�L9ڛH���m�r�@�&K. B�r���(+n �}����WR�^:�
q]C砮!�/U� br:��2�����C�i
��K錥�N�&��f����!�c�YJ��F!�vH�,v QSޖ�0�����y�.��t6��`���>X�%�S''��e�)�m��%Y`�?1φ��K���+��qf����s��Iz����gSj�*t>Am@���ۀ��ԏ\�t�]��Y�eH�W�H݂�Qi��JÒmm"m�lۦ��t	�pm����A�5���A�gc�������&�R������l�ԉ��3�5�wJ9q���CBAÈRf�Y�"�J�l����hagv�k��P���V�}��7�EF�c*���%��Ӂ�_�6;j_K�mL:ű۸$��U�Ԙ�GP���S��	�$n�:�?�]�E�N�pmI��������T=?99��r��5�>�����ɒ�<�Z�D�J�##�.�]��n�4;�I���)�`��d����fq�?�S�){&J�"�I�,��^��l�:�6��*�~6�̎.!WI��/^|���ݖ3�� )
N[ 
�tLX%\��?e���ʗ����ի�۹\	/��gO��TU��G	�J	SZb��#KO���r��/�^�e<^S��CX��6���K��D>�So{W�Gج�K����O�<q
�U'�G�R��n�R�(y��>�H[h�F���9� ��k.E߾y�|q'�% ��::�feT,���~2\!`�xXd�x-�$����K���,�B�����?�~��d����X��j)�(���St��16f�k	,��ƵU#��-t��5лHX�`��xr+��~Q�[��KNh��9�^�rs[�]���Yi�h�l��iR��V�l�#�4(�E��{zi3�AԂ���3���ԯu]�3/_��dJx�4R��ِ�������SK���u>��6�2D2r׻��Ƚe!:��� �[�@r������-7���'��m.�������2���UD��щ���p���qܶ��BM��^�>�ma�t�l���R@�Q�r�@fF���,�5���!-<jS΂�"$Q>�/�YCȄw	�P������.�cn��1R+�b���n��g�PH�)�k��\���&���L�8���t�����I�g�}(+��,�@7��5$ɦ�S�%u�����X�:2/�]�P|�\j�`$��� �b�SB��F�QY�,�������`���y�����`=qL���I�֞�|p�� ��!r��D��v�<(�|�6=z~����R���v�vc+�Z�|�2����},#�N��J���Hd�P`�� 7�7�ę���Z������F�� �K&]�����U������C$�/�i+@H�Vy�<9}zd2��<6Y1#�Kc3����K ���� mq��4�b*��&_k��"�Bi.���Af)�������1$wF�+K�-L�)��#";�a{+w�1��N���H7N�N����s������gO�����+�vX�8��P�u��B%0�M]s?��%	k�C�+��J{P܆o����B/Sn�p��!������.��7�.�02g�'򚎏�g�����������j����^O����"�� �=|���r��6�L7�?P��,���lA�F��/�z�4:;�9}��HR�`�\M�}]���V&����aI�W-�,�7�������3K��W /�Rl��vN�?��J�8 �R���	p  ��IDAT�N�Z}d�Ow��T��2%�����8�KFMP�7���;v�����sgB:�\3�U#�1�+b<�#=���놋ǧ�����C��ˆ�4/����A�����X�����j�H$���T�%�'9D�[�L��\�ڄ���l�K)��EZ@jk���<�Fg�f�R������	����f���4�,�����"�T`+=M]�	p�s�
��@�&�rAv(���9M&�"�v/T0�|�A�4�g��S���>�.Je7�h��_�p���]�*θYy�k���E�3c���t�|,^������'G����!�4X!1�0�Xi8�����ޗ$����J��]F��-��83�d��e��&���u&4}�湚���Qhp������h+k���XVA�ƒ�$�}}bx��C����Va�q�%[�� ���L1��"\T4�5#��U��'�m��83��i�F��k�t7��*������Z�,m���� A���4'k�$,5?���i�t��[��)u����A��^���bn�G"����?�R�޴��[&R9�V`Cpygb�,�f4�S�m���tώ��Nf�e�\�;ej�!z���+:5���1�zՓc�OU�T�C��z6{(�LG;z��RpO���Br�c��Q��u��9�UK
��b;w����f��h4؛��O�dX5����/�Y�fl�Et:�\�d����ヹM`�����l��B�O�d�s1_�-��zs�+���g�ˤ�U��]�g���3��H�@3��vyC�{r�z3��k�0	�x��Pw��*��o�|�'�;GM�'��˴;C�І��U�܌�zY`�='�Cz�.h���FZ<̭��G�A�syyM�7߼�����T�+���=�Sf耣��������Y�bvO�?�����j>_.//HƓ!��]��t�Ղ���$� �"bFx�˛�7����<,����� H���=v��;��^.�E�A������1.O��|��S�F���B/0��½C���|�iU�y��ڼ~}�+Ȼ��^X1�C�(�29TJk�.�\�V�5�МzFBǩ�����[��}$��m֮)�g�R<����f9�]�{{uVD��q�϶�4g��������)c�J�� e 2�o�o�"8ix�����C&x"t�-�̵XFZ���o}�\�%�۠!��0*�s�UK��Z��ʡ;�w@���G��M��Z�欍��U��)�bp��5ḡK�'��@�K�����m���>�LD&�i=h�aVfGG�`Ї����yA��$�햙�(PO�J]�S1��� g�S�!�y0��\`<c�8�8�^ڄ��z�N�U-�I�:�����PJA3c�j���fn�ȼW��Xn7s��� �����|���W/��v+:�''G���_�w����	��:aZ?�1��<C�'�[�U�
����س�ٴ�8%��H��+��-��Γ:P	���aY�w^V\���:Ӑ�B[��`0��ng�9?�f֜N���x����HC2�N�Iљ�cyHn!c��53�0GVƵ=�L�u�po\ d ��RYF��.�ia��%]�+4o6K��l���ȵ���<ĉ{AI2�I�<һ�R�`��C2%nGN�.5$ᅻ����Q17�6|�J; ����Z�ɰ�B�� p !�x�8'\` ���r`�P��7W9�]A�əv��;'h\�)�4����ﴚ�h& =`]��w:_d�O�N�>}Jq�C��������s��Yy 7-�_|A���ׯ�p��fKv�iXo��l����,r�{�٧��9<Uz��_};��;z���������c��ϟA�җJa�������˗����@t������gϞ}��'��E������2����w�qtE�@^�z�-F@�
�/~�B~��%��R����(��f��l�_]��ӽ��?��������#�����/^��0{��!����C>eY�B)�ߣ�ΓЮ�/X��d0�M�Ȋ\�ι6<��$[�߶���7��e���ݾdZ��"�f�/0b��A�����i���9�L�E����2ʹ&%�ל�]�7��Q�B�Yr�P��)�J��_�f���4#�	,�vI5"�+���<]/�-��x�\�	�@T\� ؜Z	�����2� ��16RE$I�]�e�pr�[�
s͕x8t��J[�!$�m�1�����eߠrV��$��G!��%��z>�0�B*!B'#�&��k�Ȯ懆��lA�f	*�L��L�q��R4 h]�����*s�}�&riM_kM����3��W ld�&�$�L���6:s�I������Δ=��}�iˣ��6S(�\��me܇<�|Y�?�V�,��eq�l�saa���e�x�ǋ�»3�������ɱ��ò���h����F���,���H�EBM屗�H����u�<3�Pt�,���n������>&����ë�r�IC;}rr�p�v�b�G�#  W/�_����%�Č�za�,ŭqR�.rKy�P���[W�@G;uw�8��;m�ɔ�#$	�DJ�y-���(kG[C.�\IT:�*�[�T�o;g�v�ؑ�B����s�%�~H�uʒ�i�g%)�w�9uz6ɐ��XE"���?�F������"�7.�fڑH�)&�jN��H*$ϓ
��@��1��A�4��c��i�]T��"���
4y�6��,~;�T%��G�pޮ�]H=���c�3q��J�`Kt�k���x���i�d�cd���X_RM:�"д1!��g����5	ef�?S��ڈ9�����;�#ǡ`�� �6 ��BƏ.�|5�HB��%9m}�Q۞@ '���^-؁���ߑ�����?�������L����v4��g3dR��&A�K�"��Rf���v���{`��g�^ήz����ķC��i)I|��!����U�V��Y�����r�
l%��Y�;��\(�/�7�b��	��q����H|T�ͪuJ$��?ђ2���#��ܽ8���}�0S�t܁I2��r���~���~�����׌Q�= y�.�ݻwzzJ^�$_���:��&���
w����x<ypp���c48�^�5t��v�ޣ�X��w�.��;rg_ׯ�b����s ��X�3��w&Z���D�˭N���X�@l�^�F*�X�����1}[n]܂�`4�ږh�&(�0�f��lo�@��\˖��<�VV�	.Et�-򪂫e�j]���Tn����9��-�s�x��#=���9���Ӈ��l&�2�3��G��`Ԉ�b(�T�a�q���@X� DÑG�]��,t� Lp�{ud!���SJR$�F+���]D`�ѭ�Ÿ�0`D&]��r�3NaD��`k[%�f-�_X-�n��h¡��EW�;��0�q�rg�)�#��L�mG�s���O~���h4�ٟ��_��_�y}N����=Z����~��_}�{��t���f�n�Y�]�����62�!OF�;P��p���uI���Z֊FN�;�n撙�Y��yqw�e�� �J��b��ٔ'�@�L�WZ@I1ē��Z�.\]�;p.`��9���_����e	���¼�N9��$��Z���ꗷ��z�9lN� �nؓL���E����'���"�:�Yds ��O�i�z^�!ت�:�E����%()n$W:lsq��-Ca�|��m�}�q�d��\~��E%u�l�\2,5u��b�cw
�ku�M�����y
/���ۘ7�w�:�-<{����?�w��ѣG��H|�u�N��ӹ�"d�2��?���K��Wt����7����`~{sC�u{K*΍�ŧ�~�'���?@���{n����Ir�h�^��~x�GG'�\����Qő*.�ԟ��G�899@�ӛ7o�N��1}#�૯�z��9���E����������~�	���s�	�1q�~�ӟ����ObI��,�aH���!�N�"�cm)�Z4�=\F�7��Q�1���I���b(g�-r�H�A�����c���vY|�����;�m�U����7��2�L� ������֎.u!�fЭ%����A;���E�����W�*-��'��݁��>�:�J_��t
��
@C�䇚X8��B���TV	���m�/7�&�Cހ_wѲ��;uF����Ӫl�Q�� <�D�zˬ��d�lPl�iwv\B���j��Z>��3�� ��*:���1�P0V��p���}6A�Q��H��IR�h6W�̊��q�5�>tB�P|Žh7���[�(n ����SA�VI*��d,�ٖ� s��������wK5^�٤�\��B;�̚îd�B�e	`�~�7�y�p�ۇ��R�k���Ri��ݏhw}��w�1x�eqK}��1u�	�f�s�l�|]�iGq�$�芓D�����:��nM��q3�'k��­�\8_2o�S��ˑr>5��O�f����&i�J?h'�XP�Qf��y�x��v�Sj�%��l] 4RA/�+��3�F�LD$҅��#��I?��� ׼��|e�L#1��Z�R�	tP��<I��(�9�J����4�����-~qv�n�\�J9�2��Y���Z)(n+��)�9�$�$���X�(<͘ٱi���|�^�ÑLqƨ]j����Rǽ��<��`��~�	�]�6��qd�XN�u�JP���&Gh$P�J7Z���^��#�#O��ݱ�W��^��
a�`;:�D&�.����o7�;
H� uɐR{��քk �y�Yfy R�Sr��f%R��y��}C��&�1������!q]�$M���,Ƚ ����q���E.��Dv�W��G�������d"��a	�v�Fş�	<�t��u#�}*��dZi^FAS�r�,�wN��>�v��@ǲc�.��ʜh? �'�Mw�ƅp<	T )��N��853�ɲhj�$�����_{oo��9�*=O��{�vo:��a���'�a<W��1�ذIC�-!���2YPUC�!�O�	�����U]��f<�bJ���q�~1�A0�nVMu����4Q�a0���v�]A���r~y~�
���|���kR7�������N���^{�*v=��Ŗ/��Ãٔ�W%v|>��(,
�D���
��=��H��|#F��4���h��h!�1��F\��씟�&�	�Yrwx��1l�h��%(�@r=�'�j��0"*b{�ͥ�T�l}sÃM�`q>�kӴ���!'Ȯ�Y1���E��云���0���h�"	gi�kA�r:�L�-���o{��̢���1g�V�i�h�2&d�d&b�Ơ(���$�"ᳳ���pu�0H��Hg���X�G{3k���+�~-�=�,�l�Զ��:�0l81��4���ˤAy�jG7�Ӣ�g]�P�@�#=rji٧�12������ߧ0���7_|���1G�p�'u
Բ~LZ@��n9�!�d�I���K77�GLxuB?����a�q�Uz�s��b~ra���9؟��I�?��o��������~����廦���?�M�N����/�/
�I0d�yL��0��d(��+�
�C+��V{H�r�d���4�<�;W[�d�'qZɏ�,��[�3s�]Ғi~Ls�C
D�onL��-;/^�����)4G�?tRV�J�����Gt#�pRO��ż)�o���ʕ��t�v��}+2���/v�Zh�>�~u��Cf�/Iz�\�b���]�C||�HYv��!��s��!��/u����+c��X��	�A��'#�3�kۄW^�+�(Xrz��-p'��Y+�i�4,i"��3����̐wX�Zz'StI�4U�-Y��0tڶ�Fzi����s4�-Si˓
P3��y���g�}�=��������=�0I��P�Y�FӵX�MxK��o<�?���o�_.Wn���<��q���������
<"�yxH�B��͋������r�I�8a��M��1L�m���4�8=z@f����cRt�$�Uˤ{�.�o����� A���O>������?��g?��/��/������'9�2����- ��x:���|3'�0������Ç��i�g���]`l9)d���I�ҩ�Q�W�8�7�E/=��M����u�t��>���vОD��b׏b����O�.F�=�3#b1�m}��D��Zb����"M@ܾ�ـl.}.U�n!��G�`�)�(
�h������\$��O\�t:��MI�u%����θ8�@W#Rg0�r�蓥c�I���Y�nZ���&�-���A��W,]�?$���T�p-;�m�q���$��%�d�������+w�o�����'m��hu��\�������7�t�[���y���r9�WP*������%G*Y��.�d3	[�o�6옂7=�Q�~;�[�s:�^�\�e�1�,����+Ա�����mS{a]5��r�ˉd��p��[���9�Q���NsY=�wĶ���i��.߈}���J朚��4�gvY}ڝ�uE�  �ʃO��Y�x]��eK�֥���k�_n�̌��́�?����b�D��b�
���F�ԟx{q�|kL��Ŝ���6�3�r鴔�ȫ3ا��4��<���PQ�LȌ���u������,B�+�j.�XOZ��^{Z%�3o@����j��4�W*yb�]-&%�΅����,�Z���E2�:(���T�V��P��G���E~�LQ]��b�waYH���Q6�����g?��:���b}cHP��?e	�k�5a��#���o����ga��`SSEc�(��*���@�{����5�\gz�J���G�6�<�Ɓ����$Yn�fxI��S�!K�`{�����-��Z�N?v`:��A'���J��-�tVE�ǁDz������Z�`R���9�7[Ӛc����b�P��^5&^5�!���8�;A�e/��戢�&��"���2kt�����,_����N�k;���w��zof������=8���b���9V ìj	�\�sz �d�骰�^�4m���_'���l�X��\���@�}/�ҨSjڜV��@Z��0���3!v�����/Q�A#�2��������H��T恹Ȥ��)P�;�c;���.��W�z���{�S)��;�Dh�B�fr�g�eB`ԝ�����##�������O���'�2v%]��v��u��XڜK8�X1�u��n���_�˓���0��U����B����h�,~��7����/�o*����0�MR;�*�5��D��>XyLd���ĳbV.���K}�L+��<Ӻb��qS�^'/�r5�ST��B�����ϫq��R��{Z��}fܛE@��������X�e�@�`���F�L�e�4>xp�GT�`0�"��K7+)KF����һ4:�y0`�\,�����ʯ�'1�3E���gGesG3��tR'UG��&��R@RĊp'v���2a�ד�ҷ�z�\a'�F����Hyk
Fؑ_�0�.2�39|�sҺ�9�ktVquV@u�U�:Gt�r9�z;J��e��r�'����7�ǿ�{�G�K����ϟ?���_�I|���h"�>}J���_��=:Պ��
�!o��͇q�3Ņ�W(P����(�����Y�0��N^�f��"}�xQ&�DBBn1U�.W��z�4�f	��\��-GN����z%�6��|I2��m�Xz�w^$Ӵ�h50�һ���W��:�j�4)��{��J���`�P@:#�dLG��d�� ,umҊ�+�(�R�U�91�nm�Ж� K�؅�bm
�ZL�6��>�˕�ո��qh	���V�י4�t���.q�4ah�T��ѿ���}�!��]e�2�po)鷃�P6�{�y��N{��uӏTp�l5�l�<{�����˗/Im�{w!��`��������ߧM!ߵ���y�_��|�B�E-�\������{IDQ�`�;��\�qr-0�8�����(sq��_�̡<����^�G���/�E���_��t#���_�[����,A��.��'fA��
�rM���;����$%D����L7�zC,��V�=6�U�H�E�xזVk�IP�!!�##ӟ�A�\صFY����9���K�d"�ѓ��2+oQ�v��J�:��3I����TX�hT!��s��;���胯Cʆ�����DQ����Τ^����X�\2q�`��7�:۲H��I!ɈX��s�=�9m�ux���VF{~#��r)���`e��{�+J�p���"
�@/�X7kzO9�:�qd��:��>���w�7�������Es���o���̖E����`��Y4�8#��Ѹ��`�@ �)�>X�os{�|9���C�F��q�Y���:'�H���#%�8/�QK_���a��d�)^�4�u	
���w;�U�E�"1�پL��Y��j��<b&b��K�6O�zfA,�e�$h����<�fws�a7C"��0��uf��Tq�b�(�0h�<ɐ+�w�"!Pj�c6�\�6C�+���������j�,9�#�LUY���h��F�^.�|�o���4#�%�@` �b���tʣ"�ݿp�� �^�l�����Dx���sM7�l�X�j�!.�L�)�LXM���JH��.����r� �k���q��o(#�L�W�F��d�ȳ�&	��	Iҥt6r/��i|���(��>`�,Cr�2��CU9�a
��ﴼ>�=Ɓ�u��lw���c
�:���èP ����L�s���3���{�=�E3<Aq����g�0�Q��<l��q����Y�=�N�^��AK����`Z�����\�1w;,��Út�̥t������g>d�M����_mx��G�g�ֹ�c�Yr���Æs�:��"�a�̸�e����[
w����4@0���Ztt)�'�h7��&�)� �?��nw�m-|?���ڦ��?�:$��vddh(�e�TE��ӛ|jA�D��ԓ9 T�0ڥ�a/w[�����X�Щ���
��\\\�����w5w�җ��r��ѣG�A∙��{�Ռ������H[�!�H6:�A(9{W�;|���P��)f2����5�a��LꊼKlCI>s�E�N�!��`��N^Fӿ�n�Z����L�gbj��=���al���f{s{u�p;�����7���ˮo�<Lg(HB\��Ԑ�S�$O����Ϟ=0��X0�����]
��M�GxW%�����Y�b߿�py��Ç+�ϟ?'�#��|��*dN�Nr�E�$�9G3N�=z�D*w��mtuuw�^v|����/�����Nr��y_
n��4���ݻw?~����.+Ko�7�'�<u+��Ӄ�P�ˎ>pRճ	�+3g�e2�'O�,�C_rMʣ�9������d
蚏����0��d�áE9�����D0j:�����V�L,���)�����Ļ�����n�$�$7�-{�e5�盪Nl�V+���A�Bbl�ғ|6E�m���F<���d�3f�p�r&��.m����)��'ǀmrtT�����ϘD���s1��=����;>cn�q<v��pG���~ws}��BO�q���ɓG�P�8�M$���)�9ݦ�%O�ѩ������(.�>dLy�0�,���4r>Ik+����̐����٧q��
����[3����Їl2T(E�H ��/�,�fwr�!���4�ң���a���^ Zb��g6����2$�Ϟ=#���枛C�SȔ��ob�o(���կ���1t?���I��\�~���7�?�_|x��"vz�믿~��K����?��?&�� kx4��S��tr�P�x�S>b�k�F=��9�h���r��֯w���e�W����Y����Kђ��-kc��,�ʯ���"*��6��DK,:����\i����Gd诤��~�kq,P���I����������=����b��8� ��a�5h�^����\?"D��Cʯ�	��'3AT��BDw����uHk"�dJ6(��#٥4� �:|�\Rr�D�mFʠ�U@0�|SPꏨ�?������6�}���X��1
8Xv�br�,�p��VX�z�2������)K�HyD(a����1EqX1 �0:���B��K�����%��"�	0�˗/��q��������'���_|�������ܬ8�ӷ��~ýu>�\(F�6��;]E+ވ��:n7LL��6���N�A�gA��{1����������l�ެ��^�z�
Bg����d!']V��-�Q*�3���V�*���W�m8,$r6;f-$]��u����T%a
a�K��!�8y�'KpD�$2h����B�<P�4�G�����#�d��^A�P2� A�y4g�\	�KH���u6�Z'���YN|����YZ&&�T���T*�\zT&z)�ؘc�7IPwb�����v���������kv�Ê��J$'UO��pn�t����灺+J&�u��.��#�\L�vQiMh����A�퐁�ٔq1�D�yL�D*�C��Z0SE�2t�9�ʮ������09�p>�X�����[hZN���s)1��"</���Ώx_d��c;n�K��Jb^^��;T.�����E��N���Rt"��%W��섴��~��#?tm�+?3'��"c2pN�FM�UD����.���yy]�R�!���R���t ~�/���p�����Q�����2���<žԍ������B�V"Od2}�s#d�"�w疉3��F�fѣ�+�=g0D����Lt>�y��Z���^т�z�����h䃹��zݙ ��Dy}�o��Q$
��|��EK�G}�0�UB�A������r��; #��&����v����MJF�]���\�E�{=n�k堒���-ce����,�R �:��i�l�.�)�<�?	���(m�F�7���?����-������:�:�y�a�t�L4iR'A)f�f�W�]��Ϊ�EK���#�H�5�eЖ��d�4��1}�mbɗL+��t���0j��%���~܉��]�a�0ʉ�����*8X��Wo~���.s��V1�����KA,s�%�Á�H'��g��T���AxT��^��Cf3��58��b�1IS�t	��$�y̓� '�Q��wB����š��SK=0o�u�$őt<e���}�X�e�l7j �����A��e�D�+.6���l��U��p�smo�ADVt�r}��N<�4\�U�sY�{���f��'i��J��Vt�NR�U��V��f��TJd'N�[r�NNʺ��n�p�r�F�ea�~G]��(KPPh��X�R���&���`tǼ}�����[�G��zS'�>�ٳg-0���q���������7�:8����[r�1���/^����?~��oA�-6A�
m��:6��'O�\��Jz:�������|���+��9bi����G���ׯ_����X��Ig@�aMp�P�����z"�@�IW�X,��Y��rZч�2O:�,�6	�B�{{V�sќv�@�#��E�%A[Ej�E����	h�������C!i�Rɩ�(����'zm.J����e���[z`� �"��Ag�:%	A;5V�;���Ѡb{GK�v*�f��CG_�^�%�h$��^̗��"�������A� �tH����-��%�$t�<V��<Q	7+̦�� �xyV��	]�����=J�g�~�%��ڐM9��2�����i��uH/��1�̅K'�F��- �` ��jy�3��}���d��Q�z�!�uCA�a����盛�_��_���:�X|f�ш������0�E���9��KFA~|�s�2�C�3W�����..���K&�W#O.;��V L���6�x
����SwC���9��:�C�ī�	Íg,x6�j� ��f:}�ص�U�)�dsl��q��з�2�Eg���a��*ӑt�[$Sp���d�	�i�=�Z�Q��E����z��M_E�`{}xX���BY �ݧa<U�tv4����i��v�I'!(��؍P�XZH�F��&<N�n��cHuʍ�Ůk����e)��k��})Dea��s�\p�c��W`z�T1j���X1����\i[���u|j/�(C��2�����ٍ&�W��=�/�l~��WL�2��`��%r,\���<�M�%�=�� �b�/�bt7���@E!�i�8$��Kkpsf������E�����9�(�Kw��c��w)�(W>���q��-J5uh�^�"yͥf�c�����,|��Ħ�i
���|f�DԀ0�c�Q&�ن3��<�L�x��BT�4!QGӽ��������.ԱG��t}���ӷ8�� �'$�1��Lcyv,4�����M��Cd+0i��퓫�`=|`BE�����e���x�N�a�z�k�Y�hZ�T���:�9=�7廼s���\��h�uͭ�_�\p���t��� ���۶�I�^�:R7.��b%"*��p��\�!Z4Ê��|��K܅���B��Q�c� �[n�ʤ#[��k�Т�c�)�����8��i�
�\t�s�;E��If�<�Bҵ$�N�,>��X���F=�f}�ޣB#��a���gz��
�cdL̰���!v����\�^<����-���lGs8�`�qR%2z��?�Y{���A���3ݑN�#Na|�!�-'���Q4�|��:�>�HB!I �d ���z�j#|D��w8x5<WVN�`tWv��[R���c2��"ƾ�<�llO9�Uh���c���\+{A�-��G��~Ԛ��R�8 ���Ѓ��0��a�b��0��ghU[a�W'�HI�2�*����#~4�{��}�.����ѡk̼j��K;�:��L��&XvG���F��_�Z�`9=Ա�V��	>[�A�tH��mD�$�L�\@�C��@�"��/^�~���_��j�ߑÐ���� 3�\	2Y�nS=���.O�{�c+�"(��� ~kZ�E'â��nߐ�ӬhqD�"r`D0���h�;����	��?4ߑ���*D>e@����cx �tq7)���K�\�Z���J�R-��Pga��f�%v�IQ��\�o�����d�������Q��t!�P2Z��((���$�DNh��?l��ۇ������X�*�َ-,y�m�p�B�跜آ?����vߠ�eNV-��aD�
n���\,f�MS��,+�2+ť�
o$_��!wZJ��s��ʈa1$�>��\ke��`w�i.QN&B�Db����1&t���<���S�M�?�#��(*��|�\HW �"7]�3����K���V<	G@c}��,��i�޾����^Cϗ�����G�O����?\1'� �'+��t��/����������d��矿��Ͼ=�8-�"���6�Z���������Y(�0zq{J�:ٿL(K�v-Y<M�����3���Z�x�]�/Ҫi��G��;F�^��Lumoj�W�GSA�%���LA��2����i�IJ�B��s���#�$�n?~|� ��U\���kPK���|���G��)��EUfJm=�/Vmδ����k
h�-�9St��t^\AATׄ����J�;�~����c��rB7�Z��8�΅Ħ��$wM�����6Ķ��ϫ's<2��vk�;��A������8����guu4�f9��v��= �@�c�ߥ�@��@I>��Q|b��'���|x/æ�A>�$�rOtw�itv$j=���+&�qxa%1�{�g@.LG;$v��FI{e�?XX��V	��h˝R�$>2��:�i)�	ɯ I���J�N�a�������������믿��_]]��;�!G/��qiՃ�I8L=���Vh�(":��zt���$��x�S�n�1��^��0�&)��S����k�	���Qw��6)�tm@F�s/g3���%il�0@�bB�*{ ��|{ޛL��
���	�Gtߜ�(Op��{�Gc�����јy��9��O��4��(<�EBY~��F�Qi�u$IN갘(�A�ǎ�,Ng��@�"�1�$-Jɕ`7j�\�<=b6�2m[i��A�
2m�f�^.���y��Ɣ�(2�n:�(��D���NTf�lT����f�}�a��
+���و��k�*5V�REV�W~!�(��$K,�<�2/+HB��"��`�ZD�kF䩮szz:����2۩�y��k9�>���۴��Y�zr#���'Kڴ�Q&̏��53�|�}1� ��@{- 󹖾�li8��n�ޮ��N#;>��i��ۮ� �&~&;�Մ<�����tB�!�H:j:�!��LQߡ�}RM�?d�WW�B阐�A�x�_7{���B+�F�(��Ԃ�6�>�z6R�4Z3��G��N�0�F.���b��>�}�(�,:C)��eKy��������QlF�8�8K�X ț�9��!�mje�FS�MG�LI�F� �0~�^�'��Z`j%�8E1M��6Az<%C=�yʹ7?j+�Qƺ�B	:��ݚ���m+���3z�;Kf�?Y&ڮ�\bl:�����Ft��mV�t�j������ݔJ\�>D�
�Z���9��WP*�1�?��{�	�����I��Zz.�)�uL�C+S�C�������W�EJrK�Մ�ڢFxYiG=�J�kx�?y���(�fq�L6p#�oN��eˋ�|&��ǲL�	3�a4�˾ݍ��J�QC#�1s�E+�� q���ubP!��'IܧͿ�T&LW�!�4�H4��)�o��t
������g�dj�Ns,Q����n�Ymî0ӱ�l�2�Y����˜6;�v��;rV8'�r�Y���[��I�c�>�	�uX���]L-�8C���~`�Gq�[�$��Tdyf�G�O�h(dP�x���l_7ma(����|�x5�&f�݇U-?b�n_:ܨ���<wj9���Ի3w6R�9��^'�i��qn��"ɔ�*����8Em�,T�8U�+� ;v��aR7��G�T�ƘZW�&��"�j�Q=�T�9�~4 /�8
��+�z�"v�q�y./�c��lw����Z�,�	֧1K�+�XX���"KB�02� F$�R�++4�j�D[�U���ܨHA�S�'*E��K^�!�����n�=��] 6�4 ����*��(Ǯ3���y��O�^�^�+�w�����P�DR�� ��e
�Թ�Zs�!#[�u�Z�:8�]��񒳫�L�ia3�ܐ�C(�ۉ��+�B%E�̀��`������9�o߾���Dtl�Ӳ�%4Z�^�=˕�#h2�יHr/?�~D���y
�p?C,%��ȑ���6���ɓ'ggg�<v����B�%}�5.L��̪e�x���ŀ��L(�t�/��X��)�@Z^\3$o��� ��l����섦K���$5��_��_|��7��p�P��Ŝ�<p��æ_�9C�N�נ굱nB�
�z���eg��J���___�[hł�]�v��q�0
:��i�칢���a~�i<'�#�Q�6D�ե�q:e�gU0��X�R?����6(� �e MXa��AYκ�0�O�{�
\��gTEH��\z�>~��޺gϞA����L�ͻh���0#Y�P��?�h����r��1.st�2s_C�@�e�292�E��-��V��t��б��~�:�#�{hI�o'�6���3�|���O5�j��X@(�S�>������|x;�$�Q>�	2n���"e���wf PT���i��(ul ����R�W#�e�\w	�Ū#�=<�H�P8������_�����򈮊~ ;,����]�?|��JK��9����k���?#�TQ
�G�����h��̉��Gq���g�_����x�Ƈ��vN�mU٩qi�VYjg���L�@�H���t�}B��T�rT\bjdT�w�(hQ:���䜈�x�3��bp�n��q��+9�
�6�i����#;�צP����F=V�E�����!�`)�L:P�c?6W���P\vH�s;@��}��8��fg��6 $���~�ޘ����(@�c=�NEg��~E�t5&�Q�'Y�ln3}���ƺ���e�1�0�#G�ˊ��j�Y�����]����n��a&�\���5h���%�RjK	����#��a�͛$.`�3�6h���<ࡎ�� 
�O#(iw�sw�%�!'��U��1}�R�@��A4�ӣ{?�S: ��S��L�7!��i�
'�J/���#6m��,;p�[����xWY��E�ްQ�]�ʂkFB�$�O�t�%_�	(3�£����pH$�#wN$ʨ��$�������	��z���ĹO�4��<�����'x�،QrH�P��:��I�U�0*�DE�|�)PU�WiR��>i�qF���ǝ�C�a1�W8l��0rp�.&����FRc�����:K��R�\hk��_�3���x=�|o.F$�f�sh
�C>x���EE�'�#+y�dt*�6W΄���a����l��Z���կ�\ ��$/92����/Úc��������3�Ʋ�m���蕆��4ld�y�4�����UxWUMp柫H�̠�r��X`(����=2�Nw�����ט���ii2 �������L��n���#c���èw�i�e~�9��b����S��%H���2瓚Z�&��"-��FղQ�)�ښ��>�^�r!�c�"<�w%�&.�ƍ*[�e������x� }��\RyP�>�<ާ�S1KP���i|��"�}�.�s!���]j�eA..�P����]�uBkO�d�i���"����M����c]�N9��Gux���Æ� l�E�6�z�B��^3k�6غQ�*�Iᇪ�Jyf�6�ryHz:�)�u{;0���hر��q	�Ü;�a�F��j��*�6P������/�{���$!j�,Y�J��Ԩg�ԉ�X7��x%�L�edX�qgzv�s����i .,�`�%�=j��S��ߤ��" u7zg+|=�Ǎ���^2x�}@ջCk��M�C��	ß1�$���Gt98w�u�N���͛7�c�LK"��|qhu\Bxߥ����z:AV"�����A�H'�;��l10��ߜ�J50J(��C�5��պ��P�?z|rz��T��bɢ�e�͞Bt�o�K��]o��K�_)�d~��c�OԟC�
�Fӣ��� ���ie�nooo�͇΅���ofY7���}�\�g''�'*ʕ�M��!y=>����2wL��d���&bF�릙/!�h{�S���Þ��}��5����ڪ���?y����?�lVp�y���'�n�he��C�b����Jx�wb�Bu_I����'C�7m^ &�x{'�Q�_�D�.������%�i�/���lN�$���dy�s&Y�f�7[���Nf��=�yZ%4�8�5-�ыϞ={�<�d`uu}�ݮ$���v$l��>��quwK7!26��I*���=������������`F[.�=�ꆅ��9�K9Y��<�-��x�wdniy��:���<���en�XK�POav)�l�f�@EW`��"XdOf�o+�2�������	(�ݾk�횶q=�'��=*J&�}�ӧ�;�8_3�p�v�\�,����1��TBU�X~�B���ڝD�5�Eo}È�`a"s�ΔU��$�˭i�XL��=ܓ>]v���E�w��f>�s��X�`~��d.��������''�t.� H!�V��䰧�0�U�WE9�)���^��lc\�I�Ҵ	���L�������f�Z�$�dZH�]T�5G�C�{Xw�^H������F�+�U�u*�F�]�il�t�,�
EA�Eӊc��p���Ydv)p�&Ì5��t�f���	`M�KF5�=�?�L*KF�����ݏ�����ڦ�x�T����������~��_��
S����5?��#�v,L�)S0>��*5��و�!z�=�'���#ސmMp �z��9�"4�O2�GT7#�$�"Sj�.�1Gh�4!8v��'�f>r[�Kل }�t����e����g@fw����(J�Cr�fG��II
 �ŵ2#Uk��(2\�mB��R$Nc���}^g̵� wz�$B�}3�L �Nۗ⨺3F�$.�sҁ����1��$ȬP_!#6�H��w�# ���v����u%ְ;md�}�#�u&��\�`y=&�RNm|���p<���E��G� �����a߳�D[�� �~��]��(3p�+��^nω����H�J��իW��G���䤐Q��g���wQ1Kˣ󋲨�!'|z�����5�������)����G`����#��{�ym_���SR�"+��8H�!g���_�����/߾}{}}M� !aV�%��z��Io��`���R7�ܦ?��F �l�1��y%y�+(w
�j|
h/p���3$rI�0��u�ɣس�I�X��O���M'����V���}m1�}>W+���$1�R �Y$���m�Ѱ	���3r���~(�>e+�&ˬ�{PF˄���r�Q��Q.u}�����8��tt��c|
����9�bR�?�;�/��h	���C,9�nl#��
�ǋ�.��h��K.� �k�4mJ�F���C�QQl)-5�T��,"5bW�H}e'�=��o�K���'mp�petݧ��|�O�?[���0���kf�Df�z~�z��X���Ռ������cexw���9,' �ߪ�vG��it�^��a˄3�GÉ�q꥔�8'�K�S��'d�����$D>w�䀣�w�1�6����x��!�w0�E����OyK�Rj�s2z6�I�XO�\,qB���]*a`̀Z�}���(ٝ��Zv1���'�l� Q7b.�d?�#f��8yٸQ����E�SA��B�Q�I[?�����J(��Tp2�h��mk@�I��`�p�R-_Rn��� �]Õ'��f"��LK��<z� �EaA��Q�bȇv���6��vT�8�YΩn�8����)A��*��i2A�%����8��9�ҸZ�)�Ὶ9�at�l��[A�%V~q�4�F��5��ù_��c�||c��G��TH2��������.���3��>^ኃB��]F�$S�4��+������)̈́}�yBvw��.�J�*�&Eh���\�RL��g��-����N��X�]b1�g�]�i�j��Mb⋱������dSS�xc�ʢD���O疯�!��	
$��-��E��r���MW����O�N���!Ĕp��W`z)~#�
���z]JJq��Ok��)� yYXY^%'��QA�-�DF"çX�'؅���Zns;]��~�z�b<�����y�ȋ���t!\�L"�"5��i���WZ�Ɏ��=~�X� �t�)U�'BtQK�Q
��ryyy{{K�z�큤 ia�;6~�)��ˠ��D�N��fe(Dȅ�e(dH�N:���-7� �I�#�q��2taV\%g �"O���bJ7N�I�~~�D�9�&�Z7���v�eѲ�����3�p��y����[<������mw�|��V�t�P�r�������;��ZN��!�N��@>ҵ=y�䫯��NS����H��O��K~�x�����ի7�m�T��u�'2�^��y�����A�%a�h!�FOG���gJ�P�<ߠ���9N�!Ќ�љZP�WY�-B[S��Ύ������|����S2
N
̦s�(P
ʻ��C�	�ߍpP�(��D`�#���˗��tY'l[4$�� �a�A�������{fȬy!N��ng��3���fXΡ�&���&ű2�Dfϡ.�
٨�w���!��_t����.����w�����ݻw�߿���K9���G�yd&����P����pZ�{N���FU�����2�����@���'��|ύ�fl��4�O�<��X��UR�	�{;��!t��mKc�p
�(���9X��GgP��V����������{�|����ˀ����=Y�W�^�q�r��J�d8���k�hy@5D�Ŏ�G����h�/P�B��E+)	��VM�[�/*�`+i�p ���"J�Kk�`+����3Y�vP�J�`%ϱ߅x_$u8�:���"=L!�`(|҇���Y��1���B�M��!L�߶��2��
M�:��IԄ{��4�@e*�~T���t~��|���I+�^g�����%�|����5��k=�҉2������ڃ�Rͯ�����4�A��ыmWtҴ�L8n|�EH�;�c��vHa.� ��G�6�`�tir���+G�\�1Np�F>�A��D��+}8=d=0\,������<[���~����ZV��������9#�
�ɸ2�x"�HL��^�%%�¼�OI:�K鷷�N@[ta���0t�S�3N��^�sr�]�']q�f�@�����?���yf��t�ɦ��?�ӿ����ĕ����9�ۀ,Im>q#X�j+̛�� f��_�?�p�W�G'��O� �w���nL)"c�R���r��ڸ�m�;�π|���L�E�d�����?ym�n�((����:n�A��-��X�C�,��9�#C�Tʕ	���9	y~`��c�T�E����J[��4��K��[��+��[��\9��kPM��,1ڐ�<�^QT	�!߀j�pԐ)G��P��1q�G�XX�G�]���Q�:o��|��(�����E���T��5�7��?��®������/^�W�\��L�$�y��)�v)���{�j�?wNsn�g@dj�kY�t�U�����F�/�9;	���K�5�=)} ��ô��h@H�B�����GL���=P��,��̞PT�KpQi*Ə5��zE�9�s�R;�����XN�.�+/�]��nQ�
����k�h6j�6i�?0sG�l�=4�S(A���5�jo��h�}��8~������E�A�9-"�-�O0��x��w�ʴV�F�(k]b
� �P���X�P��n�B3��*�%uA�>l�B�ʡm�'u )u"^���g�l�`q��:]� �Ԍa5Yd�yI�#פ� C%�L^�)p��^�z,��Tp�@朠Ͱ2�#S��V��ϔ����;��{t�9Wc���I�9(����H��%�'b9sGL��#z�r4s@�I-|�8>~T����H+'@��,�0��v�A!$cg7�ڷ�{�5OOS���ջQ�^�#��s�������������������?�"��c-3��ޥ3�A5���&�_���<��\Tl�>����HJiBR�<aS�}��3M�g�HT�'�-q�0���M��������)�Ӑ~=W�x�1~��w�?E�[ʹX���lT"[�Z=xˁ���$֒5p2������X���v7'�v�����W�?��������4��.Nώ�/N��v���������ѽ� 9_DB��f~�b����~�ͷ_��^�g��v�$��Lgw�К;�)����zZ n�ٍ.98�L8E�HT����$ntatb���N��K�́B ���"�wL�8�bT���k����bR~�H��wٝ���tB�C�'�;�&�i�]��Wlzq�)�7o_�ӿ�OB��< ����&��Dzss7��H�Z�E�J����V�y��t~$~m�l�v�t=S;1�T�{�)��P���oڝ�M.EM��М�.)2��tV���on��P��G�0i������D?�*47��դ��
QH �4�����w��`�� ����!��Ppr�X��$�����_�9F�蒀���T�Y��y��Q#0N� iЃ�Cj�T"a & (!�~�m���ն*���ٳ�������G<�o>u:ר钞��0=?&�˴�	���ٳg�#~�X2�q�����	\'�ݬ21�g���r�L��m�y�%�����h���C�_�f�I^�f��C���lz�����ђbl^�u(�j�$�C�n$�;���.}���3L�P����%x�@e>��62F�N�t��6��6u�Ify�Gx@�+'T���ĔAE�Q$ۍ�>x�H}f:�6©��uxŚa(�(���?��Y� ���,�+N�����z� �*�Z����y���N� �٧�9\�u\ˬ�}9������ۗ��ct�}�2Qg�ڿ~�ʄy��6 �I�~:��!�/,+Oa��6������4�uF�ƴN�4
��k��0l}9bհ,��XosT�5��a�y�A�����y@��9���c�$�f�[!�[��]�p������d|e}d s��2�iu� �m^�%tLT�����G��k�e�ln^v��/sJm=�N`6�*@t��v:��.�5�B'� ��t��ɔ���F 
zx�6f�;�s�xP*	�-8c�4 �����F�?��H�Y�_Z-j~�U�m�D�@��+�4(��+l*���/��h��yC@��QO�y���L(꨼"�A;���e��rO���銘�*O6?���G��뫫���z!���n���L����ݤfjYY� ���N�������������𞮍�h�������<9Y��Sw}�d@�IҚ�W���X�������N������Ls|\Mj:�>e� �/���o1�����8����&R��S���'h�z��k,u!u�K�ǖ�h����'Oap�:�)ץ� L#��u�O�>R�^�\�"}"�\��H�t��ɛާ�2j��EZ܁};:�!*�g&99^���m�do,���kJ�֙-�O$G�u��Ցs-�C����f��.����+6dI4We��h�"��,XۧQ�Q3��F�${�%�>�)a(��i���P��!��8VX�x��ʁ.Ŷ�a�U=�3mt:\4��ŶH\����m`��ؤ���G��f���$~|ꥺ����iɓ��ܐS��(~i��P��^�Aq~�]f�\�fY��jD��C���(��l����S��T�g�àFq����ǜ���'��ŭ��5��8(V&A��j�S�;q0T{���d�Ұ)wH�$k����d���,KVDM���_���,;ț�s ��!z%�0�cvD�����F�@;G�2����`)Bs���
K������ǆ�_��XK�h>DΝ������
�ۉ��`F��G~q�,ˀ٧��J����t1�~�0�ή7;���E?�6"Ɉ��Cvv����N��l6*���F���:��v����� eJ8Ǌ��������e1*�,jU~HW#%J��靘jiP�K��'.\CI��5A�@�YJKUX�j�a�,�-7:([d�H�N�C�.�q�O8�2E��^�	��"��1���U	�'3C��ԺOUֈ������L��,�k�\gD�v�T���_�i*ra-di s�8�Lm>��>MV�Sxܛ�f��d�^������7�|��`����W��2�oz90�\=70��	�M� �ҕv��[�f�\�J��\�������A�=���뷌`�� mt�R	~+�-"����زH��qrrr���������P|SY,�k뱩�J�� �I�\LR�+J9W��A�ȤI���s�M���߾�������://�e�KO;H�|p�t�4����X}���{��1EW,�N��z�f'�I�Da�$�tyts�wQ3����M'� (�&�+$����/�|��3�e�m�	��">P1#���	m���O�1�9w��t����3#��9j��������5�:P��@��"#gD���gh�r��:Ǡ�"���H)�0�Qxr̮-	\�N�1�}B�31 ��ѩ<;��R�����mX����2����L'K�ɹ��9gX��޳g�Z)޷�.%Ģ�Ώfpp�R��ŋ�LC��S�x6��L/��X%�X�n�����������Ѓ2�X�	�܍��ƹ;���cL�~f���q�\D:�LҚ�>��/���y���0���AkH�=y����S6�^( ���U���)��-o�r\�b�$�@w��g��d/�	`��a���6�y�eЅ������ O���]vz8��aJq4P�N��`��+6O�a����v1/<;y�P F�/�ac�Xf����"�{�Jw'w���-]�氿���Q/|��La󁡓�	��ڎ���JQF�Փ�x�Ȥ�%ߺ3U��!�~�^�亩!K-���F�,^�i�gd"9�v'�����耼{��k>�^O��W�V���>łÚ��*��iQ�J:�) h�.�W`�&�������y�)�#�J��ώq���n����n�Ie�O���\�	ࢗ3J��� 几�p%Hz�\���b�%�^�:r!��%�-Z*�x子�|���-��Jn�+#�'P��������ȧ����h�7�f�_[%H#��sT����%$��Y�	Z(��GAǧڻ�f��J��]�(u� ��%��N��ɉ5�%�/�bZ��A7b�.�?7����-C����*џE��+!A�g���Fuq˒��
E�� MBF����c>8�
��0�+W���T��HA��)����9�>����ǀ�/[ ��lqh�d �����@Έ�~Й��"����򬞻d�P@�^���Q�J�)T�|dfu� ��%�CM?W�W����dF��o?~L6��������i>| �}��#��^oe�����Ǐ����5��3����+0�����Onn޼yC/�'���%��?�C�М������|�^sm2������S��䄷���9=s*�@�p��6�tm��l��P`ZWnhQu���u�OuZ���)"�2�*2��"���'�: �,B�Aj�����#6�`�fG]V��'W|4�Y9
4x%�Ҝ`�Ix5N)�Rv�'�D�4/�Kh0'�-��?|��H���N��t����3@���b�� ��ǅ�L�uT^B��p"z�*ɝU5�J���7$��!f��^�S_#Zp�E�j1ӏ/���#�M�(\�\��љ[Kg�L�d����T��k���-��_s:Dk����.�������Vf& x�S�ʪD���Vfp���ϑu�6�[fyJD�n����y�]�����%5%r�<��u���Шe���7�o��i3�&��&,5�����Bg��G��e��&|:��@�0q�8�Й��C�ɻ�(=e�n@ri|���#lBn��\��NۥǷ��H5��ٝ��$�!��Ә�5l��2�{�2�XvE?�0���L�=;*MA�����L*Ȫ���:�ݐ��&m��O��;~�cYd3�6w�v=����¯#ga␑���!��mi�0��'���!���O�p��Q�ܳ'g�Œ�Ʉ�.��5�1�\�n�I#p^;K";��B|��wy�KŁ�=�1$��;�܊�\(B?�TY_���nJ�d��H���H�ᄤ��| � In���TN��M+Rjn>I�4(��� #_��Iַ�A�:��O����.�r>�lZ�=�ٛ^LyP)�zv�w�n�KQ���lF�1g��dF�(�M���/thW�2���	����јCW���ʅg���+s:�2C�BEB�rɫ�O'�l:e�wiN��|����:��Ӧ�'0j�*�v���H�":Eҗ>��L遼�L��- 0�vNK[=����
�/��^ms�x�]Ҽ��D�����V�韀-c^0��:>�(=[H�� u{��R��h!)Yz�Rf�s�*�	�I�7.,���v����@(+��6�c1>D���k��[��L{O�s��n�+�?u~�v��S����9���A��t�#���R����Id@.OI#熄����+�}<??_�7{�:̳��&$O���3��X>}�f�>dztB�����7�ޕ��k4��n���{�|^��8��ђ�z��q���6�|	]��b��x�J�@�I[BW���{�4�UYM�`��2�)�_:�<>��}︸�%j�q�L����B��;Z�.�����L�|zΈ�LiRf��>��n j��-f%�F�j&Z�]���擲����$�}�_<>���伂��2�8>���=!�bO��-O�.�m�y�8z�;:i�#ϞA��mv��2did]G�=Y���I}>Ė���'�����E��g�җ����Vx��Is����CR�m��v(��.�!�����]<�9,
��͡��y��~FW]��=]�l69;;^��fuss��=��>y���Ͽ )-��½�Y��w���K�WO�Ɍv��ggg�M�ż��GG�d���r�b����ّ,�^��-q�D��)��Ѣ��Fje|r�7�ȵ�|"P��vz4/ʚ���]w}�ݥ��`CS���l1i���y7�I>!c��-鎞���9��j�ow�]��|���
5]�o�W���h$�WW��Ͷ]�6�<O\��2����k	Vw���9j�)�hyR1)C����w�{�+�$���dB�eA�?��/���a��_�>~\�>X���0E�|ytv�"��S��d��[qj�~婄�h|��n82���E�,<>�U��<��%�4%��:AN�����~x�m�ͦo�m�8&�n��}��UJ=��������e�t�	�G�<y=xr�;��bz|~BB.9&W����Ǜ�ۇ�n�o��j������A&���9�3ߓ̴o��>�kȹ�<l���3S:���N)!kFW�\ϧ3ɪt���zwO����Vv�I���~6�a[�v �R��.��/i1d�CF�}!�~���-l�����r����gS��64E�����7����秛��ϧ<yf1ߵW=C��,r���t��7�ѓG���{�k�fG�ƞҼ��ɾ��kN�<�Pv}������*��,�O�B�d�h��������/��7d���9�-�{Wʙ` !��:y)�˃�.'�Y�dAKP�x���t����],��<�o��]���O��$��~��J�^�]?B?m�T����� �ytO��O�C>9Y/|�d.���16Ӡ|�92=�W���=�=�S=�f�*���q��4V,�J��#		(ٺ�6Ut�:�YQ���zp^{/���A|¶)�p���PrUȇ`Gn��g��k)�.��^�O�`��뻬�B2Ǆ�N�c�8�e�p�4ol�*U�	��F�$����\�
&b����3�\ld���0�a�Ŝ�2}5�w�Ǝ�	���G�:@�9�1�����a>_ �&���̻�c���iy�_O�s�=(�	HPbS���lp8�A�2<�+�?L�_�OȂ�����sP���8myq&�YQ�����뇕䠹)�ܕ�z�&MKW�bFw�ChZ�O�����|�.�)��j9�I)d�ȹ����Dy�[]�M蛽�s7�����=��<�f2/o�y��b1?99��9w���𬺽��{�@���H�����=	�n�Z.ȓ��)������W_}�I(�?%��*.߽~��3/�V�1.߿)J�ٽ}�����K�(�#q�Sn�%�G[�rׅ�|�ݶ��O���D�~�f}O�L:�����g����a_��"i������cU9��e�����QR4J�+NC�jȐ�3ø�
�CBǇ˞����������3�t Iog�u�Y�3\II	�\�u@L�����ؓfFr�����R�`S��4
љ\�?��^8��L�M���'X2K�F�"�h�����$�ɤ[<���L��f��!N�x("�y�n߲L,�a)I�ǅ'�l�u�S�a�I��Z���T2v�I�E���J+�G�W�<J�8�*��i[k�lCDN�̻�T&�1��^�(_%Ӻ��%3H;Q@k����`�F[�D��$�A`�|:8�(ļ\)��r�_o�M�N������.�GpD�I�X���l<�~�}���P��%Ezrn��%N�0��zʊw:-��eBHQ�8d�f��$��{+L�G|��pC&�R���٪�ْ
j-Mf����׍�/f�S����'&A�G5]L/9D:HR�K��V]Mzn��4R9!�^Ԝ�#3B�[�d�k�o����h�2q L}G��
-�	2M
� ��28&�g���̖ƩȘS&�x��ǝ���_7@�ib�K7��C˔�P;�p�7��^�V�*�{����Tu`� ʼ*�'ػ���������cI���}�CԱ]Y����&	��6�5wGyT����;\ZԚ<�<� �H.��2&��^�k>���ؗA��.$�Ӗ߱��j�ߞ ��vR���`C]ezޮPZ\��vJ&XV4����J_E����gu%���$-"��]��'X�ej�'^2�&**8u�Aj��і�E=���^f�K׀�����ܭ���*�T%#|��G�E��c�\f�pA����48]��g���r�Ҕ�.Ern�j��|�:N�T0����Q����j:MC�P�f���U&c3�g�7ʦˍBP7��0h����S+G��,�VxP���CV[4�`.xPD$^������L�T;bÓͬ"AkH�|��wϟ?���M/~��)������4qĠ����jm���}ɥe��u2�"ġ�q��ނ��_�����'S�NVل4�I#�X��U���x��$�J�v=e%z�����t�L��Ӡ�\a�����gP�m��֡�x��-��������h���'�(x[
�v���J�D"|n�tm%��Q��(	"�B���\�9�fDrU��׷מ˛s;�t�?��#��BFp��>F1g��h��j�آ���'�ѕ���
CT�� +d�<���Jc
cCwz�����ο��k�B�.�?D"� V`��i��U��c�~!�)�9B��mPF*s�-� \�lC|@�4rf���Q�Rv�H��A��¯�e��TE��
�b�kV����ݿ�?�����ƐpO�rZ��hеaq(6ȋo�_�p�D�"1����W�O�d�Ealt�<�(� s�����(��
��;CW�tm`Z̏��+V.�g�{)���[8@��B�gZ�P����2�/�t���o�e�u��	��Z�!��߀%�ؖ�~^\\@��ɂw�7�d��:K#�+$����'��pG��§ѩ�,���w+�<8β��M4C�d��끻��������Ӈ�����c�˞���	}���-�swO�b˰�������i�Z��v��3���\̘l���Z��:����T����x�Vk����]��
h�M���o�wް�?��jAF�Vr�l�t�.0St(�NNy���'�+���l"CJ�5�'�9��e"j5xAClӌfx"	��x.��t:P���
�C�τׯ_O�K���}�9پ�"�V�<3�>��{����"�h��v��N4\���Ü�ld
c6�$�"d)�Ϲ��k�gB��E-h����K�[XZd�3���p[k(6���<�ҝ�"75�@�B�a4K���889�1j'��\'_9���QO���σ�╟&��P��2 �s
u�EK��Mg���ãSF]sr�W܅EG��e:��]?�E�71��ڧbjv6׮��v=�@`�k+fn�oHS&�ES�A�0g(��+��K��7���T���N��ý���1��f�A���,����cŊ"��,a����;�9�it�HI�	��(qD_=��K2V�R��V Z�Q�@ͫ�jb <��2G���[L�C'��(�ݙ��>\����qǌ�N�͎="���`ì�;��U��3O1�ܢbIp.��@?OϞ�3���^C i	�Ԧ�n�Lv<�r����]3)�?��p#)����_@�����(��!�����m�����ej|+/�ğd���`Ϯc��K�
�a�ݙ�Q|BYb�;��M��U;0 ��	����I:� M�r��N&��s(�\=��_b��]�X��6��mY�U��T��\�����-��$~m _R���;�;J�6hj?�#�PE��ˈ��%5����D�����,N\��C�2�| �5��,h���d�ϩ��ݶA�E�u#��MQ�.pG�d�F\��s�$�_�� ����Y��Ð��)(Sj.��q �Kr�A4���؈yr�E���,��#��7Z��`��(��~>I`�s�qy"��U��08:K�����񡓾�W�;$b�
ņG!p���*�.�A����'�.�k۸HݡE�*^��e�˔!��#^��YL�+	o����cb)|��tx��n��)�I5���D�R��Z��|l\`�]�(��.Z����묕�-�F��I�y2����8=�F�Ǳ�����T'�[�Ю?�t�F��俈�;��ӥa�>ͼfyr��dzc��r���\*]5y����ًg���e1�E>����=E5%���Ky� m`6�Z'R ���#�C��YQ�p��2�t��T�D���BV���	|/."1R���/s~���p_,��?�bq�7W����f/_؋g'��"k
�3浭�x<�
F�ߞ��.��ً�9q�z�>k�;ڭ�Ld�f�C
-׋/�`S|�%�W>�z�FHT�_m�M��]͵��Ja�'2��.�q�F�ޝ2��EھD�1>Z��f�29m�(�v�_��_~��Г	�A5��n���{Z�����g�Ua�O���F{�1QtYj���u��3)e?R��vGv���'qN��ތ�����g��+OŚ�|�hϵx&�r��Mӵ�bڦ�������jʶ�N�2�m�E:m�I���P�)����{
��\)��}�����W��jvvv����v-�5!&�?B�!;�50�i*�S%�FV�"S���޼�$�1��x$��uY-G�GK�Ä"!+�Q�4p�m+�@��������ڐ�����\-kHÐ�4B ���!��x:*$����KaE/���n���'n���#L���)�E��Z?�<�H^��N�l2�O��N޿糸d�����b1C�;O���Y����D/%L�*��)M�+����.e+|1�̋�b(���'���)O���~F7%���뢮�ه������۷ﬥ�nv:a��K���sG����������Ǭ9��\�D����o|�_|�b��nWդ�f���Ǐ��uߴ�V2����(L�&��6�;���������Ų*'t�<A�i{A!�ye�p��EA�sye�]��_,�F��puu��}x���f>[����a+.�z����%}�dF���7?�#ZnNd��er��j����<Ժ"kX3��,�ya�ŝ��y��w�p�2�z/o��dtx>��x|�x�{���u�3hu�M���x�a���+BҦ���ƙCO�q{{����͎Qx�vɯ$�G�y^�;c=�Et�vBm� �,Uˠ�h��]��;Ɋr�����f������B�{YOx5����Q�@"6�a��m���G�j�Қ� Fb�� ��lI�����A�Av:K%YK�gK/�xÌ�<�[`t=t����w7�&)�"#!�	*�N�ϝ�L��W9M�%�[.�,�QIy� s]8�K��b_�BaCL�P/��m��$z���-�벀+��B�n�v������v��&sRU{'����б
�Et�9�Bvܤ�!<p��NUd}Nw��3��p�����V����������w5�`�p���Im˼���̷;
������X����Q�S�ցq�܉����v#m,^f�
z�B6=� r��a��R	:��)Z���:R?Ɓ5�դ������F���h!G����y����9�.e�<RI�)2u/�2�}���b���6�ʿv�����O'f`)Ɨ픷]��3�y�Xb�Xn"j61S{# 	i"�Ä���3�c:,9��B�c�3`��m-���%�'�05B��<�0�Y�U�0C�K�S��lP;��m�~!E��ǥ�țh�Ct:����xqq!�sk�ѐ��}��ۚ�@2E}v	[&��"��p��	r��@Δ�N���$|pk���u��1=S�41��L��I%����a��r�������g����\��q�7Y?����36���s27�:�%��|����� @!�cޭ 9�\�"��!m����C
������5�����_�2z��~/�0����2U`KL$�/�û�mќ�s�c�UM����`�3��O5���*�FD�b���I	���ڿ� ��J�ڢ�s{w�c^)կI2�]��*�tܹ[�'�r&�>V�b�a4E]C�h��6e6�4��k�Õ5Uc����	-8C,f�v��C	��(�������D����*N�Xz�Q������8ܐJ0�8ˢ��e�:�{o
B�q���^��ᤗ�(HG  )Bn��B��Ñ5��#||t�q_E[���.�рhFFӐl����b�� ���I�&>޵�aYN�>Ȳ���S�g��Ld1]3	�-8L�:������b`��,]HQ�UQِ�D�P @�f���w���(� �#�eܾ�>䐻��0b̓��L��qs�X����8Ib�a�udZ�sR�*��7� �\iOr���Ē	�V^P��ٗ�ͳ0bT��>���Y��Q�ڤ+퇚"�F�9������j���D��p#�dRZ��+�%��7��pմ�����N�#q���Gt��ˈ1�V9�t��J99aE߶L2�R��XZ�wPxDn޶�w�F��a*�4נ���P胮�r�H[��^0����t��:k�[�$h%�����	 �+�)1�x�+(У%�.�L��%�ԝ�@͏�57��gO��X�,͖6�ʒJO�<���V��j�ۭ2�+���h����a�ς�ʵ(��j�4�/�O�u�Ϡ���Ҽv����}As�ci6g�Sv�G��EL��xQ,�N��ݠ����>	h�i���YPa�E�u�\ii�F� �~~Dm�+{?$nݠ�)}B�;��_u�ͻ�WG�5Xy_{�D
����t�����=�;�;�i�M ���������
�7�k���tڒ����vvv~qL@�����p���x��"S&J&bϻyuu���[�i�ۂx��hV�eS5�^�����0�q���+�����a�X�)����+�$�A�BG"�ʼ)q����1*j��z�av!q*�/�1�I��Zф��$�����d���g��d��{ta�GțT��G�\��FSDYcp3�J	�*�����	���&�p9���G��0���i�*Hu����ŷ�[��(n4.+����䈥���_��a'�"D�,K1!DЈ-i�t�$uta90f��.��3{�z��.݈��Ag��OV�z������Z�́G�9I��Z����}f9w�������{�⮊;�y�A;EҾ�^�I�e�K?X���b�$�SH�gx<���#�-N�]Í��XE�m6���l�0�]T��`�_�c��Ē6H�u+:M�a�����y�}�\v��j�fa[�s���^|�����;I/l
��E���-�.��͠=(h3Jr�3� �hh �JxQ=�h���� �xw��şNHm�0Zg>e/�Z�@9I�'ʡ,�9BX��;@�Ak���I&�d:�
oD������^� �G��Aj_m)��XO��t
`򂿱�p~�蘿e�Ҕ��}'���ð�]�,���j�>麡=44 ��5;����_�'�z�h�Z@ӌS���e�F�Z^(Rk�<]��N8ܛ(R�������`����U&rs��q� �+=#z��pF�cN��l�4���i�\Q@|[T`�*$����e#��M3�����Ӡ���dg�������!�'��/5f\k�M����O(l��{8��a,�����(|��O���X�=�6?��F��,���2�8(>�ɆmY��ѡK1!*L ʟn��0LK|� ]An�*��˱F�ÄB� �:����bԋ`j'C�F;d��\9�*�����)�!Rr���>�+^f��:ȍ��`����6��ڰB��w�#A�L��G�c���f�D�Byɺ��4���_8]�Z�
t<��\&fD)�b����Pr۷{�"Q,�?����~���}$E��͛����9�
I���
4���R��fSΣ]ߑ��ӟ�ŋ/���Aw������������R��!˧P����� ��GQI�� !��uz19��ԙ�������/��W,�R \'������6?��������]��I7xw{�L�CM]HyR�TY:����g�<f�3�we�[%��A	I�A'v��C�ܵX75���8�5_��7|i�;�ƨ%xI�Jhp�8��=��~ �d�1�Z��t�p�$t�	�u:@��&�g�f���	�	J���E�l��ܨ�|4g�Ićpf�+�Z�h�DP����]�H�B��L���+�C��K�3-��m �t_Em��kH`=���.��X���@a���(,�4��r�wa���F�e�;$�
e��d�0��B/-�z��%\��>���?��0�	������������.//��Qp&��;X`IVQ���u=�$��v~������Q�Ru���
�2�J,s��\�Ǥ�hm9��м�l�P��a��A��(/a��=
��
	�.73a�4W�J�c�5�>,�!���6�q������ᚽR���5'O�$�F�Ʉ(Ӛ��_Ʒl^�<�e�'��#6t�e$3gċ����P	�O���ܽ�D�N�j	�Z��=�*W�&5.i"�g���h���Y{�&ɒ�\,⬹��]��` �h���kF<H��L�O�5��f�(�  f�^��֬��q���<���fJk4j�3O�����w�t��m5���~ \������߮.]�%�{%�Puu���n��>;�<��eM���#�ȱ���W�gNKd�<��<�bB�!˛������xN��r�A��0�$��d�-	w�ߑ��!f��:��v�TKHyy���hf���ƪ�}���Gm^�YUV�ݼ}'�f���r�n������A}Ó�fU�C�ߑ�NV5R	����EO*���8A�Z�m�#�3���Lq���\T��鹚~���Q���fL�;������[h���T�b�8�İO��
r��u�өP���]'�+y�������}��pp�8T�"-,�	"���L"�4�YB�d��t`k�v��%�{1���d�1���#�Ozdd=*8���2	��V������f����J?_��s��fΗ��^c��Di+�0 Q(S#J�p�ϸ��!=�3����2����5��r�m�q��h����!O��gQ?�ϋ�����y��bj��ryVW3��0��}����o��L>}��M�>�R�΃���k�۷�0���܉X��L��1���bvh�)
�7�H��������vC��"I���k�Vw�pu���z�$��j5g�T0<<�-Z��\�M�ɣz�/.�f���
z��m�ti� ����֎����qG�@�����+�������>/�zY�O��4����; MS=svqHY��?>lo�^����kiC+x��lA���vw�m�q�{�l޽c�B>����6����@������n���2p�����A�)9D:�D�n��򫗤0k&)g�������I	}Y�Ø�u�4�SGq��p�I�e>�K>l<��Qx�����~r�>�����B�u.!��m�oxB��[�����x���Z��xQ�毷L�CZ�����r�X��L���|1+�w'0�g���tѴ�g�R��9�������Qt|��\�ͪ!v�PU9_-Y�������N8e�c4+��xz���In��6[z���A��L7�фZ����g2�V�,�g�<3���B
�C;��]�eۆ��};֋���x+��%q�lAA���}V�](�ω���,ߗ݃��	�����P�¥H?S�	&�Q o"䌎g^s������4���� tE��jc��K��H��H���٣��O*a�&��K����N�(��A�en�2��Vf��f�K�����&	�l2n�!�0R���p��(J�9��:*����ЍY�s�ϫ��g�2�����l1cꗶ��Ŝ<�V�s[_3 h�0��o��\�?�Og9��1ǟ$R�m��C��_ �AR�n��t%���謚7Y�ʋEY�H)���[|l�
����Ԡ�K̬��,hAv� v�9}Xz8 �N8�S�)4J���7��C����Uk|�y�Ӣ�eý��Ԍ2��(�.u�!v�W����א���A�>��*9N1���;�
G��S&�В����v.�Q���w1�,K�L��PK� J���_)�tKd"�d��4 �t6�ך�����Ss�ӄ#8հ�:�em~��J��
�V��3�Sa��l�V�QD��l��0(D�����d.)��������_�������.G��|EZ�i\d%%|*N@+��a�G���J}�S�{�\x$>����Ġ$����m�P&rl��x:�'�V�*{�MP
�F�*���$�g�}c�(�����3���������y@"����O~���/�g:����������9TLH��U`�uf�[G�Y�9�Pe�Lٝ�f?����\��\<�����״J���o��Ɇ�g^J����������~ n������=���@D-�$�H��2��?��W�|�g�gϞ=#�jv'G��N�����KZ������D�|���ׯ��_�xA�*G�Rݿ���:CG��G�8"�E>���Y�b/w���l��vodf�9�-/ߏ�G�)|pl>�#�Mh�A� p!�;���1��;J�+֮Q����2"��
��ظc�#�X@ز�������o-F>)�-�C�QrF`Å���1�[6��|�4��<0(�z��65N>	�{\p|�8�\�,KI����}fh\]tb�QSKQ���sy��P«(Uj�s��;��)��;��n���`����$f?��t.�^_s�R<1���
/�b�)v��P�¼`"3o�^���j��$aD�����闿�կ����>���-�N�!=$$UAf`\���,��~*��z�4�OЄ�SY]���'>���G�4����t�D�45�,n�m�Z�r��=gs{C�eI@�� ?�a��Rf����dn����=&�X�QY�F�j�#`O4-PA�I��P�����`�E5�+S/��`��3$�{ 4����Q��*�C�
�m�-� �l���VTZ��	9�1�7+Yk�.u hfw�B&�Ʋ���^T	�b�}�TJ�g���ӧO���Ou}�I��?KF��d�6+�Iu�60���N�A��K����a32����F�~gf D
k�)�?SR�B��&�&4��g~�_ `�n5g8��b���'�G+�������.*���狷���n��K�F*��p�����z�
�\){�ͱ���nr��Lm˰��a�,ˎ�J'$5Մ0Oc�G�S7�cpP�0ˌ��`���.� rV���JD�n��Uy��hM�<�@f �%d��j�T�w��VZq�@djs��6]@Z�t����%b2�\�˙�Ѵl������E�f�� 3�g��Qx3r� �B�qT��U`�q����!�M�×_~�r�^|�D/�r%~�e霪@.6F�޾}��W_}��7 �Rꤨ$���s�-碒�"���<��7�p#�m�a�P��˶"Y���$2G}BNt�@ڗ��0�~@���JcbHo�-b�Y�þ��ob����Tp}2�!�B�gN��0N�����P�I�B���Ѿ��� Oü����׿�{m�&�kO�#lw�S_j�<��a߾y�fu�'}�,���Yk�/)�͡�x��Q*o��KZ&��}�I�	����s �]K��� %���8C߻^��h��Q�����>�yw��?���_CO:��1v�=>A��������Щ���,1���p�\��NQ�F(^�Jq�(���@���>���E���tF�5;��r	���dQ+��4ՇvK�,&It�G�(T�Wr��ضC+���d`���&�j�*�I`n���J���<q�|{K�������5`B��pbP���ŕ���O
4�Ch-XE͉J���ρ͡w����X�$t�'��p��pG�'��xD����n���++|� �N���H�q�Wŉ6/3jϋә���<z���a��� �_���n�-}���X��%�N�U��0�7����%t�ѳ��|W�!E���(��c�`� �ܰ�&TZ�q�m#(o�<a;�UA�h�A�4�,���@뽒QZb{h��Vn�7'm��I.��u: ��s0�����}�\�el��ތ:��б��d�s�Ve�uk�wD����,�x��;��1a�-h1�Ҍ9�R�:��ً8V��Y�>O���Ph\�n�bxv���)�d`�a�ݤ�	�A��o����gI��%�DA����(���@C�u8)���l#{�-��;������s�npq�X�oP ��>����&0�����u�	MuDm��B�4:�G���%�o�p�,7��by�l�ޒ����s���:��G?J��ܛ����|�J�;I�Iɘ�,����.޵۫+��̮��9�u��g��=��� Ec2[��޲&ִ�V������\����'�|B�)����S���o_*W8�ͷ�-t�w���	.!*�%R�ظ^���X�V^\|r�-�>����Ӎ���ۿ��������O��OK�a���D�?�=L��g(��zc�t�^�l0�R�M�1[s���R���Ng{�"��^���䙤��/�S�L�#��� �&2�
KL��1�0E;f�,u�O8��K��s��H����_S�����K�>m�t��(�r���d��1j�%��U���r���0|ʹZ^^ �Gs��&%��qe��TfSG���ʝ�P��Y�\n\:w������n��MXu�3�6�3��OgXg =�2g#��]�ւ�����S2�u}�d�_��_\^^�i�0_�oA?c�{�D�~a����qn�������F����/Pa�.�T[�HL#x3�^�s�	/�c��X[2a��E��岉_����&���i�Ϲc����3���>��-���yɴ��B�����V-G�τd����kb�h�&qA�H|7��#6ө}��V�%�/��1q�J!$h������m�M��|��b�3�q|?�Ӄ�eeAǽ-���OP����'�����)y�k{���Y��L��+OjTxǇ�����³ B��M�X�,H dx��q0�b�8c�#��d=I��0%8(�rg8��|��O�%�u�O�˒��u8�x���ο|��w����g�s�RG6�8����~RI�lN��-�wA�c�r%��f�-�==�٤��i����ԋʋ�j8~���S��x���!+��T<,�Q��AMp�g!�Kzrrb`u��Y�>w4����l��_8n�oiәi.��v��B�٥�8�N[��S�jt4�F����Uvf`�������>I��ЖR!�qX�����u�yY/�gE9�YN�0�~�S��v��ɉ��������c�`5�n�[̷�#_ed��~�y��������ݻ�IՒ>��s�C�H0�>t�8b96�M+�*����uws�p}�@7�W��v�i;lv�(��BB���*<NxVT5O�e�8�b�N�@7wc̞�WԤ�x�K}��Ho���P����WH��qa���5�:jd�IQ���[f������0=��w���fw`�.
�����|���ZO�������n�n�vՌ��j�zג���XBʬ�BH��Yn��f��x�a�9����%��Z����w��.%�y!5��s����<���߳[zh_�z��3�L���_�� �z�d&+�M������j��$��� �F�����k^�h��^ޖ����X���SRͨ�V]�m�����կ~��gϞ}���_�����%���'H�h�J��k
���1?����w�[�o���F��-EBc��>�?:��4�B�D�r��Q�@.�����-��9�����zse���猙uܫ"=P�"��yb���r�����}Ɠ����������$��<<li�Sш�9��6<E|�o7:�`�/i�����':to�������ţ�ϟ׌~���eN�/v[��@Ze,k�B���!��/2:g���_���Y!c빐�Iϋ��4���aK�,�֞�x�#+�L%�<g��kZ�x�]/�6��@����固�Sd��l F�"��ɢl#�k�j����S���#g'��^E��8�6��z�������k����	�'g�$��0���v�aN(1�w�ۓ����w��\߿}���k��u�	j�A�!����3��[J%eEÈ�\N����ޡ�9��O�S���L���`�n��9�����{,H��1R�:-�	-�!��@�t�ĤU���O<i�LF��-E�n�8�VM$w�#�q��q�w�><��=l���)�>�M�MA&D���$���	�BC�L� �x�э��|6�2u����̶�7�?�d�N��wJ����k�2K�����3�Q%	���#���Ō2���#�� QZ<u�
���?fθ��ֆ��
�1��C�!|/2��Ak�0�u���/^��UE-WcH�Af�p(�t�-�d������C<l^���FT����t�d�&~�g!�Qß�'��1x�O�1����o[J�jP��B' L=�0)FZ��3Q�s�$<;!�Dc�n&���)K�m2��4��r�KŏH�/dU���5�S��C�n�aL�Pt�*o�Kk�VvH󅠔��f�b��,Ao�O�OW�N�uǄ�I�R�jZe>�Գ�+W��׎�\�[pz�Z5��ɵ,��/$Ӈ{sH ��ʹy�r�(jb��k�2<)�n}+��n�Xͫ�BJ����K,�䑐����wW���Ϟ^<Z�HK�;���?y�xX���(��t,9�c<�9?��/��JZ�������kɷ�f�VXrGK
��G��l���b�kP8�0��nKA_�:��YC�&�ڛO��g���o���O�Kd��Dj)�Ca�O����=t��WڅǏ.�V\M�������P�l��+�ĜM�A8݂5'o�ښ�A��)�8ݭ��r�-�/���a�&4*u�d�$G�
��yy�ᕒ�0��b����+� D�G�I�{����H�L���t.3IjaPLLT�Ӷ_KT:r3�,����0�8v��Y�/��T��_�Ct����E^y�����P6S?�����ú�ɡ,\BBMx�i�7����t͢H-k�V	��ti��l�PG�r$ih���Æ}esc%�a����y�#K�6��ǒ����5!]���������?��J����������������e��ō�v�CE�*e�Rfǚk����qx��67�y�V+F$4�u��ڣT����+C�W	�a�\R��d��G>@��}8C2v�����fY���G2+�)�h�Ӵ,lwN��jkv3Pڐ�B�mM��qɕN�@?�,��O��^�\^��2f�>ʺ��2���p4v�MX'TXK�$�$�c#(�O
$M���Kv��*y��1J܍�d�ruJ:(�?�s_¦r�D��<��d\/=Ť�`�ZJ�˭B�!��T�u��U
��7����~�-&l���
%7�&w%�� �VW8��F%��RO��N���7@�SD_a���[��4W͸*r~��3&��������e�\�9'm�ʠckҡH�#�ꐋ����ǞyU����̉�6ީhB��	eޙܗ"7�#��M�u��;A
m6S�_c�ԓ5IF	fSkRd�Q�Vd�0�7��G�Ws^��Ç�����<"��}l���v�z�99�Ɏ�v�Ӏ�f§��!l>h�ѵ�F��v l2���:�,M��uBϕ��)�|��%y{�_P�sd0�)^a#��I�~'���(�n�O~:>kF�s�y8�qz��j>�w�+�-���˼ �3f]�M)R����AR$l���+ط���Q���]^^b�/K�K����k#�J�C�c���^ݬ_�z%T�wVE�:�śa�m���P�4W�B�"��|J@G�����f�E�W҄��)�~uuE�����=�Xٱ�V�R��W_�ՐE ��@;s'�W�Fx��n�9x�s�d������A�#aM�T]rS��D1���o��+�{{�\�� q���ق��7�|�/��/77�P�t}�FY��J�8_7E��pΫa,ᓧ�͛��o7;ڝ��}˙�2!�~������9	m8�I[1E��_�%��~8Ht�{aR�GM��A���	���ϣ��vS�$tC�ۧoAӱ!C�f��-��5�[Z�'O��۸�����f�棝q���tE�*��ND��Lc���q�� ��e*Z��Ú��d��BR���/pi�U]3Ҥ��
����� 	��W���^'��yi�dז�b��K����Cw�]��4��́ד�&V�!�hA����ي.�{��6(�� 8���(�JH\�Ɨs�X�y״2�z#�@	Q�
+,���2�E,K���M<8c@�������@�ɻ�}��$bAz?�Dz,Co	��):͒�jV�_*���8*xNBqqvr�ٗ�ge�u��<ij=[�mkI ��Ϟ=����ڊ��w:�����j�C=�}ߡ�DEA�y�޽{��	� �J~dL�`;��i.6������p�a4�AA�f�Ú6~��� D%�T��NMq0"tr�*j�4��G�.� �R�S)G�>DOq��E�A�-�E����j�q�zow�+æ]�3�G���шp��UG7�D���<S$jx��J�%T.���+\ �z@'(i�̛�oeW�>���J:
ޣӶ�a�A�4�u  n�"�~2v�<4Y�Ԋ��)���O 	�#�F���g�������{�j��� ��p��s�im�T�S*�t�+�ۚ�,��y�v��E8�Ѯ+�3NJ�N�/,���r�r���Ui�X�a�=��b��3��!��7#A��� �q���,T��z�K\3�����X�����*F� ~..��.��q.��#J�h�p�e�K!	�)�L�7�0N�Q��x=k�h�j+�}�T�|�{�@�Q}�t-�<@��4���W�I�9��e�_|��g�1��$�p�@v�,sI�`��߇���:p�gg�:���
}���
"�0@ a���`	z��X�h���q5���̫�&h_�z�u�B���C�Z-M���z�q�#6N ΐI�� 7�yf���G����)'�tYL���?̏O�o$�pW�T.�
�d�ZN��iR�����X����Xw@ݚ��Ap~a_p��/E=U��v
[�w�n�KBP�Ŵ|��� h�����"�G��	3yƛNY����'H�J��^J�d���|�p�]��_��a�@���h:�A�mK2O��qV��ʎ�������tMa�x�V�V��1��I��(%�I�|����Gᘇ	�� �C(����8� ��a�,�C�4M�儔��u6T��"N1R&�W�I뱛$(3m&��&�0nƊJ�ag*�%s#�,2mytj�2E�ڢ�M:1"^�Q싼f�$������Fl����$��}j��*}�t�J�<�U	z4�#,��s:���2d�RJ�yF��!=<!���Y��*KF�A���3��q�����D،�L�VI>��8�����&Z���̂�Mƈ�~�h��Y�Ia��{X�� ��^o��b��f�o��{[}�tq\��eou�\�ٍ�m�wImAk�jO�tVd�������asqq���~����]���8+���~S-��2Mf�葰V �6�42A8�֦�"���T�EN���[��ڍ�п��$g�8#%'�8H
X���7v��`�N7�v2�`�Ʌ6�D���:�%�0/�=�l�Dz���JB��v������������7��d�C����f�����g��)p��`�l�[S��2�:&~~<��"<\m�զx9G%��q#2����A;��Zb-i�PN@.H2�H�����%�xs��#P.g�\�§KǍ;Jd�ʐtWh9����JL�q�ƭ�~����ns�=�#i���-�rd}^�9xX���� }O�0Ú~��^�zEv�b.��+={|T����z^߬�����Or�(�A���Ö;C1�t�R�mv@oo���<�x�k��p�Zﻛ���%T��"��º!��⎀�V�n�?�dqr1\�"dDp��K�J��-~�b�����LT��W�޾y{��6�� ���۳���u�\�'G�i6�xSV9��r�*P���}6F�#q.�a͡'8�B�c��������B���.N�r
��N���Ww���҆;F��ͷ��>��\���{�����뻽����2@6�;�L4<i���[�r*�@�O�\6����7�|Ǭ�t��y-N���% ]�ևX?������I�?��z?I�g��@u)^�%��H�.J��v���EM`q��}�^���S y��B�2
9\\na����@Y�
���]^�ң<z��ߵ�}��R'�*��V�A�&I�O��7���$Ϟ=��K�ɢ�p��~{������%���\�t1�0��(]�����=�7�[W��?=��a��c��%T�������M��!�&i���ö�Θ݋];���,[��Xg��~��Q�7���1�O�Ļ큂OZ:���$ &�Ÿ���ss��$�)�� ���H��v�lv������[-y1Z��-��$Z�y 8�dz��� v����ӧO��t���}��y���t��n�x�)��<�TׄM�N֡�W�t�k�_��\��=>?�����n��۾|5�C��e�峥y@�viT/㱔r*�����p6�+����>0�A�!�CHC�_Kٓ��2˷�r�y��a����=E����u�,�k&�爢Ⱥ��q\-8���pF��l��x��ɧ�~z=_��`.c��]��$EH��L�9)�nǡ��y�nV���kN,���\� �p9cS�!C2�͏��H���1�E΋Wp�r������o��HC���`4h5��
��^fv1�	.�`��Ƃ״-�o؅�tu�5Y,�$8�@��gX��m���t�B�E���`�p�����4";������%a��j��{�g��B��U�	��������ѣ�D@̄w��"M��b&ܙ68H6Yd��F��5,�l��ˬ,��v�X��5ㅳl��N��'�ZaR���@�<(��r�t� ����'�M�nQ�R�O)̉[�:�u�zm�р32����1�9�K����A21��/Jt�`�I|� W�&�a��+�#N������Z�6��-�g'�iCV�kYZ����+y��Q��w�j�D$}��3�����n���~���,���JO�=�����*��n��f��/VKf:�t~�3��ʓ3��������|��9=��k���p�}��:7zr��l
H��=E�u/R��R#d"j�O��C;K870�tsT�;I���rӲV`�X+�+�l��߿���Z>�t�p�$v�\�~�����<*����$*���ճ�ƚ�s�����TȢֳ����F�+r.��o�G۲>%GrɥZ�Cۣ��٨�"ρ����Vw��8^ά8���񄴄u�<ah,��I�����'�B�&��WQo��L�S�.��-�!�d�`Z����������F4��,��L�4P��1Xɨ���\�:�|��L)^�Q�0L���O���[H&Ĵƨ�9�=�S"��޸?�����r'G�i��ն�Awy؝n��AǓ"�
) ����f�Ɏ��<���B,����`
$��a��oon�߿{Xog�
�������n*KЉ���9���C���	�ڃm�H�7P����J&�����0�rV�'x�`:+�Q�\��T5r��cRF<�\����q��>e7�A�������4�-� ��l� :D�zMˎ:g����8Hٕ�2��J:g�e��}��4����x�u�d�SDW6醶�q���ۂ�p���h��r�8Ȼ�ޘVS�{L^�7qǖQ���J�:�Y˱5wľ�M<�d.�;��D	y��,_i��ym>?�;�~8*��p��^yB<X��n�Щ���9�6��u|��=��`ߒ�����&��N	�b;�t鴖t���V$�z�*!�^/�Y�������Lx�AOV[0�KL5��|n_{R�x�x�^�0�m�fr�M���2�=�Ax@|�s�Pjx6K�Ј�P؂�RK�'�A�A���<w�,l���Z�0)����o����yB�J���������L�H#�p�r,����JƩ��51-w*r^ً��<��ʙNl8���`!3��hygK��t�)-&'e�Z�ό����fM?��	[%s�@b�����/2�d��5�,P���&���W�tw;����!��w����?�Ïn �vyy��qH����˗/�i&�j��p����
�����e[��c:jF��2Y��2�����{�߃~�G��%Ʒ-�(V�"���A'pa��_�d��9��>�^o��ڎ9�uX�%˃O���a���FN4?���o�q��R�z�G2����i��" KI�i���b�=�i=�Xt�����pR=���\��fR��`�}��C>#�g�_��n�����;��KMp>I���a<�èiI1��+ow<��	-�D��9�t�BW��o�j��'���N�7}�a�6Mn��@�� ct��v��q�<u������"^�9�%�=&����c@!��h�����<�o�:;;�XaPGӗ�����N$��f��Y^p=�����lVc���<�uO�SDc��J\���;L�tA
A �xIry��Vr��� ��DU!%�fX!�� �>5:)�8Щ����x�8?���e
Q�h��Em�E[>��o,��ϒ�-�螇�ܕ����5�ȂL�[̯0��š��v_x ��@�y7t���]ð��r^*�*0z@��J�<�G|��۠�|��(:>��P!)|��� G��u0[��y��~-ۈ3�g	1�i���
��A:��A��g.g?����δ�@�!&���������Eś��ŧ���/�o�C�<(eX��c���E�N�!5QJ �C��0�?+�nG��N1�������C�Q₩��)�g��$���彋iJi�g������� /�D��\"��X�tB&SH	~�0���ՠ�V0�^K�"�{�׃1�
�����+��A��i �M�0N;$��O��q�M��AW��3X&�n
*��
��-*���I�����$�T9j�N>aĶ(�iV���H�m�v:m���E��QpM��Q�"�-��Y�skF��ӗ�$h|�=�%�F�v{��	O�]��DBSI9��e ���SO�+�S��Ƀ9�^�85Hd �F~�ה4}�l����|f}9ܢKX�IMf^g��S�*F�<�\I�u����D�O*7��C�{N:s1��l��㏐��(r�����#��;O�#\O� [�Q�0/�rmٙ� ~2�Ұ*�Bbg�	0�苲�7��ٳ���	k�b���ʶe�a����|{�qo�����D��ΓRa������� #{w����	�8���Ny ���58��%���΅��>jg�W+R�BR}H��"�'�&;v2Ë�s8�]"�=�E�y+L��L�-�ط`�Z�-�X��� S��r;/���A�[4m��^!WӤaP���\_3;�����
�����B2h��|�
7\�c�lZdq�[H���0e�����|�	�G)5?X(4��C��NCQ,�(�&���Y���$nJ�.8��:�����\:xh�� ��+`�0��̊9J�˥�Xqi�H��R��S�P�Ǆ��F�4�e�ӀMDh����4,ų� ��K�������4s�'�ͅ�M��w�^�^M�O��G�)JHb��$s����db���d ��?;�/S�=���ma�<fo��:vl�g�&#ȖӴ��bN��8Z�@�(K�]1����|�,S�\��u�p(�����$M&���! ������vO[�e�[_ }(/�xx��YK�@@	�/J!�G�o 7!�=����옹QjqC.�m��ZP����L��V�L��l��0K��=֣`�ܹ����}{�'���o�'�U�(�a7p�vl����r7��ʢ�4g-��;:�xz�D&�%�æ'��iü9�Qs���V����y�⑃&�q~�M�-k#Q�$
���J���	Y7�n�AP}Ƀ���-q���s�Da�MCe:Y�������V��y��M� 8)f�/�ɓΗ���`�n� �'%�^y��`SB�_�G�[@��ϲi�V¤��g~��� O���/*F���p������Yv��L������4����#v����+�͸o]��I�y }d������W���s���ۄ����aZ����kG�%���g�)_�.��zX�^��@ֻ��n��8�.��pRƻ��FN����vp��M3�ۇ�l���L��'��$e����v]�����_}swu�H�����P䌣��sG�ˁ��Uն�})RǧI��ì��ẅ*~�HQm9�t�G�L��pc-)m���ɏ��n����������Ņ����ĖA�#�,�-��Jl!�i������V�]��^l�Ɏ<]f�a3
��k������ayz.��1�l�<;r'�\�u��浨��s������S�O�$t�X��.��>� iE�y��g;��%W�R�����b��P¥=��:0(���:whBQr�s؊cR���;�1�Z�Y��Ot���)�,�wo���f�=�������.,2k�%� �jP��va�F����
5jN0	F��E�/%*�����+�Y9��$r�iIq�W���0�M;��'�3�i;_���7Y>��Y���6�$I�g����G�H���t/�Xڭ��m���q�!N]��ɒS�����"�P��Q@��₮��ŧt��|�}EQ�A繍�-���;�<�"�����b΁+��c$9dQ�I�C2m�giP�J?z�h�Z8�w}� �My~δ�$]�7�m�<�R�����4� �Xҗ� �I��u=�b���m���zs��]5��}��CגK],V'm?X��e��h&ӷ�"`MP~0G�.���Q���;�ut��ӚC�ӎ�z�<�^#>���L܈!gn���c�x&���g#�9��C?�u� 
:;
{��!����Wg���ޯoH �r޴dp�䞓�\��a+�o�9ve���dI�x��Թ%��Y[�&t`n�?3�;�G���Ge� �+��V��F�4\s�xM��g�FqN����_����t���l�/3��;��,PV�}0�����&�%D������6:�&�m���z��y*d
�8��Y/�8�2ӆ>V�<����_yu�-}��ih*l ��U��)	�h�OX(�y��	
���Rmpr�� N���H�d&�Z�� ���wf�Uv��LO2I\�@y	������,}���[�dH��b��S�_�S�b�A�F帰���+� �Fm隺^_� c�:eA	R��d�P��4�J���#HNb+�+�Z+_�$k���ʖ>���(���@���q9�=@<��	7� X����\<{��2�	���Y��`O�2gVB��#�qd|�U� a�u���	%����gdM���܆�̛����j90����t|cd�r1bƺ�x�БnHt��"ʛF۩N�2OY`$��:i ����t3t���6d�_�����%c���}����q���]^m�;�X/����g�²����m�q.*(��,>�\�(`X���ME��)�H�س�$H̠��P!;- *�Μ����ѽ\J�J�q"�^g��,Z���6��$XC�5���K���Z�I:�gL*1BBC�,
��mi�p`�Q�.���>E����/��t��� gQosg���:#�Ǔ���/����.1�I�&,��nb���"��,$^j!�h�W��O͉�{�j_^^������^h7"�b������l�$Ӌ�����EEj�L��ʤ��"vH���I/�M�~�n�={Fo��)y�=�dD.HW�4�V�q"�JRv/ hK����o���	A�C��FL^.�� ����Ú���+ש�xC�d��hh��M�\A��y��	6�Ң�'�V8����
N�i���̷��i!s0��I���X�"�G�m�h�?*V�?�}@P(�I�J;��:�5���>��~��Q�	�E�Oo@�K-�
S�o�������Ę�r����sg�Q��
Ix3� m_@�����hⴤ�)y`���K���<n�y Ç��3�+lp��Y5#�9!���0��B��@Q�n*��aD-V;�6_y�N(��CS�"�O����u��&;����7P#��bw�"P�e�&lX@�2=�1���Ni��y�!U�	q1i�7_��k�/�|�\N�0[��Q�׾�!�l�Qҁ�����~�aY�9n& .�����>���L���i��K@N�Ç�|�����6�I��m�0ͧ���8��+��( 
r�Y�8�V�o��@=-�yq\��f^V2�t.��e�ϵ%��g��C�t@�O��#�-�ٿ��������U��QH�F��3
�\9�@�6jw<G���+��a�ٜ햑z'�K��@���;�{>����հ��[�b�7 }&�M֊Z��l^$*,ά���1���D@�{�'�x�'w�нs�G�¸Æ�vt̥������J�9�9�����V��#�b
� a^]%(J��:�f��7�>\�����&�N���,��v�#U�f(�cRv�L`P�D���Fr|��.42p�����a�� Ⴓ4(3	-�!�j8g�=��a�ZBTV����M���N����{t�C-�.�2L�W����W^��1*Xj|5 ��N�>�k�&@H^������8<(:�VN��z���d����Ω�ȅ�4�$�}�siS������$�	]��`�9z�Ղ$��K�~E�r�[��ȏ �������NXtYfR������O����Sm����s���Di� *�(y��~�)�9���(F��G�"��kf&�/�T�o��G҄ªi!:��R�Ho�x���L�<�9z���rC�T�M ݐ����S["����˸?pL�q�2�;˘�fbfN����WH�B�>rZD$Xe�S��<q�j+D˒A.�VhI����|�ɛ7o2A:#�9L��~"����*#�˗/�C����BI~��:�,h�� ���)CKHg�d��A�;ʣ�9�FX1��(s�#f���Ni�u���밠t
[3�OT}uX�YR7���IR�,,�kP�?��}8��Ξ�� �z�*%�a	��6�K��e|K��Wf���ä�)(s4j�i 3{�}K�$��27�gG�)�\�㤋�J�<��v-�)�v�v^�?0���}iә8qpr�����
�C�F��㴻G~�1��Z��������@�al���Q	��P$�*A�@Wd��5f�T�j�: ��*�4l�������q<Y�O�Y���)���;T���"K�l&�N�~�w'�L��h�sm��)�Ș���+ֳ��"_3�UJ��	<�/�?n����KG��Z,>s�B���t=�������~<2��c@4h69 `����?�|�`}�~�yx � l���aG���,�8+�����i~��ߋ���"�}Y��Mj/N���,��ԑ09a�"2B���j�g���ÿҕ��)��e>iz�P�cϩ����:�N��N�v{�sF�o���3nX(ۨF|��+��ݒ)[����7�`05~,�a��O�:�	�x�3���
1�H�Һ"m"9������w�p���;�������	z�PHcї�Iq"jWr�bĵ</��N��J��x����Mw K��̢�҆��^I8 �蚢7�[����_�����|�ŷ8��0􏋁���4���$p�~���@�#��;͐i�i����Z�]N{���`z��m���s��p'����Oe��q2�"�61$鑱a�������/ޮlI����R�.f��yJf5��c������	����b++c�nV��bQ�����{�w���~��l5/��&��Ud$�I�Z��wޙe�{!�Sz���،"�}v��� 0i=9E�y�jI޿u��Bȏ<�<�:��� �F��rL(�:QDI��-OŅK0	\S� !�a�::A2:�(�J�:lLw%7�xv��9�}i�NL��@�Gľ��;�XD�U�\������?�0��F��Nl9yة���1&���tfgg�������kH9N����!�d��ً�V�Ckn�tq�p���:���Р�r������\�| z�u�N���;��&�f�(2DR<�RM�:��|wk���@�vdI�������e��n
s:?~$O���?�{�DשY;K�ǖ{^�l�9�4���}揘G?�5HF�]J�n���pL��s^8����F�}v�A`U/��������|�t���P����|�����^֋�^��B�K����+�z�m���0�����S�[AK�a�[��)�}�k���QѪ�zN��g�5�i�$�,fC;�D�3�"���N<
��%}w���!P�ڭ%@�x��YA�[/œ���)��O(�&+�v��4�/�6M���f`򬚝��T���<�k�U)J7�<�=w�����4�c�
�.9}�����YΝne�̤���-�~;n�&�X�¶����S�(�D1Q^���Ö�&��^@X����?|�����~���I�,������o|Z6���E˺ٶ�,vN��jn���#_�J� bA5�q�~SV9Ϊ.��W���M,�8�����x#/F�5F7/��b�bͮ��du�_�}���"Ʉ/��o�W3F3�_<�I�$�f��=w!-$����d��n��7���Áтd�mlӱ|ί3z�D["	�jyN۴ݵ�w�%����w�S�|6�}�JtW	S�d9��(uC'�� '��e�
/k��O�v���==\j��9�$���t���׳E^��jU��i#ل�r����0J������?�Hct!RԴ�I7e�:��x&��y�Պ���adf��~���;��)��v�s�^nv���z+���;��r�2�C��1A��E!̉����i�ؼre�D�g�����g��g=;���ݡ�=~Zϖt5Z�͖��"'`����o:Z����p=�+� �QrK�S���g��R\� �wҖ#���2��pU�3��%���g�W2�f������A�41����Զ ��ŋ�G��	���:�M�s�(��g��><TuIƁ;k|�������
-n���A!���)�(�.��W%\2���d����!	{zV�9���J��ǧ�@���7gR�!� ����j��©],O����MZRa��������V�J����Xp��b+Q�U�������˵��+��J��Q�@�$�uY��f>���hP�$-A��VW��5��q�|�f�[��b��7��)�.W�Az�E��6,Bפ�|	�P4w�h}��~�%\*LCQwp"��i�܊.~R�����	}�H���������8���
wS�<�p(K9�LZ|��L�h>��ڂ��j!�W�e��>��d��L��4?j%&WP�ӂt�.*\Ĝs�q�^�����ߏ���>l����<�A�r��ɅrqzK��Mu{.ɑĺ ���_hW�����K!H��jyJ�w���֋���Y=g�ծ����u5g����-Y����+WAf�<Z�x^3�*�re���U3��%��6��j�@tdXɓ��K2xMGnyqh�Ŭ��?�	�F�8r�	�V�-E$�(;H��{�ļ��0T($$o��k�� _�&�e�s�ڌ��������~���߭7��(Kc�f+Y�eh��Y]��yr�s��8��;�I��E2JbR�����\K^;�� �KABa_���pR |FB�26��qU:��yc-�{k�a���2r�����n���l*�^q�<����f$����c��>Q�^�O���"�T��y2����tԇ�����A���U�����M�l'���Q0O���|�G貧'+|����Ęһb���"��"�)�"qt���3aY���3�!!�=ɂwz��@�fY>��pF�22i'�οĲ��FV{�Y�ܷULZ��6�wȵ!� ��p�|s]���{�����;���]<&��W_}A> ��V�tG		%�Vb	T?8�N��8�,O�)J-=�V�Z�0�	�UyK~�|�?���$1��q�-��;��~;(�;WҳL�0�����-�O��H�[#,��PY��}�&1-�1}��/�����Uz���d������b�C��7�o��h�����?\�cnt������3��;
�!F�LrC�KYd#E��!���� �6�1O��G��5@k� Ѓ��2~�K6φ^+T氚�e)�㢄`��k^�ks*R�8Y�`9��6�<�A�"�s%�p
ն�T� �qjQ"�E��9,��#͵R����'_}�md�f�
�"���Z�|��q���pk�ĎA�X�_S�b����b��+����(]ڌl����*�\��s�lJbN
��� L�o?z��>�A�f
E��)�<*2����./^|J���W__]]�*��/��/�]TԤZ;�H�¨�R�87��&"����(�3�Y�4�K�Ap��掳Eͱ�N��Vw4͞�#�mv��%p����w����&�fCy$��\��1���C.O��
Nb/�ʙ��r�?%�hh=D�]�8@�:������,��l&pZ�<M-�A\1�����E�˕�	��wƴ�5	K�U�h:��Kl��|9��������A%��_�ejav������徤�:VGc�L�j�k�)��;�bF  �X�Y��5�����p��ª�7Ez"��"\X�#��I�3�5N�K10d�H��M!kv�O2�(_.����5����YW�Ԅ%Ql�\�W��!�|������5�n�?ҽ4�[([�{��������Ca���0�>����cbJrRB��	�� -W����8���!Pԉ�ì�T~�w��B�B_E��w�p��� ��LL��5+��drV�y�Zas�����%O�\�M �nrZ4R_����+"3('èør��

;a9w�i�m���G��k�1Ȥˀ� �����r(�U�Z0��m[��%~1$��oZg�C�<3�I/�$�}��C�M�B5;D����}7`�&s��%�6b7���!�]����ؾR��H'�yA�Z_��@k��d�i=���w���͝��P�Rr?��u|)(83�{�G�l�x��	�Y �(�]	MHz���0g��'�|��A�$�0���x7)�#��+�G]'�����R(|��h�� e��̅���|�,P�N��9�'m�	\���� �\	�2E�M�;f��?�#��1dt�P 6�_�M1�
�bΠ�`�w���m?�C�Ų"ʴ��zj�W�#K?AK�q���Ц�L!��6gX�2N�q���>�꜒�H��ϔ�и�,y�;�t�XXb'��ᮀ�h��0y��7[3N����n�0�ܢ�8!r�A�N�,����$#�G�G�f]sE['m/���Hvpp�Ke�+Ւd|2gjw��ϊ�+}�s$������[�9���8̡��~��f��`��f�O�Uˏr�<�_� �)=�5�#&O���5@�����L�ɽ��O?���~���?��g�Wu��-��A��mq�5�i�z��B��N ,i3N��NR�'֦�X�s�d7�����|�ƺ�x�/i`�FO�uws���T:1e�\��yBZ���h�!bR�]M�0Lf�f��C����(梕+��bys�#;�MINi?߱���s:�|z�m�lޑ�dI��AS�62 �g�AiU�JdPy��](�4|�bs�-�#Y������x�Z�з��գ��� �N�/MU��)�UE�*@|E�'�*	cO��2Y�O:���� 1�����c�O]\\Э���x��Ҧv�,'3��!�ey=\����n�T:㨝.ej�� 	ˣA���(� ��Ʀ�M��A>}��tV����~w�k�A�ZEK^:����l\���O����(9�Dzi���ȕ3�#�ε5�}כbGoT�"9���6��Ld[o��Ä�	͔�Ҏ��k!���.��M0�vx����&(p|�f����A+�� �$��&�F���d���F���t@If:$��@n�?��;��I62*=�<`�:�Zn��(=�$|�JVx�6wmf\uA%�v�j*>gߣ��\�f�b�I�i���*�p�g>������e��3
�7�lX�J�<���B�$��2%��c��wC�sӎ�#)=	��c��.3fK��r��/���y\a�;�,��%��Dp�i����c6B`1��(������n
��d�»ĭX<��|����q2��iǜ��5��%W����A�ڦm.�szY�!���o�s�>>o���+1�iy߮�f'S^Go/
���z��v�З+��Ч+�Dʋ��� �?VO�_��A���|'}^)���	N^�A�)xd��ei��Tq��4�K��>(��
6o�1NpZ!7��v!�.��TQL8/%"�Ub�7�1�ϐ���?F/�M_��T.4����?"+����jvBQ̯����벪��_�����a�}���뢬������s�M_�~�5��S �;�� z�y�	��DF�;a���g���Y��WB�k�8����I�&[,W�_Y��22̀�e��B�i}��X<��	��F��V��Øz�%����j�܂}�2�j5�яL�*��w�_1?rv-3�f�#?BbԼ�bC��@���������2�e3����5��z�M{i ��10���u���/y��� �*$�����cD�~G�%W�i�7�Wt/�\_]qyV���j�vK�En<ұ�-bT��eaP���Q3N�yHj:
��P3-S�-f��Y�U<⹐H5��6�v@��RK��Yd�e�T7~�����3F~Ŧ[�C*7N��E^�3����a�r|���]���yyPk5;���V��������6I�Ⰷ���h�$�v}�V+�þ�m�|��8�EI'�.��v�C���S�AZ���,𰑯��Rz�-U�d������#C�8�Μ�c�s1^������<��v�7�g�i�CKK&`@�S�C�C�yri�tɳP�yK�T^ՋǏ.�aj8�|�o��� �tA��0f���՛w��ޥ���B�W2G�ppCJgM�	���V�*r���������[��A�D�!+��BF!sY@������T�����<�;�@�o�4J�Β�8:-�w�5O*x���+�e�zC�>�Jc�Z�2�o��*���u�×��{��~b�2���x�S�THs_>a�TcU�[�'�}�����&߃���ܯ��s��N/��d/�6Y.��A؎2�qh'X�b��@xH�4�i$���'g*%�m�gON�'�:�S��-�;�	�����ܑ����N
'�#��H�EŰX���]J��ڙ�)do&d3���z��n��_\����3i���p0�Q|t�c�ӈ�
	�޲��X�U*o��Ap��o� .6O�eM^ct�(�t��Ʊ"��E�� C�2N��@G��Iy;CR*���Չ�t���ؖ�LI�˗�^����:<r����GrZqZ9�g3(��҈A	������L3<��(�{-PaU�Ax2� �d�8�2"[��ƨhM����)���N '��Ch�%Ų����/'��e�qҞ�+˶Ӝ~�F�L�@�i4ۖ���;�����ɨ��0�5'}!>���<�GI�M�(?0k���̨��zm�� "���cts��6��^r}��4J��Z�����r�3t��ǌ�L5��c��������f?�R&��f>~����!A(d B��w���_�ϟ�����Y��������f�XqByd�C�K���[ҖH�0�I�F������܊|�����	%>�@�V�������ٛbD[\��\��z����dTA|LGu�wL���]�9lۍ����aO�%2���)$���$��;٠�Ҏ%h���B��-V�G�l��3!c�j%X�4�.,���K7���W8jHP+mD� ӝC�&�Q�e�%�9��ނ]�݋��6.�|�q��e��������ޞ�<�ǴD����=�r����x��b�/�Np?���	-O�2>�����Č�6�Xj��T�8Z}��H@�#��F���ɓBAܴQ�%�vDʙ2B�~a�999������1�6��^9�!Dc�����+�`C�z͊�|��P��j�aX.f�������U]r�B�_Ezl����{�l<~�8Ͳ��K�o;?�����Tq9�f�q�E��o7m��e����T�����Q�p���^!���1���}�}�<Rcgb_(aE�p<����9��y)&x�\�4��ӣ��
0τCQs*=(���=1�'R��(*��<���pIZ��#��*BRܠR� �a��*Yn��F?~,��g`�4�N&\�]�9lx�Hjd:v|�4��K�xRK�R�.f���̈ZB�?�]�`��雃��\�R�8-H�I�7*tБvf lwK%^q��p��l7oꠟ���q�)��''l �r���g�������czQ<�I呷%�BZ�?�]vH ���I�n����A�����D`�'j1�*����T��)�q�Y\�(K�<%ÐI�$
�C��d���^�ȱ=;�������w4�r(8��(��	�%�	����ɤ�^]]y���	����!��&)����T#z��7
 y {�ڍ%��# �Ϟ�<5���BĆ�'6R�,1��$ɪ��"��T�����t%�b�sM�4��'#�""ʱ%]�_29�=�hPCC��������>2�-�^����f8��c��T��QR�M\�E?,{�E�����8X��ɼ鳳sF��L���#1���d���X�pq������턪oi�G�I��;?9e�����h�i���9J$\�0�f?��~��6E���"�?L]�{-�.	����i��I� pG15��ł?% 9Z�85ݲ������	�d�����^���쉋��p����2����I?l�|U���
ykV�ǫ�S�'�D��+;�4e`�&.����d^�x|����TxvV ��WW7�l��9q9�[����d0<�����5`�>����qZ��H�5Q��d�)�J�GP��ͥ�l�ޖeR��z@��X!ӝ �%�� _�i� E����K���(xT)��9��7�}CK;�Q&ͼT��fE #ag�C��)�����M"�0����yBR ��0ς���e_�x�� Ct`��>�n6*-&����Y�I�ʗ�9�b#ľ�CE�]-�rs3�Q�){��2�GpJ#S�k�}�;����k/,���}^�NNOaq��	< kK��"�����\�zBݸvo�!w�op`v豏r^87$o{1m2�������I�A���W�z�6.�����g3F��!��6�Wө1t�En�Qd>�{Vi,l��I��!x2�i�5ᴬ�-����x�n"%����������C$�1���W�Yx�s�T;�٠�΂%��N0�&su�R�N�1Pޠ�o���v:��OPx�6:�'�)s���g���|B��EkN� Q�g���h�v%7v�6�$���M3Y=������C�=4v�j�}��y �`n�0h�IYR������f: �k/�݃�T���4  ��ߜ������¡���1h�/�)YOoΞ%O��=�����Ԇ���Q 'aRB~�x�W�^a#�0@���
]������5�V=��\
J�L � ��=\b:Ȳ��%Dz�E�}��*DW��O�<��O��'��m6l�yƞ�D	�Y�	��RH���!�@�2�]F�7m�R�K9�}Ο�~���d�~���q�n���{�3�~��-��8a�snɕWYC��������B���7�ę QJa�
M'_ډ��_�	FEؑF�C,�˗/�{�t�`�hH�I
<r��x#wE��+si����J�.�"�����,'�Z)	S�/��ߎ|�0�b��������pV��,�K�P̻ ���R���.�yq�ȁAc���Mg�W��(�,@�b���
d��n���q'P�QǈO�������N	?�r�$��9��֖Dz�q��AV�̐)���"1+��Ąsvn�d��Q�����t:�7	(������O�]%��(v��I9
Xdx�V,�u,��s��bTZ*x���x	�«���D�������)�"�6*η�9RL�M�_eS�Q++��p)�w"��9~^f)���﬽Y�e�Q.��{8C��YY�5�. Z���#�?�?�/���K7ݫY��h���RY�sf�q����_3���x�$�w�>������?�L�p��)�^D�٢6��U+-����:�>S�*��m�a��8-i�C֗Ө�z������1|�N�Aч*�d�:�FKȱn�GW��OI	xa\V�kp���C~�N1W!T{:���Yu��)K�I���ᖞ��P���%_O��[iy����*�����님������,l7cõ*�DܣX���aV���|�Ulq�gҗ�Z{�D	�Ӂ�f	k��#��o���W	�?GZ��PW��a?U��4��;�$�@H��㫭�ꤑI�x�e�i98�-�0	��V��&F�]���~�C'9�(�&uK�o�mhy��2U�2IG��Bj�.����nr�fVh7q�L�$�q;�ɗ��������>37�f-�vH����>��bu|���>NZ�}S�Rյb	��1�N`&��ӒYbz��C�O2,3�,�b���10��īa���(���"�҉-���Ã���Z��Q����߾�V�H!�]�)��`i�w�%�iW
1��X!Ԍ��N R<�`�Dd��ڹ�^�"{',W�w2K9.-z`d������#�1L�W��dn%>�a�a��W�)�� �a������7/^#YM:��b�V�((ĩ!Q��w0Ni}qNf+��<]]��͂=�NzM0�[���b����:�ۛ�ӛ�5,�맧��On���t�n�e�rr[�t�Mɓ��lj�&JM���D	<���f�f�����b����0����=p�1͗����GGŏo����G;��jfR��tSr�Ȅ86|ˌTYx`F:z�I����/!����DV����I1���J4!b����j��v*77�bzwu3�9�{A@��k���v����8��QAd���e�A;��Z,��Y/^7Ć��h7�n۷�[�z�͕�m�L�]+p�p�*qU��3�-��F���e1��r�����	�<�q5M��V8h�Hbqf�u$���v���)�S��zz�#1��pO��p�p����B�7!�C31�dCv�cZ�w�Yf�׹�캖S-�����}�1Mye�:�[n�ф4��).�A�Slgs�W7\�K+��K�r3g��/��oW���3wʮ�[�Q��W�����&#��mּ��AOd�.���/0%���ExI=1�s���k�4�۲I��m<��l�������g4�*��F��H1�0 	wҬ�����&�4҉k��j�����u�"�<3G�cc�G����[_]'�0���l9-��%uD�7�$�B�X��n/�
��+3�RG6n��=hؾ�k4�[�4�/`\a$�ooh��ˋŹ�a'MV��%,�^��@�ڸ��0^��2{mC^���!�Q��t�7/��+m3�Z�����ӹ�7�H�o7������DC%k'��Ų?8$�4���r��4�=Md�,̆0�<���ِMZu7������iu#ݝ���G>�c&�0�ۘ���i��H��Q���$ ���〯x\�8�z� Bǖ������/=|忌�=-��?�%�=�[�lVk�����8;��5-�R�p�y׍�R�����2.%��d�4����&�J������t��h*(0��SЄK����>� t�	�f&�9n����4�W��LI�Z�6�`�/k/�a��/��.�p�p4�ن�
��(_�s;��pYҥI_�2	�D!�X=Zw���t�r�hL/�6���9<�eB�Y�򤍌2����Q�QT��;�Td�(�I�D_�{2{�c|b��K8���һ��ڢ'�8Ac� }KN!kQ��i��J�c�q����ϫ<+դ�Ҙ[��5
�3��yc�/6}����I����j�����_V�!$�B��8�3��*3�ڎ����ҕTi�
�N�ϫ�K�ز����=��7o�<��� �ٖۏ�ø!?��ܢ�ˎ���zM������R�����/?���<��2r�3:��9Yh]���$?[N�����R�����%3�|���{a��.7����;9:�����iZ~��૯����oI�<}��Ç�0�z��ŋWggd}}�˟�<8z�������8�F�rvy����zT2�n�����8���0�d�6W[����dæd��V��7O�>�[>���>���
��
<)2Qw�5����	,[���˷�rA{��#�L�|�=&�Aةi윂lٸ�� ��"U�za���9��!$� �C�6}����g��E�̢�8�,	SC���r�93k�y�� ��&�sW�A�|�֐c�&���<��M��'�PxG_�6%�C��"����I���i�?�mXZ
;MD���
�5Eq��n� ���������]__����=�0��tC�...倓�� ��u��EF&-�"� ߓ	�&�����cH�Ѱ�߿/�-������@C�����o����2MI��������Yoɂ�'?E��V��.�e3:�O�M�f�V�:$GBb�����/��_�yMr ����>����!�	�#4g�dss��s�ׅ���sE�D?k�K����`�
�Z���4P;^��ua���r.�l1R�7�݋���/6@p�[�!���_H-9Ly�"��6�'����_��![;�YP�t1lB��TA1jg?3��(��ɠ��ub�Ѣ���u�(K�7HfK�9W��a�M�Q�F�m- ��@�R&a�ϔ�~	\��vE��b����[�e3��ãIV�ϝ�p����gi���J�ŻB�"��U��h/�*���H%�r#�s2'M��+��D.�@��h�l-�k	,v���Ľ�=���/�6����E�L��e�*�	�UF��i"�&:h���lz�g�Q@��N��(�"�N��4k|�iK2��`��9��A )��N{�Z�4g���\q׵��RV��!m*����,[GE��L�BN���N�<"C
_l�8�.��m
詰���W��t���C���6�F���r�j���p��Z[qs!��ƫ��4�!d*(�T�]+�U����������{�n����%���J�Z�{���i)P�nw��MgE�`J1¨�+��0β&Ld؀'��K�z*V��Ɨ�Jr�P�gjѸO�v���X�&��1�Jhˢ0�|�
�Y� ���o�����t�����i�
�;ja�����t��JD��w��[����<h͎;�&Cs�[w�2��v�Q���'e�o�ϰ��25��"�x�5H���q61r�UVX(�i
�^��k���0�H�s�+딓4V������
��F!Q�;��%e@�^_�0�L�=ɉ��EV��vG�4��4�.��A�,ƛ�,0G��=	�ޮo�a
2i�LX�h�@:g�����Bnڝ�Z�b�� �"�dH��U�l�h���R�� a�`M���>@�Ǐ����_��W�Vz�>� �O�h jh��P�z"K����v��rY�Z~xM�Φ�  ��IDATN�@f���yq�:;/5z#4*�� i���H�'	~DШ}�����+s9a߃+2��&r�;md��?d�ۄ��6�覣J��T^$�������~f� lC�DŁ�nn�b�q����1���_��g��H�F�9ݚ��'�4�=�y�E	 �`�l��C���+��!�c��¨��Z���/�Z��� �����������^�&�GK l��p;��,�u4;��=f���
���/ՠ��P2��������ȏ�T����;��/e\B#5D\�IFi�l�3jI&��^Nڿ�����˿���&Y�Rm#ɑ߱�c�Q���x���;>�b685⧪@�Qh�\�@����]�'�)�A�jf�@.^�Wu�*JS_Q�w��/v�q�L2c/8<0}1��^�QQ	Mե�,XL���4c�1�4Qiퟦ��,�Uls[�$�����S�VB�!.i�y��t�8�^�%��
Z4�܌d�ss�=P;c��BF�*��l3z���®b:j �̛�^�2	���=��mf|�t>����l��?��T������9)ʟ�ꗤ�����������[��Zb�6�b�9�bv�¼�cf%"\��\����h�͌�a�l3�E���j���}ógϖ���<�����;���˿�Kz���g4�W�^�t�2��H��l}Ġ]�&y"�W@�rM��6,�B;!�ںl�Td#���.2Z���=���%MT�aQd�\�p�%��0W�!��͎�b1k�Ҷ�v~'Y\,=�� :��,��Y�.�����q*�:~�!=��I��6
X�a��ۋKA�����]���zd��5�#��H�y<�a!a6��}AU�$3��	JJ�d��ϔ �A�<�%��t���S\��('7/G8	�� �7�HQ�� 9)�g؍0��R`$@�?[`!J�"�E�_s�,���RN1(I7��x�
�z��h,��G� �Q�3QW{�1�R�C� ��C:{��.�Ο<yr�,àk^_r��<J't�NPյK	�Xl{���bU̛�B�CV:�\��B��SHH�+��TX�� \-r�[���6�ڧ��~Pa�o�:��*�}䍹�f��^��b�4k� �}L5U�o��xQIU�Ҟ�~�twR�Z������;t�S����<E�Ѩ ���&_Q�F�l7�X�t*S���x)u�������2^���ȥ�{�0�'��+[�$��~)L
f���M�@�\�U��h�$�e�;�s�A1�M�tEK��ؤm��$`㠑c�%9���	k)�I�Q[�nB��VÒ <��6!&�3w8Q[�o,�x�*R���L݇c kS�� �.�h6[��T��wD��\S���PI�8@i�*;R���f#�6ۂf��
wQ�N��I��]L��ʴ�� �W+��3�V�ȡ�h��G(ߢ!��C#}<�2OV�?�"R�r�R�X���&�ؗ9h�U�OR�Ȓ�e0`���Y+��,\���Y@�A���	�f��9�Δ:v�m��dfî"�Q�×�~���p4utM� jdPb�x�L�� s.�V�	��b�K��̑WX~au��CW�pu}qͅ����Y��-9��\؈�CV:�����y ;c6GG��gN۸��� �i�� RdD�s��R	��.�۩��Ŗ�S�X�b�	g����� 5�D}��,G<�X�J��C�]=0�@~my�Ф[�,dϬA��Ή�ڕ̀u4�.ܔyUʍ�Ps$��ڭ����0��?�.�CS��x�8t�貖�`6`4��M'&,
"���ѷB�:]�O��4^]����2��n��O�m��e:8d_r�h!o��仴��b�pߡ㉮�2j4�VtV�J#�e�n� ������ gh�1I^^^����~a��)$�t���R���r%�ö]T6�N	����Hk��A0vJ�D6'�^�\��w��%$'�x�N��<UL����t��JQB��J1;3�E^��$Hfz|����N���Oz%p ��a���8�.�+��#�%ъ|OP�B�:q�|��v���񧟒����i��U�j]|�K���y��Z����4ʍ-*��?JZИ����& �p�'-�4U�x�
�d!�yC6��a�������] `I�����s�5]��dF��_l��ˍ��4�㏭���f+�����N�͊�k�R�!}!�,-M�Jq���Y�,m���*0� ݻwJNi�-��O�N)K�++(vŶ��(-��@�PO']��u�ͪ����SӘ������qw�o�r���=�Z���TęC��Z���i<ӞY�Z��swyk�_�6�����T�󖺶}�T5ŵ3�*���/6?�2QԒ��ks5j!m}q˾Ԃk��9~���KfuX��Q�����,�
��J����¬/��&)AՊ��+��V�
�;H[��:�S{M�8��b����U;A �FmAVY�}��!�����<H��P;$	K]Ix�p�^1`߿{���Ç�����_��?��'_}����gzn�|��y�,}�3�^�����{�Е������bܪ��r�\�LX���@Yc����3<���ч�a����8�%�����%��/��r9_�"?ONN�߼�+<��/�$�Ruq��v�vIB�4oW�7��W���q(=[%��r`��Ӧ�SI��ЀG���j|�!�^A��¼�܏�|��9C=���Ηc���b��a� XcnT� ;W�
I���p�]�P4
>Gؐ��A��ڑ�EM���ʥ�$�"_iO�L�Er����;�?�A����F��u�ek�?ҁA�B��2�ɪ�A�Br� R��4M��8�C�*ni	/�ȴE�1���NHls��I�:���˾����I	��:D$��ō���1	��i+&��u�B������Q��,8^Z˃ª�7��d�����jt�<��,4c��~���y~~)af�+�I�����%�2��������h:��7�-1�	�;;Fd���.�+n,9��l�O�)W�ߛ�)_Qﹻ/�Y�ϦP�9s1Fmih�-\�U���\�c��p���S+)�R=u�j,��n:��xF�{��vJ�Q븨�E�Q9������FѸ!܉�E��-�M�����l����&�&����ܽ�B
n��AYj����]�ÐM�ǝ�G$��`twê�<F�U�.�J���S���IX�h�H���ZNr)�`ߵ�œ��;k%)����\�#%|$�I�X���M(|'����d1���V�]�&�Y4�"����K[��
�63ҧQ4�y�Y��^ڶfY�6�29Yqw���5b��n�X��Y�c461�Y{fٌ�U��^�����{��vU�S�Hmr5�5pj9�U�F�ld$Ɍ6"0IGe��
��]������q�������^q~v�jLU���M����s&�\���a��sK��
[b�h����`����]�
�SX�����[�9�\��ʅ ��M��5������}[\5h�BwZ2��YªL8S
�,w�/���XpY��J�U&��r�!ܚ6$��޹%]�m��8�'F~���Oh�
:gA4�]u#���[oW�a���X`��Lqw�`�~��$��Nҙ0i�Jی�m\�	�(Hm�E�̌@� ����\\~�2��Ʌ!��Z.��n�ܩj�M�歴���=����v3��.njg�kbP�_h*d{7��r�RML�)v��FOm������	��
g�ITv�����$�Ty���?��y�[.�_\l�szZ3s;�C:�t���ϟ?����<��8�zSҦ���G *t���-�kl$�<ųgϸ�J��۷o�D���d胚�8����ņ~?Ȯ/���)��d
�9�2�l�-B��`S�v��d�b�nL6Р�|� Â�&� VxR�3 B�ˋ���7�y�M�@��-@I��䓏H���;�CE�P!Lj��A{�*�U���ִtK�ܚ�5H�� ���� ߁����f��!!q�;��0���3&���ku{�4{\ _���t�1�C�˺kP0��/$: 6]	َBV�"�P`��NЋ	^��cdgC(�a��6p��>n1U+^���3�V�3�V���v���[v2�+TB�s"1���W�o��(xp�:�#�-U<�n�ҳw1������ ࠻�^�qvR�Ѕb��*�*R<x�f('�JGm׫���\��`���4�i�4ְzU�^��8��驯 	����;��Y�����z�X�!��8[9����č�ڍ���t/tv;�2,IW1y���kK��,W�;B�+@f�'��i��K�D����b덪�
�Zlu���@q8��Jo���J��8`��iפC���� x�WA����N���/5k(�,i�+����w_�������ɟ��61��c{�v�������O>�B �2h��@���<}B���9�w��r�|x��4+w� x�M�E�F2@�WL~���7��;���o��I˭�i��k̟�xE���g�����0��x��g?���o�8��!� XC�Mv��k����2�5eL
Υ+�zm�l��L� �0n�k'&_r!^�]vEPAlS�V	���ݴ�Pmaꈈ�P?��B.�wl_(d	��[�?%a��'R)��<v�v�-䭮w���3U�M{G-g�ʒ!�͡�=��T�dH�i�x����R�`a~@Y��sS�i����V)�R0�L2��	�l�V+拂���[:�R�`��ƤS��J�5Pp|�;{ r�T�c�aQF_D�bU����'�e(��R�ou��h,���-^}��Z.��w�h@i�N(wpBJ�9?�*@�����%�9F�b)=~������'�0���I�f�:���9��q��3
d�+�T�Y�u�¢`[�i��pɷ�\A},�eMk��k� D�K�5(�F@d��z�N4Д��D�n<.(7Sֹ�?���`ä�$�~b�� ��������4���}�^�!�X�;�v_1�Bl�;}PM	��C�=i��8Y񝯸�,�hj��ȇ�o�i7��<��~.�����Lg���\���b���~�tGl���� �܄�a%h��ER��'Yz��}�L"��rऄ�1Ԉ�61_u�'���M�P�I�*kl�EC����ߥ:9���s�_��Ni�!���3��!!������$���<k��HFF��-�������dL�F�y�;�4�,z����xnC��`}�E���z�v}�xm��G�~���N�[�ӳ��$/��4�3��4Ln�1�=��cu���vy׮�$�ll6�fx�	7���֖n�8N��E��?�3�I��������pz�Q�X�g���Řv��K�F��1楰׵Z/ �,ew�f��w%/A��-�b�P)j��t��E���jY�+\�=��؃X��B�m����iW3mS���� `'k�-B��k�*ĥ��LkC�#�ђ,U�9/�%���tm`no����-{I���ێ��R^w�޲7���y��ł�j̾��_q���]����n$��_�6d�	t$h�oj���[��r����b��{s�?�i:�qƭT���h+x�i7���rҁ���`��H3N�)mN�Y隧����۷ggg�KȍF̡�MԎpS�9�<�eH��q͟	�<W���������f��sn�w��v.݄����Y�5���cK(8I�F��!1)�Y�Zsd�l|���[�/�6�EKoЂ.��#$5I�)f����rdLƉYk�D���������)�]�q}|t|x����1��ݿ��Ǐ~���_�(cb�H7�8�8\��ӖT�f�­�0tL���D;yA�@o��?oW�ô�Y��kX��h��߀l8��H4�t�������f���5�i��a��u7�(�Cs1s�c�I!)D��4��Z,f�׷d."& R��y�I���\ P���fY�T���zMڹ����H���#��������{���5���/_��8�|N�b1���*q�E#E��=���/���K�t^��4|nf������4	PD�(�#qB��=��jչ�T�e�����pF��v���Pݤ�+`Y�H�?�aAKD��'��9���ם4�A��i0<�ŀ��7���)����p@R�}Hv��W�����"�B#�%/l�[�h6n�x&�s����d!}���q���$3�����������M#?�
rX������~t(~d�ob7�v�lV�A2�B�R�Q�]]	�X�Ɇ�*LA���ւ���륁[��E+����W�F�p���O�tN��1��D%�&^P�j8�"h*B�"��Y�H ��a$���xt�I�{�[�@�v�E�pfZ�6�Y`�Eey#o�O{vLN�لM�*[�2%��룕`�.�@�6�On�٤�����\8oQ~�/�d��x��\�����E�[��C���6Oy�|ǯ�H�Ơ��S��������CO$#o�4�}�Y_\�&H$߮no~��:�����f�ru��\�bӋ��/�KDL�IQa�#�mpYM��NƋw�8X3�LsǇ���?~L_!�͡�A�U��i����������ϗ�l���>a5Dl���_���y���ɓ���>	�T�<���8��ef�'YN,�_H�O"�$\zKrR|���Q�ooWmpJ���'A��${��ɿ����=�5�"�V+��1�4��ԎO g@n�MW``S��Fõ$�����l�@�j��9�&�)�,�c���A� �v�ua�i�2t�q"l4>f����Zk�A�y��N{%%�l3�G�9+v�9������͉�Y��xD<���zwB��6�hD�����}}0B"�>"�0��f�G�0��$-�Ț�����VW��l�lM��d��{��A~��q�%`=�&N}�s�ݵ�3K_��LQ� �5��,No�4NdذΠ���H�fz��U"K�,J$	�-��/���DG��E�q�^����߈|��95,�m������)�oJPdlg���U�����ʞDϱ�S�:+au|vZ������P-@f���7�eH�ڸ��C'��
3�+�_U�Z8�ǞB��b,�8���>1��T���`Uޥ�K�;�4Wt�Q{�ʨq;n>A�,���w��̰�~��IT۴��83E]�-�1q�NO}��)�
��D`\f��{v���X"O̰��{�b�,���b�C�����fV)��[�]��.���\�>ⴴJ�k��4d�c�O��jYhs�Q�	8Sb�T_�@�03m�����
��ݳ
/F\�f����pw��l�Y�ZCjg�J�2i�_���r"5���S̑��qze������-V�p>�Θٵ��	�9H�ghp�$�k���/�(a��B��#d��b�'�jk�쯘[*��[����vRB����O�f@Ç�*���߂��f|R�Q��;3C[eϴ(�����M6��
=���k�>e�j�.���w��������'��m[��Y��^i#h������}	yw�����1�*���"�3�C s�Z����e":�yq��g�{s-�p3�9E|��;�&z���fFa�#��_l�4����]^\!P"'���ݬ���zh�J�Mk�ͦS�Y0;�8ad)0A�Qq�:�9b���sb�\_��p �]厜ޟ��É��(�o��>;;�Y=�:�*T����ޣK��H���F�:qkB7J��X��^}-�}�]�?!��
lct���rA�r�_w�s����࢓~yuMZ�<����8��{��sVf>��o�"W�J�ޅ���Q�Ν���{~�
W�����N��mP9�8��X8����������`a�r����r��B�R��l!]�/� m��J(	h1K&�#BM_�}$ڧ�U��sz|��_�]h6Ȗm�eO����'iI}�u�G�76��99�tK����N �	�� ��F
�
|���
� �k���g�B)!�Q�;99�ɄW�ъ����326!���A�)�I��͝K�y�;���֝���T��T@@�W��m��Yy���P�
P?#ܰ��� ��a��!�,-�8��1qm#ԙq�UZt(�ϡ��ɜ:�4\Mg2���^xzҀxnڹ�jV���fC~����T6
s���=�����"<��r
 �G&��6j4����Ł���SL��0U�I�Φ��*5
�.gq�j�mǺ��|���mϴMof�Y�SE2hQ$���[�/��Z�
!�┷ȬV��^��*U m_1Ŧ���J��A���6�r�}�&�+��Q��վf�f��֖���xu���sqV:6t벹Mw�~�����r�ߙ�Q9.�֒�*�a;mR��6���]��&f�ڔ"'a��Nw��q���vΩ���B�􁯿��y���Oim1�R�yCڏ����S.I�O�\�̰��B�4m�8�f�8O���$�5�V'�3R���&wv6�ܼ������9����s�+f�����곏?a���ϟϚ��k�2�F�FАDD�%h�oԔ06�0��ͩȴI+�C�?��|�	ߝ��?��?r��!%"Tz��j#�.�=�{{G"���f/fiu$o"�5B�L��I4����@�w#,W�\��0���ش#��LJ��+����氌��bL�����%݇P��$c��ĩ��:�TL�\,X�,3U�Jf�-��}`�m7����-Jqa!?�;S�1��$"k����1ڷ�^:�(�J�F�̡��Ĉ�n_�I*W��� ��|�
�x�ٜ`�ɿ�����,�A�|���0L������wg�h40T�����>��{��n�[��^�z��h�G�?|�P��Ć���S�)���%b�o��DҦ&jD�����S��N��fΗ�L> �5�O֢���_h��0��APt��b;�S1^ѣ�UM�$�񙐱�F-d�
6��4��+��i�ǔ��@�!��4ٟ�f��Ժ�UE���]�����7G(�;�b��ϊ3��.^ic�����p_c�'��ؗ�뗦E�\��a��{��04d�
I�p��C컆Әɑ�i܌|9�ZiU��8�s��!0~������}7�}�}{�� ��B7p��Zf����l�����ܕ;+%��~^(D�f�`ܮ�ԏg��b�tU*�*���vI ���`�-آh���v��̖<*�M���.�d⾮�Q's����w�:*�:򙮩��m�쿸˖�R����`Y��1�ńo��N=I�3њ�#����ظ_�]�\�L$I�Bsm�"D��;�`�%q����������d$�EHJ�Y��R.�{���~����J*4�<Yd�,�=�?�شΤ-��+��G�Ѭ��%�E�6�Gmr'�l�~j�ڀƪ�ǥ0vתBZ�P��v5�DM��<K�v!c�K{���.�>Q���/�}s�U��쨳�e1͙�W�邰�������;�;�N��2�2�,��Xj�[���0���3Cls�puq>����[����n֣��LW�rϮ���iX����
^,u+s����[��޾دn���ş�CC�S��L 7�p�����_\\��')|�i��?<<�$9?,�5�qOW����Z���w>/L�d�
n����\{�����6Ee4�s�YR^X2��%�eTWE��҆b�8.�Y�-�a�����jHJ��h�����R��C�b��<�!�)ng�c�*c�w:/>mWW\:�Q9E�(�����C���{�����5q�b�_�[���=<�sNn���߽����O�����䐒F��#�$����\Ҙd�d)6/���=7d�^^���o�G������'H*r�k6OOO?�쳏?��΂�//��,�Ƒ�(�)-$7�
�%n�-�I�*2~`�n$�6��_�0�����~^��?��_t��@�]�)����}�ч�4te���ʨ89<DA�M�;���������,����v��$$����V�$���m߫+)j��#��`���q��$�LA��|N��T��	��VD���������<d_\�Y� }����J��\pU,{%��Τ�7��kYh�����OS*��%lP���v��jq�	&�GeF+��M$7�MЄ�a������-�)�͆��5	͑�,��,� ��Y�V�j\	m.ga��!�e1��&�6﹞� �=��g�A��������w�co<��L����$��K���'C�<�5�pF��:HK�7�Y���U�����A���ّ �i<���tb�a�=u
�k�����U��J'+S��\u�2��r��b�,��*(��N��4nL�����[�i	�:%�������GC���OJ�_Ӡ���(Z��A�cE�B�]��捼�R!�.>�e�ހe>�rv��T����.��
�:��mYV�1���q�L��%�xR�Ҷ�WT�� �rlWÏJ��z�F�5�&�Xۍ6p;�Je�`W��>��vT�����5�M�c�y0��?#j�ܭ��8qv�aL����MU��i���ᰠ����o��;���B�)�ʯV7QP8I���'���]d�w-G���V+9:�H�U�'6c���Тߧ�]��{w%�r�;:;e��]�?_��9L\ 9��Ǜ�|~~9I?��ەH�w,�/�~>�ٛW/�����s ���V��v"�uF���I��H��B�<����`��]Ŧ�m�<5-�z=�������۟����.�飏>�����@z��˗�,�h?::�����+�U��ڪF�kf�d�LNC�V�$vH��e��;
#,�eC(K?�h�ң��I_N�	�GL��¤/z�< ��,�-Up;~�2Q$[��u��A%Yl�Nf �k�iִv]�'anO�T@�=7��F�]mљF�6����ö+y&�������,H~΄�|��}�u�aD4���o%4�Sfľ�3�a� �&L�z��MPJ }h��V ���W��j�q6�+<&b���XV��!��Z#Kp�s��9����{��2����t�ȼ�'�u�>=���>@r���G�!3���0��{Ǩm?t��_��f��������_+��za_�Yՙ��y�N�]朲z���)2�S�$1#'.��6�]l���}�kr�x��k�*��g���ߝ�_�wX��(�+&��i���Bx!W��m��*�h��6*L�eͱ�f�-}�+�8���pU(Жlʱ>�!�N��W�!����U�!Y؂��vQ�R;CʎѰ�i���|���!l��^J+���W�t��ꇔ�2���F����>�E��t�4�YS�F�.��ovAnc?A�	B�+�b��\��6jQ@�E^�H���A,dI_$��٫�6�bѿŞs���r�%GQ	��0*�b�$!%�y�K`���T2��~CY��x�崸�C�X��pG]F�6@ � Ms,RJ���m��5s�)�&'��{2l�m�(�e5�i�n��nC�sK�����ϟ���?�+����}�r�[��	B�BG1�������D�L5d4Cr�p��}/�a4�Ǐ?��O�0
��-]��LNJ��i�$����z�%��I,��d;�r�*̬��am6�Ֆ6),���e�����Ǳ������C���"�ar�2â���n>�������٠��V<j^�@������߿���=�L~��������5��-��@�%I��_׷ܪ24���u�ѣ�I�k�1ώ+F�H�B��i���u��6]��4�r��đ*����/�0�mp�\4JF�`��+֜h>sK������ׯ�77+���^Q�Pa��|Vi�lA[�'�03��(<�!~�y��"G��i,"R� ���_�zEF��@�������\j�#�/;��q�7� �^�0
�[�6s8 ����-�5>d	3� m��i�����4r2�� �^4o[튘}ci��t$I,�c,]��j����<h��17+Q����g�t�V[LB��G:g=J�>�T��uQ<�G�YJ� sz��3ԡ��.I˝F���9C����v�րCbna���Ń9�9|��A(���EӜ��i��~wI�>wh-B�v'��L�ڨ�&dZ�H}p�v÷F��I���-���(���� � z1ӽF�Jl�Xݼ�(P�V+DOM����B�7t�jD
I��T#:��n7�(���P�n�K}�i�h=3p!���&��C�y�D5CЊ'���x�l����U30]a��{.�kp�yA{�C`��ڭgך�4:;�KpmQ~(w)"�-�����'�&'����31�e�v԰�,b�U@�>�pMG�͠�$�>��u/�_++��H ��A���� ��Z9��Ulx�]�]�����#wf�-�2CKBh$��o*�<� �8�=&ܢ�=4�l�#�{�1��7�x�:2eᆤ�Q\�N�YA	%����k?�iN��P�\�۾��nS��.���t�n��L��lb-`g>��݇'��M�����, ��n����j�@��IaD6]�%�y�HF�;�b"0�����1/�R�n[�Fo[���1
��Ą����$G�IΩ��t��q%���̓��Ӎ�}�ߏ�z��z�6R�Awdp�'W��$���)	��f˖X��E�-����L8dE�M�F�{��Jc@��xdV�_���[J5%�H�@���W�X����[<��Н	!�������DJ�m�f��=���\�r�ƣ���_��WM��G}D3��L���@M�����l�l���i�H���l1�U���n�*C���ن�L u,�"}PzRӴ�H�����D��6k�\�V0E�؂��@I{��9%���a�Oz�9�D�&��/�E�E��L�@?��Ű�����ʈS.'ށ��/f*���fph��\Ҟ��$��+��狤�+�&�)`A k�2�v���!:i�bL�Fa��ae�5�;�R<;V��-��ƶ��^��a<;A\ҍh��60��z(@%!��+a�����W�LL!M)I�.�ئ�wvv�$17m�'y�!RD~HB	P��
��ˎ*�q���V�vrZ2�
2ԇWֈ\���6��߆Ʈ�*wtJ����'j7*��N���ʚ)q�߷ݢ�݅�*ȕ��\��gBU	�u���P�E��m�+f	W������)�62�����X����*t!>+ȿY�A�/�$_�L|��1F���5_�i+N�6�^���a�������ӗ{{'M;�C��c���۸���9������/ٙi�ї���W�s3��m�ہ��:<yM
�T>�iҬx�P���۾--��$g��ɷ��{ND7�]7����t�!��1�(� p��Hv��A�!O��:������>y��v˭*=M�Hg/���"��&�DJ�U�4xq2�S����+�0��mpF�`�7;*�cY�'-j�c�+��Y3h�aϔ�r���}�>����,�d�X ��^��W��8����_����F7�U�C̏�"55 i�����F�����̦���T�Ȓ��^#a�߂Xp;�E���%�pvv�]��z�����E��H\�ߣ�DS5�C2JJS�	t���*)�B���|�� ��L�/�{*�Y�;�l��b�Ra�,N�tx�ĝ��82R�t�H�ܱ �Lj�Kj�������}Lo���Q�墳�әx�����i��������;�3�U���/���&=~��DW�lV#��iE�A��)�����ENg)�GF��R��:��7g���/����q�1�T^��@k��X�=�1��p�GK2��!!#����$��aI�^i�q$ �qؤ�Tl�w��\��f�}���D�B(�t�B���4���\�Fd�������Z�-
7�z��th��q�[.�����c�n�99aƖ��+������Jq7��0l���e%��}��M`�o��ݿd�L01��(��泰\�=qG2o�룃u���rⴛA�rD5��N�m���Lf�N�$����"*�AT�`�e��*Dn���]����N��7����3�o��<S&���]֓Bkq�B�c�e��.�m�}h�aJdܭ6��f��x����Ҙ��g৿��!ϐ�:/�
P��4@��
=y�b���Ōf���ˋ��톍o:q��@��-@O���3��٬��M��h��8���&��gϿ�ޔ�'�a�e����.�z:�w����ia����{ޓ��`o���B�����In�ig˛�\��y
yE*,��7��Cbπ�	��Fhd�&	�"�v�&�9�B���t�����#�O7��{�l��5��+	�C�7��J`��O��.~}�a֫����n������˜�Ƹ���zѳIv��oo�d�pԸa�վ��܃���T�f;J*.	�(
|�G��e^6- ��I˿Yբ9���o�fQs����U��S�t��
���L��� ��rؙj�ǰ�-,���
�������-��y��./���j ��#N�T]�{Ek4����T�'�����mF/���1���I���5J�~N��7�b��2�c��Y�523
5mC��V�����'�FA^5[���I�,�\q#=Y#3�Lv�1�}����az�Jo{s��]�� 4&^K&�b�p��sw+�,~j��ҵ�ÏӐP�^6�[�EdvO:Mh�Z-��ko�4��S_(���e��i®��R�3M!��;�W�7�^.���Kf����~����s��v� �	d)mp�����~RGG��-ǌHs���J�V��b6?b;s88Ib�pT.�i�oh��ł�X4���^�x�I#M<O�^t�zsv�e^��'r�v�������;6h���O>���6q��A&�Vr,�%`潁{�ư�'����X�>���یC�xY >)�����}������!����n���K�����D��Kf�x��}�}�K��X��b�
����B&�+ܟd���u*��قlNV��h�ׯ_#x:h|����wd��A�D�[N�ƈg8��д�ާ�ğ�� �2�{��z'�	�%&�1$��F���	��.��!,�"T�2)@�
x"���>v���^[�g�:⾙ͥ/���qxk�l�����@`�"��p��4�^K�m"�#��5b������h�As�deWr��1p���(�z�3�7Z HI��<��p<A^�
��s}}:Wal�����Z%?E����I��
������#��>e���Y\�]�^\\н�	��Xs�f\����`C�3�&�<�)�V��)o ¤�2�@���KQa����im0���6Jpԇ�M^O�j̒j�JLq��7�n�XxU�r�P���m���q�"�ck�Jb��,���	ayb�foX��X��"R�D졼�O&���h'�m\��J�q�W�p�A�V���B�=d;'�ﰈm���w�Gܝ��LT�΍pm
�uo��L�pzz�6���۷o����Š3}rrB*�t���o�m�b~�4 ���1DI�[F1	��I��b٠_��"ዹ��ƃuZ�a����YWN�IN��LɒcVrP�RY;]ҷh,;D��.
�%�޾yA??xt�5Jr���Z"~g'�U��(<>Ԃ��:v����I�&��. W���:�8U��I1�����N٦�ֱfk�^���]¶-�*InXN<�W��j��OFm�@A�&�����Z�,"���$ۏs��p�����]�Ŗ_vH�������a|�^���2��V��g�H���6��H��!1ik�u�~�BN01S��2:iǶ�S���X.;Mų��&Z��]!�bZ�>�*�q<Ѡ�U1
��O��Q� �C*]WJW&���tLh��?���Khķo/h,bq��F�V���;=�<z�t1��˅<�Ǉ��?rZ�:_� j������}=ﱵ�ۧQh�Em�$�7O߉��xʻV�&�-6=# ���M~� i�^(�yy]�ZI0"��H"�g���1�Ĥ��Y+a�8ul�.��5�exm�g��**_���A�y���@�F�0�>0��2���
6��FQ�d=;����T��2��D�E�L�f�>�x/���
�U�66`�LgI:'"���*�������Ǭ7{�F�oP�9��4�`���4Ϟ=#7�i���~[�"�
���c��R����-=CާEoCi[
v������?M�ӧO��Ы�n��p%dn��C։��!�5k��(͍ ��p���yW���!�h�ڐtҪ�V��0;Q�H�`ǉ��A��a ��� �����߿~~���l�F��A��*'!�������B�C\s4���> �����{mf%v�=�i�"�3CmV�t��`.�l�P�-��n��к��X-fM�^�1	n�MR��w<�����Ym�.���IgR�e��jpHk�:8� qh��{�NNNQr������Kl-V��EF
n�<x��E��B�]��J̒��z5�L]�vʄ�BȚ�,��Y	ݚ�c�������6Κnt`�J>���+(�k�S�h}�=c23'L��*ZL#�m$lNQ&%�2� �;��!��DvR4�T�P1���(����&[�v0��L��nge�6�Wn�2~��\��8w��x�:��*�g;ܔ����d2� �M�%��R+@	b
��TAH��"����2)hӹ0�BW�l��h4�5ʙ��6`Jh��jW:/��/��"n����_��OaZ@E�1)���I����!�]�.X_=�!�|+��}����K$����
���N?�����+�px⒤2�?�6�A�氎ܫ��yQ��sǼ5��QP��(���&��_~�����=F��Y����OZ�$fڮb��CH� ?�i����6(����"͛��d���u�ٚ��~@-�M���QP�7+�iRn%>;ʈg�I�xŒ�`ڈ+��w��$�`��j�� #�k��A�glE��W�áXM'M4Δ��ژ�a�g��+7��S�R�0��{�'w�Gj�b�6%���P�@O��trr��}7(q��H��:������bY��k���p<���1��:�!�{}��%!ڮ���cc�|�R��Ӿڬ!��R	a
��SЂ�ӂ�W�������A�r�U�9��cɜ����֙�٫PKᵑ���ƍ�3.yG9����n���T��mߚH7UX�H�,��cƠ��I��r1t~?iٲmې�fCM)��+0�]k�I�����_���>Hl�N9�ZE&��|!Ue��j�\+�z*mKe�Ӡ����.���[�%4% (��]�0�4�R�#��1�R-�s^*+]�Y��4��{=�[q���o���f=�lW��c�º����� 6{a��2_�8)@WFON{zs���c���tu�V���t�3]ͱ��䖙گ��U����θ�3�T�c���� �@$O�T���RR(�⎥�|�T:C����ӻ����	��� ꯆ�$��Y�Mf��B���M\�MD��2N9�ϐі,Ad�\��mjQv�RA+!z:�7����aa�\�M��Pu ��Ѡ6N�<l��U��v�2�+(��|H 2�pXA��[1�H�0�G�C�R'a���T-��8�d��j�GU| f^b20sy�6�Òu>`��9���l����wK�A�`C�98T���|q��<���9uwML�Z�!1�1����}3�te:�&w6�� ��1�sJ�#
Nj&��riX`�A�Tl�ĥdWo��⧇KI}] ��z��"�/�]ȫŢ!G��������)�/��K,�t��F^�#�X$��7vS �$v��Q/�v}#���q)rew�BwH&�xلI��ْ�]z5�LC0�p(~d#D70����e�� ��^��NfCP̑^k+��k6�a����c���_���ǈI?um'ջ|�H��TjRR���d�0���)C#��ڤ�O� ��t�5�[��1׺)]�J����Yi��0d���ޢE>�Yf:��L�5�3y@1R�v�0N$���_��|H�Ӣ���[�0�߮�6eF̘�HK�@��-m���������w�7k���󛳳w��״V����v$���x#�c��IMޑm�o ܆-M�Mo��Ȼ�Y�`�|���ӧO�V�鼦%�:�P���  �eB��~��������-�H�Hi��x�ֱ�YOǄ_[i���ɓ��XsfӒg�n����M`�vl���+ro��[z���pG+,�� �h��d�ѹ����X�?,S�0���^s�"��_��DX�ӲJ��v �L� �a43�������Ç?~��&��47�Հ���읞>@ؑiLƩ���f,�g�kY@<x��ѻw�g�U�f���aO�E�i���r@��P�.ab�nnQ�eQ~Z��:IVÓ�lTR)z��#%ha���sޏl����[Z���I|j&2��Y'j�l�0��� c�9����~�8���#��F�o��{L���[q�|���`�J��$'���~��٩am��we������lG�-���d$���{�m��b��S���O��L?�0�2�*�1i�B8y	��|���T`��=��1�&��D��9Q�J�z��+Y�N�dA3�fny�[�Z��V�N�f��<�JZ�:)�,� ��0#-V�w�	��"f�d;;s]�$��(�J��ʅ�X�,8�<��y��Y4sDf�~̍���
�lM��'��$yG,=��u���8eH�v�ڢt��D�,�ܘ��Z�8��,y[����-�D�J��r9Nc�Q���� ��2������@3��C�e{���W��������������������Vzv�Y���?&�F2���Ž{�Hp��_�|��7ߠF�$�d�n��������?��|δ�H���W��K�?��d�g_|No�ؐ ���p,�ŋW���3���g�Ϟ=#+����ۂaې��I�.v���g��0��W���/?��Ã��G| p:��4��&n4'4���K�h�'7�Xv]'����.�Ǥi����G�x����	�����-ggoil��h�
���U*�2>��a�\X�!��R�t��0���B@X\���[Yw`����!����GY���V�Y���ΚY�1Ǜdw��)��lRD1`�ܶ�Uw��)�f� ��#{K�1	$�5��A%��I)$�e�������X�0&Yr^!a���g��b��V(#v�o�BUJJ!Zi������p���.S:Q�$�	L*��n� �zW�z'lT���6J8���1���^ؙ��!~.bn���Cu�K���E-X���p�-����s�2����?��;՜Q'��bT�j� Ԥ����p��ܤ�K�*��S$��L2���.[�*n4w�B$T'��LWZ��$yT�e�ZeZ���jz;�^i���[M�ڕgJ*�i�� �;I�\�
S�f�`�B����)�5X���lHA���nj$k0�B���,��UOd��]�&k��%�5-T�"a�L�0��^�P�!��$3��/q�ԛ�}>��0l�s��w2��5���A�&��Rn�jCo"I�n�I���g�S3ũ��4U`F:9�B��ۂ;+�h�U(RȮ+���P���ǘ���j���$i	IT���X�l��������Ҳd��e��'��ol�w�t���W����sb+�b�zga�P��Ò�H��j���V�s͖M;,a)Á4:�3��J&������n-3?���ӛ�9b����4��B%;+��\��uHQ_��DO$m=�E�{��tr(�NM��Xy�J�`[Ԯ�.  ���T\:���a.d�^y����fT*+��.S���ϻZ�ZN�i�����|��IZ��s6������#��<����L�@)�=F�g��Ţ$�:�+I�����vuCJ���i\��* �999����w]�{:/''ǢE�8縫'��#Ѓ�*�9N�vJ�\���^ ��2�}?S�3{x�Ѣ�EA(=a&zş�hs��"���ٵŘ����� �W��@!s����d�
Ah[�P���]T#���A�N�c���^h��y����y���Z�ח˄��� $Z��}�MH�@�&�{7e���䑄l�=�5")v(i��G��N|�$�n�uLgw[־`r��R_�rF,l��)���R�3B�'���^˱\:JӋ�p��T�F�,9�xyyCw�������3����4�	����9�V[��	�lV�O�F���bF�5���3r��kv�A��)�X�B��E1H�`�10?�,:b��Iz^����9"?�I�D$�� ���1v��n��8�krq�3䵾x�"U�%`�[3�\��� !�p4�܌ra��jy��7��x
��ctNi�p�,5�����㥡E7*���I�ל6,H�B8���`��EM�F�¢���H9*� �)r���Y�U�Z>"Y[�Y��|x�p/�?b�n���%�SLn�|�K���f���i.o.���[L-o?wЭ^�/�u��{���l���x;�9�>����m/�i�ľf�xMab����74���-=���L���Ҍ`�7U����'�K��%�Mt���'U/�E-���0/R+T������N-~A�v 𦀣�^V�YV�f�-�V�Z0�U����5��P���*�]5Zlk>�S�Y���߂�f�alN=FW1"i���P�&�zanM��	�."PpY�0fB��$Vb�iL�Q�I9�@�`��Q�b9Qi㹵f��*k�J�KPx@IXaU.�K`Qde����1�ŧ��G?���_>���w�?��?���oix}�����駟~����������S��{���>�ÿ����'%Bx�	�#��_����R��~��?��?}��5}��M�\��SPO�<U7OZ��w�|syy����Aٻ�yᇋ��[,�\.��N��v$��Pϴ����G��c�3�6kҮ�_Z��:a��$3�&���&a�����9�p���V�у��z�%^+�<��.gKp�ai����HOc�&��4�Tv�ap'L+2'K���lTdq��x�R���s6�,��NǌC��Ө�^�X��0sTzCO��O%�u&V(W��w��"�C��Q$���j{�)��+��E:��NG�B{�F���-<]�Je3�I��) UD�����9�4Rd�W<"��������X��H�Z|Ќ1��Y����:q�q�oߦqC%�*�(��R4 v�a�Y�L�$��f�	$����� i�=it �J8����O��a\?+��T;�mk�=������<�u�z*�m��L��+���+0��X��8M�T�v.4%zS�bNG�;�tw1��	*~�������H�w$� �_�$�~�J�j8�X��N��8U�G0š��ʹl��WBt�U��V��H���e$޵����ɔ�^�'���Bzz0�J{w=q$���m�o�񞱡I�ft��fz����5��n1g���e N,�Y[�9�rN��dv�:#��&]�J��|�Q��Ƞ_]�7#�[W��o��j��Y�u�0/�32?zњ��DZ�Qb�����nc ��@#hh���|lն(�ԁӥA��)����/��-���/�~&q<r��#f��u}���~�n�l&�IJW�jq�E�DX-�--Y��I��f�YH��ZG��Wbl�����`C?�u���;L"����q��<i?83��R��#	J�>����F,f��=|�&Y����z�
0�	[0-t*���^�E9(]��f�|Ֆ
rb}�$�㽢 �u�S��)����JdMݳ� �,�)h�4sý�e���qT���R}エ3:}i6�M
CC�'
��]�N�� �оN��a$e/v˻�f��3���]�{���k*�e������d��	K?��]J{��T�����ѩ���8�Il�شnPg�ʋ��k	��P��CְYwm�M�ڐ���͖VyM6"�t`��J%D�{�Z(E��lLh6Z����[�������=1M��T�C��0E�r�2m��!����v��[B��B���$���� zV�G�d���p�㆘Ț����޽#W�p��̬��ȸDe�������ك�[���3X�L�q��`;��m��%ᧇqVȿH��ż���\�� !�:���5>9z��tdV������95��%Am�c����0'��iI\b��KQ<K��ᖮao*���Re��mI!�P���t�i܌�6�'0�$�f�EveRm[��Ƣt�%�N8 IS��lu�Uҍ�fF�`Ϝ�D۹��Й��Jp�888�3�hd��p�JK-�����D��ƽ��[�X!AH�4n�p'�I+�n�Ѡ��,H++K�M�e�R�ʮ5�r�`��U,*X��t0l\%��`4��M����Z��3������v޹n��y`	� ���Q�k�V/����վ�I��=zD�'����Wm������@��xQ��8�Y�����rИ�����'�@;A��sҹ���p<'1�b�BA�ws�lPZ>��!�&����.��,����M��9W�������$�ꚜ.��\,8}��5�g�����[�I�̠�����8A{�dHm�c�E0�PW*����B6�K�J��*kF�'	���v3�b�A�$���2��(�]��R�YD#�, �EG�|$LӪ�MU�Βdc1�5XЉ�i�Ff6�=TD ����5�u'p`I����I�:Z��)Dv��t�z�����'e�;�W�F��'\���]Υ�F �s6��E�����9f���K�)*��F��_�>ʊ�����͚$K�s���efe�^��t�, 	ý2�(]�b�Ie҃L�Ɵ�>�M4�� \���\��`轻���\ω���5 H��J�Y��ĉ���?��Md-�yxMB:�D�C�F0n�I3:���"�N�y�͆�+��-��0�Wꌪ���ū��-��r����~���MQ�\i}�N"ň��Ω--�m�����(G9��F߈x�Kي�B����	O�����|�Ϟ��������*���o����1�bwoz||L��}���Ǐ��Ύ�I4!�����gϞ�����O������'O8v&���[���'�ʀv����/_NwgH�Q���DN���|��i��D������m���Hd��6�<8/S�1	�&��֜�`��駟޼�Y�ׯ�NO_�����WZ��8f��!m�X�X��y��E��̅�O1na�".Vk�A��ԟy1�Mhh����:�� )�e���/JJ�*���디� (�x��s�Cd69���d$�\���A�H��X�I�h?O��4�J���P���+���G��J�^#�ٍEϔ,dK�v$���I ��t�5=i��\)�{xx SGc�J��UX���#�j��n������8��J��痈t'�zi��âS����F�pg�����A�56	�B���M�5���h�%�/0_�\����'��N������X���5�f)���B��%F�˥u���D�����'w���v2KrG9G e�Ȁ�
ڥ��5c�K��b����w-8�S��F�v
,���$<���ݧ��~yw5�3��XW �`Ж��R�$G:��ޒ����aS��1#Ҥg�쒪_�)�D���ƠB�`������Q�)�Y��st�z�A
Q�m�7��XĄC��ĤK=��k<�ݹf�h.s������q<�i���{�	�!i�:��K��h�
u�*?���ŵį*���gg�ҭ�����]�x��������NEbU�T��]G%>kMf3yz�`}�%e��T�j� 
��mK_5��U1o�)<��ܲ0�.����>"+(��TxD�I���º�t	֬)��dB�A���;B<�\S���y��[��v3V��:�����`B%Tqz�&�(wE!�x���Bh�"�)[)Jl3T�è�����J���>||F�VW�m�/���Ngl�7[F!� $���"����4��㤢W"׵��q��2����=�+�X���d��	M$1鷖J9��m�h"9P���XC�-����irIx��9G����|.��#!���<q����Π'#HM�<�{���{��[d���E&��.@d�rLG�ԧ�a��q�vw$�W�'�G���9mdA۪H1!��~Z|����w�]�B�U'�E�Ԗ�݈;�h�Y$	!�("n ��s�/F � ȐA!ߵ�C�Zl?yhi%�]ĸq��D�Sn�魢�hG��[s^�D�����X^������o���~[�f׮߼yM]c�gG&09Դ��L���CuF�v���mQczZ��ڢ�3���`1�8���x��%�ɘ�[_�|e`U�W���~%ߊ��	1ٳ��y財��
�����Q=�k�6§�ps���� uqT��zb�$��aC�:���Ҧ���N WO���mra�[�>t"d20��}f� �P��w�d��E^;��FK6s��S^�)ܲا/r�m���gc�Mz�V{^�/�v����tfFm-Ǔo�u�R�r>A�!; ���,FĄ}�*,��+#d^f�����\pP���	Ĕ�'��0�8�/%�؄�hB���P��^�L`Wd�&,K��>������a��AN�ԓq����ڬ��iɺˡj�[���x";|%j����l��^�$ٝ�]�߼&��/�a�����_����ݺu�OV�{u5�d��K�� J�WV/Ӊ�b��	�eP���./��8��3�6_@���j΃�\�T���N�O6ojaE�ew:�l��%���a�n3u|Q�հE=�	�TP��E2פ��2���S+-h>�,@�҈�(Zj�ͰVj|�j1e��p&��"Il�7iB��)3 �#N�MJ�e�S̆M����J1g,�XM̕*-xgz
�ׁ:(��ٍ�-T�)3�m������pUd�MY@ޒ��������ڭ���c�71o!f�%�����(�+{��l+:���)D4�JNol������`Ȭ�­�`%=&�k��@�E!�#��IW�O�>�{�.}�޽{	�e2�jv��`	K&�جmK �r||�_h�9tgv�퀷"��o��5h�D��,6h�A_'{ZL�皯IVxK���g�qU�l��g��}��Q�c�8�cd[��;}�j#�&5vXB�2e~	�Cщ{�\�t_�U�\�+%�/?<u��3�=<>�X������w��΍v^~�4 k�`�:u�E�뇵�	��̬44I�#�}$e��Πe���7)])�Y�N�^y,()4Mh�/D�!%�4��I	<ݐ��8�<��F�x�-�A��o��k����Z�X����6���qZ//s���D�t�H�Y�˜xS�^�j�c%�N�H:#���S�|wЕL7aB�8��,����B�T��������^&9������7-��i�5�J)�pX����c>Z%�-K��54�H=BUՊ���O�5�k�E��V7���EKL��ضM�l�z�w4�������m�mm�t�Yj�*�Z����:ZS��D�m7�^{0�Lp����ZE`Fk�d#�T���$�:Ґ3�r�¦�L&⛘)�4��r�+�=�&kf"���&Z��qq��M�7ֲc� 	 ��r�MpӐ��~�����]�,n�n�LvX�����I��<=gP�y �>���)ӑ��%'�57kl���z��R?I�@P� �ӘR��Ú��i*Xo���hK����`X�����tq��*~��r�ڟl�ʤ�&�c[K��J63[3� �Ȕ38�iO~�\�$�yf��E�%��L��m+%��������Q�-|6���J�}��
�Lߠm�Dal��8*���S��NrU������U��J#5��PT���th�'Dj��^�
,�h�J��� �Z�t�I��bQ��dƂe��~��\�J�Hm�=-��5��k��bR`	lۜo7�	6�F&qx6I8*Ҷ-5D<���L�H�(l��+Ѱ�l��ڂprX3s0nb�jσ'�t|�ߵ����kǻ7����ΘWTJҦR@�4������M͡"�_�xpݥ�(�G�W��/JE�׈��ڽ��ÚD���C����h�L�:� ׵�0��~�ڢ~�oq��3���� �:�|EP	D*����@O�&ۚzۜ��$k㭷ޢa��b�;bp��Xzs���j������t���,�,�Ѵ y��Q�zň�20��_�C8�_s)�n���\�$�O'�![9mW%nǇ7qC�z�˦޸i<����$(^I��Lj���ts����F�]/y�I]����YJ��9<���)e,����+/��W��������KOa�댧�[�Ú+>�N �	Û�����8��f�%i��xy�5��l~)*\*��D�~
�=�D��t<�������D?�Z�(Cs$r� �Ѹ���$��\�vrpp Y*�%�s:t��jk��1P�y`{.#���-�C4�FEw��=�NFX�kD��l�8
�iW��5��9���D8���|�E�|I˶�^�y4ۑ6s%;	²琫�4�@�+`�,�wQ�9[dŪm���t5zLKJFJ8(S�$��=H�_�䑅Qa���./Mݑ`���_k70�����53l��#!鎎n\?�b1�۠kj���G�~���h��\�~��ˋ�W�^���X�_Ӷ�u�d�J��B;�0����ǧ�紑8�_{�cA=a�鴴�Ѿ�_􂓜����1M��L�c�,c�'8 �X���w�͏f�='fbf5R�sZScN��"W>e����ik3O]�v�͔�@��U���PLRA��[`��7�����>w_m��Dw��1'|("q� Q���	I\�[�V�
�915��H+"q�o��!�3Y�8y_(���M�"I1����JaA4�H�D��8�����L8�/.BJ��Ń���D��>��ֵ����ۺ^�6�%��q[�����s����ޥ�r IJ/���m�f8k�d;
&q���4�?��Ͼ���_�~���"\��j��l�0��Mv4��Z�)}����}`2T�vfY���톻���L�f�$\B�k
����ZhaD�3��b�
�99�X1�U�=G�f���.�����a�Z��$y�8]>����$m�7�jԍȘ�wوB �(��5"d�<���	��c��z����ٙ�����̅�3�-.�0���j��^
�C���!!L�e���Kl�'^X,:��qtt$3��#》��6ؑ�N!�ȈSJ>��j���
�"qA+�5��2��t"�R)�h*�Ԥ��Lub�!c/��?�R -�܄*��!A+�qW��J~(&Z� (<��^��6�Aٷl�?`����r��P)�#�&B#�#s�֪2�*K��\IX	���]r�ư:,O �����	�mT�h�O�<���w�ݠ5��?�+�/�.��Մ����t� �L�B\@z�YE��6'h4���,l����
;ٖ7����ŋ۷o���̦"�f*v�Wd_*0:�@�X$�<S^͜�u��>ˠ���(l2M�~�w�B�S��u+ 0k��Go�{���0/����X���(%���v�l_��g�$�Y�:���&��߇��D[�O����Uy�D��3�ڐ|���eŚ
�c�9B>d<�,��HUe;�œQ�<n'�t��t:�>0�H�[���禄l�	)�D�ɥ���,�x��ڈ-�����A����s���i�Z��A�ޣS0(��e��t�+�m�B�`�A7�}�� �4�|����0	�4�L���z�LE������c�fI`�,�_	UTZ�gxt$=zV-��jNY�j�������iu��ю6v���(89�4�]ܤ!ൖ��=ߠE���q�����b�RӅ�氵�1�P�.u�p�*�s"2i�O6��Մw������~�ޏ!�-F���+;�1V_&��CC��+ڭ��A�R6��PY#`W�Ɏ4RLܧ��zThA
3��p��Q����>WC'�� ���fa�(���������'Ւ4LL�αE��[o�:����'{�I_$���܀)�1���7wEp�.���	w�w7j��U
敥�:N��0o� ���cg�ʞvz�&ID�ª@xHTZAּ��Q��[N�ѲR�Y .3I�Mf3f��u���6t�����.�ah_��4]�<LT+|�>	��ί�ˠ}K��rLh{#����`��b ����6�r����������d��-$	9����2 ϣ�p���#��pM�^�8`Yϔ��r.2�f#�Z<Q��Vx�m�Bc�n�,�q�SL���C2��V�S<,�}�&߻�6`hك�J�V��Ha\M�a�Ѩ��lgl�靨�����jF�*臄��5`��bY�(����Ґ��\G��rZ��ZV�_șӉ����N
M2��~����4da�!��G�Z��V��WU'��Ă�ƅoŶLQ4�kKn�=�'�0kF��S�$��0ІO�3/p�}���kf6`)�2p�e�4Q#A�n�)�Œ��r{��3 �G�X*�#$6B��jkQ�z�8�m���#q�\��1N��=z��������;4������?$��)^; � �밝N��|6��j6U8:<����;7XI�9�y�ϼW3�Sy��-�����W������}�{��?�����Y��s�h>�G���{�wq�c�^5W�J���e��EQ1'"I~�.".�)��@�E�� �-^�g�ȭhƮ��/�J&"P{)G��ܛ�� мN��<�L�s�$ح�U��S~d|��\�����ԨĚaûh��4��擼�y����6*��f/7i�).��h�Ǔ�\��5A��f����ǼU��Stk���>��L5C�w~�[4�)`���k�nf�S���8;Hf���^���a��6��&t]�_4/��j� �Z zsZ���М[��1N#�������'O�|��'�V�ZX>|��)�9�ޏd-���؂��O{f&��`�0�k����J%��̽�X�.�$�ȍ����plV��#./�^c=h��0m7{�T�*.�,�s��2"�N4,�!��@����Ll��r�݂����=�1{ѐ��t><<\,VN��a�<x�������4c�|����:����A�l��T�0\!�P�k�_�>��QL�$��F*�+Cx�ߟ���]�{�L�KJo������r�	�� �Q�{a�aK�����i�%N>5�D��Z��N��6"�j$�f�S�7�OF]��Z�2?I�|�GA1x^;�&HA��s_�1��4o4*��`�8��;���Q͐�O%/��q�\
�S�� �D��͸&&��_�l"_����)��o�w�����J��[�NT�5��mn�(��H�T8E��!]F�h͇�-��L3��N���O߼9ge���nH��>|%=ܮ���|��A��]��̸��AJ���@Pv���fւ/��n��M]�6�v�����|bv-z�N�Y��!N6s��H���#'曋�06u��¾҈�SJ.hyl?���c�f��w�e�!}�Gs���Kۊ�J����6�D{�<i"�]��j�W��K�"�#ԓ)T���z��Xn�A"˓q��*�((�4/:��fQ�SdR���r0�Js�U�<s���vR6�(��H{�h4��ucZ�F{�9A��p��RBLĀ-Q�)���"MXulīQ 6|��|�6�"�w��*� �x0wף�Z���Ҍ��:lz��r����6��X!>�}jF��S9m�ÈM�@��rS��Fb����C�͒LʝI#����l�� r����Y��
��Ѷ�����PUg�B�I�����%aĆ�M�L���Q�@6��Aq"V�No+���7m2A�C`��r��5��;���j�o��q-C��Z���-���1�/ˠIx�T1m�ɿ��āg Q�$�I��t�@&Q��������n7=���_�f!������!�*�k@�U��UBʠ�A���=2i�I�F��7 G��Q!Y���[��F?���wN��״���[�%��E@G���&�θ��2l�4����-��^�0�v���N��$B���q_��Z_�Ƚ�!%�7%$�u�������t6!3��Nڃ�{�&o�?���������A��L���~\M��>�ٱ���)t��.0(�E��;u���Xў�m�v��׮��M5��El��r=�UOZ���״k�je�{�<�,��в�T7�$p�M�e<���#������^�G�lz%7�1�r����%R)��H(��^#����m��вLa�c�/�] QW�� �7�O���q#5�W��|���mz>��iK�~�ȣ��)�/5Ur��m7rU��I��+Ԃ�U����%�rXv��
i�6�z�6�nh���T�V\��*[���u�&�t�6�%n�Ը4j�QW�x~����|-E7�,�h
�B� ���;������t�H���E� G�w��ͮn�n4ޡK�B+`��!��%��/h��0�w+י�%G[_�4A�*�y���HQm��d'7P�M���xҊ�B�?�i`���us&�TA=!MG�82O�M�`�C*�C�����gtVK�K,�BO������x���$8�<�#G�A��1��)Ɯ�0맕BWzN4A��a��/I������t�Ͷϸ'��/��#���z�_\�����ݴ%ȸL.���+�W9�M��<I��ʢ��LG����w}�NY�6�9�=0��92�h���9:؇F�ow�����x��!�& �������c#���-���'?��34���P"� 9�#!9�H間�2=����իWd#Ԯq�H�n�\��g��vr���߼~�-4�j��'��~���W��4o����v̌NN]e��/��TR�?k5�ԣ1ɘ��/k�Ҿ_�Iz.���@d{T��O��?��6������|u�ƍ�����_�W����dL2����w�������<���N+�%GM� =;bRf/[�Y�JO+���\ǧ��+�8��ń�!@"=�j��TnV��ִ	So�8�>H����c�a9,tC�F:@�\\.������C�'Ӫ�86@kJ�o���X��p����]*��-�b�4�y�v�����e�Bڤ|#�j�K@������>{!;k�}"+��IҨ�˕�9�u�U����D�z1�ww����,�7BKB�09ƹW�����eb��!�X�k��QN��B�@DpK_5Eڂ���s�ͤ�˪�ߒD��Fs_��Ǭ��3-#B����eH��m�Ԉ��р�u���$>��w9�������B�PB�P|~vF�//�����Ix�ͮ���P\�Z�v8��X/;�BOOH�q��0K!�Z7�5`A��!�L���
.�בD���c�+��s�*J�D�Z-h�Q�5�_�z��f	-5JH̬���=��@�7ID���NC�Q3в=��>=�9K�[}u���볋���7���t���ȵ)$���h���Q�$�H�3Є�be-7�}�����7h��o�Ο}��/~�>��ɳ�d�9?��o!���].=>?��3Lk-I�~3�)��/_�^��s2�?>>F�H�rvk���N�Z!t��;�M�54Y��~�d���r�OvF�i�iB}@~r�;���0qea�^�������R]��l64�n��U����`�W�
���O��7I��b�;���*���۴�2s1�JȐ��w���ѡY�/HJЕ{_�F�K	����X�+`����R�pqG0�q�`�?�L`����\����Ew���p��%,jk��h�b� Hz��뙨d�|�Q|�?������ʹ�Zr��b�nG������4J�C`������IH�@��q��m����mi��G��C:5?�������9g�4go��إ�{���j:!���sP������`��*e�;�C�R߿����~������FN������%-2�N�vt���(�G4&�*x��[���-P�*�Y�
%:),f�&���F��l�|�]n��2�ҁ�%Bd��O�+%i#
��;�p�d��̱�
� ���F	9t޹�<l)�?S��i$�f����7�*+h���Ik~Қ9ٓ4
Br�� �4�&��Zq��	��9iGAz��	ՅQA9�"���'�$��d4N�!�yF�	�gh+7Ֆe�	�e�=�`�%��4� +ɂ�m�Eu�V8M���Nk�k��eyLJ���[m�:7S�-��hꔾAA|���nh�Z��c�����i5���a{4��l�"DK+�S���|�o���mN��9i� ����l����S�I(�+��E�s���ې��%��`q�^;�m�p���6$8�>�:3�{-Y�¡j�Ö�!�+-�o��V����C�O�������OkfB��,�1�Op6Hq�fJo#����w5ES<h���3,��#��jR����H�ܾ��ot*�Q<;������b%��ٻ��,`h����p��hlҜ	NTY%�Ǩ�'�;W0 ^�\�H�4�A��䘻%0+ ��j./[}�Q6�vmnX'�fEKOF�����ڵ}n�:�Ȗ:؟H��9w�Gd��k����e�k�x������)i��8s�y�X��47�bkс�;_�_�|)��9��XR˒v��C�cRʓJ	Al0Y��BȜf��(R�Bۘ|��#�,5/s�؄�,{�xd�3�" 9w�6=:9q�����V��xe<�;�������k�x��X6�7��M.��v���D��U\�$K��\��u�(ʛ�g'���Wٵ+m��`�.*I ��a�r��%�֛������G{l:�ڙW��w��v��g��Fۣ
�D:4��1�dNOO�qћw��a��舮I��I��U�4Cʝ��d���5!�>j����U�v� \àtK��b�Z����0G�����ĵ��1�B�^<�#�j`���}y)?��r/�y�4��Du�Q�i����r'�{W
K7\��It�LG�BT����Q��VgoΑ3��Z%���h�.>GG � �L�$-��^1�����7oޤ�8��6��A�t7Hervv����MS�O'���<*?F%����X�.m��tz�����~���>�oV���jI�#f&DA�d�)�f$v`�W��8�ڡ��4^�#m�ݽ .h��ɟ�ɟ����������ÇA�͚� �W�/>��Ë�<`��H &5x-ļ���Q;������2�"��\h�C�]�5�y�[(M�o�~Y.2T�w���
qB0��c��8� Ғ�/U��Gpx���S��@��N�YWҴ���f*�"� s]44O�h%��R�[P r���b�D���g���<������|`^�~C��t����Qg��9�4��K�<�S�D����e=(��e�I�z�
35�ݏQ!N4�ML#��$܍GйXA�g-z�Z ��^I�q���m�z!�GB��$~ZU�V���eǢo����nMߥ�lP_�+�|"R@��O�޾�=F��I��V�`���� y�Q�5�ųl��;(��L�inp']�ix��I�D�`����v>/�K�bM$ob`c�>D�OGO
k���4�VX�%����?��Q)�4O��c��b9Z7xn=�7�_`��O2�>��#��1��>���������������B��'i֒�8k��o�8�P=,��mǌ(�4Q�t�z7e�ԓ�N���i��R��b��.�
���îa��3�e�í�x�2���F�y�$�3���h��K6J�����WDUT��7Ja�2.i��F^I���s̄C�޶��7N�P��7�wD���ғ��pA�`���=� ;X|,թv#| 3�d����s4=8�"�4F�-#��`3�>x)/�v�Ӻ�a6Z(����O�k��� 4��=�T��d?B�dx�xp�M�?��7���1������4�ޓ��e?X�$�NJ�{��y�5p��������Q�l#�N�M�p ��1��x���(_pDD���h�83Oʦ�pN��є2����T���_'sMƚ��;pK>`�-�h��Zi�S��$���������Չ��<n����l4u9E��4��]FÒR�36$��msd�I��#_p�h����Q���4j�˕�Di��#SCTɞ���6��9�ub�[ѱKvL�_�:��µ2��4tE�˽��-I��ŵ��K�_+=��V|�"綂=�-ey;���r0��q�t�J����β�;�H���\����"��3��0s���.��ar��7�&K��i����7	k�(�rˇuRY`��M��f��A�v$L��^W<Kc���ta��{d��em�m>����lsܸq�dg�b���u�w+Zr���?�� E�v5R��֧q�!��trrB�}��b�Z,�����A̤tBr��0����L�9����c{�L���^�k�r�#N5� {�������N �Y��G���@�ﱞ,��6QZc3fv2��6���v����n�<x��]v�G���w4����f\6��"f�v�E706����x�4(7�/:Q��*eR�5�&[��Yo�VM�@ ��[H;4��5��x��[��)gpW�3e捭O_�rz%��� o��i i�JJ�Q�����I�Y���뙰�\.΢�!]�tU�R����B�����;8���ѣGG���N��:�ye��5��Х	jܔ�(�趚�#��|��E8?�$U�k��7�]�m)�+��-nNJ��S�>Cn!��XSDp�.��l��"K?_%3k̒h��1_�H����[%���֎��AJ�+M{�ޑ>[6���¾4a���
Z&�{aY�ʘ�	�8b׮]����$�Z�֢p�qw�-0��e�@d2�A�wFOP�7����m���ɳ����J�U�p�f&�Q��y]���7-{�䆁�Ѻ�7��fԱ@���f^2c9��n$����#%P�Y�����xd�[Q�i�zE=����$<#�H�KD�1�ms?hK���Iy���q�e������������hg�x��}�6�ZV��ؤB��Iōns�(��+Z���W�ci�YJ�����K%����t��O_���������UMvv���_��?��wg�t�q5�ۿ���ã�#��I8��7�i��t=4�e�A7�M��߲�0.��~�HX&�3h#�[��HwuI���p�{�="�C�Z��Ĥ_��]�8TT�5F/����Y����J��lȊ��N�%h�h�I9fz��5�h,r���I�xe������;�#�#=���Pq����,+��M&tR�g5_He�d��k�M=V�l^G&bb��tg�n��� �Q�iD�6��@�ʅF2O�+����K�7o�{��vR3���ՅH��$��QIoKUH?�tA����q����A$���b5�6b8C�G�,'�M�kF)��A3�N�Vf٢6�*�)V��ł�.�;@qC�#�c����᢯<{��n����ZsfВ?��O��A;ܺu�6 s�z��3`f�{�1oخ�N�b�g��饝�^�w�܁U�$����^�dI����2�)LE2d����� n�>�h �׎��Qe��ބB�x7��˗/IVfS���7���
k�C�`�ѓ�z;>�R�}�1=�[o�E��?�����~�[�y?���ׯ�hm]��M�k�Y�^a��|4g��CL�-i��^@g��'��� ��th@Wt؈�>Dl�ւ|����2w�����H��l��O]�B�\����f�b���mH=tW�K�r�5j��mP���m�:��v���%{�Tdy!���+��|M�d�Wvp��X���J&��z�(K`
����j��D�AC�Du!��[���)�N��bB`R�bD�9�̈́�����,�h��a���z�F�/^� �EwGz��G�������'7o�O���|�����G�����?~�Y-��e�&s��/�\�˶Utj<'�+��k΁ϧ΍-\�{YpTN�C�ü�]�7��d{6C��`��X5�
�j`�M{�(/Q�~�[T�b�FW�Kt�Dr���6�`:V�+�/_��(uV[���4�\1]e�Bh��&�>H"��������T��}�i�>��Φ�Gͽ�'W�#���N��7���O�������6E��uY�P�hRſ@P&Y>ò��7����呂�=Y8�;E��s��-@fs��_�XNQ��J��+��6f�bl�_i拍���õi��l]S<Z�EwE��� #ˬP�M�r�|�j�d�M�;n�jآ�f�]l��|޾N��e!$�]/,Ym��4uU�����4U�4��(��6,:G�t�UYhl����-�i�����D���2�9)R��"�+ �lO�#��]�U�Wa��}Rv㝎�*���|������X$k�gjL�K��Xj�Ͼ��,�x��.�h磊b�*�b'�K]"����aYv	+g6kP��g�Y�W^��R䱈�K�dY�p�܋"�ycx�n �@��(�3�H��x�ty��ܑ�v�p�q���d��ݻ@T5-ט��^��$�r�k#]zI��m	���
���Q�It��mԨ�I&�˥���LٮP�L�����zX�Z64�6$�-U�N�f�n�ep��F��_@�hA%b��de6M�Xo޺�J��X͝a��M��N�>�_.sD�������G��]�W�.
{��Q��$p���$��Ǟ�;�ۇ좬�m����
�]�{m����}�L����&`�"�5��V� Y^Ă�4)���o9g� H�2�������A��:�|�3Z�vN�/N�:GGGN��#����jP��$����R�Dݖ���A-K�+�V�|�N"G2�S���℗�Ϧ{�2*�n޼�����/�K$ˇ�{�š+�"L�J���<,v#t�r,���e�8��{\S�c��+,�>`k
W�KҥR:�N��B��x+�ф80������'''7n�x���'�|@�2�=�&��M�1�7��T-��2P݆zU���:Ө�����J��_Ԣ�J���	0�N�$l�gϞ];9�?8���(����.ds+�H�\n�L�sB.��D����!��?L�����k�o�4�4]�<�y�����룧�|IC��/��kǣ��K���X�7J򊟮G'ĥ�������A��s'>��T��D<�>Ӵ�ПhKc���]�Q�1`�#�PĸkŤx���	ľ}�������2[�rlG�|��� ��<�|H��	1�/0x�h���`�73�V���CA��5A�%Y���F�-��+�� �q���4߬�1C.�E�X!�ŋg�̫W�?z��4�h�ڢA$<i`[h-�Wp�VO/�r�#pǡh���9~�ᱜ":���A��J���Ν�,��<<�fGgoP�`�Q����;�T` M%���=ǹ�N��!��j�����H -���H�^k�]��>���i:�	@��~���r���2��h`�?�7���&��9{�p�S�&�2�i7'd���"��ҺJ-*�G�q�ha.����L��Ik�MY:���!�$G�X6N=�5�,��#a�i'�h#��vg�6)�ב&��Cn�%��e!Ҙ�:�?i̟~��~�#���y�:#4rC�sFЍx��Q�	e�$)�Ci!��2��׮�[fթ�i�ώs��B!��W�9h�R�NJ}���2
��+��*cχ��l(V[�w*<.f�=�b9������z����� �;
pr����$�q�Ep�.
�\��&ԩ���4\Xi]��kǔJ�Ԝٽ�w�L�:�"�<b�(�8,����OT 87aчo߾M�I��$7��X��@�hf�}H�Π�^��B��q��(���z噟d&I;Sa>�E��w�CO�����?�������������կ~���ӷ�b�I�t�������	�����LO+�su����vOv��%e�2��c���g�2v��w�T��Nasʦj! �}���^�

Ě���4n6'���yZ(�i0)�C#�m�A���63u�Âۅ"�DJ���aة�R�\e��No��ip�lT���ܓd�b�	X�)�2|Yi_� �aI#�a��gs�m����'��s�$��ֶ>(=��P����nֹhTA2����`e��qh�L*��U���"1s���H�L��Crain*�B�=���,F`��+�Ė��t3`@�Ӷ�\ʙ�BT��.�C�z[Dg��
��=���'����;��ϓ׆%���ǭ�qo�th1���9%������CnN���X��Z�L��Ib�5B0%�\J��v����W��zd��ƪ]^�A�45��E�!��7t�d���������
&��Em�*���&w\].MB��|����}P<B7�?fZ��N �n)-�6���&�"���x�정p��>rg.�J���G�(����Ѯ �aUJ %m�.�#�_��޶5�vÆu[8�՟��)֕�֫K��E���43��.h�wt0�}�̝7�ݼys:t@�f�n�(��TtXl�Z2p's��Tq�x5�4+���Rd5\�4ٝ���T1��j���$�����]��/��F�	达mF���Cv
<�ӆ���0W�nۄ�ʓ�ѝ���R��<k[%�hƉ��˗�bm$�,��"��nV���-V�,h�Vi 	vZU��+���R?9<��,�>d�mf�\^�H��	udc�!�ӏ�Q�w�;R��1���n��3��w���2o����i'��H�Af��do	TGyUT�:��N9�i#F���4K��~k�m'���k$$�խL� YWI=8t4V�$E�1�+m���K��΍�Sr����g��pv���24!*���
aG�W*U^�J;�;	Հ�0��"^F[����R�tΠ[q�!� H�j������\
07�`�٫�����ݒ;�D�}L��|��&�$��Zp�����6������H@0���?(mR��vl�����/B�/j��j����k�ylz�29h�՛7���4n��3F�B�~ �H㈜S&~9}9����Z��t�t��-N�2����$�;�R�*�A��&y� ���4��;DI��Łd��v��'��Z?}���F�ዳ����~��_\\��l,q֖�+�%�� �"�L/MfZ���PMg��[3������mG;
`vr��a�����擟���ݺY1iC�ͦ;?�����G��y�o�+�I:y$��W�l�	O#��o���h"�Z�������0�]�Q6IKw�E0q���˗��}x��OR@�ړ��z4?*M�UN�rz��+KL��w���Q@y8���ޚ����8��!�x��ܕ�,�Tf;\2�&n�%bJ	t�t�K��bJ�_�N�풺��Q���^����� �V?�Y�^M�:����aLz;C8;?��Z����^�B���)d-D�3b�ZXl�P5?��O�]r��g3ۄ$��b����wq�	ք�q%p��삯N?�޻�y-�X)�3h:
>�d2� �z}&�g�a���d��50?Q@Fpt-.��he��2���ѐJ����Ң�S���J^�o�>99��D��#M������E[v�a�s)�RI��P�((���}�+���L`'������О<y�Xg�x(��\s�@9�v�g"/d:qBiҸ[}���蟝t���cGY40�9L,�9h�VG>�����/�O��կ~�ڵc��ׯ�D/p4p���A�����͋~�Ȅ�!x}��֒�^[� #�(��:W���IjAW&�D���C�EWQR�l��VEZ__]j��841V�1�ZKڢ�f,*0�'��9�E��<��P;��*�x�� ޶.��Ҥ7�	99�F����m�+<���irs�}Ѿ�T$�drЛ4?����Fi����i˜�m�w"�ND19��,K��ryD��������0����ހ�r61�� ��������>��O����_3SA��_�����rԲ?N>����O���{�P�q���0���iԈ��j)���a��'�M����3��$8�e�k,�R	�~Vpoo��)/���V�x(�O,���ͩgw����Edd�F���Ra�>ǣ����Z?j��qn�/\���0��H����u�R���)�$}髣q
2�Jq�f�����O�J�7G<��k��K
$����խ|H�ZKi�f��0�\v��dz�픺�X5NK�hol�(-Ja��	�[����ɞXtf��@�W�d�YE۠�eG������j���.2�p�]Q�]�~})H
s�ЬM\�.9�W�2v-}*�P�T*%�s�\�&%��:��]w,��	�^�9�Ǔ!���Z�жv�&W�5�okڝ�3M����Uo���\ԦTf���	
��6ñ RCa�|nV��QO/h�^1��p�zm�&��A�n��At:�~ĉ?��q��KI� �1]���~������ I`¼3/�<;+q�g@$,H��̪5�,�
9��ʑ!c-kli�w�|��s|H��+�:֙$�!!�1G��$J�����G���Z�J�s�nԯ�dQ5ݎ���lV�fJ�Γ���NYܼq|�Νw�Ẽ�)i�Ɉ-?_qny*�6������"�3=�32͢�+xp��oZDw%��ߌ�{xS����H��#��%Z"^�P\�����i�5��"Q�Ae�_^���Զ2�+��=���-{N[�4#m��4��������
���0.)��/���\5�m�l]Mau��4#��BU3�l�����Y�Xd�����m���Y���i�d��,:�h��_�4D��/���*N0*����ق�l7\g$�JZ[�N��m�Gc���Z�ьSf7�_˴��T"��&�9zBw��;G�U*@��>�� / ��*��Ą��!7���r�N`h��\}���i�ah���e*���ׯ�h+(�&�'g�4|�<s��qqxbQ�m��^RH�CH:W��m��^yE�g�l�/����E5Z�#3�)좖�ut@�*���蘠�L�A#�3�M�Je6+��\f�\֎c�t�>�U�%k��9��j�����C�#��st>��Y�p�����%�δ���=W�dP��ǏY�M���_|��\ޙ�O�2�����p)MUif��������'�a0�0�k�'�TO����_��{|��w�]GFc=z�+���i�/N&s�e���!���J������������8�7�gDaMsы���#�[���鑑R������9��V4Y�V	�2�8�v�b�!��#�\6i11��!X),�$������P��K����>����
:�*�8�465jn*5�9V������.��]1S3�[!��}��~�߿��G�a=���ygiB[#�e"��b2�G���� �ZE�-O1_+(�m6x�I�������GI���B�ݽ��El��(W��^��,e�f��vXJ�s�y6�!��D'�B�&:؜��L��mI�Uf}%E��R�T���n^����Y I��JЊ(�+()^�x��zx���|������|z8) �xA�A��E�<yr���w�{�����c�ļ����<�x`�����sd�s��Np��Ef�j�k"��a� ���d�ؼܑtyBr��8nzV�����L���;��<?�<?_��#��AB��K+�s�n���|D�1eDykz$j����S�8(z���Ic8M݈\#Q(:�Y5�!�v$E����؁�-]+�R����0`�U���I�H��N{F�=�UC�"4�r�)K's�-�aQK��{zURU��^��Պ�6���2�9s��t��#���Ӱ�0!P
d?�."kYZ��軴���J�O�Mă�8�a��@fm��栖^�#j�I��EQ�1p�V�!��c��?��?�C�����q��O~�� �����\�h�gə�d��48�1����P	�W,^:Zl���Ei�N��"�x3;2�}��`OTV��<)�`��o� ��T�l#V���}(�����7M[E4����5�h�WjG,ac�y��X�I��C�s�T@�l�X�R�#�T˩dֵ����^-șL��z���C�h�X�y�Q���)�$�`0l�zT����rK��R�Z�<�2���NO2�^k�,�`����W)�R�e��%[�ʠ6��X�sW��R����b�Z�k[��Yl�-��U�z�glm�F�< �R�9��#�k!)����zw�jXW ��X�#�Hmr9�ʹ���|�sn�Q�-����^���F�p�"��Ħu�P������y�Q�0PQN�Ͷ<���Z�D���M�����@�����7~��/�L��$�n�0��B���e.4$���5���rJ��H��lxβ�aHH��P�#��8;��x̬4MI�E:�Q~�h�����uS�5��2���Y)�yEZ� y7h���g���vlߋQ>�|gϰ��
<����M�a�aX߹y�q�w�yx�Ф4�u�;!%�3�.Q��fk��&�.֚W�w�ܜQ�pMnT��w�2�n���F��Z��>��%n�������s�v ��p7�Z��Zk͜V�ؘE��Bz�|�INkl;m��`���$,�>soi@d�E�&o���5#F�F�!����d�h�!�0J�ؒN�®�����h�C0{��I34d�\��p�BS�C���w�#�/�[A�x�dLv�r���)q��K	k{2�!ˮf�����!	�-M�q"�l>2#w�h׸�kf�VY��j�����7���xb�=	��zw�90�h�'�ʬG�Z�})彽�˗/�褫5ܑ�G5������S���Z�! -������������~�}f�w��z�K~)�F�䯕�k9�C^9� ��&3{���oq�ǖA+,H@%�05����ϱ��i�wm�)d�����74ip,��2����CZ#rli�L&�V|g��V��A�:�ߤ�E?�Xܾ}8PT��CGI���0P���k�q�j�F,��.�H$�i�H���]t㝣�~�`���{�͚�������r�X�/�͐|M6�lw��mp~��pHCd�A���v��Mq�LvǳQ;�	پ�N��e�� 6��G{t�H����^O��/�]��������{oߣϿ�����G��|����{�k�B�f�*&<UGK���&���T�՗��V����e�`{ԕw�a�k	�[/W���g?�I/��Ӫ��+�����s/�,���S	p^�BR "�ƃt�k9(\A?��9���K"�O!��+�mn�>?��|���P|�����Z�1���7�^��a�]t2~�1]���!���(��+�����]�MZ.Xݼ~u�vtp| \<U3}~���`�k��"��7o�jI�Z���cٻ�����	���_��_yh����(>d�g�uy�@����)���2�+ݰ�ޕ��h������G��u�8 �_�|�u�-\Q3D:�{!�V� �lz� t�2_��&3}�2�bP�y�)vdn�R���E^�~��C��b1�k��z�&i"D�Pm�jM�S�9�v�&�-�Cf��V��ַ�_�NG�,m��l�����[�� ��ʅ=�+�]����m�%��MY\Q��]K����5'�Mf����)�PT8l1r��-�b�^,�"�霸M�B'*00�8���n�D4���C�`!�%�^AAX�4C�A���ro
���n<��e���\�Uf��Z h�I���&�?ϕ��+�ֺ`x��1`��KE�ƆvLN�� ��*e��*��Z�s]�5��36ɨU �oZV@�Ӑ;@�Ͷ�p��6�����P�3B�;�B�T��ܣ$\C� �������>*�xW$�O���s���������`����A��r=��l��* �VT�m	�Y4�'�6t�;7�)��OF���_������ˏ>���%�N�f��gg�`�]\�� ܝM./����_��#[l������i�l\�R�/��YN��Aw�!�p���X��m� �_��!HGA:j�a��a�k���E1���_b���_w�N�V˪Ë����e�\��cQe?h����U��ߑǃA�>���d�s��䢅K�_]mbOP���󵠿M{*0C�(�rEd�|��.?�%qx�.�^�LM��0,��N�9r";�$ޣ��$����@��`��S�-���r�T_r��t��H S�h����B�-x'U��B�"�+A#2m�ك�6�kD-f�d
{��4�j��/�o1{�2�Pkۚ☁�>�s��@��-�����^$i1�����.H�J�����Rj
�v��d܅�m���	p:D�nR�R�L&<̤%�8�>C�	�(�g|IK��F��0�a4��ϜOK%a��!�L�Ci ��Ƀ��
{�4�Ǐ��"�<����2���Nat��qƱ8�W��{�/}������F�v���`��+m2�*=m��b*�3e>0S���"���{����}F�P�7C?����L4nQiJ'�)��E�\�{�<���Q�4��kw3� Y�8���tB4$����@9<<��7���U�L;!J�#�IOD�!���[� �)'�Y�8 &���اV�n���13��o��Ta�t��_1���8���_��|v�c�U^َm����і�|@��-D%эl�|��E�)WTR��q�Iy�8�)i$�R D�����g(q<K�I�hw ���Kr�{�o߿g�٭k'���z�U�G�J�퇾�#;S�ʏ������u�'�,�R>�mQ���L������'��B��v�&߇q���1������B6��Л�2���1_�WQ̈́���eH4�Ur�p ��	n5��&�4
�\/z.�QOO_E)I�$ ��U��z	��P�  ����Y��th(����@nxe+�����I��#�w2�=+�,VF�5�%�q�y�2�iR3�6gc������3���\]���;t�r� c��H���E�Ƃ���tA�	J����9?�./=	��dǬR�8<phLN�+��"�����~�R�
��=�}�j8,����>��1j�Il޺u���_�� `М:CEc�(�eD�PH���GÊ�`w��D=��88b�� 7�����}~ɒ���58��֋�������#4Q�u��������`��$��(�
��}%�
���;��e�O�Q����.fR�)�N�\�5R>�J54���w�RI
I�d���&��ͧO�^^�J�P����BaU$E�?�F� �q@�=<���8��~w(�ld�A|Լ|�m�P�z|rh�N�kJ ��D:�����?_�xA����~�,�����df3�{X��a���-]�r����:�K�BdB�& �B���X�yQh]\��K�q� �QI)S`�;���!�UC�+�9/�Τ~ܷ��#%�e�v����E3B�B4m��L\s�����B�C���7ˡ����S�՝2��j���q�ŹN����I'�u��$�h!�`��9G�A v&��"|���d�=���������׿N2���?��J�KPB��:sb��#(t�����Oq� x�A;# Rk�hP&>��8��|��;k�:C� �ׯ_��Җ�a�а?��?|��/����o7X�0}%�g� �8>>�yI�:�:]�v��i�/R�Ns$<pQf�p\i5G�w"Xl�Sʈll*!.̤u����U�-r\�˛����e���8�xdZCL��A1l�g�FC�4H�VI��QK7p�6R��a���ׯ�i	�%�u�cHI�v�AzeP2�g_�?<�Ӫ�X�Ub p���P���a`����A�"����q�-g����pf-_*�Z!� 
�\����Ɂ#�8`���00�db���M��~��?������(#��o޼��M$���������ga녴���԰د��:���"f��J�|��O%��2�X|��v�V�A��Z �k�$��\���AF��.7�E@6Ш/�l�����e�͵��PFū%���*�
ߵ]�~-��h�X�*)K�
����#W
��`;5���]E��g�[�2��ʴ(����+h�E����;{٩����W�����N�#%'��1r.��6���M�%���9��b�-x_���C&;��.�q��Xiz���ʎ���	��[asK�����ѷW���Q��N��-( ��ΜAl9%j�l���$Z�0����D�P��L#AS�Ѽ>X] �_ӵvڝ&�L^C.�oR�Q�t�����6��V����6sQ�h8Nfz؅3� �l6��N��X�.A��N�0l��ȑb�Q�E.-<@p׮݀��ΧGGR�!�	��J��p.���&���,K�M$-�6��e�y�V�Ӯ����v��4�M�yѕ��i/B!lQ`t�M2��
^��mOj�Ν;����#�.���3�̔ q�Z;�Y� >^*Jݳ��t\%�G#G���w;mh��M�"���)������hw��6��.��޼q8�����NG;�Ԓ�qYǏ�I>�\u�/ϓXZ�-L�B�@�Cg�\�4�]�Y<��u���U��F���HZB!���1��|@kt��< 3&3�r�k\�-x%�K��4ˇ� 7�o��"�E�,0�4�G�r��+��Eח��{=N��?�)��HbL���q�V�,�s�7����r$����U7�� �����ٸ��zu1T~Cre�c�V�����.u�)g}��U��(e���|�<���-�C��W�g<�ue�J[|�
t9�w�B�"*}��-=Q\�$H1�r�$^"����L��@��`����_�9E.����ba�P�<a��ܽ{6"��q��!W�@�d�maOb�"4��x���A�+�
��:�)�,�{�$�(��|�7�D=w�����×�S�X�h����%x�2s��F�j�PhH>�'mn�Wo��C��� �
� ��x<1ȇ[�&��L�j���=wqq�\�A�(��LI����Q<p�ϝ�1��ĬYi.痡'�C{ۃ��F�nwo��ԭ[7NOY���{�� ���ק�E�\����m����&#�ғ`\,/�Hr�aM�\��r�R&9�+�3])�5]D��p�Ub���]U��vw��{��+�tM��g���[����g����^J�9Sq�:�~-u�a����<�H^&iE_o�Ig�1���xzpx2���X�y��b����|�.fFK3@q���δ��� �Z@@�|��k�0r�U]�%�Hw�bѡ�v�?�Q�Zx[���*�J[�K�r����{��??�������׿VF�����}xί_qD-��|����C��a���W�P�=}��͛s�)�=D�b���R�-R�e�SH�+b����i�<�~g�\ �������ߗ�k�m p���x7jf=� �9�d��D��M�'a��~>_,.ⰡM:�ݹ�_�(����X�7��d埲R���]chخl�+�� �l ''�t��[�≃�U7�S&b����;Fr�.T�7��6��P��!m֫�A�w"�VIo�2D�n*Uo	�I3����`wUڒ�� �ʒ^�C�8���E����F_ ��Ɠ�C�I��[��̍���Rq^�~y���s��mz�ŋN;��f"n��'Da��I%��n�`Ϡs��4ut��߿������ס[�MgI�#����ʡWjB	�7�v��J^p:��ᬕ��D�'�#h�46:�����ꅕro�������~�����򕯼��W?~�o��w�>}*>p>b��G�z9[+�ފ���b��J3����F��R#idO'�]�͒6����1Mt�%]FJM�.��!��@����2W-)r$;�1�������"9�1<����.��;6�Y݀/�)Z巁%l=��+"r]����N���j��-\�M��<w��УT�����D�s$zy)*�-"q/\]�84R��j
�>��0��H���0xFp@a�Ȇ�G^qN��Y�SsF����Đ�bn+��ԘÕv'3�,FH�j2�~�����d"q9�>�؋�/Q}B_�8�O�P5����5����Aj��ay'G~-:��]W����/��';\�<�r:jSƲ!iN.�v<�--� ��$VgH��˥�^�Z��Y��U�`�}8h�|�/��Zu�5�M���"�T�#I���$˾a�H��� ��KT����4��Qj�dbe��I)e5ݾ�F��B��p�2}yeMu
g��X��e!�@�wRy�P;��P$��Jb_)ON^���s�P������kK���Ym"C���F[|��32*�}�=���c�����vL�۳�UѼ�$#>fEy�����ީ�u�IL����p9ᰱ��CrͿt�P&W	!e�t�l �rW��.�$�?O]@�]�����.Y*"&���-�a�4�!��+�IR;�*�,(���z�Ze�AwF��X���7:=U����@��E_<JpP+�<y��U���?�|��E��E.0~�M��8nkpo	��W������(u"��o��:�����C��x$A^q����'	J��3��pԭe����d:H:MB�tc����d����DT����m���� �T��w��.%�O�@�TQ�S��qZ1w��ܹ��7R䑜��P6^ka�fW4���[�p�QٔiHg;^k�~r��tZ~n�rc��"VQPՓ�+�;x��/�FJ�4���ik���N��d� dX�4�m)@XѺ��>(A5"��@�G,�E'x���Xw��t@�Zά���3����V#�d�p�J&�|`F����|��}R�,֛K��g�⬳p�8&�!;,Q�3�t6�IJ�l{�1�4\R |��W�O��yd�s�	dpM�1�~�_�,��Ч"g���0G�^�۝�����J��{�����x����驜\�fjw���{\�Y/9��Oۄj#z�!�`���.n����4Z�����+�,��Եk�R2F�?�o`�1�&��>ə��x�z2F�Ą��FJlx-�c��?88@��Jc���l��6B#*�;�Z|im��h������,s\^��xn�px�O��\;�v<x׎���F#����T��]$�����`Gm��� ������4�@��OnF�!�m����텹QH�t��r�=�ٷw\e���XS�;j�$M�ans�=�9G��4��5.K�W�i�v�@�ަ�ť�v�5��/V�4?g����!#Aj����b��E�y[���T bG<+[Z۩p |����Wu5Qgv�������	!�=>����7>���k׏��*Ӈ�8�uVˍ)�"�+-�Ç!�hK߽{��'I�?�#��_�������.}�c�P��������`�@�zX20���%�M�-;�3��8����/�L 1*H0�m$MF���;���ԋ�E/j�D��^�_Џ�RZ�MYS%�.3P(�r|��������L@�U��&߻���������_i����[���E
jӭ�P+ʘ�}���Gg�73Hǳ冏x��v���!���͇��B�(n�\k�l��l��������&�Bf3����=$�;[�����,u���K��ś������"E�k)�*Q�l�/}'�k�;Aʈd�	¨Z?�%��(
K�<>��>L�+"d �|�9�-(�X��S�!Bw���S�^�Sط�����"&h�l>�n�S�◿���R8�_�֖:q��<����RD�oh-MB�V�=$�Ü��/2H�--rΏ
��eLP+C/�[ ����
f�1�A�@�z�h
3Ѧb�����|��׃��d����K��D�Zm�'O�xV(�(��p5��ŉ�4�G��QV)/h� ExX$ ya�w���3���`�i�;���0��h-�8��hK������� �E�.�MYY�0�7�:-Q8 �W�L7VNT��%�׫<�k��U;)����l_ql�� z���N!F�g#j�±�M] ���y�?i~{��J��� -�\݈��iL4;;���I�ٍ�j���`�s�/%�n��T4;�|i����k�Q	��Zs	 آ�(<&E�	v@ye�Yd����5�T��s��"��_�G�B�_�������S�3�э�.j��dH��D�*�U>3k��F��P�����C��)�)j��v�Q�_IS�e{��v2-ilyޕC�GP.dty��Z+iܲN�������,?<�����*e;b��ُ��{��j�}q���3��.���/+���Ҝ���rM8K�����m�2�PP6l���l�m`���ˍ>�r#�7 Ak��*v��sxg��/*m��5TcF:~�2�lʠXDo�Z5D���0:-�橚d�N��G�e8��U(����t��Tl�QV��}�Ӓ���8>6t0�X��@�ϖ�m`�\��2n+վ+�b��v�0u%��R���,o�璜���lf�pytְŜ<���W�|���>��C��<��iL�Tc��ruE����-��rZ:���@���ɠrHA�}���pоl�>���5�%�ΤHx�k��,Ğ+��d�i5ҡ��n֗_~Ik�|8z�J�;�	�0�[a����,,�!osa٘���.7�	$�y�f�@d�vK��L���냎��7�H��L��fݻ}�ڽS
Un�< �󨵯�+������n���TqVz0k@0�>�����'��ښ�2(	.i ��a%z��Z&ik��6�~�cz��܆��O���5y ����f�4#q3\�v�a0�(��3<vr��\�Ӹ԰<���2��ŏiL�����K\�])!���S\1S;��/J��k�Xe��q}�&�+P��w�ܾ{�/����D���D�8�$ʱ(&��k�2a�|VcgZ�����dE��J�{@/���D�q�APu� ��2ݒ	��5
��y�l�-��͒#C`���[��(>�����=B�ʩ* �!x1���Ed;N[��JR�n
�+N�D��%�A4�����(4!	R����|�5�<h54����m6��ϔz��)E� �M�:ٕ�Z��9X{����5���ƍt�d��|S�ᕝ�H�KP�(�8�2�h�~7��Wʌ�Cغ�n)7J�Ħ����ɍS�t��la|�{�����)����i�H��7z;9�H��Ą2n�<B�gϞыY�u�-�>˛-�"���D�Dz��>��	HCf����B��7��˯��_���w(6����g�s{/Mɤ[}ذ�֞!�f3^�+6�N��zZ�ϼ��ܬ�;�H�jR7�T͖��rծ��� ��N��?g4yv��U۞�b�"�˂�����ލ�[�j�-*�{\-s�a�:��82m���Fgy#�ĘRƧ':������Wս�����M�����3.on9uPi�ѕϦ.�_U��x���ûwo>�4���;�����׏�z���}��b1{���;ͷ�o�Ŀ+_�_��j\�2rbw{L�x�����[7N�x��������a9<`8�ŋ3:�ʖѶ�,1� B�@��xq�Y_��_����O?���v�q��������~%7c���D����������k�1@�(��E �e�jkH۠*�z<��i�n��+���]�}�ĕ��?� R��y�� �.08)#l�����?�"7��~�G��v"��|~W�U;e������k��,\�e#�j��!*��.6.�Qi�E�z�H4z�?�˿�K������`�U\d|��u��j�ȫUEN�M;m�s��f�k��ںZ�el�}Io�^���Kp���V
�*b��	Ү���*�nH��W߼y��������?z�%wu��}
��I�� _s� #��%�}�#m�bK��N�z&��ࠛ�R鮯�.�pl���P.�ѡ-d�������Z���!���6�@ā�dǢ9r��!�(F,�a]qm)&�P�/���k�l�x-+Yz�u���o�6�8h']A��obH�&2km逼c���FFq�!QG.���P�ܠ��ӛI`G�)z�v۟�o��&}��_��?�����������QN�4�A�� �l6�eyD���{�JĲ}X�7͔� ���;��&��6����l:_���)�n�v�[u:�����4�6*��/����2�]9�c��:)ۑ^sp�����G���E�95�'�Pdj/hW�3=Kְ3�e�*��بʂAW`y!��{��͋X��2�!Ch�&��b��� �!�a���(�ے7:������t� R�d:,��Oo�52�0�ֈ�юXνȗ���:t�TA8A9Ί#���TD��M%�@v�粋�c�SFE ȼι	+2	��/(k���m;V�5�m����j.�Ӣ�TP-���(�j���R�x�^(2-Ո�������������PJD�_��A�d{ �F��]��R���]����0N���J�pF�3�����2�q�%1��z�`�r0�����I���iV*t�Ϸ���	aLS����L�`rA���%r!L\�^���|W�e�ģ�����LV�/��;�J}��A:D����c���0��A	�]?ʁ�X>��l
���4�~�8'�fEkr���vh��ݙT��ş?��K8>��HP�(\l�k�
W���v@{IY�`6d�,n�I�p_��J�+�w"_^�A����t�)�q���\]�����j})��dC��{[6j�R* <3OM���[��1סV�_s��j[̾�	�$U��/�yl/��3�Rp�KË�0�pZ��v=�*eq�z�ѪΠڷ��Sh�v�mU$�{-���F��x����|�"���P���1��˯�Ǟ_3��tab�i�@�,��=y��LQ0}��y+�Ȉ[�r�mȊ�c܎��A8*��	��0s��s17�E�&*9�ԗG5���,<	�z2ۃo�D=�C�T��|�]n�b��f�
�$s+��|�T�s*� �{���(�sM?��.2Ur6��a)G�"�b[hH\��7
6�\R4KϜ���Gѓ(P
�	cH"Y$��3��]l6��t��%4=<<4	�7�N\p��o#37c2�d�O�n.�M ��'�'�><!g�"J��Jɧ ��J�%9��%嚳A�@����|� X��?�6[�`������ǇH�ҵ�8�}�a1p�j1J`3��Ue�x������
 t��4#:]h_ps*����*	�'E��y��B}�͊{�R�QU4ısvY-�X�ݪ��^�6o�0nR�ڛ]v �RH��1��TE�b|Ͷe�Q��l���~�>����]��۬��^9y���/{��2[���"�\���������8LVDܽ{-0�D�+�P���k�c�$��J^��^:�9���z:��y�:��~��囕��x�ܿ�3k-t�m
SY)� �W�;��:��&ծ�di_���9�b'��_QM��k��\˦�Y8u׉I$S@� ��O:�I�0���s��������_~�L�Jh�V%�^�O-���H>vZ���2\�ЇF=ٰGMs��֍��K��6�SѽQ��h��^`+X�%k�kP�d���P@M�W2�E2" ?~F�����4��aĞ�}�Jp7Ў{_�������j`	�`�RA���V���p����gO��� j��Y���������o�%Zb@����NzظBM�cƑm��F��{QiF֫b�1<��������1�����QS��J���@��K�̰'�̚�*m�3NL��I�p��] ��*�<e%�7p�骵��|l��X����0A8,�����ЈR�xn2y��00*�����٩�T�l��ſ�F���N*�m{�b��v��
ABr�:n)XDIh��r���'{�;��;^�d����'�gN�+���"_hr���,8I!ȉ3�׫���	�]��2�3h���*��?B��2֑��ጕ�$��0��s�(gϛ��v9̱��0Y�j�9-��������
�+@��2/�9o��]��T�HY��2+�w(j�5DMX���WЯ����M#�P2�R1�V��b�5��r��Ykw�N.�0���bv[vp�.)��)�����WPK�1iC�gv�	~L�b1t�ck���)b�&��-�g5eYR9v�K���<�dG]��[�R!ZajR�Pt:7�#�+g%Eaa�P�Wf��J��`TP"e��tA�Q�nhP���MP$E�N�2�Z���= x��Ù����An���
��������+䟽�~��w��uo|�!/#��8�^IB�a���@]A�<��W9�ٕ�6�M%��l���=E�uooM8+���v��0���[� v�����w���փ�w��eʪ"q�R�S��9�f���"���[3��Z�v�$s�l
Y`��+e����v��N�G�Ѧ����L4P0fY�����ǂ`���bB��*��$Z9��P�=@ +*���ٜ]���7N���9b&����ŔΧ���h]��GN���w��=�ý�2,ƞ��v�UU-'��V���N[��E�c,�P�'���VZ݆/�GtbB�CY �3y�]\]^���8W�C<����Qw+>D�)ST�-��ɣ�Y����U0	a̝��sJ1H�+a���(����@6v)bo�>z�0C
p��l��E��Q�Ɋ�4S�ǋ[7No߹A���!w�kw�M�f�I�<�t8ׁyN�|�$��x%��{%=-�x|A���m6[WP����:/f�m�S�,!��>s�7������Dnk��EfxH��F��I����Z��>I�ϞJ�n��%=��Ё�f
l�x�\F�f��,t]��YY\X_K��#>*��3W,k�b�[�	�r�0¤�r��|3�H�Zp�����'��f�(i
�k#�A�s�b7Z�f�ZR��k�?n����[�3��]֔��~���Jt�֮�4!4n3�Š��W�%=&謏�r��(����֭[��0��d�.��z����C��E��u
�FF�#�迌��=�,��J�w�X��łB��-�.�Hْ�lv�Edib��8�۱�������[�r�m'�l����]��]��.��ԝ�L��DAw�-o֧�F�E#��tlaB�E�¦��-�x���`k��=�����	9��V��m�e�B9�Ba-���.��$�]�����w�wI���ƆlR٠
���k೘��~�^��",	�ɩ�z5t &��p{�`qrz�%]s�������_[�����[i2����#	�9��"'3LC���A���U	g���H�q;��ż3G!�;�Ev(����R0 C��.�dF��roV8��ӥʝ?'�v���9����ܿ��G���@���;��w�	B���L�'Swv������m��9q��=x}���xA[q�}�ꡖ�)nV�ͦ�����v6��~�Z={��x���OCk]�i#L�޽ެc�E�'��Jz�z����!�G�����Y1�V��MZ�i6>�D�Ǔ�b-'�=��>ǉ��K|r�f�(B
3hG0�� ,�*%�H~��J%'�߰M{��)=�b� �;0�*զ �.��`a)�?���Af��sZ<DX�N��UqX���T�,�|�a�k��1��g�u��Iq���m�%V3���hA)���J��Z<����C��hߏ�ݦ��Q�ڄ�v~~n�B�Z6�6��>���mq�����}�N�E�?�%M�(��z�(�@[|,0&�pL��2Ns\�e����stx�C�k(�H���6��S�hL-Ӝb�M2ʯ�i�:b���
e�A+��Ȱ��^���Xo���e�g!?�V�i�K��G,�8Q�}������{����)�?�����{�>�P-�T�\��@ʀuJV�*4���z]��x pV�گ���.��m�E9���E�&��̜B���Ym!f�˺�ߴq�op��S�7!�����Č�;#����a`�/�q��hm{Du�{!�Jw��r�h�9_�d8`�J4�?*  �LC'J��J<�0�uZ�l@�h���U@?G�-���%���#�,��5U��\��(�c7��x�S�
n3IVW����c�+6h�`�7�MCQ;�8�Ų��YG,`A��;Ů!8	��PÖ�B�r�'fCS�������!��������(ԅ5�@%=�)D�,��ȷ�8_���JrF��^._un��D�O�D��"�T�af1]��sJ�KE�8yUV�Úz#7/n%1��{r��L�sy������r����m�b�qh�ݠ��>��r �z� ��][��0�<JPu*�����]���K��KQ��2��2���}~�AtI��5���(|/_~���F%.�V��3�4dqkf��,�o>l�� ���L��Z']V�i�Z�Rg3+f.�{���� d+�RA�r�^�5�\��(ht�_ �����2��3�V�X�II��'M�¾�0�U�}�i!�����ڟ�����>Ɗ�9ܟK�S� �C���e���|-�!U�0U��c�WZx<�=H_��z��7�T�TGdl�&V1oO 7M���ȬੂA�V_��c�n�e���̕k˸U����/z�E�4��+h-���ҕ;�5@��d�+_�r�&(%�+���0|G���?0�L�{��;w��)�3Y��כ�	�j.�R1�յ�b?�Vt��鵛�z]c=���b��mh�/�����i����%��������Nso� ? Es4&N���v��4��klw�lBIf
������-SmX%clޭ���"/Yh�����ZO����(u���5�Zhf��Gd�hkx���I�#�{�*]�N%���y�D�l��<K�8 䉰3���P��@�@�)�p_���3�]"�E��s�E��Xf�$}5��vkH{`�`̑�����I�v,#M�]d�80�&`�UZ4�����F���,.�f<��>v��i��ĹGkQ�B���AiΌO8�%�O��UMsqv���_�Lx�
�v�S�^$�������[��s_�"� �0&pv#�x��XidL���l���&}~t�;�1q�\H��I��Q&4���׉�_���FT���0kN~�T��~�}�6�$�dG;��h$�4�k�[��Q|�oP�Gޚ�TAښ0&�ފSY�7���R~��["�Z� _OB��L�lט�[�nђx��w����l�e8c8�����=	 �>��3n�ɵZ��o������_�!ͅrl�F�V|h�bQ��8u-h�w�za���N;QȢ{�n�B�CE� -�+��$��7LmP��AK�xrZj ��9��z��8��8�����C��
9WKB~]�v�AG���Ф����\Fق%�}�D��BQp��#E\���� =I_
<T/���?^3�a��況>,�"���E�Q\hG9 B��V�	H��\�� �W����	0��O�����V��
ئM�t�jk��8q 9%Ac閱�*UN7O���Z6�	�iE�F:���	���Xx#b�(iNt��)��Ȭ/�-vZ��c�J{��������Åi�E�V��ߠx��U�06T�X�N� �� &n��P����j3\#3򽶓��
7nE�*n�a�0��-
N��X�̠���`UB(��T��n=zT�.-�����?�9�#�Gt|�sJ��^{�W���g��� ��k*��A��"���J�9<�&;\3�k!�ڡO`\r�Cd.��_?���E�ϊ����F��R�5u�@0��i�ie������ɱ�Ar��FUm� ���a��S���3����2*ϲl�!Y��������*)_��q��9�l{-��ͮ��-mQ������� 9�P� (�e�>H�e����m1{����/�h�����jƾ(���N�����Q�|��j	�&�d�5�C�����F.!��g���"4�����%�䋆��h�lc���A�I$:WX�8$l}�󮴡�Y�`Zڕ�B	ER"�0����Un�?[�2%#�� �BYa=pLE���lI� ��ɢC��V� �^�����B;��ѕ����E�ʿ����m���Yg��s�C�x/�^ۚ�b���&ƚncE�k�+Ws(Je@d���&{�{-s��IY-7bw�ru�<��r��>�V}��kwaǳS�>�2�h\t�ж�'Y��nT�Z�[U�u��O�T��z���[L�\'Y��䢠}���S��IDy��V������Ұe�R�RFx���';+c�$��,��)w	v����ō����<�8e`ZW�9�XZS�^�胃�� d��X���]C˯���ʨ5��3&�Ll�
�b�]oxtN��7Xz[�h�e���N�7g{7&�����`�]�}3�z�蜥1��m=f)eqy`��A�R)eD,�0̀��R�����b!Y���ҼlTA�f�Ĥ6#�ءϠ�
C���{�ۭ��ؿ~�������K�ϻ�:�N�Ma>`j���V������KEd�Wz�x5c+���eE����u�TD��1U�n�gD-���Aʺ�27&�h��
����n��|us�7nO����%������>H[�V8й��F�t'����qUQB��5�GhZ�2sJ���vO�,3�V]X�/��)::�^�����,є�Ç)̣W>~��;�B��E8���.	̜H��B�k��v�7��`m����� �V�R��b��ԯ�;̑H�q�5�]��h�2H�6b�⇘�lG"�d�Q���+��`�#>��������� �e���W ����Se�۠d� �i��׵�ag�t.{�v2���}���"bA!y���@�%��od/�S6PP*����!�^z--Z�4!�(fTb��mQ
�jZw�7Co>b���\}�&�ٗ�2����q'pN#T�6��Is8=�+�$2'�L<][G���lB拢�}:XiG4���,�"��?��?��х��?~��79�g�J��j>�n`�:�D�EC3
�<���M�E^�~2M�j���8]�U-�0Z��g�_<ߵ��Kn�M��.1�{�kᖈ7o������R��Qu��j����?x���j���;��o�PMm
���a'7`��F.�
�,E���^<��a�vm�O��>�r��4�3�GO�KG��hs,�n�8�w�γgO?~�q��`��FzA��ޯ�op��H��2gF�1�o�}�6�)W�L�(n��v׵[��{a�H��!=�4C��jtR�wx���}����4U�n���l�f�"����Ђk?����
�&+�"\�`��j��OX�ڸ9�^눭��41��X������� ܲ��W+F�� 1�����Z����/�9���,Ŗ�꣣,�����K�m�˽��ڌ��N\P�赞׉� ��Ѧ����Ƣlp� \��r
��&z����q���/�݊u�����	"���kB��j�P��O��gN� ��P!08R����������|bЯ�^`��
A��iBڢH`pV���� -D��%}�� �����щv�Ś1�Y�J+�87��R��˂3yЀ�*8�z�W��k�8�?� E����%T�-	b���z�N1�I������%��Pk��k"�wV[#q� F����4��0���$�T���a�������DG�=؃��PN888�Ý���0ST� UD������z�������_���駟Ҙ�wa0���+�� V��Mtad厏���^ohK�wyu�C":�Ь��/�??��ڶ�Xq�Jp��s�v����I-j�O� ,a����|��E�'��$��y�J���� �B��f��B�#��lJV�p^B��Bј�kK(���!� (�l{]~��_	�5�R=��X,�kJ�.)�/3G(i�{ԊI��8 nr�@'��\(������t���&<��^�v�*#���-a@˂��M�:o]��A��Daoڸ媫�P�������Ű��Cl��I�*��&�b�e6�t�6���rge�=^8Y���	^u�,�O��a�U�.Ѝ	7��}�D�0Y�U�$�~��@k�Y�h�#Bǩh�ѠA��] �	�MM��K�i�8��8�������羲�s�J�u�ew���u;^���(GE�m�!��AJO(��+Gf���c2���d�Z�����t���=�c��T�|�;I�%�0�NƉu�8����y�2���y���fD��9ڴg�|Ҭ(���?�[��&���pb�Wt��Lg�na�v ��H��l� U�R} |���Fr�ڧV�J���N�aYhJ�_TcYsa�Ty*jS���b��-���Z[�T,������e]�nܸq��	�&&
C8^!͕�0S��|4kPZ�J��{�VsE������ �'��n�/h��|x�
U�A$:z�����WO.y���W������?���?�ųg�pr����nT}���Go^`%���_���g��|Z�'g��H\-݇��s�=J7M�%�6i>f'�s4����LW�G�� ��������������[�ܱ.�%7�L�NP���`@�~(�3h^7�w*y����"�k�陼�Y*�2,�� Ñ�c��f�5>f���p/��զLO��n
�n%AA�cԜM_����q�&(�f�¾"ϟ/�P*����П>|Ho��9�ev�X�TS��"hH�8TN�N�z�-�W%%������ܹC/΅�;�1�N��:�R4Y?�dg9���c�/x���/~��4�dz��ӧ��:���X�#��̒s>c�"x0wP+�[�� ̣g��O�ª.� !;�bHaI�]җ���|gDi���E7E/{��Š�aTiѓ4w��:N��Δ���t�ds<j��]�T�\ǂ(5�f��4�����������{��'�Z˯�?vvU���5a^�ަ~Y+9�P$\1td�q=�~���n�Y��{2U�.��aB���1ڃ6�>���X4�6;���7t��y�޽Ko����eZ5l^oY���&�z�-_�5M+��V��\�Kh�~���@����/ �d�e�	��{��1����j�{�w>��>v#-������4�Kb��~Y��΅�H�ӆ��`�ha9��=Ё�FI�h�5�h�=y��`�y,�#��k �׏C!����m��p�B���ԩ�B^�[���Px2I$M��ν&z���/�=��\�A�B�~�1)���ITYU�7p?��瑰�1T��;83�}�m��p,n?'>k����X��8o��n6�"t��>�?��sZ�����T0�p��bջ^@C4���}��A�m�:�NL/19�>IMQb���:���l�Z�Ŷ�X�Y�47�Z���
L�G�U��9�w�|�Ä���N0bri�\��!(���gQf�_�~�-��6�����M�a����]Q���Y�hX��������#8�@aR  ,=OwGo��U��,��0�hg]�l��jX<�wXT#��mR�l��������Q���^�`j�/.eU�7bu*hԖ��*<�+c4����.�7�ƕ�jS*O;#	���G��[���+�݌3=j~�BH+��WB�o��0-\X%��'��9?��Oh'ҙ�vd�Ma�m���Y��F�4����{�7�-�<!��/��qO����3#�0FK=�I6�t�^{��(��Uˬl���1�~,1M8� ��,��-V>r�'�c'�/,f��CA�e�t��BL,d�&c;��Vm��9��x 
�_���R_�Pd���R�4�{���`8�OZ�݅�
�\V�������@��#���eZ�P�THLhԐu���� �����r-pԎ"w��ʭ�y��8p�g]��j����
/ɔl��HGq�+��j��&h�п�H�'���:��L]��w�t��6������t>W���m��ݎan'ݐ���]X^��߶k��W�T�3�̡Q��E�E�8.�6m
�r���VT�o����b@���o)�T�+��7-l~Y�m� 46r'@�/r@�%N��e����[75}�c][7��S �d�L��䇯<��m�qu���qM=�Ϟ	2<"�d�쭐�c�7r���|��+6a�tE�����g����0gXR(��`�
&񌥿j��� ������6`�	t��l,�;	�?k���@��ެ�!����#�$+�V>춹l�B�-�6T_�j�Lװiw-�~|L/��鑋[y_��ojVڬB5�<y�������������͛�)�����1@�\�-{:�Q�9��{U|	��3_F�̈́F��Ƞ��t7��NS�������)e�N���'i.����L�N���X+4�M����k�[V���xud޻�pt��px@��|1=ݛ��7o�89���D�����/;T�#*/�e�S���K?�̙�����e��U�~!ja*m�sL����>�-}Bk�v/�����6��4'�w�j�\nv,<[4���f6?��gK�q���S���M�_�֫=���z
:�s01����eبL:�l$�@�5�8^egEqg�z@#��Y���N)z�+�51���i��ɓ�q�A\�4���霂�7>�wz��`���l:��<;�i3��N�;�8��6;��������_K��A����*������X`�)M{��R3�����N��kѦ��O&�8�dF��E�f��σ�$�*�8��bu�⢮�H{�O��+�|��
���r���p�*9�0� �Dx	����.����)_�o9}�Ve:k�Bԍ
;���a#cF����T*���i�p ��N����� l�"�G<�2��V��ٚ��G�I�O��ڝ;w{�gd�vo���������G}Ă�����3+]�$� e��$�P䂭1��gc_��o�I5q���ӌ�2z�q��;(��f����l>�_v_!��MW��u��ǫJ"�_!�%�(m6+9��;�r{��e�v6�N����0 X-8�g�OS�,3m�h"7K�!���lB��X� �T9�A��_��.������ے�::ڛLhn�*�����]ۑ�>��]�^^�C�H�@��	�"�V9�G�ڮh#��0�m�Y²�ͤ�K�ɟ�aI+�vg�7�ͮ�/|Ǖtt���*��Xq�Kg��)����č��������y'�m�Yu��FI��W��[��KNn�Òu�o�8�Iւ�A4�$�Zw����<<8���iap���=~�83���].t�M����0�l���ݮ�������	Ǉ\vѐ�[u��?<ݰ�H�?<�.ϻ���szM��vC�+���-b�P�)~o���nC+��7�|����!"�i ��DJ	ʪa���gAK�s+XĄ�U��G����t���
t:���ّe��>�w7���@3uF���;7i�i�M��E�"nvkr��|*E@t��-�JZ��̓� ���9E��\[uͼ�?޻u�ƣ�������56���q*vG��4"'�[5NP��� I��DC�|�y��^X�yu����G�R��I�o�������>��t���ѧ�g��1��u'+�:�c$j}���D�i�\=Y�1-nh+~����X1z>_r�GQ�M@������Щzi��i�q�u[r��ԠH!+���xDK}�Yc�kU��kyG%ؖ@�A阚�n�8aAg��8�9��٠h�-}8�����g�}��~���bew�B����-@@�`��%eRi?K���K�f�y���Xc$�`$i9���x  ��IDAT �Ϛ�=7L�cA\���J�Cb��gdm:��͚ܜghy|�O|X�6tLT�@�-f�	/G����i�&��}=-l�n�^h;��P�0[�q�sQp��6��dҦ&�&�L��榫\��o"�>�ƪn�B.;�j��\�xb9Y�Vx����lڴ�o��?��������]�YN�c4hC�i`H� ғX�K�#�6��4)�:Y�9�I!{B���(���W.+�8�ԄZ0JfYG6�t�����Cd���0s���jX������&��x:������=y���-�����j�ڶY͟v��J��=ˬ�YG�i1��d��i`F�9��P�/��i���$�;t��
%l G-���Ь�ˮ��͖���j�T��>�}���8�,(Q�M�{%��T���3+���u�q�A�"��wqbW����y9>�_%�
8�>��$�}�=�g��h�@����U�s�X,r�ez/�gtH�7~��?� M�hO��^f,:Fu)��^m*.��K`@H�TD�����Ҹ�g�`/�&��_E���Ǹ�v�2C0�j��A���Ƌm'G�^I�ţ�z��4�d*�vO@s&�.8� A���� �T#�������CU�h��Q;6���i���ȴ
x���)~�ؙ|�Э�0��!���@?�����A�Ǭ	��ٍՊI{��������J˹Z������*�E�!(d[���g� |{�Y�հ�J���[eR�v��o�Y$��Oh�(itr J{���iQO�F�A��"v��޴����dN�8��ɫ1H5�\�#���R��uŘJN�(K�ø[�UpkU/�Ul�0ZöZ֡��_Gz��{���\�}e������C���������ϱU�S����Jnq����"����;U����v�+/�
�!�7�ba�0D����	��M�ײ��d���i�sԮd�PfDmc�
f6�<8�@��J�AN9�H�a����T��P��k�VsMκמk�v�a6��)���cؑi���צb��(29>��
�p�LH�YG?e�_�(�P�����4#߮�����{��f�H�$K����� �	Y�Q$��tN@�����ʡ�fy&=g�.i�/��Eʴ�,w�:�{p�Ҝ�?��I'����<gV :fBYc6���A�=�M=�-������C��|K���֏�C�n����>"�I�:�K`M"��B��t&H��C�_�����_|�Er�eY�����Z�����3�9��������	�fVH���q.Lv��-��F	��df��Ľ�y~i/�Vz@߼y��]�U��`��KTV���ZM�4���,�a�'F�����dű�{�)h��	\)i���e��u�7���x�>�@�Cn�͕#@ꟿ�\KA�*�*�d�̔���J	��9tIE����YP��^�4bm�{�I]�����L��j�aGT��p��T6"�;<<�G����MaI ��06��0}�+x)�ߍ^��ɳ�ʄq$�)্�!�C��l&]!�S\�Vk�\X䮍�$�$yi`d��2��vw�Y��R���K켳3%J����K�6Q=8ܣk&_�.���D��gQe���N�{���($��Cn�̠�ΘV�;w�/�&���4�@��J�D3�4D����A9�Xl4���r�8�7p2�gNgF� )�2���)�+�p���6+4��yV^[!/%[I9�U�
��Q�<*��I̌pJ�?pa5�2�W�E��BzeA��`qB�v��͛ǯ��:����}-~P������Ϙ#��1�1��h����]�ѣG�+���4ڐ�k�A�6���̣�5E2N�<O�>�ާ#��&m��?}T"�����b�p�c���5�*h$�	"�ͦD�uStʖ�(��e�n�Qy+���JΜ^3�48}�9��lP}\�|Ƥi�gϞ�}�C��<�������|q��gb�F�7k�ܲ��X�q��1��@�p�I@Ir��X��j� �%En0��3�>RP��N$xҧ<��mg�0ġԎZ��S�2�����	���З��is��9t�b����8�[���b�%��A�rp�6�p;9�+��v���~������?��O��O�d��{��! t�d&6��F�z^�5�0�NB'8T�?�M���Qa���<�n�}��ӓ�V8�Q�[6J��l���#��3�ޢ<V�1~%.e]�7�D�B!�^�����b�=��<�6�T��Q��
4�������;8�<P,ئז��3A��Q�T����&���'8r~pG1�ҿ.7'�U$�K����Y�Q�rY��yM�^�똅�:��"��jT�G���5Q�a��=��O����_���R����?����Ĥ�c� ;-�Tl��d�B%p�̳�FIƛ��]Cx+ʲ�0�
KZWEQ[�՚ʊ�Apb��v�f���� �?N.�/%���Exb�R�|�d:k��y��	<+�A���Wn$�EQ*�
E�_3����78ڸ`�q��(ؠ�0���X�t�tB�̅�h�q�sk;ׂY���\�u�e�3��g��4�dQ�@v��!����z?��a�D8��2� �Y��}�-*�@��0Jx�+�#�Z(�-N+���~*�W04_��28{>}B�Y|U��Z">�XX�A+�%:��D/;&L��vT�򱗊�I�NU~+�::���'�{�]���Z��1���F�z18�j�=�g��+����Q6�T��+;ɞq�����1�tl���0���jz5Ζ}~�U��I��R�r!@^m�����m󍄱F���>2f"+��V�*�R}��Ii+x(��ج�`�80F;��k�m���7|>�X[6�>����ł�%[�H��|  A��OE9vM�l�ht�����u�.'fo޼��?[1�|ת���wt]4�7�f
��6}vf+p1��mG�l�s�#��-�1�lY��#�WM�b��1h5���+���	u��Ȍ�HI��>��O���2��y�ܖ��MM��Ew~�b�F��5��~x��7��]L3Š�y눹P��͜�M�ct��$!c�2���Ж�9˄BpZk0��͖�X-�<�@7s�C����F�;�e�깤dyͤ�n��r���4W�|���M{���`�)��Kf\=��a�L����r����^���`�`��N�$�ck�d�%D
�IY`.oL�Cmw+!�c##�T�hxIݳ��BP�8������a�N(Nx���ӛ{Gǳ錬Y��x"|�Ie����06Jrf�lryLb/LL�	f�Jc5������8�=�.]��w`^#a�*&Sp�Q"�����=�7D�|¸���RVD~~	)���0�kʬ��K�%7�µ�����/��䬑Y=���e���D�������xD�1>����R��.��b�0"+ye���S���dGmUU���R��Wj$ߋ�_�(�msk�U�]{�U�҇���m�(ȹ�8��`-��(9�)ڭ��蓘F.ʹ999�oC��rIk���Ļ�*�\�(+2�!�`%i�>�*�b�Y_�	aR��n�O!}��Nw���)}���>"'
�i�ٮ��F���k�(�句��5��Ȟ߾}�~}��9�[FQX��B�]��ul�i��R-p�#���J�,K*���h�|s{����\C��Z5����1H���=x8Hà����ʕX��jd��) ��Tu�6ۍ��O��A�����,.A�m�^���ZiG&[5za�����(�i&�N���:t��������TS�n�=����r�����Ȅѐ"dj�'�Z�`<�&t V���X�yC�I?\-�?}�ڬ��8i̥4���������?��G�A�L1��v�?��V>�ĵ ਡEo�z݌�'p�hQ���U�j��>Q����`A4�����4hIi2�V�0�����Z���-�4*��;T�e6�|/ PP͙��0�d^�Wכ��!K������Z^o�{�������5�p�{#�.��P�K��LLV��5�裝��X%������Az��0�Xh�Ӟ#_ʐ|�G)l^�[?�����2a*�L+[�3�Rz�u1�胸�kX��l�\�;u�=�(��f�/�CΔ�F����2�����yۼ(%)]�i����&|���5<�OiA·�/�Z��:�P��y4_~�գG�X�,ޅv��Y�`(I* �F�X��1�*C��٬??oIV50�"��P�GW�~��<v�RI����` �I� "Z��E֢ߛ�W��r8�x�<�[m#�<rH�t5��C��(L�J��!:mY㽖N�9j�c<��7����'M��Z"BW�Lg��ZU볻�g�;�:K�+ayS��B���Ѐ_zqq�����_�M���wY���2�!������,�w�Z��s3�ڹQ|��
�{Ȃ�tɫ�5yI��Mjk��r�砹ms�8�� �4��
� ��L��;g�J*E��Ї�FT�-`b�b�ا��c�0>x���^��FƘC���$�n�@H/>::�	�v.�)�xgu}��x|%��,���R ��<��<_?�x�������<d^+�l���#n&�nW{R�T�Y4i���d<=ROr��E�4�L�u���KM{\ш�_�@�c� �rX����B3�;J�9�煦cSn`P���Ɍ<���<���i�ys�)�3رR�!�	����mZ�X>�
҆��X�`lSHiYU3:T1�32,��ck̢��N<����ҺwP�A=ˑ�5�C`ؙ/�oV*E7(�� �<�6.6_<����|�w�T05icb��mMD،⍠����%)�[8c�;Dm+�i�WU��U�E�*�y,!f��E��K���(H�I1_@�Yѩ
6���s o��Ɛ�E�2J����^��Ze��⿰˽I�U�W�-����B�N1PK<:�V��e�ٴ��k�+CA?@Z;͋N�岰�%2A�>�$�W^1"�<J��f9I���l�EuA�&],T�E�&7��E�� �B�U��C� �=q�C���\�I�	�Z���؈�(h���c+�*ڛ�tfت4�j�c� s+���نH����}�28X�����/�>���o���[ǋ��Q�`����g��3[�Z�&e���;�y��Wj^�ڧ�
���94Vo<�*�;��T�`���cz;�H�㝬^v�����qL|�h�ܰ�5���U�1?<lݒ`7���v4�<���Kk�M �Ȱp��T{�JMYc�I��(G���V<�Dj�"* J�A2u��7O�޽���Ȼ�"mZ��^���I/q��J|`]��I�ɷ��� &��lv=}�������N;��q��r-˒/�f����v���e�w[.|���r������]7�6p�ܗm4Q���*��4���Jⓠ2�����7h%@.��(6���IWh�T�eXc����B�0�I荒�g:�t%\�.>���9N=z��N���Yq ��@a�,�܊ѦN6m\�A0���Q��V7�R��e�":&��)�t9{mV��,�x�𨏌+�W�
�;V�'��ȷ"ch�Z��5�dk訽s�.���韸?��a>X�qd�W��~�z�JCǘ��3�;��Ԏbʎ�E)�bmu/�R�Ad`4��ʎ�:�:U`!�
*1�c+�뜋��s�NH��'O��]�T�^O���HfTv='�6`<�*��^��2�tИ���;ת��C@�����b�p�K6~R���_��B�v�Ƭr��:t~봏g�
����{���b'-t��Cx��Y�c��R��ô�l����(��o�ܬ����|�����V�?�ΌC������k��:�hӇC��� )��|e>���x�MMx��,&A@�}g�n��$6�������
J/Y��LQ�𱐻<�����]���}Qi��Jj��Hx�l����'��(?��������4\O�p�8��@cx��n�(��M B��g�e�����N�G���w^X��v��I���h��` k�o)s�țG���k�Ǉ'�����5�Ȼ���J�'�z]h2z)Ej�7�`E�&�H�����`�J�ת�U��"��^�#��d1@	4�o��6�>� �(0��(ˡ "�o�[?��O�����]ϟ_�М�����I�cBf�g/�]ZT���vs[/��*��)Xrd�%˂��Q�9�����Q3^pob�Y�?!dG�Ֆ�8�.%_�G;Z �Nυ�1L3����k�)"}3��׮n�0ݘ�F9ŝI�۟��Q �m��] �	�n]-/0��dY쉅��ν���4�e�-�^[Qc_�E`�gP���h@P#��l_�0���#7h7a��:�=���iXcWX?eˀ��iC��xA�A
�ñ���g]�pҽ�'A��+��}F�eæ��:&A?���t6�%�h`R],���'F�����Yi��(8�Yx���� ���"�Άm�{��O���.�e�j�����/� �.@���r���?��h�C���.:�?��#�h4�V'����+��o��������)c[<#���O���l?71�m��r�E�/P*�_i��U�M�9P�L������Q�j_H��;�-�^�l)ڌ����2Rp
kDEܰM\Q�z��Ҩt�+W��֪Wb�:� �\��B��cDթoj���+�$I���q:J5hrA9E�F�_:-Ƴ����`�)����b8��(Ʈ�t�̱���%�F��� ڜo`��|��"KwX�R)�.)[�Q1�^��yğ��+�=A�X�Zǅ�r�M��KUԫg�)��ݲ�_�"��&�����dڂE�0����d�池=eA�I�r�����ń�����C��2Y�[kScw:���6�9�����N�-�3!S�z'G)����p�@+��� ��?�R��$'�'ta�}���\���*��ۨ�ɒ�tRw�����믞�׭Po
�ևB���wWW�B-T�sou5�1]N}���"W���-J�c�:;��Y���+ų�B��������ds���gǨ��<w��>=�{덇o��ڍ�a�麝H�U��3���O�0��`��jl�]��t�R�b�P�Zz3H�H�����Q�Iuu���ZἙ͛~p�9�^�;t�i�&u������^P��u�pD�pٮ�k:��<}�5S�(¶Y������$�v�T�Μe��0����o 󀿢Ql�*�x1���LvS��#�p��Q�LK��N����Z�,��H$��kM����1�Uq;;\�wpp���~���
d
ڪ��W�%!݂�����̵�2F�*���ZmF}
�^��W2˃��Aب���I��Nh�n��4̑y����'���M˒+�m�}(�`����)��o<���ꫯ..iz/�1�ԮkO��hd�T����z�9	+�BT\i�WI�"<<\���ϥ
����xfH�P�� ����i;�\$�;@��<�A��B �17YkP�Y������)z1k��e@��|P�[����hdfV��8��s&���X�[G�3@�J�A7'?dk�%q�Q�S�����05�HQ$�!����Ԃ.�e��v2ihN<xp��M�rZ,h�<}���Q���!]����\n(�`v���vf�Y��]�� �i�!���;@A({�ql�p��!`����sN�`谜���"���ɳ(	��/��u�f?J���=�I҉FP)WX.��t�-חW��M�I���zA�R-5s^i`�8ΜT(
��7S�H�G;��6Wm�83�w$�_tf�d��F:�޽{�}$�'���|�{���9zˏ��_��m��������FrROe�ͽ��=��=�dJ�.�������������)��b�w||9]12�b�E�Z��c׺͖pF��NSV�Zn�đ���B �u�&�6�F�)�z�����u��9��^�����"��K��̃mp+���0��1�&�E%�,��.�q��X�;���ӵ|Ŝd�ټ��!m�h�o;!��=9��m�#Z���Q�O4ݳٴ����uUe�����lxIx`
��=�@b�^�J��̇����l<���h�u���pQi}�'��_�΃�^7,;�4{G�U�ڰ=�/��0�fp��C� @\23�Z�C{M�	�1|�Ь����㤑F��ݶk��d8��Ƚ$�Z��� �D}@�h�rZLC7(/�⑺�mME���~�3TY�mR����w��ݻPr8����/	�7B��e&+��Z{8�-@�~A;����^�O d���t�I��J�/u|MW��������=���|�	zj��ț�R�	�ڿX�k"���r�]ף06����X-�r�Dժ�N#��
�oqy~am\���n��T[RI9'�\���)�í��*9Z�`h�UǤ��FH����G��3�opgk}���1ڃ�Tі��;�iG�Z��E���c9����ъ�\���1ŸMԱ hyP�)lY��򈅖�M�/�5]]]�I�61r�(���#� ���i��cN���J���3���{�n��V��j�N�:�<������{�T6�3������7SfA%�N��z�	���iM���>�5y���
�N6��@���O�<��O������Ept7n�X�9�Ev�c��g�&��0^!��yd�����޿
l �ȼ}fr�mf{2!g�v߃���Ǚ�J�cB�g�O;E����adAC.z$��D�@��n��k�|�)�1D�ƾ�N!�q t��|�Q���v�f���\�-�T@�%r4�zU�P�_�íڬ�^���o�/�"�2/���)����./���A��Y���~�ؓ��\{���n[���E#3_0�����{��»l�º�Qj��2d�~:\,���l��(��D��k�%Vڐ;s� s�|W,LɐW�6ݳe�v?$WЦ*M�%�Q�PK6����}�Q�d���n��b��ű�.�l[a�3���-O��~�tT��W �rG�p�-����נ�@��X �іJ _��1�PIۊ�#�B��e�_�+S��I��z�U*����,��>��݊�&hE�J}�~�/��ɷ2��$1H��1��Ӫ��N���e��_�X'���/ ��u�4r)�}���8��?������ۯ5G�e������K�4�s�0�Ϩ���#�+]3ᑼ�>y{P�h�˛�b�kɆ7�ŏ|^y6c�E&�{M�F�0�kl/�B&��Y\�-�xQ?�[0t@ؔ=�*����U�N��k,6	x�W�-�XҰ�G+�L�A��|�G�q �x�P�{L4��I�v@T�$��H�Qa���>Ph�
r�2�3��O��TK����b����Cޛ�����۷n�P�M�37tV�^���cT������o�G)�+�0C��^ŕ�qB۞zU�>%m }�����sFfQ ۥ@{������%��}@�؟_0�s*<#�׫K����K͵�*��C$��M����//7Q�U!+�i�0���uC��#X�N+X�ȴ��E�1B
�N����J7� �d1��oݺ�$z��y ��U쵿�z@���3�B H����ꊋ�4�x[�m;&3Rl��L���ѴR8�3f�y(�{���,���B,���cTEɏ���F� �D<c�^h;�� a�|�!�"���l�p7_�'�d�%"�V|t��� ���sDz��Y��J`���,�j�U�c�)�ï�'�)Y��Y���D�9���p�v���Vzv���;���%��?�c���
ٵ<q�O��E�6�_��wY��c��x1�QX4P���2�[�>�&��»�N3[_��lV��m:��?�����ߺ�.�et�������{������յ�[p,2dsE���Mnq���,B]�� �DEl��bUD�n��AS��3�im�,8��v�������\s`d��+�]�fb�eR9W�zO)���L�|,Gw�X���%$�ֈ�O;I)���\if�a���
	3y97M�"�5��a,�0k�{/�f�(pdԙ���YQ�@��3�����BI��A�^���_r=�Wm��:iqC?�&"c�rW����_�;E!:m��" ���5ǀ��潓�2��~�s�s��}M+�vU��B_�w�i��]yk�m��P��]���BA�(����O?].�����ҵ���?�ۿ�[z�w���~���45'�4,��3:&���>}\+�����,�\�b6�Z �d3�"��=zD�����A����2��?=�!��5���/�?d}z1��~�z��-t����_��_=z�$r�'�o�G���TY8P��&;�iu�iSAA�J�0��ߢ��������W:�R.@XI\�6P饏����[���&=�Zo��ñ`�viW��c������9�8������v�P9���}p���:��f�{�ɪqa�j�0Ôp�C���!�)@�U�n6��㳕iQ�Sn&��T��?Zll�e�Z �s\w�iE�o�jm���Fu6p%�.%�˴>��ذ��y�R��TG��} hh�l��ƾ�|��.b�V[$�ڷ�6f���*��>�<� F;D� @��cAs�������ﾋ1���Tt�������gt��������k���5'}����Jt��Se��@~�,K�eؕ�NFx'g� �O� `����C$2�p�2�6�>9���7��HA3�l Z����ȷ�w�p�X�m�+wm�ڠ�^�g-��U��!#-�$~@A�(��2�:2�U�ޔ�T�e���:h���)�.f���X��"�s�x}d�Nߚ{���U�>�}��:�S��tJ��B�63�bw*Y��+�x��e�F��mm�K�5i���c�Ь�M	�B�����jC�$���J�H��P�N
�y%-"�Tz�f'�~��j��������� c�?�����ٖ�|;�0�S� H��G�}WU���%��L6�ѶW���Q��D-��UZ�<��
����g<dP9UW� NUtBǦ.1�EY͋�f]d�	�0Q�e�ژ, �յ�h$)ʛ�i	�}��}������#C0���<��i�(
hq���)q,=��e8CO����
�Fl݁$Rk
��ٯ�Zz1d�Aׇ��޽{x�O���_��szz,��n�Į���# ���ޜ���F�TƘzNIۿ������x�w~������j�kw`�8�2�
U�G�Ӗ8QS1��T��A�Y���!jn�s�n��\��ѓ����C��$���G׳�wU�붝�\0����3��;K�	W"^.�Ł[ N%�	��U� ��_/����ջee�i�g��1U��銗�5�8�a�1�F��H���tڇ+�֚)��6���^Ib6f�������Q|2�&��I��X*$5;,��|�maL����GR�2�&c=E���f3z�0���j*�<V/��E�K�j�ًti���ܜ��9�F(^ �F�����44�%y3��5���V����?/�@<+�*8��t2�߶��zo1�?򗫁�<�n.�_Ф�}`8i{��d���i!*�aLm.�QP}#%�ǡ�5�[{�� ��S��N�D�$mɌ��@��4��ʠ-&�O�t"f���!u�E���NR�]��X0(M2�Y��2 `��}��b��F��K�E�N�`+h55s���4Vۈ ( �7n�ɲ����Ȩ��� '�y��A:F�w�$`��3��ŐA���̅�>^^]�_��-�xg�bL�}.�r`Mb�b�&�+Y��U�@���aL��n����Cl�(�����ώT�������4�Gz����b�+M�����P���M��!]����9���B��*��+ٮ7������#t��1-�n��CO&�)~-�C��)�3:#�YC���P��k���-���bYR��|$'����i�cq�������x�ޭ��AF/�{�v3������:�����I�M�N�M�2�n>��>,f<�t����*��������t� s1�흞�t\����<�;|������v�.l>;�o߻��=�l�ݤ��W�mV��R����'0�T*@�^L7��|�*�݂�1�F	�@� ���R+�����sb�/ˌ��C��Jv0�L����f'��h�M�uxy�����}�4EȚ���|>o����y.	"��l:��ٜ+ևԯ6˶�.�f�g�|�rH`�hK��$^\�Qt�"��Q�� /��s�MeD���a���=�.P�Vd.����x�%�G�C*���i��ly�Ɏ��t�li��(���d���<6���U�"-��wn?���M{��9u#s��޲c�XP��+rz�Ģ�\��	���Hc!TW(�����Y�m�q&�֞Θ'�;uk�p��,�[2RdH/���F�!Al��o��(���`��a�XB��F����Y�(��,Vխ;e�9�i��񭈳�R�}PU��<g��׊�_���E[e��L�=)�O>���ޣ��;��;t�_���߿O�B�Ȳ=����@Ʉ����}��e&ׁE���7���[�X@Ύ?�-x,��U!�szƘ���]�#��SC��/WR�Ș���t����}���|��bA��fZ\�!S���.����r��(��2���/��乶�w~��P䐿:�l���r3r�V�i��ٳ��|���t0,W��o���P�S���T���O/,��h��?JqPj�S�g簀tL��׵w�l�Xκj�VJR�yQ�7iҊ����ـ3�d+��RQƬo��#�J�T� ��X+0ؤ�q�7�\�;�JyH���s����~H�-��*}���Pg@���D�-��o5Q��	�K̚��pq���ٷ���eB��C��0�.�z�B��᩵��m�!(�u
R��
�J4	���U�,&nǙ�Z+��Wzj���:�(;�k>�x��	]-��O&[&4�?�W^��洷�����*E��b���O�h���
��m�S5]%a���e�8e�nă%Cz�l�E���ػm���)���7�l*��68>s�z64X��������l	�M���أN�c
�R�lwڶU1aK,zR�"�)W�̧M�����hj��D�b�!(Y�IT�K�L�
����^S3V��X�� ū�Q��� M\@�1XY��^8V��.��'+�[8	�D�V
��-J�s�-9�i#��\R?����Z����������y�fl0豛+���%j\m���������۲���q1 EoL���fN+���If��G*h}�2��0B���L� ��f,C�[5���w�z�f�c�,�aˈ�)�n�D*�ETZ�p�ks7Ni��Vr�}��Vb�,vFwZ |@x�R(d�.�E�p�g���kZ��r�v@<�)�7˪^!��|�^� Tz'''����|K�H-re�]Њ7��~쁳����(�|q|�2�:��9�F1���Y)|=S�+����}���:�<9��V[T��9FZ�!�t<4>9�7o���׿J~���T�I�/y|%=�-Rt�\�i��&3��u�(s}n �8��֡���J<!Z����?~�x~�D�E�	f@�8U�;q~|v��
npd,��	<�ժ����$���ō��jU�%�����`؎&�3^��d`Y��0-���Co�j����})�'}[[�b�H�����5yݿ���ۣB�BR��Q�ib��>��S�)H�����>��]��j̰� .�h%r�鏳�g��!�*�J���\Ezr�A�9�։3-� ��h:2��)/�p�\��`�����E�t��RitS���s��_I��pa.!���b��/���5j�z  `��b�+��A�
T��Ν;w�ޥ�~��E�m�x:��޸q.r�l�����_A��X��K�������0;H+ٷ�{�|�"�+��pX�����)��n�g't?����pBC�+$���)ˈ�e�}Fo��üB��F�C�P��Dl�U�j��y��@�G�� x˹#�H�#��,� S����%ܙm��ˊ[YOOι?�I������N��1D�Yol2}7n�؞L�j�U���HA`�K�&�?���qN�$�(�j:�l)P�A���M��R�|$"��f	�Wpl T<Qtͪ�䍮s�w�X@!,��	)}8�g�]H�l�N�0��#W��t4�<�t{)A3���X1�A+���7�O��]y�D�>
c�����?����՟��>{zHJ�[�%�i����D����@
�=�g�(�0�k-��gi���P$h���^P�µO��w�α[,�Й,�XH�c�����4��B���`P�"�z�sba@��S�,$�f�dĥ�B�=�0�%�$k����b��f\��r����p���\_�/��{lt��RТNၝ�^^D4�ݘIB"�dj2ڈ��@�����w ٠�<��֩�E�
��b9')��i��g��mzS��QǵB�ClVcG�nC�� k�/�@�K�A	Ƞ�ѿiQ	�s��0�W `��JMQ[%#�9����#i�w$���iz���Y�
���z6������K��і���[،H���C �ʌ�h4f+�F.#"'H�����"ő�u��Ç�>}���}����'��P��WZ��3R���YN�|����\�����������M���<{���������`b��
���m�X�ed��O~Q�7V�^���C�������r�붆Ko�z'2;Vp�5	��b8xP2��@��6�D^ꋠ�3c�v�d��jk���Ȕ ����)M��5U >jiC�B'�DQQ�5��7�b�ڸRb>�;�������k̖z�6���2�s"�zd^P�2��:� ���0h~�t�^�v*h�B�~��D7Хi����Fg�a� �d�aD"��eә�}��-���8�^ف�������B����d"�q��nç��C]�I	�=Q��Ͽ
G�l�����&4|�#3����H~�x1�io|(�gȀ��6��?��,�X�l6����z��.��4�f�c��W7Qv�~����^��N�-�vj���(�X���0�Lk��@55$~�}�)^��9�������+Q0J��mס�[0b��d� E����b�#q���r�݂�4,��m�m�R���ƈj|�d7����+t欙^��b����^]�EE}���=.O'~�=3���*�l�b%����u<Ҟ�.M��N��@d���O��j��r&ۦȝ�U(�Ħyȫ�k��91$�8\����H��a��Z�:��/L݆�ѵ���j������[ʕsʩS��c���If���ٲ;��9�����@"R��C&EF �4%a����)VZ��}I �^�S��܄�Y�0�,��İ�D����˯W����#צ<�y1``Kp��\��hҞ�)��hv��r�ߑ��6%<���4�Y�|���%J��G�?~L�:3Q<�1X����[�ˑd���e��Ӥ�Y8��Y��{G�V|~\�f����{�=|p��ݻ��9�y> ˶G�3�й�F8��f[$%�iS` ;�֌F"e�|hG�+#I&��%�ʊ�O���̼��5����j_ �D�ttTq��'uH�������������w�-�Ǐ>���vm����T����b%3���ȋfU�?krE��fí�+�y�^[	�6��%�^l&��Q�v$���i���ټ��13��~�@d���;"؟$k�g���Q�_��b�L8���ۿ~m���}}o���k
�drt�cN�ffTR�X
&Q����e�"8?+x��}i,����T��&�xE>Y�+5&'�,��%�N�z��d����'I�����,���BMà�D�hT����e9]7�`�.9Mv��%۠��*.�����I|ڲ�u��AN�^dԌ$�N�p��dn�$�B��^ȭ��"��N�r�*����ȁe% ��7���5d���8@%�H�����q&Z���Eib�	���)j�Z�����6��89��Dk]�"p�����)h-z?Ezh�"@l��Zq�@�WH����k5�S�g���E��a�{x���SXRs\�ꊧ�R`�e��{�h/����y��&�l@9�����M��w�*>?("E=��Y7��ӭ�l{*#&�WH��S�''����7����� VU�.�1C���>ߟ0L���'��X�+�[���R��
�UΫ�#U�>l1]�sv�SGBP0Y/֫m�+}�t����j�]�����uU.dִ劖c8�;���u��c�?y(3	\.�cq���r�u|�����D��!�7J>خ�ttG���W����׮]�v��-ڻ�k�0l�>\	��_|�k��w�������1�d�����H���4[��L����k>}}��vWt��:��&c�$�`h���e����9���)e��F�CF#L�U�OQ��[�'Y�o!ς�W��`fDR�Ы��:�B���|�y�Gͣ�o�*41�DkH�nM�,�Ra�)��0jv6�Y+$+Š�8'?��e6�qx�g����b#�\�ҢM]�0��ٔ�<�>K���j]5��=����c��w��.��ݻw����x�Y�����w�Y��ʎ%�d�zFt�)���4�K��Dd����ݐL1�S�J�h���yC��X�,����L�	7�p)7��M�1-��3��r%)N���h�����#��l҂��2����b�F�mOEՔ�r��Ƕ��ঠ�k��
=�����!��$��<|���7_�����?�'SĆ8��)7B2�L;��J�]�X�ȝ	;�3�$i��r�pT ����&y.��0�	�0$o�6�R�e���h6W|�����NQ���_�w6��ۿ������'wmU��7�Ȓ�\�T�#��݅���
t��ã�?�����©M{�:A��,i0ZF����pF�o�����K�k`s�2i݀2u�)�k�g��0/1bByC��88��V;������V�;)i���S�M��z�E�k�\���9BbED0��?0s�Ad��J�ry�=�)CuydAC�J�p���'���>�ߋv�h��ak'>�8���H;�a�+@�9c��~�� |9|;�'SH����&�S�*��F\�~K����(ey:p�1��)(J�QҞ~j�P��8K��/�2&��>7��< �:&�9?�MI�:��H�Pe�۰��!���.fq��"ʓ�����]m$�!Q�O�/����R$D@��C�"^\'�)�&�"c��F�<�3&Q�P��.�v���Ȉr�@5?jc�tk�%qY��)�W�!1WkUX���k����Z�6˴ս��ң;�)�4e�#5֟ޛ��v|Z��W��]/y�Y~�1E`�`
��\��y�]%������':���H��^\���X"�P��>���bU�LG���d5�Naf�4u�J?�Hl
x�x8���B�䲭ی��|�S����e�!�5�n�2{����;��2{io�sG�rb�����3\H:c���-ў����^��Z��g��! ���+!�ml�;qv�u�^�:��"�v��E��Q�I���n�N#�Cd�c7��T�s�2N�Iu�K�n����tS�u2:M�S��|��rH@� �ex��77�Ҕ���ƣ� ��LL��x����#�lA�&�����Aq��B�08���h�M�t�v'q�f����~ ��a� �Y++�%���f���Q���F����%Ϡe�\�g�m��x �	���rd*1��4HVQ�W�V�BC�,��o��oܻw�Ƶ]�#r��-�gY��`7T�AS��bB��6VƄZ"�ϋc�e�.��l5�֋�I�c&|�8?���L����ϟ<ea���rH:81d&S,C���ךT���	Ih�F�vF�J�%��a�|t�f����l�@;)Vx�ѓ�ǉC��m0.0k{��H�h;0Kb݀��󁌏��1B��on�,;�>I~���Q��J���x�eT��/������G�GA�i~�a��m�Ĺ)�c�,������[C�M�3��y���upW�Ƨ������I9;��/}/�T�g"{�֥9몔�F �"��>Db��:��}z���G�W�'Onwo/Qf�@�lL\�\����i;p�Q~O�@*j��2	���D�P��|wB��N(DP���!e�&��}Z�4a���(�	��C�����
]�u�����c�x�E��� G�Al@���d-�Ѧ���V���B)��x���L�l_tAL5�����D��^�Ï!'p����N9�kU�Z���d�I��*7Bt�����8�]c�"�A�;;�B]0Ӣ�h�LzM��h=f�إ�'"Ƚ�;y!�w.)D~2�YQ����r�Rp�� �,�`E�	?�����m�Kα���� ����@�i�H�b�+}|�rչ,��h;��G��zş�W��_޹s��Ç�L&��y�C�nU4��AZ�o|��b�g�gR�Ć �>g��L�޽K1�i����"�f;��@F0/�[D�|��e	q�H7���gjĴh�3�8-�[o�E_D�����:���lb�F��:��{�b����=��q�l��
J`(�IK�2�<9�7"�4�W�J��ԠI񭎹��!��iS�V��-���:0`�@�Zs:�y%��R!���˂}��Eno�B��sڗ�^MY�j���8�l&H*ge[q���u)�<7�P�%�hF�E4@���B��Vk�̀����ς�6�S�!�>ơ^��{T�dX	��b�Dj6���$:�tp����wߥA�T�t� �x�e�q�	E�I�V�DE-�ѓ�޹��e:O���C�b��Z�h���L�� /Z?�6O��芲���g�}F'��?���sE��$m'��
i�Dq�(�[t&�v� �鴁������:�r˚�e��{���L^�E�/�����3Jt��_��Z���(t2x+�1�}1D�.18!2�tگk�\���L[����L���kw�ב�ؑV��80�Y���s?��-F�2�R��E6��"V�D�P8%Q��FxkR+S���O�%�����c극.��%Cǫ��T1�Ա�v| ��H�2x˙Rd��E��i��m�W3й�=�ø7
�l��o�g�
�$�m�}ؒ�R�]A�1�̾�R����AJt��a�p�}������qf��!=�믿��"7�v���C��98���].3�@��B�Y����rf����зhf}�,C`2i(D:~k<�tG����G/�?��n�"s�f�)��z����\;��xx[���tx�8�A�����~�S�7�~����M9�*��=�eډ�Q�v�|T�і���Gچ���h�Vg!X����kmo��«і|��s|]�m|�ԧ�׸Aas{�&�e�=���&�{,��/���htƐ����1�-�����/�܆>�BJsS��Pi�
�8U�έy�^��̍��w�
��P6�{[E1��N���O��$������z^@,p�]���lך�#��RP	�L��;����!Y:W�~�R��]�kh�#�g�DC�eUy�٤_f
�{<�h�)�2��6r#��ǩ,5T�g���v��i$�:Mņ^��y��D�'��X[�CX�=�F�Z�w�^8�{]C_pΨ�����#W�j��"���~�eI��9e-i�v]�5l�4R���7Ӌ7p3��(����d��a�$3���/��@֓�L�s	%s�	��TJ_���*���\�"#[�K(�=oR�E� H4X_��)0Ҥ��8��7�o����n^��P�InZ�	��p�ǉ�ƂտE.sj��r�h��s�Q�ښ�8N�X\�����R�>����O����YZOO�NN�g���G'y���;w���|�	畺X��#��l�:�C0a`�פ9�J����V-�T|R\2����p���)�ǣKZӆA+N��=�qN���ܥ'���Se�&!��������ŀE��l{��\[�L&��I�$n��V��9���d��u�3;�A1��ݾ�s}{g�si�x�Ww		�� r��$Z��������l�Ȕ-�6l��-sA��ٸ^PL��~��G���&�?99c��G����[��0����;{�12�p�4=:>+VƂ��`���Е<2-�4З�usrv�����m4��F�D|N�'�|�Iǿ!yE���O�Jy������eh[�:1w>1|n �ra`;n,����d1�s�F�ހ�0I�AP����R$��Zf�x8�8���$5r~cGO%�5�ԥ�V:�Ӭ��j<B�ZgsA��y
E�� �����Z{Rk ��z~&h�&��ΔQ�*H��'���x��B�̂$�R��������m���	��x4�?!e�-:�d׸- �6Z�2���~e���6�!y�Z2-
L��q{��I&)��C�	��Yf���1�l�n~�m�!�I{��\��G/s(�9Ib�D��z���7#���a��U������;:�����&���O�rWm���b~F�DO:��Ԗ�j��j�H��*G�^�K�#h���n�d����a�a#�vc��~�������l����v���Պ��h�M�,�.)��ٖ�nѢ����g6KM�X_V2?j�\Е��g��U26H��$29o���dt ����sy�2V��X	�g �x2��ds��x4i�7d�&����%MU,���vww�ig��_-�k�es��ȏ��N��O��"׼��w:��=����l6����~�5#9���]^,��xv�|(�R��1HY�~%�SҜRm�.�8�,���k0�p�u!���|�\T������={�=
  s�v����ud|�]�Q�
Ĕ�c'��[�l����."��m�0bn2ĸ�=������uRjM�G��/�)H"���ц�c���q�����bI�\N��3�uhi�y�555�λ�cp=��$�}��M���I%������P��Ds�%M��H�v4b������w��BQ�(o��g�>�=�/���\�t&���Q��>�+����.O&���Tpɋv��[���Z��<u>���Q8U�Ғ���k�˥3!n�,f�_,��)Wa���R�ֹ��X�<<�ୃy��`+��g��(ޒ�3�Ĕ4y8dX���Lg�ƺ{�.y<8�}�,gF<:��I�ӧO���Ȍ�L?v�s�^H���Xwa��]q��y���Q�֒6�1�R�(���l:8Z(z�C�hV�tY1z���/���H��ĩ�L!��iK����E��h��ϊ"�׫fP�|\P���~"`V�%[#��HI)�N�%:\���L��	�u�;�*Մ�	��J��4���u�&'��ò#����`��L������lΘ�f�Ց��"[�$'���8�(��"�_���i�^=/��j$�p:���N���H!,�π��Im�
�L�2L,�cy�Vq^�m��$R9�%KAnѭ[�\d�Z޹u�5���YtP�j=��y�=����X�¡�:_Z��X�(:��?W_�M["�d2�˨���a!ٍ�Q\, �:!v�t��2�3]�?�� g�wh�j�	s6N;�OL^G���2$�Ω����.M��tMR}�{	Ґ�<ɬ�E���� 3������ܩE��o�t):\t^��$T	:#��d��.�����Ѕ���z�*[
(L� #�.w���E���[?����%�X�n��T�-3%��7�1�8�!~�=F?!�F�������
3�+��d�g�zX�L��I�6c���e� �#t�ZQ�r�[��K<���%QG �#ݎ��=0�P�[k،QGɦ�65��s��j�Z�b��Ml�F%��h(OM���^B ��uN�M�(Ү�=�|W�`I�Li�R($!f���J��ҥ =�(�������*����ij�W�&���:�mb�����������Z�,��W��+����=�/��Gd�sq�q'x�8K�9d 1�z��(u1k�~��#r�����?Y��2�>��4IH��D:��i�ɞ1���(u˨)F���h��<�Q�П�T�=��'-�g$��!wA�τ�e!I�F�Reρbu�
��H=�=s����ei'������P�A�HXa]�g9��&��rUx�r"7�v���u��e7�v�Bh" �L������XdD�5gj�i��ϙ������y���0�2km��(�T�=ٲ�1Il�onp��[�V��l<B~�5;	�"NH�ܓC0!����M�c�<��:��8c���k��Ś��9��nR�Ng�	
/��B�
ٰ]g����zJ�sLN�Q���Ir:cDpj&��a�g����l�h�<#���l��0�"*�:�u���x�W�H�d�]?r<ΡI�>I����R9�pM���aD5�6�v
��]�V���Jx� Q ,`�)�]H����x��o(B�� =���e�\�a�i�p��H���},V��Q�,����UEʿ��^�m��Lt�Y�/��8�"�7�0l'<������/��ЛL�~!��D�Y�=_�D���c]�lt,$z�,c���
:]{��{@�>H�S͐�!J�Y�����XNY�9�ҩ䫥�<����Ԭ�� ф���Z2�d��	]�&Sw�	���̄U��zlM@grx����ƈ��"󜙊�1~\���|�yUG�l�-�WV�g�D����o|�������/�q'�O�@�":.��ʃ��@"����,�����܏�f�#SH%ܻw�[����o< ��[~�\�6mc0� ��?5��]��w����秧�g��tct�<�J�)���m7� ����1��'����ޚk��*旌^��O=#�w#pp@�,�%�LH��[Qh��y\]�"�bR�m��9��]]����v��T��O~B"΃w�-�Z�fM%��X��-Rt.�L�'#�uT�+Ls:9>�HV���>z�O?��0�i}� ���FM�=��a^�<m��ۯ�wF���*��})����X�ظ��XO�����W��v�;ҙ�fϏ)T~��1�v�/eZ�3�!�u����Ħw:y�+��){8�q�����:�S!��D�|o'}E��������>��牽�Xd�kx���M[���cK�,��V\����0�np���q���7��HG'�+cX*sG����*R�KP�����$�N#�FBF��b��
!����b��0N�'���`�@�p[I��?�
����d�ĐG�r�������o��o.��5|��,���#�<m�c^E�Ƣ�n���r!�a��Q��%4q'0R!RIn�@N #0�A�Z�4!��kG?�!(�[�_�3�=]�;\���H��aF��plR�9	�Қ�cYY��u�v%�V	�\9�漠�++� ��''�X7Dܩ�=!Z!���C8�on
���ǖ�)dZ�I�AF/��l(
0N���Y�:<#�ס���"X������R�oJ�Pc�\A��
�s�W�zErY��k��t 3���!K�Agq6ݾ~�:	6�
z���AnY�V����k)C~�?#^���C�e�0��n�k���mv��ѣ��
��jכ�!gJ�K�pJڜ#�����=��D��&��F�[|�44��fM�*��2�n\g�m�I�)M�Y;����}o��:o�VV�p�1�	L��mt\U�V�n�i"�P�;�E��%���*�����ps��V�1in3���Jy��敺~Pw'�)���y�0��U�+��+� j�e%���芙�l���6�V������C�!	=
�Esb�1��s��g�rR�� [H�& �<�/���!��0w�uq�9�L����"��f)�)Csl/�&�����$	���v�[e�}�]���lS�r:�4ҡq���Lכ�*#��9TC�e��0o�t��۷���oSl@����}��G�v+�"'�q��[Y��Q��t�0�!k\ʃ�Hl$i)&_�%�_�����X�4ܓT�L��Ԁ�79d1cVS܅�G%�"I��D@�b�h��ô����^$�O�7�(�I��՜���Jz�d�\��w��h�D�➡��2BX���0�z��YcQ��&I���D[�����65��Wy�O�j�����S��ķg����=?[�8u\Lc2n��IUr�*�iג7C�+Å����FW�-��@�KV�2Lǥeݵ���6�c򳳲sm�V|���B�x����"]W�����I�Wʝ��CuXj���P�@0A7�o��_q[qf���,TA��)�mM|[6��H����ޭ�ݹ�5/hebCt:�D?$�W�%����1+j��ܼ�$ې08aݢ���m��Ã�gϞIb�\�����yyvvI��g�-��8CI��y���:_���rܳyF��2~�I(AM�-��X�("���|~��1m�r��Y..��#�9}��lnA(�ျP��w%1;<<$w��m{{f�D�l ~�|��j�$M+����Cz�A6���T�V�y���u��ޜ�	c�a�TV��/�O�>�;af���JJ3����nʭ)�w3K&ޢ���:����z	�&��Df��Rn�(��)^���Y �e4��p��Z����gz�D��hg)�� �$����s.��Ύ�꣰ү�Zz8"u�y�D�r�4��J����&�!W��]�L'6�As������E ,�أ�ܹC�'�x-���j�2�^���ŗË�Ǵ���#Έ��P�8��I"LB� �A���N�-M���c�F�<8�#��r�#������rB�)�jgP��z�R�0����.-�����7���/>a��N��	�C��g?\��+6�;��4ʒ%�s�(�p�,��Eg��d�ytC��H��N�9��7��K^�Ze8ܺu�_��׿���}���1��I��v8�f�p�L����8a�w5�ڡ/�s�U��i��+�Q̪:-gf�u%}N2,A&? O�<;�,[���o����ͧ�~:�d��a�灞Ið7ޔ��gL��I�ce�sm�4oHz��r���h�NQ�$�Q��ȋ�'J�z���j%��i�"�l#�t
�p�H�b�D�[�VarT�D��,��6Hz+���i��ϵ(�b��ʛ��7>������a^�Y]E�pvv�����	�
���%�e<��qab!��/Ig��Vh���=�|�X��#�5�pge�.�Ab���Jf�Ur5��7ca�N3����z��fʃ�z�D�"~����鯿������SHy��5���ϟ��?�poo����{�k_}�+�<�����3�����*�al�S�Ő���5<m�q_��;����H&�����;�$��	�4D���g�� =������9`�����:+�;�ʹ�����Y���~#ϟ�<��N ��XOC���i��uU�,�q�E7w�d�q$�	�Ueo,l������>z���;������O�%�1��#���8MCJ�;�a���P����э�Ӯ�R�������4I�Q�w�`��v.��G� �4ҵ,c�1�>�ʳ�ax��E���+�`���3km��e�I�f`SY�2��d�2F�uP��K�=��� ����ȥ�,]-�g G���Z���W�/,��&�����.dL�J�J2 Wv��,�jkʃ��L"Q.�t:�.
���wBc#�0�4��6�5H,J��m7�>(��{p�䒐^$YF�ޝ���\���r��XLצ�-儣��\�Н@�z��9���Ğ��4�r:.��ڷ������6�vQ���"w�"d��],c��׍43�'���r�O�@�ӍK2�����	��H);�s��C[8�*HRެ�
�!i���J�n�q���3-1q��H|�+0|�:���۝�A�H��Oz<W�G�fRjg�ȄG.����	A�T�m�O��u���{��P�N;��'��^ޖ�a���M����k�������!9<\f���s�K�D�|kV���B[)�Cp�q�k@	}m���3t=hO�`�`Ѿ��\�"��zM�u
:�
��E�"�B}�kF�˄��q};�N9�b��>g������R�I��X���7���)�����<'���[��&������@�P$itDf�0'����L�%�9?�Ta;)6�n�0\
)��d�)�̃�|���0��ohwH�Y�)D��:��Ai%�^9Q�
Q���_� e���l���k*�����B�����FI������:h'�\(ߡҥ���*��E�`�JVsI9
�Z�Dx���2h�i�F�����Q��9o;KRIV	օ�0
�c
> %��Ɲ X*t2XR�	p��@��#]kl��$��W�&�z,�)x��<:::=�`����OA��s�3��i�V˄���v��G	LX�����g�%���+ys�=`�`�|��������끔���\�@�cƃ��3�G�UQ��3��di��qtA�6��s���R�۸������7o�L3<���������+?�O`��Tn׫�A�"�	G��ϟg9�E���
�d��$��|Dpt��k�BGq�&�L��+av#��0�,�]���Ko�Y�r��?rxE�A*�k��YHȇ�\[��ɣ����a�f���
y���@#Us�}oov��p$���gA_'%�I�Z�8�{�:(6�x`��	� i��
�~�)��6�޽{�b@E��]��pv����:�2n�� ~Zp,2�9��8��0��a�.�C8%�����"]X�`5���уS){d)"�Ԛ�"eD�i��'V��{���(K����E��|#�pH� ��D�5�4�îu��2T��DK�V�滒	�A�:ZҜXI'�=�QF!	rШ;i�Y3Jt������0ǹ0�D-b=ؿr�� W�v�DD��cf�4ƥ�l=8 �����^������������I��2�j��5xx@��3Hc ��!)������u���pN�`~��GE�}�_�����c#�)¶a��:���	��(��!#մ�ntL3�gb����I�xA��ܠ�Y��mc
�7*v�����y�����SR+�W�I���`j�
H�6��jH[�\�؊Dat�ր�0r�aú�%�e3v��}x�F�X��"�����$:y�e��T^��Ȟ&֗*��FZ>�Px�t���֙rY����42)��4�Xa���{[��^:�붖�%z,X&�w�_�F��_�>Q�.1G�6 zF�P�+��<%5�Q�2N���O_SE9S��|#B�>q�إ��@X���Fb�N'�J8(W㧾{��7��͇�C����s8���~�B���k��Sz��^��/���Y��#`�$������o�=,P̤���t�>�sQK�W���3�0BE7�)�u�,ɲ���F�1�`Ʉݿ�+_�
�p�8��~����gϞ��~!w:3��=H�lMe7/.��k9)P^�+ې]�Q�u�����w�Ɋ�|��Q"�D�v<��Ӂt��#�|#i���S�	\�T��i��̉�RVj�U,�(2#S�J�V�}l#Z�4�e��"@7�B� ��#ގצ��ɒ8�2B�r~I��Y�����H�=��`���0N�Y�&��Zy�Y�H�hނ$�ϰJ��$K����M#S�6ۚ�8!E���'ɒ�G��Ff� Lp���e� :�Q]��C�,�N+�ϗ�����2S%j3�@%�p��4K�Xrʖ��d�.����VF�LJv{��$�$��T�^�d, HcJ���L9�_zJ�{���s�z}���D}���z.�fI?��t�d&ю]]�W�5���};f���������U<#�Bz�]y勂6Qm8lf�zn����/���e�M�!�)�]�
���&�e� ��D=������ ��Z|��v�C$��/����CN����qʸ� ��h3 ����&�^�nv`l!B��n��f���B���m�i��꘲h�s���I�C�+81����OA�dKԍ�r��,��g�ō4��Y��FF�ry	EKg���a<�Q���Tq^s�@F���T������]m �z0�D���,�P��QN�~��X�с*��V{�pI�GZ���~6'� 4&0�,��=&��:��)�T$�0���j|s�L�t2	~�!�7��/^�E�a�H�ŉ�K�����W���tk��Hu�`�A\#�I���� ��k��;�lם�َ���x���N��/�P�A�s�ߢ��������0|�g������o?�� ��ӥ/����/O����M�F���t>L���Qda{{v��M�'��	ƻ�H��'�m��7ܭ۾b�E��f��*I�*�\$A������kP�ݪ������˓�SZ���K�B�ʶH�A���� O���e��{<����ϣ�A���O��
LA@����p�i1�����<$�+t��C�x���Ca�R�:���Y�Qڴp�Ҡ��-(�ř�-5�ˀ��0�+��vu��Y~~���H��˔�Q��җ�t�U��"O�v�t/R��0��l�h'������xf#�q���:m}���x��/)n98<�,p�K�6��9?���.��@!����q��|A�7��"�9}��x]�'�q[�����ٙ].�/O���Y���[23�|����&��.�v�4��)<'�"ٕvҌ�<*(Dk�01ÍFNO_����).�jH�|RhJ2om/H�u�@WC���I�,�e.��[�n��N�A�	��k��f<]����b^	���VaN�J���%%א�Ƶ�.���L�z�#r�R^6��)�՚6M�$ThǦj�)���2>3^�A� r�)�����J��.5��D2��`���B�797�Y��L'6�ܺ!��LH���y��Q3�PJ�]����-��6]֌_Ֆ�VX��YV����<f|гLﹾ�I��(ÚX�ƹIgt��oq0��b
_��-��s�r�҂p\W
��5�
�j��<I|A�:Z!^X��0�SSdE	��i(�?98|>���<ݿu�����%��}vzv<���NzV՝�^�~�n�:�~JS��1�iY�����q���?z�闾��j��ޙp�R��A9\��1P��M�xkzvyQ5�Qa-��CRr��dLi-y�mR�@�0e���#�eS�?<��B���KV�q72���(���痟?z"�Y��-z�m���N�|g�6�%�s�*Z��@������k��3��6���g�y�L��-Y@b��n���9�&bP�N�M���A��۴�R��!7���	�J_פ�Uq��M#u�X,��k����%r|	*H���i͖�5���0fr��b.�|�5��4/c�j�g��m|�-�Ca����_F}�
�����V!)&>���XX�41>J� 	�&Y����
b0� ��;���9G�o>|���ocf��t�[OJ��LR�2�#���ֵ�/�w�͟l��~��?}����3�Gr��Bw���w��l�>�G�|�}L%�<Q������W��r��Z5�V/_��<�@8:���y4M5_.��C9(�h{k�g��U�&W��stp��������/��nBT����|�{?�����O>���D[#��2-���9��%�@vAPQ3Q�(��� ����x&>�5&�1�p��)aY�:�E�d�Cu)x�$~5��<Sg2�D!x�G.��n�x6��~�W�3^�;�cW�놃P0̆X�FCC:�y�k�e�+	�x�;ze���T.���Z��r]/�+y�k�m&Q=K.O7`��Ŋ�J3)�@t�
<�"4����@�.h;XdR���X�6H?1�P@^�����t����9���g�:q#��?�]�V�J���_z���²X�gi�F��=<�N�N!Z^2d�ɰЄ�X��_�*���,Oh�Hӳ��������N��[Z�K�ye�B�p�ʴ��Xi6,][_^p�`���ԭϖ�z�s��*K�bq�#z��lc>���I�t���o܆̔/�K�Z�aC�,MÉ����'�d�$c�iwkzzrB����H�rjA������ĩ���0����1��x��eA�V�U���,^�S��˿��'57�S�*�[��4 jH��i�~�:�D�t^N�@h�\��@�f����W?3�WGv�h'W��M7�^��Ν��]���ڠ�G6X��\���Na������̂D� ����nd���Y
�]OB���i�F���{�W��c�נ)�D�����^�$۲3^ɞ���|!-��y;���F�޶v�n8 f<_�*��Q�Fv)��7D����8�&o������_mkԂ�P')���p�2�g��B���$�2�8Qt���+�T���T9Ԡ�}A,�|�5��_�(9�r�s���-6��#*_>�*���!�M�L��\]<>�фQ�g��E[�����rs�aw����/SL�+�b�G�s�A�V�W�`�1>��X�Jh�<Z6��o�gP�yM�cq��XJ<�� ��P��P�ǅ���on%J�#P�v��S�����o��2ƪ�eU�AC�;2b{k���޿�D��)�隶G���X�\x��\[?�
"wnP��sO�΋a��'O�t�{87T�-���������@����N"\��qK �Lz���<f^�i����_E>U�G�
\�D����w�2M�//����A߇�:|�Q�y�È��$��Zg�Y:~8t:yi �sk�Qk��7:�nmM�� � !��/��Yl1H��SD�� A1�+z�J��!���I(��(�s��O�P4B�g>����Ϲ'�1[{B�9�C, H�:�]��xYl"wƍ�^�p.��n�����ժ¦�	��s��EǍH��& ���j�ׯ��C�4i�7�J8�<�V�K�� G��Kݻw�"(�����:ण�Y}��S&(	(iZke|��6��j��p&-�f�����{��,���t�!���t/��N��&:X������cg:�O��~�@�]F�.Y�T�|�����_1:4��dvZ�bcڴ�m�Ǒ��I�Τ%���/^��Er�o
�����V#�B��u�t�O#�F��ʁ/�V9#�NA��q��覉Ls�i��J'�� m�;�$�l�JpH�:	���U�̉�)sr�<i_ֲ�H�"C����e5NQ�3)!w��>I�h����_S���\����NX�x�=�+)�o}�[����?�eǰ��锬BN�QT=���J�At�z<B����]IO[�9�S|o�[P�Ky��&�X*ң�����P��J�v���nݢ5��s�H�6���!')b�Ԅ٠(���W�\Yb����՚��ȏG:^�2��v�Z���r�6����<�"�2�>[mŭ������ж��6�&D΅k�=�1���dD{D��x�3�o_�W�������Ǝ��:���J�.�b&Y<�1x_Yn�0��9�O3#R_@��6��]D~l��%�<��)�b9hNsr,*�-����l�c��Y���]`�E�"),r�g�	&�.Prb�k#X����l���6�����v!3�n�e�<��]�����w���A�0L�l2)�6�6`��V
�,�����~�m
���Z���ѣ�ǻ�����c�
�=��?�ï~���Wu��Át���Z:	G���?�s�9{�q�'�|�A ��>��9A&�8���FX�<����+�n�}���x l~�@�Ma�Cq��/���^*��������F�IC�^�lv�S�yq@�g�Z ����[ظ�tާ�I�����y�zҟ�&a��ᐓ�'��Ij@k��.H�'m����͛�K����W��1�� �Ԍl�N;�l�:� �y{J������ ��5#aH��Z��Z��F�3t8�RQG��JƗ�Q�X�T��q�����	�-g\�хYTˤ�	�Sc: �8b�{�Z�����̃��U�J��-_1 �
|'+��q��+ŀF����g]b��O��/a���x8���th4��~��� ��g(�vZ<2���V�D]�1�#��&�;`���-�6C��y��)w�:	ʸ�%�-��b��UN6���t��6e4X���&K��:��UR�<�N@JKb̮�j��s��RA��}!|O��)C�����y�vo6Ԃ���ve9ˬi*OguĴ����H1�ʙ�7�kO�s%�� ]ӷ8ɦ�4�F�+7���4eQ9g}�e�&��a�n<iү�Z���*��;���u�09��x��^�@"�e��kL�ۅt=���<Rh�V{m��hu���.�M�����F�6C�����z`�u�m+�I��+�h��l��[��
'5�JH[Lึ�� 1���Ƹ�Tڼ���v&�xu9�½�em
��ϲ�ݵ���̼�i�c�"��@��1��d��:�oH�z1B;�qʑA��Ԓ�m�f�:�=�e����N* �~�x�b<(��&?�H�_��W[�e�p����eC�4-Z盲b�φ�V�Р5��Mp�g�A�2�oJ�,����>�!��<���s� �5��� 9�,�a�����m,������:6�>®����("+R$�D�P��ғ2�𬵁NEn� '��	�i�nh�ʆV��ٕ'��I<��r�eL�U��vk�qln<̳��+�� 8�^,IRi��x2a�������\&Z�q~y1�ǪV�x<,\�7����k�>4i��K�gٔ��&��I�^^#���e�/�3�if�o���!9���|�g֤D���c>�]���u��zM�{+FT2EԺj�����I����vq�TQE�����ޕ-K�U�j�L�|2Z-k�QW�����(�ԯЬ$6�h!-TmmH�CH�aA��:�x��P��hď9?�g����d�f�Яe���>���u���.�S�0�/#���K�P�_q���jE�:�����&��� UÔ*Y���HM�
)i��܎N�Z_�^yޚ�oM�eVt
�O��|b�xp�t[�J(JM���Y���)9B#�_�kwv�~��S�GB46oD� |"y��P�k����C����3#��^�� 	�L&���������3?�M�t�����hTv䚵ň��Re)���OW�:�3F��1	;;]��1�������|1D�X0�Pf��B�����!#��l@H1m]V�gH#��;�mfoY3S!)�����k�XN�3�H���W���!�9���ř��'������%q�U�IAr֤��S�/9�2b�����r! ���Sي?]O'#6(����|����޸q�CGGGp��xH�����ꉖ��̅a�T�Ւ+FҭIZ���,�J�g�oڍG-'����5�x7���Eh|�rYO��N�nd0�S�h����K�%�b&K��S"R/!��˗/��u(�$�L��C�9-�g.�7�'�)/������H 1�"�9)�f{�1��[���2�)D����Ы�<U	�w;	*DѦ�&\��L:�O�IIՍ'�����B�+[G�&Y2�L�E���F��褾��=���G�ɬF�ZQ��|�SV����xDԵ�ьLO%䠉�a����.I�����g:;=�w�����$�_�?�h�w��lgwJ�;�i�fBƳ���x�e"6q2�|Xj�AN�\���h�f�}	�b�<c�{y|�SM]��D���F�#�
q�H�Tm��k&=;!-<i��jSW6!��dJ���G��OVU�y���둓��d�']��K�G6h`nt+�/�^�죊v]���Z���\�g�mڻ�����r�mڴ�rM~�7�7�1Ojy�;׵<_ph>'�.(�2��NV��lT�~ �^�v�?�o��!̿���o���G?Bs1ϘM>�vvH���?{�r-��{���+R)9�%�Q�5��u���N���O���/g���g<]���R�Ir�ȝ����<o%O��&)!y"T+;`l�kE��� �',��Z���`�ق��/R8��2�f�YV
'�m�Z����v�wvfs�1�������O���.)�$[F)^��I�{!��
�	�@4a��/�._��Ӎ�a�\��\J)���!yKɻ0�q��D4�!���X��ş^y����U:����t�{mw8�g�l�W���aN�@_����������bE�����'Ő��ӧOI����$�C��r�x͒�����/PV�7�,��rU��ݝ��ru~��T��������1#���h�,Y�W�^al�$O�a	��i6��[I��~���h�;�}��l1%�;��$E�`���P.W�����u#O%���b�VRϵL��+�.=��X���<h���%��J�S��H�ۂ���f�"�Ӣ���}*LLSo_������s���sQd,>����hl��ii��.VGG��yɖ����dQ�d���/Θgv<@j�N�R�S0�gs~qYL���O��7�}������?�����g?���������|����%W�&SnXI����vݱ�8��狓�sr7%��dY+���uz~J����_�l3N���'O�/YQ4k�aq�v{w�L%&
v�/�(�o|�u��-[�|��#�|�4����	��B"s�xxtDƅ$yUդ�֟�-'���ݻӢX,�[��,�̝N1ހdx���h�����<�\"�ϸ�0 �ѵ"��/yRR���dO�x2s������,�
2o���rbaQqF"�3�=������/��.:��Jѧ%� �w_q�#�e��D�bt�p.#9�0�6��K_��G�qF?~N�I��X�s5q�cb�4�0o�e�Z�+�*�o	7BΜ�-�6D
���K��C��R�䌀����Sp�I�㋋�tJ�����Ogv0$5-�����rp�#�)�"o�:�d
�a��˓��tL�I�谉݇u[ed��	wLﱳ�5��)>����w;̤�)h����6}��)�f\���ļ%W����e���	SɊy'`^ncK��-
WH�6�		=*=��F�);�Dj//�_t�eݬWrq��D־��C[���puw���D��q��N�L�����y)�91M#~Esy􄚼�A��(:Hdlo'9�T*-��{����d�^3b�ϥۙ�-�U�Ӵ@��yi8�S�d��|q'�9yl��8ʘ.�evw�G<��cCj�	��m�Į�*��Բ�,g�i���0���+6Ǡ|I��������
�7��"+�!�^lw�Y��o:`H���;'c�ҤD��t�R[FV#�9� q/@�x�R�J.�Eмd�Z��tC8�^ZE��Ø<��VR6ڗg	A+a��*��<,�y�D@��l#�{���Ҕ��s�v`.X��	P"�����dqP��a��$�,����\�IE����[\�D� ��H��:�Y�+�^L���eO���x��sh[4���X�� ]"9���JY�ݙL��9��~�:�g��?�8k�7»>xA�YY�<������D+n��Bz�֢����v[�h҇U��
����/�7��y�w�ܹ��
��r�9��F�ݝ��L?�ބ�D�{����M$�Ƹ-r�?~|���gϞ��+p���TrF��	l>�i̒�6X@x����R[	=�iê����Jρd�4��'
���g���)�-w��J��3�HT:#;H6SptNd#�?V2��+2��P\�FDYl.C��Dbހ0��2exܖ��������:ӭʔ(=�r9��"�A�7�� 9B�=<��G��b� �u-5R�Sa�$Г�/�E=��^��(�=Ý�����J��#��/����E_�::а1>
��Y6���8�I��I�����������9��iWN�,"�PZf�%�_�`i��b�Aa�/^� �
�V~k'�aȌ�D�<�h�2���i�
�bÂ���s����I�x�����;�%�w����5)/\ot��l*���c�8OP��3�ܥ��7 3{��K��Ɲ;��r��#��!���[+�9|g`U �D��M�pO��G��ӷ��=Y�F�AOУ�AXAu�|��Mzۉ F'#�bx��0��Ձ,�!wظ����/�O{������a{&阮ʕ�ӥ�EÁLE��#��^�0 ��s�2�T��''/O�^"z!'n"�JGջ���\:L1�]<9�LgG�j�Vs;���lk%wH�ԙ�9�#�^RE=h�D	��ю*��0���
�6���oP%#��n�G7@橮Xc�d�(�������O���K�J�n�D���C�]eyn�R(c��4N��N�<�`:�r��oP���Y�e����J�Oѧ��Q�Q�a-�3g��˫rx>�L܏�:��Iﯰ�P�H��J⅊~��6��L�^���|�ⱦ��tK�EsY��ebA�4<�i[�"%�̉ua�5����HW2�䳖�����F�Mx�	�6Q�4m/FJ�Ã��%�X�*>�+�
��őŴ�nm% �j�	��&%A?��O�����P�{>'?j�`����בx�w޽��_���t��ӧ�Ҋ�h�l]�P� �t9+^��qJ����O�_<�i���q�i���K�b@7�"��HP�ۑ�=:zQ+[:+Ó���m��������{����{;�sz̐��Pg�K`ۡüJ"@��ð�!BS7�K�)M٫/�]��վxqJ����w�{��`�m�lYʊ�e$���d$l���ɐ;	��v�������wхz�ƍ������W��������������c	�oއ�1��u�ʯ�O�V6��~��靋S�o����ko>�%%ae�r�{�w�����/H��?��������Rڅ���nt�C-��E��[��_�^>yN����G�}~~�
n���n�^߽{����;w�����b�$�qt|��G��<#�\ݹ��ϝ{���#���~�����_�;�y�������ÿ����򂙎�#������'��p��P�UIW���8�a�������訝m�f��C(ٽ�=�� �m���%>���~�z��O�굈� ���� m�T#_!��>|H�틋����o{ꕠ���R�btd�L��TG*(�.2��Ü
��{�^��X:��\���Qh�r���=ge�3HS��)�\Q�WP�^I'�d��%}T��Pʃ^/K�lP��Y?F%n�D*�¢�~̢i5gn�
�Ė�~B�<R5�)4��S�#9�L�Wt�%�,[�9\��p�tv�I�v��u��>N�i�����Q�#��ĕ�<�:ۣ��T8�	�ZK��2xt��3'��d��rRP^я*t�	�%��&�	D=�G`�l��l���m�o�S�&v�ʤ�$�+�z}��|皎d���RFF���7>��T��|��hǮ:��X_����A�]:ߌ�s7&�u�	�%U�5��)��i*���������z�}��T�l��Z��_1�b�m��W.�L�s�N0���2	:SB@;�ͷqP�uN�L��g�촉�N��g���
9$2}�/(�4�&nI��T�em�yA9n�-��i4fwU�},꾲�[���^]����y�5	ɶ��y���lOe��L�x��i,+y�ٳ�-2 F�X�E���X.�Հ�M�wn���2�&�'�BA7rl�X�R�hA�Y��	[��S�bd�8��5�д������o߹�co���i��<]{@�{E��b5�C�<eH�q��>~y��'O��^>{z���l�&c�;X��h��4RGmEV�n<��'��<�{x]*�L�;'tH�Q�_Rk���Ɩv`�av���BH�M7���w\>��GQA4��q��s�d�U� ,	.��KJE=���[rp+�ʞ�����M�8�$�[P�k���������;�� oj��Z�E�s�f\MC�� ܷ"��]PR�urɎ.P������������w�-�AY��򤨈2e��j��}1\<B�F�S�ƃ/!A�]�SyKJ�D����/�2t�b����8�[�i[C*�)#�)dC�]7J�g�*8%I���j��� �A����aw�o�)8*�C��a�88O3m"�D:���� �m7�0@��u��M��B����
��}MO��Y�)�!�Z�� hu:���O��=�"�0�t��uE"<n�2�t1�KwG�Ow�36" ��;�%�0�����̮B���/<ZC�6�j!+��@�e��Oz��� m��*0��-+�3N���:��tL۔ɜ� ��NNO��i��k���kHB�`u�.�Ѻ��*E��Zq5o�
�k$8�ʬ|,��1c��MܾXØ�a���0�1�"�K=�t$K�7M"sq�,��Y��<���gOX <�4K5=��ɋ<㚗�1d��aTK����ild\Yc �eCh��Ro�r�b��i�����\�W��x�9,t��A] g�q�l����I��z�&I��J�̯8�<��k��g0�. ���%vWH���O�_(X�@@�Aw1�3}��u���FU}�^��!-�U��fjz>}:�I���0c�yq˺���p���P�c��'���oCC_v:��� R��Z�zH�TV�Vdqr�B�@���#2'�-�� X����b�zU5�P�/��V͒�d6T�W�4T��Xs��Cm�S���$S�n��-���s:E�x��fC>M=xI�d�^xA���5h�<�Q�k\!D`E�Pđϕp#���9���}u}�D��n⹦�a��J�բ���|��LE�GjkF� ݉�!G�c{��⥫&H�o&��w�b;eu�6*�\~����F�m�
�l{������=u� ̻w�އ~���c��f�� �~�O!ޡU�-����f^�YŁ�����5�T�>��_�wY�����_~���B*�J��3U-��W��a3q�s��9���A�c0E���������8EBRʕ��}�����	���>��0!�<9�'?���y~~���goNO�ߞs_�}�Z0A�6fA�r�w\q��0�t4��e�	���n�g^}T���}���Y?s�6heX�t䴸���*#��v�hj,�q�M)]�"�*����˗M��"�|>���b#^���Y�0en���|�H�ŊF�vv���{�w����~������'�^������qqq1ԉ왐�5�b[ˊ�п��� ���W�������o��o^>����M=��26�n���߿�]��)D)zt�]�h�G2��w_�����ַ��,�O�����cҦW�_��M?z�?����t�ۗ_~=��_�M�l��o����)[������㓓#Ү�@�������?�������k��b������7�����k�����Z���]�p�f���ɿ%c}vy��r����ϯ�}K�4)��FX-,�+S��&�۟���HX8w��!� ��9�G8����H�~����uK���{ �G����Sz}
��2��Y50 W�����H1ϬI�E����J��{�B�`�3CN�Pl1J�d��rZ�W,����a�=�+�ގ�C�R�u;��$��7_IB�t>�ul\z��%��)?
�l���N�"4�u��"}ȆG�t�@:���Xiw΂��k����E�-&R2�AgY�"3��lZ?8���2�� A��_��gBD��X.����]���<��oSu�Nd���$�g�N`�e�xv�v�����k��S&��d!�d��tq��<s�X�9q�����>�hE
�Z�Y��k*���^��!� ��}sA�M��Y3�ބ [�L��m[�Z�9�fk�b���X�NQN���Q�;��v��y(q�-l$Y�m�4��>"�R���(�:[%|o�!����R`�0�Gv�����Yנ��ZyFM�0������)�8;5~\��Ɩ�Mtl�(�δ�3�7��P���<c~d�xNs1��ɊR��3\pPD0c71�̔,ll9�xۣ	}�D����JL���@S�.�V[�p��E�cJ�S2ߧԫQ�����+,9�F��$�o<�L��X�Th�W:B~�`�R"�]��"|i�"چ�%�s��bU.e�/�o�,��s��*�E9ɭgҝ��dt�^X�XBЀ���j��)�����5�7�,�C�����
gM��7#sieN_�%� $��9�4?�����٪U�Ǿ��bn�b�m �߭jX_@�쳠��K^�|k��N����*<�u�O֏[$$1%�1�h����դ�B�S8����A48�Ź�J`H� �����[�d�O��2�?�Ȇk0�)��s�9�KeJ���ogil��^�.e\o�]��b�g��M���b�
iZ�r�RDR@G�l�nѿ����M�t�9N�ვ��Ht���~q03��$�k�o�O��	t\� hk+p1�S��`�vw9��/B��E,N��S0y!��q�`6�Υ��s��)6�BÇ̅Yg'�M&�)1B��(J�c�.i{.L6@T�)���hs�D�s3����!�\��&�b��RHh�2^ż� �L'�ag��B�%m;Rp���{�'�A�"�Fg>h��M��-�t���;�+��YC!I).���� ��4q"�<2P`�0�w^�6�?ѵ�hs(d�֐j�	j~�c@7�_�H�Jۊ���:�$$��c�l).A��9J�6�8U髯8S�8i��w�R��_�x!Y��Z�Z�-����S��b��� <|�K�K�e�ӟ�����W�^��a:��'�[��$E�����#�����ᮐ��2�j TՂc�Fe�F�s���y&ht����F��l9_��a�{L�8ePIf{Q�{F{g��f�ÄV�!Ș�2�x.�2d��n�r�������N`g�5}��V��X1
��+�F�|٣8�~B���Q��Z�����g��4 2������0�1�� d��>�Fh�Yq#���D74_�vt�ФaDf���_�ʌ�A{�)!'�e��	0�w�P��b�3뽢��tZ|kY?�-G��,�9�J����tc#f��jer�?���ӧ��mw�%:g�+�	�L7���E�`8� ���(菟��g���/�o�H��d5����E�C'��q���<źdeK7��_|��Oh��O4���d�?���Ǐ����y��h �?���������djp��i��ۮxp�%�>~D������p�ԃ���O������<zb�Fʩٺ�5T:��_�L�-�O�Npn�VP��?�B*0�6@�{+�P��~-�#�sp�q)�/цdB9�_,�n�t? =~�p�d.����1s���SN����l��7B���̴57פZ��Z0>�q|��9�!�mx�,m����'��������'''��_����X�.���I�...�d�T�O�<�կ~E�D�~����hY��������/�4�G'�f����|ن�aF&�w����I����ඣE#mu�������ݥ�:��g,�LzG�#��rS���)��/~�קo?��Ã���/���D҉���yUM�A�7�=
6��BP�7�E�Ȥ1E�"Ӊ�ggg�-X	
D� �tq52}N��c:k��o����=/y��R�8(��oVv��H�(��
(H8Z:���ġ��g���ކ����ɲ��''��L��5$)��ێrU^5>��}t+ @�B�2*�29�S$�E\�7�(��(��)u1n2���u����=��������Cc�m�o�ڥ���$���0X,]�]�+T+�;�����i�*/�ﵫ�=�G��Mmg�l����ܰ�b��σ�7G�`/o�@#H����O"�X���'f���+ ൘�UC{�\	����B���2f��Î��H����	���r�͚Ɗ>1v%�uך���g�$���i�F�Q�^3J��x����ҙJ>{rr��J�sl��o�F�G ���l��;�~̬��Lۃ#���A�Mzܠ��z�H���dg�$Yi"�{�B���Tҿ,Ua��cy���Թ8��J���C�@��]�Qy��TP��5;�������l�AeCܑ��� v����x�{�R��6az��ib"<�ţ/�k��TuMa��}N�>�?�J#!j�r��k#f9����C���Tbur��vww�g�"O��w��G:d2b� ���0�(��}����]_���/G"�B�Ӵ��p�=}�pw2ܛ���D���왩�0t�ͼqJF�D���m���V��`�l���g�����t�����~Ƙ��<�f2N�L�7��i݄MٖU�6̻]��TZ�JƱ�)�\��U[��Yy�"�(#��-�U���Q�c~�����xg�d�(�S�V0�N�YN��j	mj�mVJ��Y� �X!	�Ǥ�I�9�!BYୡ�L�C5U�\��6R�h��8���=~��d:p�§�7��ھ�� �d� Y"r��@�@��I������rzz��ٳ����_~wqqy��I�f�:���qӾp��P���7<���?�� j�X��#�)�cJ��b���$���/�{{c �}p
���U��G.	�*h{>�[�Ϣ'{�B6�}g�\���ő͡Îj���rYK�ЉD�>D[��3�)nF_䐹��K�{�eG� |�\����c��c�x�e��c�% ��ؒ�� ����9}����vJ��崍��K���8[���E�%=+Y�֖^��OM�H����l4��qԥD���|"�'G#Kf���s@��s6[X�[����������f�K�1�=�18�ș�l�A�;�(}�Y#	k	A3^X�YE�s��*gs���C��6��)�7�MӹA^t#Qrܠ)�DӶ��h 'm��kwO$!H��=zԕ��<i����dDvr�Y�I�V��K��tυ�*�ng:�Ýi3(�/�},/8����U�Ȝ%�%�QsIN�͔�gϤ�#�*�'�� Z3�x�9��jv�`t�$���hi��g������G���"�BM� �6=��� DMY�I�&9�	2]�{���Xa�%��֫���k�d�0��Gs�GG�L�p0������Z���$g`:�C�9S!/W'ΑגDJ�4��{��b,ۛ(�آ��# ���u3�1*R�-D�J��1�r��uDuMMВ�G�WV2%�����/<�Dǐ+�#�r�Y�r��s�w���;xy][5���j�W9<�Ji����|r�.��f�?6N\�������m�6tnty����;0��<�c)\��%�>>5��<\X/uSJ�~KՄ{D6�K\�qrR3و���7��V�
6$�M-E}��|-y
�-P�PSNcWd�-��UB)�����$R�+F#�*=}�����ѣ��)�D����-���Bxm� ;�,hs�g�d��pېƣ8Z����{��X�y�������_�����|.�I������C��dT~��7t��G�J'G?��[2�>�O%�Ԋ��޻sr�z��_r�&S��[���b�^��첼`�Q ��Y8o��i���|rx����'�_��V���>�]緘�|���R��ԻDKw��<`:�'|~I�T%���A�[�H�.��C��|�jE<��j�?��P�DZ��*ud��wR	q@NOO�f�=��^�z��<�S� �����b��͸��est��L� <w�b0ٔ����GOvw�-,Jdv)I������ݝ��8g���ow�n�F`HFӧ�E�ج��d�H?̮�(آsA�KGM�t�I,?|�=Oȉ�#�͗_���^�/��bsx�Q1��IJ&����h��������\����]�OB�2 �3�磐������zU�Eć��/�!�����^�jڝ��$�B�I��ʳ��O>��?��`�=�m�v�Ql]��p�F�>����<#���v\ �d� �0�&5�k������ɓ��EBN��C�PɃ����i���T��xL%��ts_�!1&���v:�#��j��yMf3��e��pؠy���@�&e����9Z �7 gw�q��w��2l"�mIy�[R:�5�F1�x�P�����mB�N��A�{Q�z�>o�0-�ztI1���k�R���'�,ˆ6�~B��l&�n��XΜ�5`-p@�L?����_�	��h�h��	���f=.Z�@P+��u�]�\n\
k�Ԅ���i��]�[�j�<��'�uP�q�yT��49֗�0B)�uj�E�~���VqL���ۑ�������x&?�seSJ��(�+7�\�qڹ
W��9}
�	��z���}0���� 敒؄�* �k˳��V�p��U:��@:�1R$��1ei�Y"�pl��Y�g�.^oy�
�D}� 1\�{7·K���,3��N���8!K�d;`�ܳ���b�^x?1�ǉ�^Q��{��k7�e�s+�1�y%
e�2��/a�@�k�H��&��A^�lP�G~{;��r����I:�:M���_������:ȵ˄E�id���d
<f�W5�#�UB|��!��U�z�y]I,�{�s�ʵQ�ry8X�v��r�5�	ԉ��,@$�N
�JՍ@s�ɘ7�ڼ�qa;I��Rݚ����z|/kO߸ؔț�'t3Ϟqi���R�Y��Q�V��@�g�M�3��<#�?�b#������~X��cn4N'њO�'`��3�2�1	�p�7=Yސ����BA_wү���\��gX���콕Xx�3x-R��
I`7xӫ��\�I&?��}�
XeP����{95��50�l[&�5���h��۷o�ϯ��8;;��I���ZL����l���6�A�G�!@*gk�E! -Qs�],,��:��IP����y�qp<�8�JG�E��Ǵ2���&Zo,�2`Ll��aF�yqZ�m�k5�zf����Naa۲���a����'Gn+�@�&�}{F�h��8��*��0���F��IW:f�i��Hڛ��1da��M�@Ȋ���# ��[��rcA���e.�:� q���躘wΔ4�� �
��B�w���k�2�ͼ+������Kh6˽�'�kL;$Dl28������y��߿?��ү�� ��y0�>=�T���q�F���3��C0�ި8���ʙ��\�q���a�=6���9��{�$4���fqnؖ�n�5]���ٰ�Kn��.��\KM��y�dC�����C4tx�#?yRm�0>��J�z'�Ux6�F'�o���ZZpR8!�cO	z� d6��-�Ҵ7��2�)��8�;��\iR�t�����l9m��;R?��Z>� 	_��.9:�g��fN��h2�������#��g/�a���>|H"t�歠�V� MN�@A5�PfR�p}�٦��G�F�R7���y��+4w
��]Ñ$	�֖e�ogʔn �X���4�6&�6���޹Zn�p$$Α���DJSx��7vJA39Du!�&��Ai�	V�n���JhU����
9����N˟��lztT�z�*��@��2-�VIr�T�(!҈�d�Q&�b�>j:I����S��
��x�?4��k�D�`��G}���#�(���<??�������w��(�n˨�F܆�(j3�����ۗ/_�c@����:�$��|�|���͋zz�cm�x���AY�> i��>��������ݿ�ۀ�`
�}m$tf�y��]6����Y_ غɬ�"�H��ɢ'��Ew��pP��N �L�Z[αJ�e4<YN�с��+���sl��"� ��-{��|�����i��٥%��7��
��0� � �N�A�t�y�����;�UC�EO&
�:壷y�0ּt��[�8�Obcȥ^����`I�=e������J��HdFk%����p�b�䙌�LȞ�������'=��qY�I����5˳W�t��ŋ|�\��cava�ReKb%����/I�'O�Ԡ��DA�gi�)7'''�f��q�G9z���NG���r�����J'򆞤VҦm��G��,
��� �%��@?����Нs������mt�[���J�`%6[<wq��H������A�X/hn=��R�e�$/F�Yf��=fE���Bb�j�t���a��X��<lcy���������C�mf�$.Q^�6�DmJ��:��\�g��A����z���(����=l���S���K���wY�,;���ado������D�^���O�d�`F��\/^/>Bo g0U�������St�Zc5�]p�-�����c~,�j	U�|]��؃�U�,�3�V)���l��"���
su��ZZ���d�p��1Uh[�k�ƣ�J��Ѓ�}�_8�恙{�+)�	�-�肋�w)%��B���[�<�F'���Ŗ���
��\��L9n0�$D�V�Z)z��<��A��u���a�T�?���w��֙�����c��Rۉ��I���D��2E\Z���قg���5�G~�@�F{������2�:ʒ9ͼ�u�2��Ds�T؅\	�k�՚g��l��QG �%>��t0�w�\��r0oRv3Zn�*�+�d|�2Iq���@�5�IL�;��Ó��s��"�cS�v#����Aݵ��.�5l�?�U"dؒ&w�JMO&����L|���޿{��;!.Kȑ	]Sw��6���"cg�A�cQ����,7B���fyVT%\�P��o^|��V���W�O���E���^�˓UI���M=_nv�'U˞�h<��v=�R��f�I)5�+�rL���g'ha�S�4$�Rޔh��#��֤m}�/'�B���f�uK[��S�EwI#Xf/c4���V�°eH|8��p��9$7$ݗ�AH"ήiX=����'�߻�s?�ڵ\!ρ��YJ3���*L��S�G�|Ƨ�1�ݮno�]��4�����mH&�a �Dj�[^�$(r.��l��$ag4���)^�Mnډ��%�2j��'�4#�G>%�hNIc	�}��8br�2!o��A����뒔�~�� 3h~̥���o2�����)��%�I'�	��ݻG�݌�ݨ��D8� ������dLG��F!�w�EF8T+���9�(�kt7�1���SH����S �e�& �D\2�(�B�oc�	{M�hh�5��^���ہ(^ �"s�"k`�*�-���9.�]��0~,]�:S�$�K�9�����Ǹ�z�K΄
�[��p��Vp彦ű�H*џ�D���W#�5�BE7F�J��|�����b�1K�:���9ldM�[�*Yj\G^:���
gE�Og�Ժ<;;���&#��t1َ-�r9�P��5�c��qɄg4-6�͊$y�����x����<�]�'��A���xRi�<p�>cc:t́�9�`^^��,�ed=s���:j�]^��=�hz'=�۷oa�h��n��i'N:ɖ:m-��뛛��7o��^ݞ��]�_�G�]�X��&�̼A�Y�9����)C�-;WdE�6S%NF��p@r@.}���aU�'w�v&�2+Q��#������#��˗���4?�J��Q�9*�Jl���i��U�s�e�n취y.�1����!uS
�C�҅"Ke�6���j1�S�z	�z�a���F��)ީuӖk��6_r�uhKòѽ�A���jS}��s����,��l6

���g-Ȝ-���(g�Z��m-�)X�"4>�ѐ�mS���Nr(���������d���5���w��d�e(hA^{><���d�*����Ձ�Q���_�C.��Es,�i����"xE>Z�b��Y�D�b:i�G)��}��V���?���P���-�����o_���j�'��}a0����A>%(�~����o~�Y�}�x�ػ���h@�ޑ��.5ok6ޙM�F2U#f��� ?������������G�waq����-��$'�L^�e5�妜-�7�yݐkʞ!]v��9f�!'jCo���[��������ÇOOO/�n�D+X��|z����Ε\�_���[*�6+�������m����D)D:��`X��iݛV�4�?t{f$kB��2M�b	���@S�5o�Yp�N'ܲ�'���'@F�uݬ�����+�+se����x4��<I�н/H[jd��)ui� ��\]]5
h�sS�U�&f<,&��7Z^/g6�C���eE�����eÀ��|&���ѣ�p!H���QU����zO֛��"�J���H����1)���8�;�̜�!���mH1H�b�\xn�ivv&]S.f�7߽&]��G���c�E�׷W�wN`X�L#���Y��4Kk.�I�W6QΰKZ��'��	$ �T	�"�P�D�al��-I�b��.�i�����o?��#Zj�.Í$�yX�_C���45�����{Yo�9Y^���i6�nY520����-m�dAJ�.��p)X,�8����Rs#�=�^��ZӾC��=C�C�)t��B��s�v�1Kp�=�N�y��!ؓɀ�ǂ�hV�-�8�^����O�:mˊib1T�D���运y�g5��Z0�[�(��
��0�A�8�#N=�DI��n�.�*:L�	0���G���t6ڬc9����B����Z�ۡ�8��~���{�yn��tȔ7�H�����w�+�(Ҝ��#Bϩ��@J,�$&p�^�����N'GH�,�v����!��`�۹�2h
/Q������YN4�}�m��1��o@G8ݼ=��q��<��.bm󜦄p�A;
+���).ò����ڏW ���3fA9��0�]��2����B+��ʳĴ)~R)�)��8�����V�V�-mJ��@�N.���r֣�e�������S�5���t]x?�7t�|e������t@
8>|��@'YsD�'���O�SR�~����3�P4�tK<�|��6϶�W:	w��	�<2��Ж��d�,(�YeK��`����r�5S��#)��$�q>B)VĜ;�\,��Ѹx*/�ཻGܷR$�H5��Aq��mٵ�|���@{#�!��\�"��ߔ5�P��e";�I~'�J��Te!��S���\<�ȷ�aӕJ����U������:���
�8I^��L�O�킷Ò{&��nA�t'}��q������!w��z� �u�<����t���\�t$֮���1)"�����L@����G%��3��<�+.f	��k����e�o}yy)ٓ-��S���L^ހV±��iv,C��S�S>� ��ƕ39��L����{1#�&}C�Cw*d�n4*����p-l���í�J ���>���赙�֙?N2�̥5�}aҮ�X��)��k[�#�A1�mo�z O��XO��쀭���6T������_�C1I��7q���t��駻w[tWh%�oA�WN�OcHJK�=*�o�	ʮ�*(��(� �9�{Fu� �;g@�p�.D"$T%�D*;����`��8 ���R�lev8^��Zf9�Fl� i��qh��g�d7ҸJ����z�:���V����~E�X@] �s:[~&�D�'�:+���~N�T�,�k�	B��,f'�HȕK%�*���^^�A��'��i@/�V��#�yQ�92ś���H�.o���j�����橦�O��v�ڸƴ�4�C+;���|���P2�O�<1�=�-�C*X��w��F|��W�}����65L�4�&&9<]J�d�J��NDX�"���\�jb���vr�>��$SڤU
K��qx��H��sjc�a�V��=x5̮�F�DkE��b��XZY�u+�P-��H�h���<��"��W�#����n�;���C�r0���7t `)������
�7�nreڡ+��y�"�f9b��W)D�~K	a�ܚ�l^�fS��LN��w:C�.7������0h��,(���l�v�|��-'���V]��`�0>�.��H"3X�蘈h�e���j�0V�4��L��N�b��7�I��@ONN�ݻ�e$/�:�I����l7Wk����M�v�f���L��z���R--VVS��a��1K8�?$��H���+��a\,T"��h$��Պ����[O"�����z���3R?β��n�ɢ�]\���O�,
�Y2"�7��4�wh�':��J�n;S�3�]�`�|H��O���\'B� ��
�éoc�Ħ!mɲ��i[�g��1i��9�=�v 6��N��"!��q.�.�5ӛ��l9���Lfz�Il�	���9,F�	� *�B`���_������\�,8�U1^U�X�@h��d���.v*��$��b��O��f��p�-R�+�)�fC����8�\�m��� ⌮x�=,�)�A�(��*ǃѦ�0��K�M$ة�/�F ��:���ua�a��?Gx��a\hLxx�p("\���o��7�z! �8�Z�iK�����b��Y�́��"����H�5!�$�ء=��t�oU|�Ckp�gݦ�����1͑1I��Ǟ��<�G�0�Ql�����|N�-*�[Av��d$Or3���oAY��7;Z�cŘVY�»hxS��p)���9EL��t�9�&�s�{:���c����~�f9D���q�ߘi1����n�gK��M���&�3�Gipf���28O�T7��@o��$���� ������ħm�
m8o]�5��=x$G�Bo[��d�)M���Ff}fD��iS=���QL�;�Ao�۶��-}����czx���"�ґG�%��/F���1���4�j��*E�'<�:t�9�2Ɋr��/���B�-�/5�N�q3^�N��D ]�a��l�b+�T�!1'��)J��OTyl����I͋m�I�>��Z�����7h� GY���|���|0,�BbY6�CH!���cp}c�P���*A��V��e*8
��A�zw:}x�><�۫z2�rg�UՒ�ia�ᦠ�w�WUEl�6��DN"���
24�#e�N:��'�L#3�� &d(�#� O��~ڶ��O��Y���L���ɕ��-���ӧO���M���t#cr�
o k��.��5J�?�NN��dL�'�TR+�2������H�����vy~~=���+��]fx�n�.�MY����^Y1��(��A�	�6z)"�F�e��H��wEF�T&9��8ނX$
�a6*aS�u0�ae�W+� �3� j4�TP�����:;	��[����	 É�C��V�I�E�mo�\9��@\ö
���"�|����h������xR�)� E@�z5�ǝO}�N�p�+�t=@ٻV��=΍d8��\U�Ey3[��WI:��IR�됆F���bo���9���3�y-jN0��l�\&�ܦ�tuz��]��!�U�&
�(:���2:��Ʌ�n����8<�;�b,#9/��vU��Y��r�%�YU:���FǽY��ck?TD�D�H�Z�3�t'0�����3���$�Ǳ�!�h�h2cdz�N����̀.����E+���ˠ%G$Ugke��:��=�Ώ¦�" �pI�%��(�d���p��!S��9���?{D��ɄAy�s�W.���Yˋ�|i0�:��J��Q����7�]
�#� �r�t�[�� T����pH�@��ҐŒ���M�N��e@+��'�P��QNt>�C�'�N���8��׷��]~����MmP�����¡��=^/%#Ã�72A��c\���+d�J� ŐI�lB�]��>2[0��߬X��[ո�f�MC�u����f�X~�I�w4ޥ�&�'�s��,H����~1�-��ں�E
�?�k�O�c$��c�I͘�TA��f��眠��o�m���o���g?���Dv��C�V����}��W�����{��eᘟ�_��p��P\Ճ���C�MY���d:�ɹ��Eh7�I�}+�5ZZz xD����y3��Q�l����^]�Ov&L��	]���������:�i3i�÷�RL�%��rh*���Z�[�i90�S�#��.7�z��&��ԛ�����o��0�4�dw|~~Y���^���&�����/��	 l P�i�)���)ɂ-
#�*��������j�R���`��݄|&� ���T�� �����b��"K6����z9_̚�ޛN�l���t��3� �$>�jn�$�e���i�Ô|4:3L��!Si��+�	ҟv3�,�O�M(�`��݁B�Nw�� Aj�%�����=�/�I�Li���n<BX� �{x�ޝLQ��n@خ���~e�b�d�U3�/_�|�Zm�Wx��5i":��8�M|3��� b�Q{{�������4sڏ!)4ҟϟ�|�����uM�tͽ��|�4o�O��֛�?R\JD��g�y��u�2ցs@RtI飙�ڊ�Ʉ	�h$���0T�%A�s���L��i�I�r�b� g��橶:�
�G���Ј5�LT�T
�?ժC���#
>���S.iì�)8d�|�Y�?�c�l@Kʄk''�$����֠
�٭Wܵ��_�3��A�ۣ3{�޽��R�t�{��L���t�OI���6���ˋ��������%��<`gՊA��ڌ�8L���\�{�>x�)y�;�18�I�%�;��_͒�)#��ɿ���tJ�ͅ�"#��B��F��fV� ���o^�spgw�ы��p$�V��	y�wRl +��U�,�"��ۡ���=y�	R6������ZR���;������|�
������D�
tc�~�����IZ���5��h<�|Rtϳ1\�+r�d� g�:���8L^t�u�!�9}hggb���΢W������}$�Q�����#��IO��40��\0蠏L1�A�p�(�1��4���<.�BM ��A��:�c�c�����`�xE@KR	�c�s'�B�}�J<Ȍ�������&��!Du�,;��r:�%G��)G��T�h�ɇ��;B�g��kѴż�N �&l�����{x-�u��hiV��L�˖�J�ȯ�7���\�N��,�����u:)�W�g���qz�R�B�Y�����!M��̒0�����p�F;De�eq.(߈$I2�lN�,EǬ�ej��Y�8�Kl!rp�⥴7$$�[v���ֿ4:Q%��H��x]��A�R,����{�R�8�n�:�r෥���"�o�m�ubOV��f��f|�2�n���3ݵ�Y���lm�c9��"[�2�����"�dc�&�X_��RV"�<�Wت�IЉ�mt*�������q��C?��)w��6jH�&UV�W6��2��\琠�e1�W�")���ʄ;��(�T�Cp�0=�0�KΖ��NlU�1��2��+(ŬLj��d�~�vB֚���5$�HuK��7��y) R���^��&��7~CбEN�ǐ׶��� ]���N��g�_W��Y���BK�䑥R�~����\iJ�%��y/��U�)7��V�"�Z�-��9�����o޼!���?��o�ϒ�U�<*A&l�M-��_]�����"�M���~' I�3P6O���Ne��N��b��N�v4X�PS*��Za�^QAT�c���
h����X�Z���\*<N��K�A���6�L���9L{�0QW�!�1&QD�����<B�Y�j�o�ڙ��ӝ@�,뇄5*91ܵ'�h�a Y��9v1'q����x'�؉������G���܅�� �d�u�Z&/���|,�i�s�����;w���k#��2.Z����X��/^�@��N.�T��Ģ+O2�[�N	6�wtt���8�$�wyy4+	)g�m���	4!j$�0���?`��0k;R�����W���Z`D�v)q	��v�$����P��R�;�
p�+���G�δ�o��c�S�2�X]�z�
\�U%�2(�n(�UPQ���Z@�6!t}7 �e�1|nఀ��:@(���<�~ �q�U����������=d�=/�8q��-�S)Sɣ�\��dE���V�[�D���#��Hd[W����m,饊�B�&C�F�C���7EU2�a��+!9b���	3�]m��g�����~�z6[I��3��#��o��z5А=�m�pۺ�s�;~~~�O��O��$	��"�K����r/�=z×_~��W_q3f>�Z�P��,i�����"���+y�Tۡ�! D2�)W88(s:�Ɓ44�k�f�T�+Y(��������x*����r<>��-���'�s�[�&7��r�r��T4^m���X��zq)�{�S�У@�H�D��@���Mc$	7�0���	�z��f.9�P^����ٓF'`��	��]AE�Ġ��8AG:��$�F>���a��<-EΓ}䫉�B=OY'�p�>��%��ݻwI��������@�b��'iDo X7~�����'Hx".R8��9E�lc�Ȭ��2�L2t��
�\�&o��n(�z�Ǘ)�ׅ���㖠�P������{�O���kzpz�yDA���h�Z�/�	�A�C[��4tY	c��ƑLx]C��{F�j�`��L6�mFn�`�5!r�P�lO�=rV݇�R ʭѢIB�h̹������i��]�HK�Y��)C=���,�S\�C��0Ξ=��wv-�b�+�knO�à���Bѳ�:��k1���N����FV�1�	�iP��d��=��x>o-��h��i��G�>��Ӎ� ��'�裏������(��ҟ�z{-8�1�h��0z ��hQ�H�l�՚��p�B��`�c	��Ͱt�!��z�왩PZf��V�ɞR��\�t'���8.|b�@�y4ن��>�ك�'cv�a�=���1٫k�/>���tRFHJ��g�{��+�h����d/�@�;?L�JR.-ʬX�D�P���	�K>,2˧7��~28W��d����x�+�+*��덳Cؽ��E(��!�5HW�9.f$��%��cH��kc� �j��X4�G�>��s����{���x;�3�br���������	fy�Ī|�����(X��+b֐Պъ-�F@��v��0�x%}u�	j�Ϥ}Nȷ֑?ʛ>��f��D�]��S�B���ȸ�zW��v���l��j�+�ڡ0g��v�����:̗��@(+����]}>q8ȲᵹT�p˭G�=���=�y�f�P�`�ou:��I�%d�#��=�����fr�P��{��ӡ�V�2�ipQ�+1��^Fj��f���.B�'OQ��j���>l
����ոs	�ek���]�̼�r���X%Ҭ�ne+I��Vb6���b�eB�4h	9N�����H����"�{��E6�V)qͦ�-��0a�6;$��-�J��?k��\@ȄV2 ��3^@Ҝ�w��=��.�!���e냹P������6������<�2#����^T2M�;�`1���A�B�T�}��:L<�N<!��	�=�3�C�9&D`�������G@`���/J�R�Α�3CWJ�qs��w���v���`�@�$���1K�K�����U��	r�x�m���hg0@��s
��A1�������v�Z���v.-�*��ߴ�r�Z�7x�+>�,`��*��Y�;'�k�-_*`[^�(H��1�����J�GVGB7�ݶS������|Qb�?ޯ�LĠA��-أ�*�`ϔ���/k��.U2�!�B /Ӂ�b1�����̻�3�+mGO�2u]�!1O9�����I1�- ��v0ɡI��y�R���YjN��J�1������W߼|���}ߚ���|�壖�5��v.6�I$#��%��%���djh����0���mV�@��(e6�yHZ��2[s*���-5���֟�0ㄞLFxL$�p��+n=G� }4�ǁ�·+����$�� n:V���'/@ϐn��JC!�=/9���m�D�!��>q��Å=�۷o-]蔓�,T��3l ڇ��?�(kܼX(y�:EʬF���C��mPD�}�7���_�"[Z���������0�rB�U�׮R��rCD�V�J��FB١.M�	W`;g&��,qTɨd�{���Z1����핕�R��2
�(��w�����3�b��h�h�fG�dڅ��"�d(u#'�A�bi�k:^n���\_�Q���&��1-���
dO�Ft��Q�"�%;?�kʭ��j_W����b��l����@B��O��-�q��ɪT���Ú��n�[���vY�,�L
�!e��@�� *r[�
Z2Ҭ}���:�SI�����]��.��ߑ����8D����+�^l[Z�g��6I#��vg�C��X�%@���<�wr��<��3A �xL�rhy�l��i�\˶-�m�r�G���圴���zI{ty~A�v3���L,��h�(&�[��Zd���\���x�XaI�ElA
���X�I���LOa8T���o��O�ggo�����'�7ɢ$d�k����B�'m#{'.|]mF�bor��N�㔓�������D_�tg��N�r3b�Y��#h��Mt�E����8��u&hX[d�!�h{ģtJd�
��+ ��,��O�3[2�*[ɂQ��/ȬP�����^2���[�>����r�\��͎��dj��=�56y�Y�I�%�|�+�+��9f������R�̣^�xB�J���
f��0xu>��ۧgs3z�����=_�~�tAa-,]������K\z��.��������v.���i /&��X�������dg��.W���{W����vr�#�O`8u�`v:��bH��^�/�b����{�-�s���D�}A�)���Ő�c�G9�9iB6�Ut�:mk��J����,�;�&7�!3ta8Dhfs�/�h�ۅ�z@��Z�(!��7�X)�K� L�'����gWί���������)����!n�l.�St���3�N
�pGb��y}�4 �v�)�A
˿��o^���?����,��&1{���TL0m���\Y����*�����.in�/�r5OBsg����b��6����X�Z-�����|q�p~�,��p��z>x�0<�n�6�T���������gw�m���Gd�������$�Ao�]AZZ���L�ѵ���|���tҵՐtT]�� q8��O���P����3oE�$ӗ/f��=�a������{�XGQ�*��.L���:9Y��بW����:2d��f3h����i�oӢ���������C�@�J��z�p��N	�*K]V��Q�6�C5�u�p���m��b!�z�L��)E,��q�"W����qD�mt��*��!(�ĊL���'���]*�tu�FD`����a�C���2�:	��lSf����e��/�0x��^�,hn􅤟@����-𗬇C̔�J��U��F?�v=��}�%m�T��'�o�B�qi=-��y�,�07����\j��m��<^a|N]D�y3�qU]쎍tl���/�x���0<��elM|�͛چYF��~���������xh���N�D�x	�"$�O�/
Pk��L��v�\�MFRp���Mxu�˕f�m�oI���B�}�iP� ^4�N�?�7W�%k��*�{ؾ��ʋ�jWc�� ����d�x(xo���NuLs��{t��r%dVx�Lp;��������p1HF��N ��@R^��g��)Y�[��S�v�⟽�����<f�F���4�ә����@�&@�DF	�2�mW�H���\#m"�����v~~N�b�$�٣0A�m�w2L "�G(Hb�v	�J������/Șsp�D�/3]NXTP}
3�d�"�j� B-�����{'|�����>�]aʨ���
�x�@[DS�
&B[}�)��	y�_}����<%ÕՋK��23�k���#�"*H�P`��D���$P�w	�
9��O�9;�� o��=
ua��&TS����F�3��N�L������O�є�|{ ���`�8�L�2k8���8�Jc	�2w�I/d'dm�ΓT&���a�K�AJ��������2�TS��-�9��b�"���ￖQ \=[on�C�ǳ�WP19�&r��.�&�⚍�?��[��9�6��%;��L4���J���a:� � 	e� �}����قV�>��7f�"ü:,Z��uI��>��Gg�>`?AT,(�P^������b�0�@4�B'������]�W� ���6$��<r%�;<<���>�u` 7�a�5��b���Ň�����5�
��T���{E�ڻ�_���Ȭ	�@x�;c�a�Y/��z4_�fː4�x�.�3ݣ�����#L9�J��Y�;�)��-�Sz?��xA�%`�"�i,'6�D�n���#�̳�ҜN��+�[�/!�y��H�?�z��s��'�� n�d`���^u�N�)���ǹ(��F$��K�e_^]`4*��]N�<j��Q��S�]+~|�<�>�����ʼ�ÞVl��o�mm��8���v�G��u�'Y��/.f_~�%� ��L��///�8�%`�n�ec��ֵ�_�`�#�|��� [�@��H�U��Z��'tΜ��7���l�@f�����53��lq>(��<b�2�4Jhc��d�F�H��`�(�Fp�������Y���t�'O���WϞ=��`P���ݱ��mk�9�N�qr��\p@{9_W�E�덤��DG�QS)ȳ�CX����+������3�� I��R��_�r|L�3��<��'���B�9@ĚVj�]���K�[���\�V�0U�'1�%w�k[n�D�8�,�E�\�nkz%s��t[Y1�p����˒`��A=�l�wrx��{�2��������v��-��3��)3]�s:���hVR'�%l��=��>�W�^eo"���	�g��G:Spv��k��!M��; 7�;9"��͒��2�>*���R���D�BUJ�d6��<kH���P�`��x>�4����$��ݻ����5�"��mZ� �wvvFws��"mj]P;|"*����灧;��M/IkE�I�d�>���_��g���[q���~*�,LB���{uu���Kѧ��)׳�O�+X��b����'���^�ӳ������o>��'?�	P�PD�O��Y�G��φ�	Z�mM��!b�蝴P��u�c2���b��������Da�i[���m,���
%���=�8J�7*F���h��J2A=wJ\�	c�����!���EY�ı��f�&ڰe�K���&`�B���TH~!�(�@��DŴ7�����c��?K��kM1I#�W(�6�	�ȺZ�8e����u�{c�/~�)��W���o�s�i��ǒgo+�͗���.����T����*�s��%x�m��y�r;�]
B'����U؛���@�A���G��{c��{�EX�RpZ>
7��	2>���^6�j�kB�����#S�A�U
�c?5dx�9D؂DY�"�,��:-���\!�t��Dg�)�u�����w��m3f^Q����}']�k�Δt�����߽�Ї��7���Y`����_��-�'���Q��cڢ8��k����^q������f�T� i�Ċ��I�+�í�$+��v�̗c+K�\�}el����dw7<iw[����:�Q�@͊�����i��(�������륱 ��$� &x�^���_��2��m�Z+6��E���mLq�/)4�S*�R�R\�w˚����l�ß�x۵��!m��_�FOJ	,��'�l23�"����[�w�p�͛7�U��e���]���f�7�զН	j��7�yu.���W3M��Y�=zDo ������t�$V���?�da�Gw!�γ�:�~8�ƃ!l��j�Ԙ����o�mB��8��5��w�9}{��7//�V/��n��9��"��ץ�r��EոM���ҩ�1a�,�َ�9����<�y�Z>��Gt,�@���M�5�b1���9-5�N +��q�)/���O$'^ŉ�QWXP�8��!/z�ꦵ���u`���QF^ yQ��ז�DB�f��ԡ�� �'�|w\�䝕��˽���n�G�W��[Aכ��[���f���*=�K7�����/�}��볳�9���°]��@���)o�I�"A/FE'������x�L�La)mrvP�׳�A��e�(r�Z{e��<V��40Z%�i�������0�'|
��L��!��cW�>Nk���t�Y���`�ŊсecD'�]P�u�Nj&LՊ�9g�����!��H�Q%�����K�N-/�8��/F ��2�M^=�)�
�$�~H2�q H0b��&Vڠ��"#3��8��T��P���kuJ���8��p������֤�5�,�ӑՄ�B4tt�ږ<��'�p�=z4�#��������wdh,��],�<ϝQ{yt�%E�-�!��/��ٵ�U��9oD�@7��18g.M@$�-!�D�-z���Q���"\)e�H�Ô[����B�֖1��@]0a.PB77W�x��8=0����� 3F����e)�x�b?,'�w'!k8XC��r}�~MRY���h�OzBt\���_5��<II�BC���\&�<�ũ@l�F�:��&��q�pk�}�s�q�/^� �2�g��:θ�3��Y�@n�Y;�Vѵ���.�J��
���I�zW5i�Q1��'�`(��;_W�k�<[wu�'���	UI)�+ت,�����RH��jյ�oE&��>�f>gRHXD&2��Ã��m��h���zMU[`#ϾMv�%�̠�f�ŋ���WC�![�bd���;\,o�[ɮ��O���� �"4绪ވ_���3.��2���I)�ٛ1�w�YW$�$���j���(x��s� z$�Ѡ+�ɕn��B2!zk���,<ꚧ�6�,	��x|�E�m�a^�'Ca�c�X�ã;E&!��t2#��?�:�%d2ⶦ�v<S�\-y)���Ȉ�R�8���A^�c�fLx��y�l�hY��i[�*ȿ;�L���-�:En��\/��Q�`~����/�$o�Ԏ���Aa�Afkn�E��4l�$k��gŀ\��j}s;�:��W̢���3D�~�\��}}��+��C*�4ޔ<ɪ%�e�Dc������aS�!�8r����&��\Z�;�Z�5�|���N]�pH��6�ߺ����yM[���p	�	��rb���r�V���Z��d4I�<~�������נ{�X��Mg��t4�a�=�}h��U�R��>==�͹����U催�tz<L�ܥ���d���bͶ2+�m�����������V2�u����z�d�f�e���pw�w�z���|B�"q{�\I��\_.���?�����פ���o������r���ͫ��ö�Bی��,��g>�:pnNdo���K����_�������}��u���~�t�YW\�#���~"�	}�����7������Yjr#]^�e�>9�Ǖ��+^�_�ab�|�7�vv׫���jJ��$�Hu�0O�w��.���W����]
|�|��h�7 sJf ��,�J��Abe2X�1�&q:�@iZ��+s��a?1ct� �(O%W �e,�`��N� 1�5P|""����t*�" ���Q�i����nїxkr�Z�- o�k��i'�L�I.|�����1���W��������x�G����X����(�@�� x�T�|4e��p��L`J����<w�4�	�&�>f�:���uȻ�L.�)^�ք^���l��7i��Rh��\K@դ
�{�,�a�N�u�q�u�6�v���4��8��a�Ast�ߤ[J�m�Le1�op
���+⤙:fN�[�w�N~$��Dd]�;���hx$U�-������ՠh��	n���R��Cm����kz<`[es�,[��\���:$%n&Y�-���Vh�^/sбt�I���j���O�G�@߄b�  ��k�d~bLk��3q�e�i�<) `ے���E޲`r�mw����[X�Jp?�������[D�e�ȮuƦt��I!��ֹ-+��8o��,�P�i�5(x���)��r{��'T��b���to�f�H
9��@'1O��Q��4~S�":wm����&��܂�x�긹YR�?�'-	 m�=ʥ���[��y�cB8�)W6�����0>�c��x��
�99"LཷwyyI!��1�[�ñ .�m��o'������j��>N��,7(J������ѳ�dT��u�P����`�?R&B�$��d��I]PM�V� �/���5�B�μm�c��fs����4��Å.0,>��*Wx�TLvn� �"~g���F�>�Q�Q=dx���I�!�WI���Q�{"<&�2}���C�A���4�8-1%Z7ׁ��#	 �qggJ2F.�\�3hH�HJ�'����0��ߙpTO�(��hAg	��SX"@�M����߱�VS�b�Kq����}���˗��gb˹n�Y�f��R���3�����iiN�{�\s,*s��� � K��@�
��=b� r�j�l�Z!�����<�к3���d�PAũAD�d,R�7�(5�����x�Ç��,���s@ϰ�Ȕ����q�����P�T�Y^�k�\'�d�TG�A����%������(Fz�\^�et's�p�
<��?[R;�HDȃ81�&�D�Л7oH}1�^2$"�{!7�b�D^� 9&Z24#EסU�i�
y"�43�+1O6�5�`*z{e�j�<�UǟY͝�k��JS�@]�A����I$؏��Wػ����NG�����8Ԁ&#�BB̭���O�&�X3<�ʦ����kg��4�O���%� Y
:�io& ��u@��O���f�4a��X%��qB��^�$��=`���7����ˤ�~�R=kE�`ߡTc�uS�0i�} V�#hnE���Ѩ8e��ƛA��{8�O�bɳ����quum���?dQçR(��)�M���JA}#�h����r�7M���*�������/F�!��ᗡa�1Tg2�n�7���[+A��T#����z����p�鷳قtS�J���o��m��a��Hj��.ےb'�@�׃W)3*�1(�A`'_��$:Y��3�% md��}>�`k�촭X�NB�,�# Ё���9�OE�N�u�\��SyA�(��y��1f�ьB��Ay�P9��:K��!��pm�/�T�PG�x�������.�ㇹ[R+*���E5�R"�(4�&�P�t��,z\~�b �-Բ�#�=+�AI3���o9:�C[ ��@����X!���HS�7��|-�D�C�x�CK�TQB��`��6�0'�cf�e!��*�5[v�����&:�_i� �z��9&z}��O������+���[�?�ǩ��\�=�AAk뫜Q�^�*3:�~^z'9l�v���,%<I����Ѓ	�_����Q�K_�ܔ���t���0�Zi��{��M?!Q�	-Y����p�w�w����t� �,��/=>xo!�t�_����A����� R�(=�%����������R�G������݈��Zd�M�DϞ=�������B'b(�s��k�'�������Y�eyf�pT!3mbn!�P�N�)�s|�yP��v�I=8���YI��+�\���NLk��7T����@�b$��U�D�C�",�k!:��N�<o�*\	�
���1ٲ�F����'�&���e�B�j�~b�S��(��&���sF�4��8�:|����%:�|��D�ay$;q�b�L�ZZ��(�BcN~?��?�)�O��_�Ϣ�w�&�hoKdY��{8P��L�+�.�^?�����-�?���N/�/����',M��O,��_
:�v�f��/�7����@R�y~^	ڿӊ=��8��1ͪd�?��e�f:)8U��F�!���WAa棘�)8�����$��R�䐞x1���)�}v8�VhJ��Q=�6��x�':P�iKo'�pf
��{i�do�;(VU��"~LЂ@�N[>�]ɰEV�i"�I
2��k�l�	�EZ��8$øeģY������  ��IDATA�V���E?y���`P�D��	V6Q�H��Rj��~�Ĵ&�����ͤO*�J)�q<x1��z	�{ n�)f�v�W+�h��QF�䬅������R6k�#������gpo߾���OR�c]0�r-	��'�&������I@��N�o[�%ֻw�1 w�������N
��������V��b���Y�N�,��;�h뒯@Z���M����<��Γ��>������N�fI��2��vMԻ��,s�}GE�Dy��vܩ�m��痌�j)\Yҳ��Ζ�:���	gGӉ�`�4���w�#�����^F�aV�i1�sy$3w`�k�2P�:�y��C�����9�^{�ō�W
�$8l����:(x�~�Sr�y����"� ��E�1��4b����GItx�>�� >�����]�=��������{���w��<F�!�(	~O���|_#u>f-a&�=;��j;�
�~H���� e����\��r��G>r�%�����)��k�������A�r�A�bG��+�lXN��rie�K�I��g�Ͷ캎k����d�@�@Һ�J�umʮ���'?���z�?R�P��q��*�zȲ$E��	�h �	dw�ݭ��sE�J��3((�8g��׊���$sH1��S��!�k.>]gVq�:��!���KS
��D�0�V�|�ⶊ��#�}��'�z���h�@�/�"��-��
/$��1�v��ೋ �a�����)#ח���7�dRC����q2�m��'2xf�\���H%ϸ#L�m�+���"DԳ�q���)�X5B˥de�,��D-���W��x���'�h*f�pf2k2��|��7n�q�L;�аy��6�`����cʭ��?"$�F�+�2��N�3*��Æ]����Y*gȒ\��!GCs��L�k��҄e�),���#��="U��R��zM��t�haC1�, �9���z!kLo�i4}�s���>d뗯Y���뵲z�d�$6ˍ��}�8�l���^Ϧ����;�(<{Mpn��$G&ou����<�i4�mHF%���]�q4-�,�-{�"WMN����K=F���O���c�5�\'��|$�V�ZL�Q=A��͖Y����8��K|��	'W��ΘO��D��B��J�=gA��ZՁ	�QP�����q�Ц�V���<zU��噦j��!WM�QQ�y-jJB������u!-Յ8�GG�����X�W�E~�v�<&f�G��1)���byu�\1o�53�j����
qL��Xo[��[�:f_���ŕOS��3��7��R��}��[�%���M�>���r�����(�ɫWg���ʊ����Y���<����߽��~�ϖ��n@:S5������BYC����^:%��L�����zK]ϤC���7¾��%�Hp)4aa�Ѹ�&�!����x
�M5��� �DT�z�O.����#j<�M=>,P�T9d��<,�Kz���1k������d�6��d֮�e���ݤ�%�NҫM�|,�0g3����nݺ%�xv)"u54�������E����O�~Y�����E�H�|�N��Yx��8��"!t�D��&z&p������g�(o���M�Rv��y���a�������9��A�|��_<?1��҉m�N'm�X
R7��ӓ�ޮ�d�1�I�x���3Y��?�я�I�����ɓG��{�.|��)��T[�ĭ EX��8k��M�."�����U?����蓘:W��!�������KV����u����i�ſ��_�y����^.Ө�~�T�,S�!��(��̧�r-����������/�E����YY�w�w��i9===�5��Z擶R{������߸�O�����|�@V��ʮY�T�yp���e�~��_�U��;oi{f�/�:2~R��K;$(I��ȹ����`p�iO�>�9��0w�ry��ZdL�N�C�s	��|�F0�t'��5��9�r�#���6�s�����G#�`�saSԙ���*Yr�|�`�i�q�y�F;ED{�gFO�7�U=�o����Z������$e'������� ��p�Z����ۿ��b�\˦�4g�u%9�$\>���);j�x\�r&�5I�ڰ���w�X�����-��ᰭ���xǡ\E��H'8}D��!O�}8~My�,k9�WO�6  �3㮦�u���d���#���f��JEg�P�H����x5��x���T��Ce���?ї��XzK�~�:��YF֘@��k�h+Bz��̣��xL�2=��|��0~�9��F�o0�M�|���Ʀ_���W+��ca�VfH]�05�L��	��q�VS��1)��M��3����@Zc��R-�oS�9&c�paK~9.;�G;�Ԏ<t��T�����pzT���q�s�\�jT ��?�Z�|���Y]|o�%��*��7��f�+�/v�����V��� ��Q���"=ݬ�m�����y��|��_���?יJ,��z:��6��(��(���WB�q�:��2���~��)Ke�K}�َ8jw�ܕ-�P�������!!�Z�89Z���(q�8�*ܹs�a9+W�8��%/]�H7JZˆH������,��U|MIۙh.c��|>[�\�Z�f��b-n�{��TB�l8Um��}y���)nY�p�辐���J�#����uyL ��U�aށ�(O`~'�u��EJ1ß+-ٝ�^�Ni� ʳ̶ФjC�'݋9�.x�X�\��=��"��m)�L�����̈,��kO�)X�ew�^L�Rff<.�6�GVճ�LGJPƭ��j@!�I���b$<�j��@]ߘ~�S������<|�u�=�<;;�F_%~���(�>/}�rB�'��dV,��r����f���j���Mg#�<C5ϛ�,���)�Ǆ!Y��V+.0�G;L�ɲ��GI���#qm�Ld�;�IЌ"��u��27��	쎎�#2K[S���"�+�E7n�@*r��-!K�y��Ra��<��{�G��I>+
��I�I>�56Cd�{[9�0.�S��-&K%��fi���l;1�`�I�ڦ42;��~�W��[LU�U*��,<K��EB|%�~�UDVKT&��V>{��c��^�]�^b�lT1��qTDBP�2�_�*����N>"jP��+�oy�ݽ�D5��L`G���B��ʕ�̈́c�b�꣹b���0�l��/,)���d����ne�$�du�t.�_�8���b��D9G�sJ&=����Ժ�� 
c9�\3���Me6�Z�S)If�^o���m�m���DCj���~�"�U$�g�3���`&��7�%���=�j���q����kEQ�����k\����q^��p��kZ����1�u@��uD�Q\�R�D���`��(H�n"Kk�偍�#n��0}>�Q�Q45�q8���ڪ0p��-�UYe�r��Ĳ�$䆌��^/�d�`:�@���6,M���٣�"�0*��>���������zumr+`Ke�x�Q ӑ�[�ԫ��Y�E!g�O��8u):�2h������+�N�@�����7ni�s{ٵ׭x^Tq�Y��� D�O�bXG�>,~Bp��߾	��e?��O��(N�Z�~>E�>Lz�+�|u�� � ?`���٨!���_��'�)�ﷱQHW�0I{L+�Fl^�|���>{����NT�Wo8+ݙ���%��B�b\@$5����#O�c�F>"��[�~��_�O~v��:�E����d	 ���A�]r.t�������?x�x

K�V.�,�:��� -�3��`�U�f������	�4��(�����.�*���Ѻ&���裏����W��Ki�T��ɓ'Ϟ=;>}��%��J�9��<�Sy�Ȳ:f}�駟����e�EY� �)1���ӗ���O����O�����|&��|�|�g�}&�<�¥���jyy��˭�*5���g?��\Y���7�>|({:?i�zy���'z���v(�?��?�G��HZ�Q^I0�iV̩�Ը��NT*j�Z�?������ꫯ����+Qŗ_~�����\�k�7ꢊk����a���믋�G���oЩP����>5��g���{&{� �g#��8xZ#Zs�� ����%�7LI����Ʊ�PPo���`̞�G��^8����"/����@_c����҄�������w��7�#�/8뼨P7��<O�,�7��-u9�FC����hWQz��Gu���#R� �,b)0_���4FÕIh���-�/�a��S���v��8�@!$2c!�����(�F�П��Q�>Uo����_*�����(�0����<O����mgM����f��;��d{T���),��C�ێ�9�I9��]�z��j��$��i�:���~F=-5֎�Fq��*��8Ne6�x�A�{Z�������K��9��Z���LV���"�r�e*����,�N�N��\S������C?��U�hP��l�\���h�g׷)f��ժ)t��l'JyF�g�g�Ǉ�e�^ޓړ+t'V%2��)��;��o�S#�ʉDf��_�$��I�N��\������?oБ��1*q�Ԁ��3������=5̗FNDIP��ڂ��j�'�@����-��=;�C��[���-�r�P�s��V���ٰWEAO����^��֛J������oܾ��;o�5Y���ԓ��b�@����ɇ4�w0��/�4Q�g�0_�3*�Y���03�"?���+˄K�C�F�L?� ��U��`gU]!�6�OV�E��2�Elt,���jZ2zd
��J�|'��1Ux�\l^��m6�f��l�v>լ}�r`g7U۾�����ݙ�'�j6����O&&x|��G�?+�݋�(!�D��i���W,�jú�����o=z�����\�b��������{����Y������R�l�l�hP���Z��\��E�Ot}�z�	
�X�?fu�H߹��)�9u�y�	�$���g�? V�$�8<T.�^-,W�rZ �PgV���?vgg�&��7o��QJ����UFy�[� �"s�����DG�jѝ�~&o�"��l�W��*_m�/�w�����N1���]Y�A�VV�!���
�6>]��"�xG,�j�.����I���j�R'+|S�Ðǵ2����D?�V�u��7n��o8IV�e�RwU?��َA�ֲ�i5�@����q��Kof
8kb:�b��_B��jl�H�,�r���x�d/H*��L���A`}(m�xl��y'�h�1�0�S�;�0^��o��S~��s��-��(�%���|��q�1>�U@;���N�t�׊_��d�0�Bn;C�Ik��8��mr?�\	sh��z�Zq&n�0��i$J98�[,����65�b�s��b�Zv�z����
��4(�#���&@���D{�R2M&ס�O�94��J߸q�_Gp�SD�鴺*«s	��z� jFS�@�N�����k��ށ:�0:�D�[	�0�A����'���)�پ�{�,''��j`|x�d�j�,����WwM|��R,s9���{��i8�
Ңe	�'?Uݬ[	U��+⺽ES�AT`��^���u7�f�S?��k��^g��J��Ǽ�F����������"�� }�l�B`�|4��46t.Ŵճ�r��ά�Da��г���8�+��mz9��'h�P�y��e6���NsR�əϋ�h�����M3�&�YmR*�:.&BqU�es��kJZ�WߦS�ݶ��\�ܧ%1�r��{u�ڶ�SM�I�7��YH��t�Ab��;b�DՈϠ�tݦi7����ƥo������B|sU�u���?�X�:Mq�+�e3]���o��hT#'���#:NFb�H�g�I*[E�w.�XJEF����o�F�u=)�~��3i򸷿/����;��((�I΍�� V�y�B���M��yY�Yu�${py"g]s��CE�fZ��f���P�.M�����"|��_��G?���������ןj5��r�տ�|'�XMa��9/R�?��Z�4J
9!��|����oZ��T����F�=1���o����n:y[�+����/�,ҥG�\'��l��)��)�]=�.���|וzwU1��jI#l+���9�+6� �a��L� �F3�(C>�EV�u\y�S�=`�-P��P'�j)qD�����u�n�w�:L�x��U����x��w�d�ݽ?8�yS��B㩇�!r�&�����a3��l:�	�X,���=�VgK�|�q�8tZ#���&ƀ,dJ�.f30H*TɁTb��`���r;��X�UAɎ�E}����˿��O>��w�~&w���&b��.ϧ��LVfӝi�o����wm�=}�<�_�0[Q�ĕ��XwQ�;;�Z�����Q�h0�]~��h3x��s^��T�D�_Q�H���X,zlBޛR��3�,Q�k��Z؛TT�%�Zm�hӮ��!�^��T:yЁ}zL�ؿ8��O~%D�΍�ܛb�<�Z�T��������[U��q~��l�w�{����Y_�8 dogW��H��Ү$�z	^�ϊR����♕H�L �=8:8�u,_�˟�\���>���������z2��~0ߙLg�Ur����ys��t~V�ڃ"����g�5�����}~���Rl�b5����jy5]�D�Gd�D�u��?��?�^>WN��j�$&hg�@3Yռ����~�G'����,�lv�Sn�lGZ{y��"}~��T��
��?�b�!̭�#��h󝙬���%zC"4ME��Q2�A�YSl5�e���L��&�QCxU��\��0�\�����֬��������d��|�8z�t��X>�ڌJ��YB���[���ԮQ��Y��c���Օ�\�@��C@������#���D��th���2r̽�0a�I���1{���r)�M����j)_,��(�2�������Nŝ̚���S���r}���w7�|�_u���������d&��ZD\)�T��W���R�j��E�h�]�{��RL���:�<�G�g��Th�ʩ�[&jFf*p������O�,'�PV{�!� ��\�QYkMֳ*�t�`dz�daX7�LE`��2�Ô~�O<�)���跄]�� &;&�|t�ۤ`���OY�-�q����Ԁ���4$K�>��ׄz�1�!m���N��%q0�`@6D#�m>
���S��3̈́``��&���v�ׇ.c9���Pr��Bqo=�Vu�Y�
�C76���A��zk�b?X�7�C�m�v{{�S<��;�7HHO��֋	�S�E��g����i�����Ec���83Ol�����W�A��P{�'�n���Q�>�����h��6B���l$�8	;$���ɍc�ɔ̺�yq_aQ���=I������ۗ���F��%��^�B�ͳKK�a4B菾�ë� �yˍ�X�������{�=����|�׸�tV,������Z�?ie�I60����`Q�`������y�~d@�A%|�I��`<����������K=I�ÖO!��,hͭ��gx}FL�<��*'''WWJ�t�CB����аaH�I ������;HF��������D��x0Lk?�M�A;8����TJ`M$���*��'d9hB��XW�E�� �J������L��B^���Q���:����a���9P��JP��R3�ʡ��0�$��3��A����J�
�ܳ�^����k������b��E���x�^T�W�F͊79����륹A2�"�M�4�I�H���:���*�����#&�z��؝z���8'V������7��� ���\��@�ΛF�>޸qCv�ᓜD�W�Mi�dQ֖Ȫ,����~R����]��hV_}���d�|�/�O��]ͰL�T��(��لb�F���-���>D2󛬗CB1�/�$ާ��8���
y�<e@����o0��[��';{�r�Y���VI,!�G*:V�������Z{�NN{��͚�~QؖXI,K��Z�U@��3���j�]����+8�o��5q#r�5G�P��-�p*�%ZAy��xF�`��dq�+Ͼ$��I�1���64���<K"�w�6�Ԫ�m���w8o 0KBF.,�e��*[e�vDG�.4�Kd1�of�Xa����Sݻ�!M^f��1�E��Ɖ4�����O���܆�#ÒP��z���|P�/�)K�`L왺��+*@���g�/o;�V�T�k��|��j��\�C���z�ؙ���j}��Y]'��z>U�x����X�v y8��'�'C�J#K�<��]ۄ�}X*�k�&�CO��U���0���0h(Az�"K�y?�5q��-|p͖�S�\"�P�R�Jߨx���Tb�����ߊ��*~��t��%��n����PV�H����41b�,������C����&���|i��ɢK��t�>��/�qhD&�����z少�|�-�y�6+1��#� �5$�o�ؿ����B�֐����Ƀd����|�%�~���jKB�����}���D��Ճ�Ϟ=����Es�"=�yg���<�.��%J�eQ{m�a�׍��k���&��u�z�m��q�A3��������B����>z�ͷ~�ӟ>|�\�l��'[:J�v��ɺ��D��(=�Ѽ\G��Ӕ���<��m�gf�1D��g��s���Ľ֖X�8��X��{�x6�t:5L��D��R�)�-8��dmI�������_��_-��p��ǋ�e0,�`MBue�G�!��&�6�@�)"A�V&z㛓}m�D�E�7��"���eZy�/�����l����%p/S�:�"�����o�}i�G,��T��Bޙ���CW�|CZ*w�����Y��0�C:\\(n����q�8E�1ո�l!mB^w����nv��@�j͜^\䆠�����a��M���B4���,y�c�,G� �]�Ҙ����Ȧ4��g��)Y��}�^��%��8d烵B��G,��p�"����b�l��;HlJ�������_\]_p9�{R��Jp��W�d}�vEd�{｛��M\^jSB_�RuT��˓��3�����aL��ՊSx�⭸�<D'׳�L/:��	��['�'=�������ќ|Nw��Mu��Ճ/�v��w�R0�o:��&їS�*�ǳ()�'�){����#�_�Q���F��7��$0҇��@���͚�^u��W���Ԕ��b9���O҇�(SGz�f�v�/�4����\K����`�>��~H��LG��� YNf}���1j��5�e!n�������-o�o�Q뵱�Spzϩ�p餣OE\��T�f�խ�Ԧk��D��"i�-�7D9.�X����j��a�`Ĉ�".�P�
]S�R�Q�Zm��ܰ<�0Z
i���J>�?x6�w�b��a$��,3ܬ�6��#��f�6���`s�s?K���訣�1�,�{Z�o�րt��ĔY:���r�N������y��Gy���87��PR^%��N�>2���,8_],�"�p7�������G��m~EH��j�k>��hx�Y�Ǐ��o!������٥lB��R�{�IL���yk�5��V�Ԇ�Q�xk�(4�e�pSˈ]^.Ř����iz��b�)�q�����v�bD��^�}� ���ZR^�kT���乑F���˦M���*�jS�/�O����w �I�{d�������`x��>jkz��P&��k�T�N9bu;�K��+�'SA�mw �'p�yo�S�_����l��l���jΰVI1vw���Ĕhp�Z2�ᝃѨ.� �A�0�h�Lggc#��Q�󿲏5�y�0��έ1�bd��n6{�
�_�[��ȕ�|���m}mQ��g�M?�i�,/��jET�j�J�]q�<M$��2�e�߳Q�_�&R<��r
��3q��Bƴo�-�~��C�]i:�Wr��+J�)��I|�)9�r�h2�T�9	!����=g�ݑ{�[̆E�Tț�1�y.�*����t�ʰ��my>���V'H��X���	h�"[�+ɧ��0�h�/Cog�8�*E�yR�t��5���[���w�SZ���g�M{*|�$�M"js�J���ʶ��5��'�]�q�5���V,W�s��П�}n �e�e-�� �t��h\F��_끺%\���/<ϥ<�loOG�<#�����`|E��S���_���|TSAp>�_�1`W����R)o�:�ʼ��Dx�X�:y��C612F
���	X��Nl#�a�A5��d��{�&f�ؚ2l�4��o��Aj��|*��l��m�*}��[��^�����)�C"ac/-7.��ZR�Hw|W�E�r��a�_�e�����b�F<u�$'D�szz*�%'}�:%�o:d���-��Y�oVV ׼�ұ�m��yV�3��OԳ0t���3�%�z6K������E�F���1 m�տ)����9۩��z����Z#�s�\"ѿ[�l;f��t�c=D?�(���z��kEM�� =�*_�Y��W���_a��{�aS0�=L9���c~�֭�?���?��7�s��|P����3���4wYhV���"�ʔ�����AK�b	7��Nì*�D��6{��x�U�ЇS���o������#mv�˳jr�C�6��|�26}�`��u��^/	ր�DDLQ�k�S4�~�ͣǏ߻wogo�lop���	y�m��2�����ߧ��~(����酘mlٶC�|@]�[k'A8���%�b���!\�R�$���ϹP��\gw>�}�L�'\�|����~������������N&�wo:Q�@�ʝ��wn�8��'�gƪF��ڮ��9��H����o�0�OPo����'z��k�`D�ZV~Z��r�-66U2�zF��&�)�4X��r;X�`j���1�?R�43&j�Ԙ�2�$�DY�˂tf�\�ggV�G^��iޭ_���m�O��h��B;��|�v_ƄNP��:e4�=�-���T��C
��'7���)N�t��^Q'�?Z~x��ܹ�0� �^2]Άh�R��l�$��y]D'��a.1�SV�S�����O�4���Rdᨌ;����?�a������Y�/S`�^���üY{�r�
Sf̾�V��f�v��6Njzkو&ȍ{o|m��ΏV��m�5O��F���Rx��]�fU,�QS8=(�eqǞt
lScfPVB|q�&:{3�
��.�	NЮ��%FDd�X��h�`lSH�G_1E�rM��1�	���N_��$�}�7��5[W( I��<��?���g~�?�C������3�8J�����ݟ�0L*��;3Մ����v%�l�t�>�G@�8(����t��(��O�>��/=��Q�`P'71���A�{��}����ƙ"�ܳWft�)��Z@��I<M���ԧ�ː� �d�˵�#dEV��2ƥ���5d�d$�:�Z~Trb#Q
x�Xe<-ö�9��,m*��5��7s������F	(��6R��ZW̓�4F��$�Ta��8Ք�\i����V��%�@Q�
c'i�r��y>��iJ�O��l�{��(K�a=�1O8ߦ:���0�:|�QjJd���<�@�!�G��'��ۢ�\8�"��l���������+�P�I�X�4��ni S-a�,��CB$�L�]I����HT>��:�L�'c�5=��l�d��?>�x� �u����).R�y_}��&���(���H��D��m��`���q��0�%����Zޘ&q�U	땂��x1�vW6�A>�|�� ���aT�`��~��7��C��qR�lA�)��,�0�a�ͤn_�V�9/�^ו��T�\�`,7O���X�z���΂Ch'V\N�� ��Ƙ�۵�R#d5E��1eFi)���%׏|�b�@�9R�)��SnӴ�aC24��������9E��{�L侙����v%����� �i@�k#�|��~1�M�9$m�[�H�G�xio����;G���
�'R}q0m��ҙ\��mc;���j��Ȓ��� �����V���Avr;�R�>�U �J޿��|�#}���i �5��_1�����O���F���?��#���_����&xH��e^�ۀ���}V��/�;Վ�zk�;88`I`�q�D��}��ȋ���HxL���	9����4G�`;U�7����fP�oic(�nL��0ź�d�V�莻ظ�l¤�,8S	��7��v�'Y��Mm���ߛ[?��S��ܯ���O ��e�S�|��L����G P�yY��m�E����:hz�#��D�Q�/�����l
�M3+�ɫr��0M�%�e��SSH�4y�Z�-a�/�"�}!?,k]]\2#��01#=;��yn��I���FL���O�V��(���!i��I�^A���`OY,9f���&m1�	}�1s��6�����k0cg:�e2�L�Fl�-���2��
%�6��z{Ӧ�ܺ�W�7�_糌�V� Rء���7��v]���zQ$B5c�͸P�I=s�䎐�����ӳs*"�r�Cwyy���� �@f��x'1'����H�Za�W�j<��nP��Ru����-&���%g��c���� ���h�}�#?�k�]�h� �5ֿm��r��&"�La�����~*Z��?�?�����J���̌T营��	���a3J�z�.	�����`���ĸ pe�Ʀ؉X,t�9�K�PbD�=����Kqλ*I��__+|���)&�.1L Yf���Ca�����F�(� T���7�<S*d�D5e)�$�ӟ����8����u��,_#���������T7�s@GN���� d*�Ǐ�\�X\�L=~�w�YJ��w��/_��Gۤ���cф�Ղ4�`C+�z�<~��>J���7��:�-ݼ{�_��_�wvŎ�:;c�B�vr"�������osخ��PV+1n��u+���$3#��W���A���<����s���ݱ�yl"�!h�Pҍ�����8�SX�}c3��*�1�.�}�6H�Z��fya�.��RW���Љ���T˖C�m�o�34�\"�3�J<&�ɹ�����e6��V>��#˖|(�B��w�Z��FQ�i�0����Q �F�,7#"!���_�C]yy(�%��o@Ht@�ʟ���kKVP��H����l8���Ҷ��� tB1����@*�s�ڲy�4����hlH������/����\���w��Q�57���̞V.�y�Ƒ��������Vmɀa���j�&�4&�ߞ'H{�D� 	R��k����<ͣSǴ�?�k'�'�}�씁���yj��E�2��꧿�D���js7�e�D��v|k�t�F�
�v���-�A�h����r�{@�/K���F[����c�d_����s?'Z��?�7�H������|���nA�(���j�
M�`�5.o����ο`}�<8\�|6d�u�X���"қ����V�\qcE�q�m�ͯ�8K4�%L2�@#���`Е�?�Y,R̠���d\���9rK�u.ս;�:�:��S^7< ��0G�=��]�{��T!�O�X�T��צst�a�;���+���mb���h�q֜+o��*6!ᔳniSr��N��E��n�v��ь?�egH�nq4B����a�t��@_�����,�m�)�힫�(Ի�����q4{�3�wCqfS�MQ�� �?Ėy��B�n�T�'�ם���a��&d��h&�6vJAD�������"�N���Ucd����]��߽{~@<99]T�15-�25�E��(�gف�������
����,n��*ur)� y�q��mG�Np��Ka2Uռ3����z�������ܼq0�(���gN���l�29��U�d�I[dC�/k���g�_>����������D�79��A�uӲ5F�y	�D�D�p@7r�i�$�e�$�'A��:.�gdH�u�i��Ԧ�:��+�+J]E��|@�R�3��0U�F�TGJ��d#-��������#deL�9 ��K���O��U��Qd_Ϗ�f;Se�_I�\�"�qW�����,%pa�m6�u����h��]�������٩� �Y�4)9X�9�D�iH�4o9��gD����TV���^-{�5���rqqq��&��L��4m�JPrx�lA���8N��E��gϞqe��(!j��!j*� 7�LZ�1$N�&AYM�9�Q��޽{��-�}�ـ�tFk����[��h��$���	I������SRIiJ�5g�ܖ�h¨��� 0��V���< ]j�̷�Y�����}?q� �n\2�)q�'�i?b�|i4,��`/s�`�:t����wp�f��V��^d�VB�CfN_��P^������al��Ag,�+�RMSղt=�&s� �El�:�n/� @/{"c��S�{A����;�{H�EEM"�P��֭[�7�f3��$n���������n�lT��������0�;f#�&P �ףp�z@`���f]��[���*�H^��mM�k���S�O�d�o�X�C*l��{o���qU6#;eC*�YLX@*����a�i�K:��2?F4�G�H`�0���5yL�E�B��Qg�ԙy�\V��U�j*z�?�{���G���#�`�]�g�M���X/��2��6J���س�Fp��.�fC?�^^-��]��
��5e�T�K��,���lj��8b5��k��o�0���FE�kM���&e{��ߵh���+���cG,��0�-]\]Z\��ΰ�4>��/~���c��G�"ĕA�6��I9֌Y�1�`�A�G�#ņ=�E��0�H�1C�&�P��Y���"�V�[�����������XPE�
t�4-����4 sH�?�o9R��
j�ZB���_��Ŕ6��#+���!3��GWS���>���?����MLݝ���8<�O�}��|�7�|����߮m������G��K��#Q�b�OO/��?���>6g��ZI%�qyجM��O�����8Y�v��/O���T�M�3�f��ɓ�}����/��/O�>{�{�w��/�]Ok�?}�TNM]�"l<���rl��ꚙ�K���^�bX�,}�n��d�E�o����Ypqj�TN+m�dE��3�4^�(�6՗��E� �N�L�&{�勶�U�=��R`xK�4�K#j�zm/���yq�*S��;�����eo�	�=~� �2��� &g���{_�_��K'QS]_�Z���?-1����'[�*��`u��L�u9����f����=zr�X�ޠ��H�4S��m��(hD����,�J��'%�m�V�����
��$zP>ƀg��������S����[S�h�xl݃�5���>�q"ƍ�[�0ʲ�Py���O�p_�@�������&�����$�:�4j���8�%GAt���hS���e��.r<%xQ�ڮCԈ�O��Qb1��A�Y�Z�f�V����a����R��e�x|��͓gO^����\~�����~;���~�g���X���/���ݩl<}�A��֍���\-�~��f��K�t�/�{G{��iݼf@e��H]��(��g�=����m������B�Ծ���:ÈH-���Xm.8�S.�����s�9�M��נC�� ��m��k�-c�4W#��u�kˣ�N0��,t1TI���������-V��`|����8K��=���S%]gpn��3�E���I���@4��$xf�����4�h�-�)�mR�����<���p4��'o8���hH`z�C��=d�� m@-��@�s��x᫥�kb�R�#I2��҃��F#({�_z~JG�ؼc�*�<յĆ���*DTEbkcq�!:�x��ۄ_Z�`M�\���z��y�z�YA�Gӳ�� ��+j>�`������!:�f�ro��#��
�)�1ظ�¦UR��~(W�D�����7�Ӄ��r�h5y��OW> �nYf�1��[0&6�H�9;�����/1��vͤ�P�4��/�)�u�q"��x9h_	\�n�{۱ �:P�%�o��s�I1ʌ�U���i�������XK��`���4Ѧ���܀T`UW�'�'�Σ��D7��R�Y��o��� �#J�XTi~���X�(��l�VM������,[��"J�aZ��g���� ��K��ƽ��(��h�A�Qӓ|U5I��VG����:�O�c�A�M����|U%��$)\+e�Y'�bVƁ~iz����$qĦ����uM8d��F�rk�hP�:.��«	�9��tކF��XAm������F,����Xo�)�.%��C��n��1��%Lh�^T���!!)��z�^��b8�i���e��_���ʟ�)>]�@B�+���dsP����T���cf�c$Nc�ƨ3��֚Έ;s���h\gN��n�lغ��Br����Nאu��X3W6#�0wkt��<Na�UW�M�έt�v��q�|�T��z��M�qU�Q~��ۦ�;<�E�~j}�W]����;���Ʒ�>YPI��˜(�๏����Y�"|�{����E�!h�mǝw3�k����#��:}�o��$ȑN� ��Ζ���A�v�$���A���,�v���� q��K���8��:$���#UC�e�u�v���wRQ!���Ω��(BЀmHs*���'ڝ�����TF���,�(;ryy�l^c^y�K�mZ��t]�F��S�n�EXo� Ҕ3���o}�i�P<�]�Z� y���j��]|��$�
���p	'C���R�����+*5��ļ��72��G�'b
v�}��T��%-��>�|��+�899�����bOv�Ǯ��v(�mE&����ӧO9j�����j��R�O&ӱ=�f�W�S9�rZ]EQɬ."Zyհ���&�A�zz
�,]��	����`~��TV`u����+�6�\�����[Q�d*�L�h>�#��Qm���-s7i�E*kN����7�9:>$��w�aFԸ��{�~���~���r�<�$u���G?����N�m������S�dK�we��<� �S�����~ɩ_��v�@YZ��hwB�����#�Y)www@������ �#�~�����z�i�C|���H,Uk��\^&"E���NF[���q��t�S8���v�ſ5p�p6j��^�W�$��X�;k���ݛ7�e��`���z����&�1�z<KM�j���|::��V�W~=���O�I��E�y?
��M�F�}-ZmD�0,{p�˼`�.�f���݌���Pݡ��ހy��~\4�' �ΎD\Rfi+��i��J���HWf!��I|L�F�2��u�+\]/y{q��,C���s;���ZG3+�Z�i* xDLg 3�9��X늨�6N�њ����� ُj�
����#�)	|1�������j��h�/%r� �&��`��Ս#���fh�S볊ʁ�'cf�"�.�L`3�q��W$֝7n�f�A���[o����㯾�* ��S�[��<�ڍ���f�ͥ�9�ZC����s�u^��G�d��d�!v�w/.Z"o���C��M��`@��
=-A��!3��8a��F�T`����7�{냿-`++�w�˝����Fz�a��urZxR��^Ke�T�����HBJ�Z�$�N�B�j3Jq���8��ÝM���{�#�~�1��Q��:�DO�x+z�y�Κ��\���B\�%Jl]Gb)���icX��{�Kc�}jMj�.0�ț��*j2k6d�V�&�x�Pd�^��:�1���`�WI)�,_QCk yl{l�:LI�v}k�F�|T���L춣'خӅ�u#n]�~�@�I�����6��d�g\kz"UV!K���0�|e��a�o@�4�1�����|&�+����;o�d���T��mT#��Z\L&w����w�������]5ێ'�?/�T=����iH�"�[">�Q>F�2�0�cc4��F�l�D ���bþ�!�˵h��(Ģ �Ӫ�@�c��%52�"*��ll��lZ}#���7��f���ذ�`���H޶c|\!��L��\�&�|y���e7��<z�e3��z�G���k�C�Ǆ�R4\�L���@�r~��$-���{b-qfE�R#gn�]���:�Y�q{�Yw ��k���H�\g�����ڈ�-���@zQ��X�K��b�#"�\��IT2�h�P���l�������������'�F��fJ'�O����x	�7�v&�����F8�&�  �bKOy�,��)��r���p�������=;�Nt�'Y���Z�A̔�%��",��z!U^�M�Tk��?L�2����g/��&��tv���Rɵ����^�CP��Htش*%��-]\7��M�"�|����\�+���B�|JA�ŌI@9}��=4F-�'y�tn ���]N���!�ZX.E�_��E�����AR���pA�Y�&��U�IFM�%@�/�Ua�N�3�5�ț��#p�4:vcJk:�L�@�~X�/�||r{GЫy�eT�(��6t�8['$�a�F���8�"��wwؔ��	��P8�J�B)J�i�Zi�P���?݀�(M��!����>��z�՘�j~�� S�Sj��?���ԉjȪ�4��r�Ns�h.ZOG�9��yp�Ч�RRQ��NM����嫳�É �ڈ�� t�٘g)����d���q�.�S��Y1,d~|�8%\� O��hέ��4������TQS��te��Ns��҈o*��M�B�<������i�W*�e�§>�
#w����������D1>���?��z������OUT��s葉8����⇦kqn6ou�H�.����/V�F��S\��bF�\n���WKI_�+����؀�!�a��A8ji�����|�$����y�a7�Oq#��B�[�������m����t���%����1z97�j��.���睝�(�z������l�؊�^V��S8ty��A]'�E�*�r{i]g�v�S{��U���ЖI��5I�pn�s�Y���aG4IM�9E����L���������g/�N���l���I)E5N�3�Q%� �LSB!T^�����p�2M��뙸���Ĵ�U3�"���F�/��+�ͺ�H�+IM��ѣ��?;:8$z��[��N������[7���k��g/t�'�|��(1���٠W�ճ��~��b�hM�8��l�n��!d�$3p�i@w�����nh�wf�"�8�:qW����c��{{ڬp��]���|��������ݻ7���&^��#��ZmY��&V���������秋�Um�񺻿����n����-+��b�K�5�OXY��_0�à�x<�CU��
+��)l��j�)G|��z���	
me$V7g�M�( �40�."o����~q"r��U�S���(��x&8S����|gݮC�i�F��� Tc%�� �Q0Ǝ/WK�R�s���$\_����x�\H���R5Zi����b��N�b�"�F�+��
)�T���3��f6³�I<V��yy}-�S��ɥpz��$�Q����Mb�J��Rj���
���{э�"�(��Uf�6U}�3.���N��~^��s���b�a�4�b4 ����,861hڔ�����g �t�"�UA[�!��)k��GΕI}���+p���W���&�*qG�y"A�S���m�P��Zn�7�<��5z��d��o���nNg�rbd����{o�y�o1�e��Гm���5�=A�z�s*FN��Km�ٟM����؇������"ک�R���Ҳ�˧ W{	�Jo��8L&�{�����C0�I��Մ��D�"��2_%7��(�_f�9� �9_3���2��	��T�w-����Ů�;���DaD����G��7�s��E�����~���;�z4�	���ڰ(ڱEр��y=Rfi.|JLN5Q�8q2�N>�,ڔ�����o0d���{�4bi~��C��A���6Q��,\�#��~4Ș������Y�E^&`����.����Y̌��f�e(\*�gW����G:~`|�ݏ_�8��Vb$my�57~��*B�&�2cT�B�6����K"�/��Z/$.UM#��1���F�Cw�TG.��E��b�rle�'��=�c9lS���V��F&k�ٟh��?�,F�F�!T<�[7�y�*�{�Opvv�H[>(_`��ح[����2���}����N�`�Xd��u��a"��5�$P0xҘ<L���gt}y>�^��I]�
�I��B��o���/6Z;��c���~��SA|�G�^�
���`k��B�SY|Z�~Ճ�r��m 
�S�ef&V�3Lk��R��!�t���BL,H�VOY"�'W$Ӂl��8�4Cv}�)q������X��
�����εaP����3��4I�������vH6e]P��s�g�&M� vN{�8�DBu"S��h��z4�j�!���V��Em4Ƀ!v+k0|���믿f>�%e��^��&��#�+"��*�"�90cx��F䪔*H�v�ΑsK�I(�s	P�ܹC�9r�܊]��������|���|ſ���D���E&y�bH�T��I6��qm��1��	�DTɷ0�)� �"%�(�J���X��TG!uz�ޥ���Q���c˝�WP�zqz���9���#�s^j�w���V��6T�(*OC ���A�1�t0�Y� (�nUF��=�h�{ZC��x�,��,�Wi�㮈���(�n߾�w�N^��W-2�@�m�pc2��W�m:9�-|��ƨyq���ViD�H� [�]��!K�7
0��[u0�5]vzT̴�m(5@��z�D*����T�����}�P�W�<�&5W���n��hG׺���'E|,��ўO�8jud���7�-,t�ݻp�M�Ig��Po����T TI3T���Uj��c`/�%x ���o��7�7������+G�� ��D;g�
�����UJ� �{_�s~j�^A��r���8\��QqDi�b:Q��,Q���{j�-��n�s�둡�z��S���	x��)]�p$���PK�	dX㷈���*E��4}�Ⅶ�����_�����(�����Ŗq�wU�Ф�/'��Æ>�<��{��1n�\�RӠ�Rr-CaC�6Ϣ(���Ȧ���d�6:�(�yx�<;c�Pm��,�Di_"Kѐ�>	�j�j&����>l�4��cdhBb}R����ѤuOsKPxx�����)�8K������o�EJE�8$DW	\�TP���u��7��_���wѨQ��	ا�,�:bK|I]�jޞ�O�V�ҏN������5��)�#��֠���F�'�$z����ӽ�Kܠ�xӬ&�,��>q�#�OD�J�[����B�H���̟!���E�ϖ&hy |���3DEZXJ�%F���Q0�-mbI�ƶ&�E&?�u8��]O5��z�%'��#9�9*Su�o1X)�H�7��j6�zO���ݻw���f?>{�L�t��:�[�8?*%,>���,!mZ�ΉD&�/��a�ad�-G�A~��@�@īc	��<2t6�MX��cΡ�2����d}�{�O��1F�5�Ҡ��`�.���F=��ն	6���¡�F(�[�u�lV;5 ���s��cl��ٚ��}�`�ޛ$�.W0f� �٦*/ #��=�KW�Q<�.m�n�d��	��S-���|]m�����O��q�s=Nt8 ��D$�0�˰߮����@�C����Ou,Px%Q�0��i-���ۧj�_�(T9{DO��#������Pr<\�x����R�ۆ��0d��ozH�&8�R��UO�̭�Jm�q��O���!O]�zC�|�\\�Pq�6����@�7Py���^Z�����#���,�E�[�@;K�t� �NghYݒ �w:�p�}+r���潄ي��!r����R����X���6ԁL��̊��y��c�++q���Q�:�9�q��6�&���&�;'lt}��n0E*Uq�5�ʆ2u*�k��Kܡz^:�'���#v+�P�|j�\s��3̥��Q� �l>�<�]�Zڮ��؀�ͪ�DԠ%����Y�;�/rM1�������}�9���)��Z�nðy:�V�9��`�.���pO��Y��1��.G`��R���S�y�%5H5����R	�@����t�6Wg���K��$E�V��*g�B��H��BL]���&�Z1\�fF#��������UW붑m醀C+o��$�O(7N�qV�wԏӹ���p���u\�B�9�^yQ;hn�z�u����W��%��ߑCL>�e(���ŷ3�E�yν��iVh��I=���ɬ5��:���K���I5	Ct4��wOzn��
Q�B!���]]r����K�;��Խ.�2I=ƶUJ�Nr���Fc���PU�5m �X��IT�"j�	��X}��<-|�t��q~E��ӗ//��X]��(�qC=��P �'�y"3n��̽�ޠ�l��)�"�������>tij���$R��Cq��ZK�G���*��[,�V���bX�����?�l�逈0�J�+:ȣ���=���p[I��T׋gg˫���۷t?�oU-7����ԕ�ພ��ND�%J��bF#�}�Q,tp0x�����XqĜHĄ.b���e��uB�Vô��WH�47M�^��r�k��5�QA�S"=�3��y�Tt��S�1�z||,O��K�LqY@�)>�U�b Z��?+�"�*���SoH��s��ˌ��f&��Q�n�z����6=z���x�P��9��yZ�Q����ke�l��o�Sd�8U�^�1Lg3�Ft�-�P}%h�'��햯��<&{�{��p���fEGYMC��q ��]v֪L�"����HM*����b����lȣ��/���m��t6Av �3qyuq�����]PpF�����t*�ʆ&�㫝��:_mQ�BN&IP���lr���,�Ѐu�\��JY�D�M&��L����-���ϸƀEn�Y���:U�Ib���[���>Gx��e��!K܅\�1���m�������Ș�	d��{�Jkh�~A�UR�c��]zh�q�@�K��GX� �"�/D��?�&�M�Y���5�����#��3+�j\FU&@1��R���B�� 9��{�
���Q�4<��h�l��B�SE��x�L�bј{�ɏ��mp���tU�������HwN�K{�]��ƪa�7r�⤔"�}�l�Ao��%���n�ԓ�ޞ8O?Y^]Syn�ZX����= �T���Uur�����?zZ��vU_Px�]���=L&2��6�fC DbY�ԺE���j�Ν7?���L����6�['��f�%�>��	��N��e���jK�PiL+zEl� ۝2�ә��o�̉Y*L����qڤ�/��z)�,�<����F�Kh����F��ї�~I�~�ρ��r�n��x�����H���/>������i����7ߔ��k��a�#�_��+47�����7z�QG�Qw8l�l�`iqK� iY�a�l�|3�˂D�����N(�&C+s�E��_O4���ܫ�����W#������2�(�$�S"���?�!��;;����^�<�srrr��}�%p)эK9�Ķ� ����͒�h�r�h��$����7���KV�\dh�Q̲� �Tt��A����FD�͈��Cl���^��9��'c�d+��Ÿ@k��EI��mZ�o˻��#&�{��PP���ї���\J~�w�ST��{�:9lYP�&KXf�#�Fe+1O��	w���*9�7��I�X�B��AC�-��U�eH��FCAi�e�cN����!,gu��rd'�Աib"?U�5�J��-Ec��lC�J�6�,�臭`���l6&����fo��b4�4M�7XX����i{�fN�wE��#V�n�8&�O�iޥ�CA�':?���4�ڵ�+ͳ�Rұ��T(�2��Y���e�6ʉ�^�2�5�Lsz�9�o�D��Ə�i�� ���|�@�ʧhZ,��������E=�#!!�5���T/A/&����;��Ng��Z#&R�i@W'�U?�-�'�OU�W��`�hӃի,=��U�� �˞[R̓q
s�~�È��?6��otɀ���R� p%Ŭ4
�,bm�:eB��F����D2��)�r��d&-���E�cW-�>�=l�)gm%���?��Jʼ�D��`U�_��J����g����Kޥ�.����ٹ��@"��AI0�����O��ҸF���M FN����1Q�'�����ER�k�P���@v�N��Aq� ��y�u�S��A���	� �gY^+�򮅋��o�9ZO!��73��s$B���`�i�+d|�zj��Nȶz���cg&���8ը�X��n���pz�)X���5/�G� �w=%��3LFf<�î,R���q�?��G�<��P�?M��m:{�U���Z�;;��a��@�*����d���=��d�>pB�A������m�o�g�#���z��y�,Y���Q���ms���s�\E�@)���*�8tu�c��;Ub"[W�Ӧ�&6��]�1E�DVP��hr�+ �sv
�yJ�6φHO��S�  ��py/[�c�ht��4���4�<Bw�l�����?��a3�>Nl�tґ��Ƞ�>7��c�T�)�]c��LI5�+��H�>�g�]i,�y��M�����%�y�Z�'��$�J�C/'Ӳs�i�A#����?����9�G�8qe��2/WKA,J��"i%t@�x,<��?�gJ��傡R�)�$�L[w�Q��ʄ��+� ���cM�c�Ptj�=�#���[�4z�ؘɒ'Ȯ��y!X7��m�����پ�x@��,����۷nݒ�>y�C�%�G���e
�8��Y(��y\���?�Ѵ!�b�=�#[E��`��
��dO}@���f���nZa|�t��H(���G.#U"#�Ir���.!^I^�#��Ҽ�ޚ5q������t�`L����*�
f�5ҵ�<S䚔o��u���'`�M��p�ӼBG0����O��e5�ֱ�����kH���lMb3`��t���� 6(Anh_�U��J��S�,�	f�c쉬37��&���e�`f���G���y��ޮ72�4PS���E����{v���F3w,*Pki��vЯ���ϟ>}p�����e �gqYrG�>�2�X��y缠����y
�jp21��BPU�z~~���yiQa`$f	�����'k��CXX7�z��#�����Wk��\�&_;6M+�T��̠.r'�l�j�Ƨ�i0�lXtd����L�I�ُ&B�pi�R�	��ݑ�����.PS�t��jn]2�.:d�˸����X��88|��ᣯxބK�l+�!	�"���U%�XXk:>�QN�#���N��r��EB������tk�#�d�Ld�ez�!;kQ��a_���:$��&/~���t��%8� ���?�{�����;*�<sPC��ۈ�sfW�š�a�d�C�U�K�.W}�8�|�X1h�S*Q���,w�q���B�u�-�{�^��ӛ7��W�e!�=��K��[7AG�1Q(����� O[c⣡��ӃG$ b
V���ҝ��~)�eF}��,������G�D�ҹ ^�w�ІQIf/�')�Ol[ntT�ScnN~C�bp���`U�̑�ɑ��r�B�<o1��N)��,YɥH`J�,��5~���+����;\.z_~X�R�2+�OM���3}�@����4�~��z�hV�#�yg0L>��@4a�1�D��dR���[�
Ƅ��_y6=w�+՝G�n�<���s00�~r#]��ͣ�`s\��O��P��:Q�� }���8���|QK�'��|tB&��F8tV�D��k��RDӜ�$��L	��y�@O�T�&�?����mv�K<Nd�D��>Xn��u</@P���fsEQq����cg��N_<��[��Ӂ��Q3pp�3��̶̔#إ�+<��a<~w
�0�*ɭ��s;�Ϡ2��lD��u�#�G�O��o�G,����pq+�)?�';[ؤ�h�u�Ъ7�F�A�U	���FM$�~r*X�[��8S����Yo#,���Z��< �v��F6����+�g�,y6T����s7�z���2�(�%�]�e�SO-�3,��/�:���m����@�Y�,9�Ab�"���䐣@T/n}����[#�Ŗ)����y�{�Xa`|�fq�qOe1kͻ���	S�Un���Y�GX�y[y-ފlZׄ�LO�X��#��j�]�fz�"��D�f���^D���1Ր�*���d�*0T��ܺ���,��A�~f<*�G���݃5��:��4b�z��;66�VJPí�ޭ*M٨��\�D�G���f#�:u�����@@��ge;(�4#�"��X;����2�X�R2�5�pg�XT�]���K�\��~ .19�pJ����f�<1^���h��� h�@�|�_eI��%��LJ5"0D&��w�jq���>�Y�P3D;�r�w{���ެ��UB.]Nmߕ���t@����8T|׋�F���f-�Hd"��
@�AI.{H��d����^	�\hj&�(�H�Q��<5l��	��H��;��3��C�ԣ��>S��U?����9�pQT#���0�B+�σ)Y,N��w��xţT8X�����p�(9�J��|һQ��PM���C���f��e+�14ɳ�]�E����bRϡ�#�v���sUO�={yz�!�ܬz��Q=�����^.&�p�����6�j6��7o޼s�����<V/�ཷoݾ}���G�1$뮵͝i]����I:��9:�GG���^��BU�rfQ�b�"��0& �u�0P&ۦ��&�)�Н$.����_>��'���yT�Ny&Wc�'X�/>0�Ae��L�����m��O��A¼>� !Ђh����[������X���ǌ	�j<&����e�,��~�-;��6-���ݝ��}<�\�<��(�y�~�b8�=o��3+rhP��{�&Ɏ�\0"ΖK�ݵ����KRC>ʮF2����yF���l(�#�$�@�X@7z�-+��Ƹ��y��L��V��<yN�������Cb;��	�Ц
�UNq.-�R�t�DI&�pl"����
�>�X� �Ě�v���٢u5�˴^��У�y�~�&b�!T�a���
"�GP'�-������Mg��zg-��z�H�6�%�It��)!438g];�\/���-6W׷\X6��Ys��+;�{����L��G�
��Rm�-�Ҍo�"^iɤ���Mu�H?��*G��*Eb��aef8M��H�����)��[g��V����2�?�K���r����0�L��|�(���G���e�d���C�jQ��̓a��Żc��z�-]�+.rx�1dxLm�H��y��j}Yd��ә�5��ik�qnhU�t܁��&�@�3@n�c��X�j�f?�)��>��������2����,[��$$d (x9
�_��� -4�����%ۭ��
|6%���xf�U��3���jO������D+��N�2?��/�ܮWtjh���lΓD�zx�~N
������ &�jn����~:o%��;��Ҹa�4<}�����e1)rZ���k�!*/��a��Nb�v�殤�VmB&k����91����Ԑ;��w������ww�wu������G����N����M�d�ݚ��U�*�v���������!��x���˗/i1��ѿ�E1`�+-��Ǐ�6n�t��/_�y�b�G�����u'��8��j)Y�%t2��u�����D�4?)� U�	�Y�u���\�-nn�VK�eM���Q<So6�DnQ�g7Ik�C��ZPo��.qF�j���-����A�X�����(����n����" ޮXy����� Q��)��2�-Md������DvPJw�ل�	m��c��m�OH�1�dY���~���S�hP����������ŋ�7���ꐉsR-��nfd#[s���
�O���%����5va:�����h��K�4��%λ�
>0�XƌKE�5648��I0���ǁ�熖2�3����X-ӿ�WH�sd�ͭ�Z9e,5�t,;D���%�9ŋ�(&(�ٝN�f
s:OߣV��_[L�����x�A!�^��A�킦z�B�a��l4��-�6]�f��)v�����e����~�(x�Xm2X��;������*���j�Z��S�W$�s�=�f��;�Ϡ/�RȹS�$ǅ1���r�n9=���+��+ұ��đݝ�&���œ��75#����B����9��":�o2=lZ�}�.��0�9��§/e���V��J�����l�mq��2k���L,�n��%�@�$�&��0/(���J�pB��$��~�A�S8�KN�fkQ_�d��r�~x0�2?��xC�rkxf�}ʔ��
a�1��yp�rI���W�A)��"a��V��42,�vIV��p"��csMe����XV13�h�A��|(���+ b8(�A: �d�d/�ȁHۏ�q�s�h�1V���s�)��n6+���\�,V<���(�:N����9�E��^s��X��A-�VCn�4B<tŌ�S�kT�H+�������N�c9�I[I!wF0�V��>��*e)q������'q�#�{ h�+o���w���.%_7 �*)g2@���̲����+�S�[5�x��-���	�_�2���Nz�y��Q�<
/+�5/3"����$�_�59�1z��N���P�9��ά\��[�DO�2��v:U#�Ŀ��t.5�b4��l���ݻ��[�����y��d�҇�נS�Mu�BY��ذ�c
�?O�\���_��&C:��}�
�!Be�Si���ì+�Q3%���=(�J�:�	0.Z59�Q��ϟ���1�2����a`����U���⎜�j�p:�uQ��v?���V��ڙ�sμ��HvV�5tW�Ӡ77�OO��_� $(����m��RoT��t
{E@*��
�ډW�d���#vǽ���g|�O�.d�X��oo��O
t�'������˿3&J��I� �](Ȥk�榏!�&�2?W���!$t�����7�]QHc3a���N��'����[�Q1mФv�$} ��HBL��Ld:%#!���0�7$�
eY���i
[�����w��i�p:Kğ��=�99��km�5��c�ݰ��ܓ�P`�h�!������O�a��S�\.�<�j�OR�����D"�ߧ	�i�)$���$�	ҵ��Y;02)�C�I���S�I��w���e@���TZ�[9e��Ga��6P���Ҟ��DR�!
���S�7M=A"x��ɥ�����N�w8bAҝ�V�+͒��B_��D;d<x@���jN�iϪ>��LE�)��hpnWH��_Pۮ�8���%������h��'tGb�d[wlq���D	*�{��-ݜ)�W�x�B!S�����\�3���8P#����gǵ�A�k����'g',i�rЂ$㈉2/�l�6�:a�yDX.Zj�]��L��!��:��9�[�]nH��)BS�C���P~DW�ewo�Fb1�1��6����*vS�(��Ѵ�io\�s��du�+�	aU%VШi�^�Q=�/�$��:��O^��"HuhYZ�'�4���@JLky8W�S~46ѥ	?J��§zfiX~���o^3�yZ��
j����@9Xh�F�k`;���UY���ߧc~��R"�j�gX��3{OJ��cgr)�)�8�R!��X���n�3�>6�崶�����������^�z�H���G���qb"��5#*��h�h$ÿ�����+��i��R Ѷ��::d7z=�{�G������o���T1�+��iɏ�ys%���u����W_�e=z$O�߅�-�M�d'�X�:�CQ��Ț�-��$������c��[y��ۤ	Z�*��T�hl���:O�������v��g��lm{2��W��(�T�w�&��%�RmL��Ǘ �1{%
 1C�	B�l4)"��VN>���8)dB��U߅��t�m`(�zG�UC���/�8�G��	�a�xIP��w�[�R����������FS�pE:���{�<�)���^���pLl���6l��6�`�Q��.{�4�7�K�98CR�+�<���LdkB�	yn��$BNy��5��('����h��da�ø:etɕ`����#�\-*�EP �)��	��A�V�쬆f�TA�X����y�;��4�;j�Z���'�-u�Pw�I�*�
%a�Nt<���?@�QF;n&R���qŒ?� �`�2�^�s���� N�v/�6��8�Ŝ塬�u�=`�;�@��2!Z�h����co���Կ�EX����Į��,�g�ʏ��(��k�-E ��.��U�e�7zY�9�/o�N�
�i&躎�28�u���Y�u������(��t#}�t� V~^�������O��9/դ�MȇI���6g��fRV�>`O�~1���K�@I;�#��z����hY�=~�p��SXRU���v��!��<?c6�����_bv�����(h�.oWn���$ZS�?w:�Ż�5�2�`�̋�eAwK.E[��o���i
�Hd�	gWr�w;�dd�$ax��ߺ�qD�[2��E��F�}�<���RT����A��(��A��	��55K���+��W��Ԏ�ߕ
qrjv�ip�P���=�nP�!h�n��iY�L��6� ̬���=�����T���Q���9�H���Ԉ4[���W��떝iӖ��MO�˱:��f6�tܝtvz�jF�.����,3��"��Q���,�����W7�D�-$晘�<�|m?H�i�L;��'4���`�w�-G�>�P)�2�ڽ}��g8�K��Od��;(h���oS^�2�n�+4+)C�z�( -�t�&{����݂�T��v��!��xtG�jڱ�7���"����hĻz!���ϧ"��xю`��fӝ�I�7�*�D���<G�?%k��+Ӑ����H@d�L�:MI>4
\ڣ�xȡw���(�>�]�J� ����N� � �����خ��$���u��7N�1#�q\	�:�6�� �5|z��{,u���M�g{31��ݞܟ����//N����w���3R_]m��8:<�k?pK��<����>�b��%�W�Ŵe~7�6�͚�,�O��7��Z姟~����|Z4M 2�u����Τ��N�Pi�����mH�Dm7���+h
��t�m���[p���a���Ų��;j9N�I���O��p��[���0�Ob׍��֬�N�u��ٙu��(�;==E��r�wtļ�/_"Re��%���4_����s '777t��W�4���;��(80�'N=�\<(�#�Ȥ�C�I�f]������=3�u�G�z����:̤s:��rޅ���kƹX��B?�>/������Z؝���.��1���5M쩡��0���>�C�&]���,�K6�����<�
�!���穰��K_�m��a�l�9_��H�e��PV���N9��ԍ2E=�c �@��_�M��bП�Lj*9�9�vA��QË9)�v?��dv�M���3�z�nb��	�ch�� b���:�M�V�
��2k�<Z�Պ�� ��87c%3���Hu�|�'̦��k�L�Y��;*��i��VՖ=��"8���6�����I��?����R\^8��۶��fZL��)��Q0oЪ��ۻ��V���,��6�N]`�~;��,�U�^���tl�]�l �ɄY��0���f�)/WF<�qK�ˁRY%��!8���Ze��|uuu)ٽ*�C�9N�\ݜT���{�@�9����� ?o��z�!�R�;�'×��r2H7о�y}�]P�?�WAJL�����w��mߚS��Nt���Z�((��X�Xm�4��"&�	�wO�>�������gt�~���N�쌗4�ك�A��9yzx�yw��a�:H|���H�"gw�r?���x�6�~	+����|೤Bq����KIw��7��N��I�������"O@�R����z��-��?��?���)�Zw~~^�};���>����.�98�t�n@;�����RK��t�bG��U�Ph`�
t�C�!3�����u��WLI��ΙV�Є����7�U3�QKAX@It�"�eQgJ�$Z'�����5;��ݮ!6$��"2��4�J�Ծ�b�r�AC�Y�B��V�~�I��%ڐ)K�y Y�҈�b<�`��H;�|��鉝�挋��d^��gɔ௶�N��Xd{�7U1�@c1�kۍrp��̣�����ܼnDl�+��ƻAs�^��
�A;��9$!�(j���bh�:	ۀ|\aJ :�l��A����zD�X�l�����d���q�$�q�łv������{�Q|6�]戜���K��䎔ȝ�7�8��nЍoǿ)0.$�0�R%(9�[Ӈ,K!#oN$E�<t��g{{w�;�=�[�+L���ޜ�z?��'�fAF�������,�zR�H�,bc��;ʲA1��te��nύ�!�m˻y�2ߍ ��k�i�J�^M��V�g��=#"2AM������#��	�}1�20�Oڼ�B&&�T���O�g�^��t�|�>�ʠ'�X����0��d�'���mbߔ��d�^�;�(��l|b10�� È��i� ���f�p�W9eH3���HAˈE�¦B}#�O�qS�@Z��<t�EnN@�8�`]���-A�!U�5m�t�����~�f	h.��>��z��I%y:�5J��I�/�T�<�$##+���.Q��d�?�oDE�ԖSf�e�Cw��v��˞j�v隓�;�h�FM���1�� Ww�� ϔ"�⁨pV���7M�I�#4L�	�8,̼o�T�eȖ+�]��tv�~���_�@���}!�H�Kb�9ρ��Y{\d�l��IV�<��eY���R%�P��}�A55��s�����0eƖ,��s!�Q��ִ���=��0�� �@�����_��d �a��ϙ7?"S��Ӧ����$M6�����s��!�6^M�i���L���<�^��.9�Hdg#�I!Ӝ�UqʢW)У=_�C�|���K,���=������#w��������{zV��9��R�<|\dv����:Eb�������EB��Ё�h%��~j�ɀ[̟	������A`��� *�teh$��K�pˌ{��w��D�d��Q�8��B�b����/��E
��c��?C&�R8�w�Is�TOςvR��pF����t��
kȵX
�8@@�U�Y����duqq��7�����h�	ܤ�/Mm\�Dfɋ%8�Fm|�X�G�c Ƴgπ��6n;j��љ�Ҕ?:��6�}Py^ cseQhu^0� T1�����,�}
�E��%�o@�(���)[%rI�P��ҹ�@�p�(��""�@pSz=l�rx"�6��V��#yK����	��a{���"O�Y�6��3�d�g��CH���0�	��wݬX����<b{o6aD���ϑ��<v�7: �i$E��_���!j���+'�I����Q�:^q���z1a�u�?�<�Nq	�>��:j+�k�(�O��ĥ���ҧ��P�o���,s�M����,�
df��.w2儎���+z+W,�@��0(�k��qN�N��#:-�D���p�����|R�^�H���:��,��~)�HLg�ɓ'�� �ы�t�r� ֕���CW�'��"�Y�!OKjp۸�	{>�����?<�8��T2(�۵S�_;��x�U��%�hI/�)<`e��@�`�qN���������{�w,�t�>�/^� 	��\�a�	�jp��G= �x�)eQ��K�۠�����G�֛��f���A��
�Z�?S�/X������PCp2��d"tT�S���-�W}�'��]���K��^9��Y��u	���DgJ�Ŕ����y_�h׸ׯ_�o��/�zi1?_j�!����2�����Ri���GW(��8�L6W�X�2 �A��f�������˟�����͛����絠�f�_na ��!�n7���,�,D����d/ BP���no��>>�d��g�etȕ0>�`���j��;�>�^)���F"GҒ&�տ��;y�4�C���������f~�3�!c��[�(gʌ�]�(�q� Ƈj2	́0,n���6�!�i5������I�B�`�n��4�`�y���j(��Y�"���L��٠u����%
��txƃ���w�ӧOIu�N��&�u5��`���w
`#g�6�L�4����h^#���d[ɿ��Z���V	�g� ���d�u�5��_�����v��M�nH�!��� B��4Fi��t�2�I�R�i�:P�S�%}��ADf�c�)�8X	IU
����#�E�e`�-�%Z�g@6o˙a��
����m��/Ȫw�� ��
F3�%��=���H��Dv�i�_�]4-v0J����0hCg�^������2��BV&�3�j�m 3�Nn�9Nd��)���/сdɎrЮ8D^p!�f�"Q���S�����)t�ᥜ����4��G����ی`���uz����d
'�C�����"���=�\\�R�G�K��U��L2����^�@VV2��h���@A�{���"������,o��}E'�̐b��.�E_xF�Fq�[����]=��ѽ޻w '�G���ЪN����t�g�4!U$-��A8���bt�R����t�di���خ�6������V����m��R������;�&���O�9p6���N�;��ve�c�2w�Te^p�5��Ҹq^�|aBP��8/MeS��i���)��q��k��W��Xe�}�sPL�`)@��ʁ�U��1d^�tɷ��2j�'�0�Vȫ�ј�ř�T��J�,t��(f������ou#����X\L��2̽������`��a���Lj���Y�J����)=�=���Cq�Ŗw�"�v���M�kn�ʴ9��'mA8yJ�QiKq�w����`*h=)G$I�E �>D��g���0)r�;m��2E�
0+n�,]7[�ȟ��>�n�����ʶ�H�>%�����o#�=�q�)�����K��ͽ����\
�=�V�^e�p�-����R��L�L�oڦ��۝/��H9���d���G�M�i�����Ȥ�"+���B����i�-u�3K���DC�I����V�	�piA��Qs\x����l���Ag�c����d A�U*����c�HǊ���P�a�V�i6�/�����8;�Ѩ��x�tv~"+P`=�����`��M95��"aUq��1�Ejť�=��o�1TJ�nPz�5���y	W 	�fR��-�z� m�Iz���Y�ʱ���Bg$�9Di�͵y6�)���a`�!�-܂S;H�.����8ߵ�N�x��J��	�q� 28�ze� M<�L9J����D,�}s��������ُ��^;� �X$�a uW���C��q]���b1�����j\M�Tjd�}T�ru-��sy*���o�w���Fo���o ���h����rc9�ɠC��$���8�����+��dl:e�&i���]��,#�u�E�+����g"�*�0KBb������;��۾�l~s{WM.������ט��H�(�kmk�hS��;fY�̄H瘽0�p��9�K� ����@xf�7��7܇a||`�ǉN�
_H=���4϶�}���?�T���e l�%;��2�c�C���Rb;�;��iF��\�(3>�M���M&���?��c�ؿ]v�Ƕ�������ڱJ���&E� ���	�F��3�L��:���1���`�I�<x��g��f-T_�{I1�ysyw��(����6�o�P2���̴cb�P�Vk�E�x}�U��
���x{��p��I�-�g�N'1.YL)��7ʧ"2�����A41��8]G)�X�g^��^4���Cn�[,n��=�Yϊ ^ɔs�s��t�8��w�r�t1[`����S���ߧ���7�ƈ/ym�Ot6(k�,�1㐯�%}ZR��L!`����8�k;m�t��S�W����	�\�!��o~CQ���O�Ҧ��.��n9���]l�@���6��Ӓx3��`��y�3g�ہ�������Bn�}j�(�^�p���+Y�Hל̦�ɼ��ɶ�p#��O�
�� ��#L�H�gλI�|���덼d�X�|�����޽���O>��޳��:M��:ˮe�Ԇ~.��	���+y�S-jG���1��7#��yP DE��}f��G�i;$<u�K�p�j�z�
mn`c:)�|���aU�'E��!Sʹ�w~4�|8�`PfӺ�����UE+����Ƃ�)�
2e��[wsH ��1W��kТH���� �j�	����<�a���h�:�-�,�ş��Ė�C�
���P/���M��p-pʰ&^JA����rJ[��\����6;EK�QTn�kF����;��h�p��@�����+�#R7J����{VC��LTg��N��f���ޡ�Ac�>
ʻnhZvz� X9	��d����T�-C8�Qэf��W�g�~�S)��q.tu\�u�)�ï���B��<
:����ٖ���m�V�Y���gH��7�\��53Y}vy7��I��q�d2ib�.;t��=��T�/�� 2���R-(�f� qU���B��t&O6}$��	K�S�O>;H��4��F'^܆�YZ���:�i�<lh�U]tҝ�rr�S{e���äQ��N�f�`�5��2{?�уp�����^���E檸w��AR?Dkq��D[�B� �N��A$���)� <6�匂4ZP��:N��Y��[9�w6j��z-g!�������B9%��d!k�ٔ�Sy��n�w����d@�d��ۈ�D�{f6����u�֠gq��+<i�V��ꔌ�ħ��N��Ei�!t		���m57�&�6���1me�6A��M&��Y��u:2�[s�z7A������e�3� �ڛХ.�Ds���W��߽���6h1=��H	�7(7������-��Q���!�{�q7:)���m�AEEi90�V�з�U)%�ԥ�K'���i���K�W8�GB��q��U1H�wK�A�Q^��A��`#N��S�2��oߺ��Z&�l��>�k���F㌕���pX
f���Zi���<��fvR�I�I���MgB��j�,X�b�0˹�1��"|<�d7�Y��ۦ��ppX �Gቒ�Z��A��q�V���/C�9�Ɣw]T����z��c���^�j�I|r�ݬ�AM��mH���"�'(V1�<;�������LZP�X��d�:ƚ�[��^J�r�M�V�D��ɽ��uJ����`̍����H2�+3�� ]?�"�����}�zU�1���D �)͞U
$m��_�@Zk$�te���.KUQ�fB/��i��h*F�ɐ��'K�����q0U��J?���r�#C��<A x��ś�/^��0dV5��
B!|.` ��Z�5�����"��� �����#T�x"{FDD�� B���D@�	�<lm���[�q}��G��6�&�SLX�4�\H�I �B[�(���'#(��D��刮+�I��Aq��Դ) �24@LP�Emjl��Ҡ�
*�J!:�(���  >˾]�ZK���q�K�v�#�o�����f����+0�8c�O�~��1ٖ/�x����E�ΰhE�-���a��� ���k/Q����s+d=v�;����	��.K���^\��cP�&|�����.Eb�d�ͷ��%�������!(�/VWR���axiH?�+��u���͝���%4d7�؊v���f���Z�+B�V1�~D8�t����>�9����7�y�.E����,.ߐ�X-��_��F+M��H�3��E��v������N*��}��ѣG��O�<!!D���f�p�`��yLSP����ʈ�i?j5��N�@�������K��Ea�eZ'�p.)�(u_ $�A���+�܄����g>�4������*r>}��u�8�z������7��P)"��$ ���cad�"�0��w��[ǖ"(|a��q�B:��I'��n6y��_�%sx����4��NXZ!{Ȇ�� ���$�g�(^j���	2"ay5E�T�M� ���NZ(�p�%i{�F:I��W"��2x�Dn����g/H=�������OI��ɽ~��0����§�}��e�$�u�~J��P��Q�s���̴�R�4쉅 Ǣ�F'��J��4'�=o���c��H�BM�$���ɱ�
0�.�;���[��b�a;�Ih`�E'/d>d�"��l�Z�]c0f�� ��q�����k�㜕#+�l+�
�d?x�M��g�^z���B��P)DQ	s�/���_���h�S L��G��B'ݯ6kX
� b�a﬽��nB�tr,�J�Kp#��(��Xè���;�+@,�O�_7"v���ׁ��	�9B�Rr�{��n4�H������S:J,Qk(�R[��6�؁s���y��%�K����J^O9�c{��ǟп�^�%���+<����s�?�T��W(��N$�I��inXj�J�hK�4-�wI8�-�����	`o^_�n��&�r��f���}*�f?�7h��' �	Ɵ&��N�S�3R<��᰿���F�
�F��N{Gz'�D����tuȸ1'Lea�9������Ʃ�'�fX�'��HQ��s��k�oX�o��r�����-���$�|��	]��f3��1��.�󽰼�$E���>>Ȟ<zĨ�P���Æ�&�-o��S ��E��K,W��딲&�v��M����|M+뵣p�A��ٙ��K���w��
�����5�t��RU��)���t^�y��|��[�ю۵UX���DP��'��r��*���-2r�H�nRz��k֏Y�!�W,�aV-�#�eRfnt��w�O�Rw8$��bdt�`Pi�(��|)/��{٣N�z.H3 ��F�3N�:N^�,��eN���"Eδ��Lb*��C����t�$��vr2f>��M-��^��d,}Ws��h��b�]?��[��2t�p�F,��+�J�� e����R��<���nC�pR\�\��_޾-'�ݫ�t�"+����0��΁���D7�Z��o%I?�����r�di!}��=$4uR��!�<�Li�<z�$6��۵�����iy�Ih��H�����z�준��6m�ظ�Do�wH���!ϫ�#���A&��n7�gkAK(I�������;� n�b�s����"��|��D!�O�ێ�zE[<>x>,��n��C?7y�<�tj�@k#]*%/r��-N6�w�UƬ>d��]y�2m^��9/_�$���Rk����!��>|�NXx��gL����]��G*���c��D���%��O>�&�w��ŋ��������v�H⁚�r��[-�o�QH�@X�	F��(���Mˬٮ)� ��q�JRJ��8/4R����J�_���-Р���2�[,�$)���� j�	�����0�U9�������-YG�C��GG���2� �O:H��z�H4�c��)�w	�0�1꼟T�IE�S���vh�v��ȇ��?ک�"��b��ۺ������?���"a.��p�!�o9u߈.=qeN�9�|��ɿ�[����h�+IW�i�))��acB�EO�@�u_|��rK���m�F9ƴѡ��佬�z��{��Y�8�$�:��^d�i�)��MRtv���юnyӹ�����SÌѬ��o^�NvS��K��bE�X�t�h_�7�;Fy��g���=���l���̋%�SWcC�_��*=�����"D" +2-~��lry}�tM��m�V�t�n�I�߿JK����^�"U���,����X+�:���t�e[/�8�(�U�Q�g��5�������ȦEEf�&��Ç����
�ĀN�v��)��C9JMQΙ7�Q��r[�������r�x 5[:GMW���{�r�
2֒U���9��-��}�wғM鬬������;��mٮiZ�Q<d�"�����zRL�v;�aZ����t��y�����td7"�|ӑX��G�gd�͊ɤD�!s�V܃����t>a2�y�H$�Z�{Ӭ�<���J�"�\jŜwY����W�����5-��g�r����S�I�Z?�� XwЪ*4�9B�����OCŎ5-)~6��ge���2ꊕ�4.]���n1�M��Շb���gՑ�r2��Gi���'Ɔ<�ؒŧ���	n,֓�mGS��P'P�������,�V�wxt 
BR}�S�$�}�ެH��d:�#=�$s2*�{�}@�| �Y
�W���X�Bւ� XE���mﺦ}���'|p�?����
����o/_��Zw�?W����Q�I����ٶM10��m�@�nV��:t����ߟ2�������N�[ܻ��bqs����8�q�)܁�:��5m1�-�����=dR���J�dvx�\��S�m-�|���-w0ƍ, ��O������Ml�i�7-��������D87��9�Ӿ۴�wr���ۻ;��Ȥ�]&�!�c�7��&�e��|��ڭL�ȋ*��"����A8�<̤N�<��رf��~�H�L��$3�1�_�i�]�@ij�؛̥�^<{���0�������_�-�M�7�n�\#������f	{m�rÀ7���1Z@�k�cia_/n��U_^�p��4eeڍT������� g )&�޻��Krþ��[������>�ơ�ˆ��yG~a�u����)�{g?�V�����/����a2G;���eν)�φn^�,�y�/�c��!,B�7�Rt�9,>z���]k�5|-	��A�
I
i ڠX2m��d�ס��m���E���n>���s.����t�C�Z'����P�r;��� c��X�#�}��fف��mGw��S�)S�},��	<��:���(d+vB��������j��]��D�uu�7g���ma�����]��<�R䓮W[rOs�|��W�"��н���y��m:G_�3���{�a���jt����MY�A{J�n9�Ɏl�K�lj�'��TR@�|6���ΦN�����3���2�$$]-�k�!�j��I��3Y��R ���3��|u���Ҝ�̉&���<8�ZJ�5��N&cd�:dR:���r�)�����'��<�V�}(.��������7ųGU����'<��-;RC�=��j9�M7]���K�I��̪b�,��fZArf�̆�k��q��q�����~g���'G���u���Ϟ������K�o�}:�Z�y"O���o�[�L��rLN�|�ȁb%��}��YS�Z0ŒN@��V��2$`�.��2Z42�d\�¡#����|��Y�-��Κ���⼕Bb���bSw�  -"*�[\:5�N�!�r����o��� {�ۚ�����%�@Y�#g��h.��8S�6��&��I�s��v��l��Ym�����-u淐���������y���H�6[Nc8��!]�2N�a��"3K�C����fqyu}��a��pPl/��!�t�772���;��x4Lǀy�v�+���02QRe�J��WX�a/whm+}�Z�&��(�iR��6����D��^��{� ��3l����W��s��{K��"�h5�\[�쉜V�e\�j��HC�&�F|��*$�b�r2��c�`����+[��ǲ�֟�@��z���`�M��D���/޼yc��&�X�^IO,?k)v-�%M:.�8m>��L�d�K�;�
�;����c����_�'�;���d˽Em������N^���H�)����x���$�`а�X���δJ)��U&S��J�s
�ԵJ0�b��]��%�`�SȼK�:�������A��LaV3��G}t�p
MT��0���:��{~�~U��Q�f�����#:�8��u����`sz���SȩD��5���J���e|����mD�v��L�=zؠ���J�d�R<��� ᨖJ����6����W"	�uSrD��	T�<��t/�y���'?�Ƀ�s�I�?IT����?�_D3�#f^�������w����c��T�8(�����܎|�0OTY����U�s��^���d��@9���h]�c�lux,/�^ �ԷN��R�?'��.
 a?�cn*�6�p(r��m-p+�.��T��lg(H ���w���Cp��
�o��/�|N�c:)���x��|������g2v���3�BGk�+�E#��!7KF�q�5�O3�g2FG�>��O�.�PmP�1�N0���g|m�.�^�\ǿ�1��F���R��^I9�\�&��z��1�X"y���p*�r��nV��-�� s�9n�D�?�s}*�7��	@.����>@��}����$���	4(���
��P(!r; * %YU��jR@���Ar�$�� :�^���|�(~�4� ��`�t .5�%�:�7�Ij��3�Q��0y:�v����Ŝh΃L*^�rƩ
���P65K�xn$ ��`��������VS��f��M�UI�s�C-i����;����t�vH3�H|ڃ��f��lD�o��N�>��豏N�/��#]m_z9�L�,�E�:8��po�2h6�bQk�š�T8L�2ioz��>G����N��ئ�n�'�w�D��P�v�_$J���,S�#�d��d#��5����{�?O�2�5{���&w@-n��X	��r@'�q�� }����lԛR�`��jZ(���#��^;�$��B�d��8?�U`��uG�?َW�x�{�2z�\��z(��T�@aT���8j�W�mp���Rt�?���"-�נ;���F��	*��.�~��L�P�s�;������&���:k��_����V@�g�vr�[1^]]	�nM6�L����@�B����_�:�`�{�o/q���T*	�9+ғ�)�k�F�U���~OH/@dvqZ��o�~���_}��f~�����Ch�$"��ܿ�L3��߄��5:}��V��u
E�\�K�.&��.�(�O(��-:��E��S^L�khY0s��t�;��1x9�D2^�vD<7��+>N"����p���&9K���؋˕[�V���d6�R�-|�����?��!����̔��2/���v�A(�����0�W�?~	�o�^�sQA��C��?��J�%�,L����H��aצB�7���%5./0���%6�kc/�L����NHZ�I�(µ(ö���-N� } ��qx�+���
� w�еW��A����|�Zh�Srr�E5�/���<���	-�(�Y1�[�2o�|/�<�Ǭ�&���8F��AmbQ�F��v�X�L�@�G�[S�cH:ʹ���ڧ�_��HG��,̷]���mK�T;���"e���P��E@�|@�����?�0�t�.��ǅQ�/��J����
�"��D��,.���6����rJx���tl��ۍ�1�]��Ŷk�׍~�x�H��� �I�r�4p+D"��9�s|���Yy%����������r���t�<'�Rm[�Iδ7�Nf�;�&�A�2��	�L��Aٛ��Ƈ�a�&�xMյJ�cq#��up���	4:5�.�B�`���#2��B�h�XV�|42�I1�哖��3�"S��yI�IV�*P:))aq�
��D�m������|���π�!�ߚWm*>�2�e�.K ��X���cr2�[G)�͆�Y���)����9Sm�҂z��B���9C^�3�p�p����^���ǌ}�:E����-Q���vB���>�dLtԋ�!t�2*������.���@�m�Dvkh��G�ڔvR��$�r(��X
BSp��ӎ �
DL���"r����2Sg�0EA"��j�l���r��� ?2�L��Ž,�6bE�*P�#�`���ڐ_KB1J\��%����f��M��B�°�ܘ0�lGKo�	�OֶCo�紕�6]�r�藆U�����Qgn���6�+fʺɴ4�V�si�(�͢�h�z=_���X����#�=�i���r<S7�hS���.ܟĐ�\X�3�fԪC�>&Y�����M��CT�H�����&�*b�b�����i� W0��K!t1�������Sfw�:��eH�<�/`偯C��� ����	vT�Eŉ�Ks!z���r���[	7����B8�i����v��$�V�dЛ�����G�/y�������."��#4ОkA^l'S�Jr\���lV�!m��E�vE�̗r�΂)�PzZ���32��~��g���6�J�G�:��%�T����Pr80�`�:-+L�ha[��4�$jR�P��J�D넪7t���
:�t���F�{{8�&��t3H"�޶6m��L�<C�����RG%�],���5�4��f4
�~�[2���>}��}�o.�����9���[z��Ŝ��4����p�&�*����� c
"6�7��v�����[dgк&G�sXRZ� t/�'�Oc��0): ��Ja�GH����5���G��b
CF(�l�	���t�A�t��sL9D�G�eR��Ov%x����5ޏʟ�U,?b�2��i���}����[KN�7f� ������[|#�0������+dcS6�  p6��'4$N=�'�9B ����5����3ǁ�r �3�"ps1�Q�4$�@���P�����
�Z=x�#���j�Z�%N�Sp��jJ�(�7��{�w}}�2*�y�m_�!(��(-�<a���� I5���h/hq�(+7�2hܹpäb鸇��ȏ�1�!o���|`�*z-�s�*J�3sê��7[�%���O9VP��R�1y9�T�`Y`�U����#���#P�I�=��~���|B��ŋ�~�-����2B�e�m3�9I��`2�W�(�se�F��\	��Jds��5-JA/�j�m��_���w�a�;���ѣG�Б<WʤCK���	�Q��U��2��� �36*��7�SSo0����*�-.�Y�+�$�@�����iL�Ԍ-�@�(zY���5����������/�����:K]ͭ��z>��Rk�2P=���"B��1m�r���_�聖)��q��&x���&/E��L8������!\�����j��e�oҫ]8�����0�S�P��N�6Y�@d.�R��_�M��g��S�� gW�If���O�F����l����$$����dk�������`������?|!{A��O����Q����)�J���?7[l��ؓ���W���^rm����'2e2WJ"\bc��B�^�����t��r��k�����J"���F"f���A_�K8M��Q
a�UO�l�<l�t�n���Bg�
p�tߠcI�s<M$����K�����l�M�$�U�����>b����Cii��E�ǭݬ7w����9��VZS�9f�lT�F��B�tL��sSG�G����*��I���LKp�V��(��D�q�[�g׋�^�[�Ri�F!c5�,P`<;t#ڡ`n�dGze�4����v��J4[����iלp������S�N��'�4��g�`j�<�M2�$�0���Dn�Kp4!w�9�l�b}v�'�"����N	F�)|��k\���漘��	�ѭܿB*��#��'�&���QI�s% �۽���ek<�Wm�\�6��;��b#�;»�9�lĥ�5ڇְ�:A|���	:l�B߰�^E�*L����ܨOua��3���+X�s���<�'�H�Wݗ۟�0�����+�t��oo�fy�G�<�v�c�r�7V�@j]��/����N��ho�+j6��)P��IаpCa�sᏰ;4%9tZ����i�RE��A;XF�E�矞��4��D&شO�>�[����xf�$ËA��8���0�N������ٯ*��}J���3����t��h��"A�L&���7eN�0c_(6k��r"i�5w{��!�m2QD�=`2�G��96-���mm��s>$��N�A{���_]����!{M��>���$A�k93��M
ݹ��n�R2���h�`��<�h�^���UI�c>:7rf���JEԵ::S�A��jPy�0 ^K����
`�
Ɓ� �Z�LT�&���v�|���#�]__���+��on��rx�<�n�#G���Q�4��};�cu�Fh�蓑�M�q0c�΍�q�����{n4%���������e��9�����Nr+�L��>�r2�(qcZ�K��s_��D�5�QO9������F2\�"�8*4�D�իW�@� E��(ቄu��H����ȅ��HMF��s�����anxa_��7�.�����AO�;鮐�D�;���-�C��̵o/�}Ƅ�����W����P����g!�;7���s�p���
��f��Mv=�Z\I�_ �i���q0	2�O�-��XX.=�}K��҃�8E���Hc�z�))��$��} s�I��R����i &zky"�%ыn�����:�<;�`�f�Cj��F�tp����!�N2�wt�t��t�a�NB�JF��J[C��=���llw��,L���Ё�q�� ��Ag��#�lF�!5L��y8-��[$��O� �%=�c��T_&%�'`M�d�<������n����m�s|�bM^��w�1~�ʫ�^�������)���U�r8N�|����|,�����3��CJ���7��j��b.�$�J���Җ�ƥ�)�Ff,~Ԋ��6��a��錙�0�*a��b" aT��;ܦQW	9���N{+D����q��|eY~������"M���'F�.�qT�#u�)}!P�΄�w��Í�p��w16�L�!��1!���I�P��R�աq����f��:�Z�s1
�*;�e�(S�?~�"Ú��)@��@WI%#��͊Z�	�`"�M�lֿ�֟��ѣG�s����� $*�����=i셋یh��3lJ�[��ڎdŊ%�R���Je��/5�-'z��_���r`��H\��B�Qb�"��M[ru��a�=u���Td��$���0�Nr�䜃��I)c蚭)�[����?����>b��Պ��y.�O,� x/1Q"m�ߐf���kz�o�[�l$>!��\��و��n��>s� W�e.Ei��\��VB�	���XЛ� �U�
~�K�Rܿ+ !QEJ�Gy7�K#j�v:#uR��� ��y`���XFF,2��.����ѽè �Œ�Q�H6��&���G����ӟ�����;�t �3����R��q�e���6-gΤ�A��Aያ���+sX+�l4L�r��5Z�J���פ
`8H�H�,y��,=B!���ܩWWwggǿ��/pe8�Oɰk��~����|s%�����,h�~�t��W �Չ3e��Q��6a
N��k�XX�A�ҋS��
�g\��s���8���4�0 �+�?kǀ�,����D���#��������~�	������q�L�J��
rYIA��+�+�Ҧz/r���yE�-jo)�v�+�u�r���*�@ܼ���4�Jd����"Ia�5�tj��Le	{E�Y��J�n��pʗ2$�Р�ōB�]��+�b�����e�R�m��s|5����a���-E�`������s������r'�������r�d^<x0�=fZ��/_���i0�L6�V<C&�S���m+� a�{[Sp{(���B<Y��wF]�9�[Y�~�jxd��#!��
��M�Y�]��8�t�s7��M�ǟ�K:"9��=�G���ӭ�Lr؛�W3���rh����otn��A�ɑTq/m�!��BDW}��s�f��0�U������*�^]<�fn�甔獔>S�6���"�t�oS1��b�8:���(\w
��3��b���ކ�"��k� ����LP��q2h���ua��e�-�1�)b�nŜ���Iː@����W�g��[��uyX�M�^�:I{�x�H;�\��.<��-�G������C'��ã��'�tD=֧Ic�vI�R�j���$�a����2�n�f:���M��@f��Д��a�H��Ȣ���K����-���&���H3;d����R���٤1��S0�3p��WK��(�jl#�j����k��\����0i'c�w��Y�dd�Q�
�\I�:��/�a|����a-$&�P�Q��Ēď����a�y!/�LL��#�u�>��{{����Y�{�R�3�>�dOں��5����)"�<��(�\Ԡ��G`��5]g��#�K�Zzh|�[z}��cã��\�A�m��RJO�k@R���Uɮv�d0��/����]��Y{�I�h��&��b�� �2���u�`s�+�Nk�� z���DP ~��i�q�|&��n�Ia3�g�	j�HV6�Ȁ+H���Tp�(��cc�=���I��;��N���F�*vS/���G�5�g��W��g³^*w~ԩY��0H��U#=���5i��h:���K�H"U������ҿs��:Ō��S*r�p$ĺ�w��)�����z:�9��҉��PV*u������g�$f�{!S�"����Z2�i��-`S ���?Ć^\<DK8I���10\������"��5���6�b�Z�@�ҋ�T%	>t$��Hr�1XR��8�W3��Sh�����d�_|ǡf��u�V���א��Еy�D��2��p��Nx�p��F�4����c7�d�5D�8�N��&��{��Z�	���i��AIN��)�d��̿�>���k$vi馀d���ջp(�(��°o����Hy��5���ED�����T�ATe�m�e�p�L�Z!y����M��Zja)nn�H�O'�H%]�!bאyy������O?����;�����8�X�M4�O� ۓȝ��`��n���!���8�"�%Y���y9�u�B Ə:��6Cg�Kt�.B�E�"q�4dno2C��,��P^
�/%�cI�tm\�B�v������|��)�'Et�Ϗϡ���p^8p�|�i���="<^Z�s�zqy�Y�^d�����HN[�����a2��l082V�������h��}���S�o���1��.�r�H�9۰�85���luׯ�0���A��#:���� �C6�K��`ȖK8o�'�/a�rh*��a�HB�'�,�5�O���w!��'OY!����_�}���߿�~r$6�1��51�NؓHsJ��������������ӏ��?�CN�n�`o��@M���J��E��ﾣ�B_D�K��\��.hMH�@Z4�+1�"n�$����%a��f+R(��"{Kkr}yIo��^q���L�#q�r��>��i��'/�	=���៮���������g?�OKQ�X�( �`�C���r��h��<*��E�{���\;��� ~�����	�pq���SdJ����k>;E���#��|��(N.TraȽ��D�:=>]��¯~�������b�U�=:QG�[�^���S��#���"��Mx��iuְ�Ғ���G��QB���6$�ik�M>@�J�J�4���E'g�1�Ӥ��l��]��޶E�B��0����������f��C�xx�&��/��Q�`a~C�"�]~���Ȉ3%��Q�6n�+�g%���.� q�Q
2�( Nu��P�i��㙇Y��n���Êh���GS:J/Z�|������2�S�<`� j�dC[�f�|vp����_>���f��
����Lʍ8� ���ZG揶�Ei�����)̌��'S)(P��`G�n�m���Y
L��K�3y������?3)Ixؓ�'�>�0f3�eT^*q�6(j�j����[s��u�\����"��L;fv�ܻ�ql�ߥ�3��N�ۥ0|E�Q�*m��J�Ʃ�i���B��:�/T���u�Ǹ�ߎ�q �߁H�H!*$d���bD�����C!3�� ��d��s
��W�O�#~4�m��i`&�*pLѦ����)+Dh�O{��;n��w?b����I�t���m�|�O!�`�b�c������H�PB��y�B���n�%R����k|��=0��!� ]^���^_-�N��o��wm�k�Ł0�5d��jἦ~ ���3�O� �����K
�F+��=	�Z��\�,I����E�8;�aT0I�8˝VEPO� �@2�(	_@fRD��\T���Imޤ�d8�݈�!�e��4��
��[��z����6��
�״u'w��E[Go�Щ>�Gq=z[�b�)_�8W2o�׷o�ҧ�߮��7����p�(0O\�Q
d����i��q�g���n�f�i�J����I�V;�#�r�������X�y& j�wDH�)�@�-��v�(�0jx�Z%3�i� �x_��y:8�{h1��/H�,n7<���mZ�ex%�J"X�
�f�P3h�a/�BXp��6h�k"�7A�#��PJ�:�����K�y�-W����O���	_dcS_U&~���F �z�
Q�ݸ%����Jd'���<L�T}�,m'�/^� ��K��)p�
����D,�*4� �zH�ƨӱ��hM5�Jo �T��:$�t�t��|Z4�H�'�hd�ץr�"�D60Ϲ'�M�q��! �Y��ȧ�v6���.� pꑛ ]�\r[1�2����fw$�iD���꬧:=���W_��:���'ۊ�2��g�<c�C��ǉ��L�FҤUZ7Q�yļ�3a�!/�G7��Y��dPS$��u�q� �Q�nSo�6�D�t�R�ņ����_ OAϵ�0�;)b�=8�#:w��-���T�ƍX�E�G�VᑱSc���$��wN��F�n����t?��t��~�����9�~�-�&a�E3{lP�s�SHa�}�L:��t� �¡RZp�m�ۙr[�3Ϯ͔����9ZG�<����X2(�Z*���naJhG.ΏOۘaA(���{��	�>����;��Ĕ��N�H^X4�Ak����;��r�0���t�?W�,���U��Y�Lt�t��'M?O�
^0t�l}2:�
�k^z�����40�c�y
�(���V��͊m%KR�S�T)D�2����B�m�'�0N16��
[�(�g��	r�犊-�y��C+�"������۫ݐ��Nc\�j�� ˔���Ǐ�=�4�8� �A�;62�
�^14���>�?�QǢׁ����a�ΰV�A���c���`#P"���Zټrz'�V�?�������煮�ݓ�3a/�y��)���=$!�������O>�ۿ�[��<?���H��[�/��A壘� !�,����\"r�D�u��Mb_���,QSt5q���-���z���W_M+�����"���&��_7��߭����iP��&V�P��Xm8� Ŏ�.H�����	5�9I]H�M�Zd�#�UB>�iu���n3��'�u���XN�9tl�V�uJMÊ�0���'�8�js1�����3��;�nˠ�)�؆����O��д�@� �#Q+ͥ�Gm@.��t���-T��6�pW/"�Z�*��'���ɶt����h���1�x���3�G�����'t�<�D�H�r�\.�b��e�&:�l}$Q�F�) S|�����JZ�=���Ç���� �� 4ասWg�����NxE��xg�E��~� �"���q#�r��C�����8b���'W����!�X{(��+���I,wJ�4m���N|ӽ���@�&:��Ъ��3+��S�t��pUe�0�dv9��H�"�x�|����W����2���IY,�5�lXh6��(-W2�����дLGDg~�O�5�o������'��i�3�Ȣ����ޠ#2������~ԯo{,0�n�o�ݿW���e�s�l�-��N�HE�{��W�ʉ��Lf��"�'�Jf�t�y�&N_�6£�UY��4�h���5؏���1@9�d����	�ߏ�d�۹��fp�"m�d:�&��fi�g�h������	�?jQl��]n/�S\�mYB&%^��e�Gc���D&� �H���Dt#v-��<p�	�e��'�m�ă��� �؅B؈��R9�h��>��HL��J-9؈\P��1M��_Wi.�s�١p��ى�x�c{<^�s�le� <;p��������D�3��
B�Ʉ�K� �;�G�Rҧl�( ����x��c�aY��l�+�xs����e���
ΧՃ��F�@�)�@�\ƕ�ȗ�[g>:~.FTzN�� �-���v�Ȍ��B���J�e\���[�w�_��e�-�2��%:?���`�ظ�b������}��a2�g!Q�rK�
y��A��`�j ��y���y����-|_z3���v���ķ#�$��BB+|���{�=zDo~��%�:�1)�U���
hK��;�+K�`&C�����kG"	Y6E�pbh�Zhu7��e�y�#P���_`2 ��Z�f.;$�$8�?�� @f:
�?\rp����s?TH���X(��_�Q��K��H�O#R$@��F0Dy�!Kbn�J���n%�0![U!�~%:�n�I��l.�`��-��=��0ň韯STM�[ p� �+ӠO�UyN1̤��������!�"�Cfǃ�e�s'�Uڬ/^l7z�����#�Av8��N�� �HN~��Iv�Y�)i�A���$�� �PI�F'tɴt{sK�ؒ:;������CfW�<��^ja������(r���'e�5�7-��=�5�$D���+nӛ��i����)��3��A ｅLf/�0m�G�J�5�91��8�	�ݤ��Pne�2�����N7�ƽ���{�}a�;:������`2aEq�ޑ�R��X$o�VzRe�p�iQ�j�XI��_}���2Lx�y.�=��_a-Ȑxe�IG<3�x��䧻�J�Z�S�h�i����x�ub3�&�����3��^8+�Aߐ��Ԓj>�����G|���s�JWE.�>s�9E2F�"-�\^�`��<J�J�E�+$d�����iڴ#�XBS>�S�A����j}+~>�X��0\-2��zWH�H�ôM�ړ'O賟~�_��m��26mM*p�+cG����%���K�{5[vYcU�{�ms��4�� C�$�c^�?�7/�2� ��c�4C a�h����M�2sU��~�G� :n�>g����Ү\�ʍ��֟n ���+���f��%]H��Uj!Z��|]�\ϗ�t4G?7���<���a?7z��[��J��2���G�o�jcD+�CA0��|��P�
:d��9��5�r~�4|�O�K<<>v�<D�o`e���X1��A:��,��)�u�n��T;��f�*����5 [ 3,�,��0���>:A�#�I7O������;w��1�u�!�~���B����~��_��-3�w<�kB���J��F���9	pp{x���{��'�b*�Z�� �/�sAK8�/���m�k�g���{R���Y����7���Zv](a뙭�D[%S�L�ͪ����K��j	�*.A�:���*6[�Q�n�����[lq0��A��1L�T2ĵS���$���A�YA9�H;���bkaqE�w1��ܛ�Hc�ݳ[�W��a�s�� [�z�)븆/�+�4�*m1E=�'�����2i �F��p�,�fhk������0�'����-�<Kʕ[4SlJ�$�Xۨm����#�C�Hw�)�T�ԨH��u�bB�(/>��­幐@ϋR(��W.c��MD[q��-�F278P�v����������������Gӌa4L��n��z����M}}s�,�M-�����<�ZZF��<�(sǀ� �PxB%���K�٩1��G^��N/�Mޮ�v�\�n)�,3�6��i[�B�F~�]��!ݦz�6�7  s}-�a�M?V�ǉ������V�^�7W��%!�J��3涾�Y���޽}K�������蘔������Lj��;
h�#�m��:�w��4�A"�1zG����L\�x)�1Gh�|�� r;.˒��)�Z�di1��r�Z-
rA޼yC��!�.�ZRk������d{D6��s��XG��D��`����yr���W����6U���+$
e�v
��:�~��S�{ȕ����,!�~,&q����[�.�z�u���}�$U��RI��wF�g��υ\��YכK�Հ�b��VY����\aP(�z<wZ�O"��A��^K`�Vi�U�sC!�PQ�X��my��@�)�����K�y�D*4me��)a���͜�y��R�m3+���I�[aFAƲ�����;���VJ�*3�p�>(k�&�t2���V�5��Br+��j�D�q���J�U)�N� Hg|�`��I�C#�n�L
�q�r��������\\V!�K`�<�1]�ф��TQO���Þ�*�Ю�q���� 2�{�:܅#/���f@��2xWN?ǵV�aq0N�;�� 5 O �v@�!�f;�N+f�r4�9Ak-��:���1�a��sC�h��K�I��������Ҫ�&d�߇�2��p�ԛZ��7�Ac�о�˹8S��ι���~ �i��a���5SP�U5l�E7����ĿzY����Qs���i�H���	&#��%3�����Q�{x��̐'"G���hgo�իW''�-S8%I���I��r���?�����$~H�vi�]�J�O��y��������v'�wR���JĹ��aMA�9 �9��|1O\�#�aMd��޽K~?�w�N�)��V x�y�P�bŋ�z3�B���Ν;�$ f��byA�h�29D��@{CC����5y�B�=���d�����#��O?����W_}���;�PH.w�^iJ�9bC!�"]�8�������R���w��FW����p�4�O��#%a���T�"��t/Ws �8�!���%b$����r�x||<�q�-:�^����\�H� �e.��QK�����4������nЦW��JV8 �$~:� @J�^��w�{���ƣJ�%�'/б�+�^��<~���{g���>��٧$��U���_��+�a��P��Pf�N	;|�J�BZ����9H3�G� 	PSN:���b*��5��v��&D�&��Тa��H��U�\^ДA_�I��6�s��� Z�s��r ƕƜ����1���AH��O��Ve�k,���i�K-��[B�dU(>X��6���?����=۠�߶��7��D�U�|�d�Y�c��1D�t�ph�<yBEۊ^���@��.tm44$�5���_sPX����O���8�̐��u�Ϻ����g��שnA7�����@9H��3� ���\�
#��$�����;�ȃr,�P(qM���m�F?��8v-�i���7H�)��vZŇi�{Q�R��k��)����ѥ	�"���� ����*�C����#��KerkjYH�gn��@x�s�:˽їJ�2e%�:2�ʄ���V��R�� ���%�×�'%��{T�tLBٮ���B�s'�A��(.%���~��wò"�!sI������,�){t}��/�˧O���wkk�<\)����b���!���4�5=��:i
�uö�m����g�������-/�g����&�90��X����zR!�I3s�
�h�2iP M�6T�|)��H�^�_�X,��4�$(1<8!�d f��Ǻ��k���/M�A�:0��uǣȚ)�>�i��q& G&N-[������ ��G3򰰪��*�r�5Q�_��8t��NNη�'� � o�S���?�A�:��[�������[�7�<�&N��eL�2�u�
B6$�1e(�~|#�#Ȫ�^
g�1 �)\� H�$�ٲ�����!JR8v�E���[�ȝ;?�xۇ���@I���y�6~��%6�3�SX����8fdߡ)��f~��� �Y��	pp*�����5�ݠ$sF^}(�i�<�	m��4��#� ;%��8(eT,!5hѥ9�A���,3���>mT+ ���F�s����I���z�o��v>M����J��UR�CQ�<ysx�y.�PZ[��y�7	����j88���k�9R�W<3 �:r��i'}����ʆH��	��0�<�י��$���l��"�纂�J��p�w�Z,j���Z,����2O��D;�Yd���lM����/��ϔc?Cg��E�i&��EW���<+6G&���9f:$y֙�f�aAq�pxҍg����\.���l���������N�ojN��aDQ+CL嵬�A��I�+���Fʖ2�J��5��4j-��Hv�8�i�7�yk���[E�W~2��16m�4ϳӀ��Ւb O��l]��^!��6¼����U�rh.g��n��y#3��.x:�P�1���7��xT���eɃT�,V�9�)+�:�5��КYV�EE��P����&��0����<�e�d�P���\�M��ޙ�违�-&]	Qv!"�}��?�ʉ7������ H�O�oל6z�n�[����,"oޠ�a���M��&�t�����ᰲCZ� �\���>�Dp��A��MRl%�FIA,>��3t��>�*� L�Ӫ��t��`�	k&♞�*�m����Ld>�ڐ��Lb��y{ɝ&���CR����Ң��%fYgJҽ��ȳL��Ƞc��f���{�L��ge��w��4�,�٤Z3A����M�q��0`�Gp����<g=���t�ȟ�Q�E�#I��Z�81u3���0����SL�j�.1���9��D�Z,t��0\!J#/|�Fyv���t�t����	I���C
�)`g<�:��'�����)��H�΋�d ��\�<H%��7=f����(|�R��L��Yntwo񛤩yq谷:-K�+�:q�.�^k9�	M�c�4n/(B���?�;;b)R�}���DW�-F7�hx�b�l0�B���2�D�6k6�棻�g�p��Fc�2B!�o��&�7��8�'��7xl'�g]˞���i��`p��D�p]���BC$�K:�	�i!�'��~԰w�P�m�8�| ���ȡ��Kq�������\��n~{yzL��F}TW#j��9�ڣ��^_��v{zrQ�?�v����?���G�w�ٿ�񇗿�����7�g7d�� "��B��m�-�TRSտw��p�3_�^�c�:Ė�"��H�aCj��JJPe�j��iIT�AF1��ziM>�����1� �^���U>}yJ�Nxz���wt� ����,�&��/�Z�Z���$�6�)�D�mt�����k�d�+���/2eć��}�{���>�u3��eg�$���YrX���M�������8��G�[��ۙL� ^OF��$+xM�TB�0��i��i���\K���amS��E!�\�ӟ�={vttT���-J�Kr�A$G��1䇳�5����vN������Ǭ�×/_"ѿX�)�.�f��/(����#��'�:��C������;~w�ߒ7����,�t��Y����8���P���R���'�K
�����Pbf˘�5�v(XO�p�!���WTL�U�[�l�}�Q�Ɲ��A����Y��v�D�<S��\�f�(�/�+��5�B�m�q�����WcW�V����_~������_�A`�@j�����ޡ�K;;�Ғ8�Eoˀ��A�F�S+��r���:Š*�8e-���6���2�?��k�aL��$Y�2x@�o@��z��?�p��$�-�������'�]�|0:��_�&�Io�vә-�ā��,{8��!%-�Ç)���@�kH������B�ȉ��a25�S�_fJ�E�&�����(3��5�G��%P�#D֖��iS̼fM�U���9�� i��t,BN����2��O��ْ�a8�jK?���:�Af�%�%�G�S�):�1�բL��+f�D����	��n��j��/�/���|�Z,�-�*����X
��ׁ�l�<�S�exfW�@fݴ�T��J��pG�F" [�5^��f dW3-�n<��fvpJgk���X��J
�Z.� N��Zd�C���:my�B�,����W?�tm>��{��f��������)��UdcH�&t�Y�ഝ�Ȋ��!�����G�s�k�/���'^E���ox�f�_ �jhͥ.;.���D�������K;;Ӫpw����$9��#1����X�c��9oQ���~�%��A��-��+9f��M��(	�.%W<Of�+�W�_���޼����Զ��$g�����+I���fe%$�1��w�ϯ����K�p(��y��d�!�8ŀ#0����ڄ!Ϣ`�����`�@.�Jf�ճYKjG`F�梅����0�H�iZn���!�?��u��5��M"di��3�bQ�Ɩ�"�~`��\���Z%�������-�嵷�i������8۞�l��{]K��SŰ��rf��C^�N^�=¯��7׼7S8�����
�7 �t����S,��\�-t�Y|lh��Tm}�&]��4Q
*�k�TB\~. 䴒�հ���X:�a��&����C�	��-���Eԑ��Ulᗰ�s�
�8��ؐ>���e�gǘ6��۷�;���3w~~N����#1��
VS�a�̿!OW�tIBHd�N\��]"��+a�l&�9�,���7�̈́�Z��B���f�6.N�6򳸇N�2�/&������9J&� ��(���!�����P^ҵ��CE�#<�kU����^�d�4�E����B�0rn�u�<�]g��@�Ͳk?z��p*!����R�{-��������\���`�f{I��С Hw��*=
�G�9���-�"X;KA�oV2 ��M���WH���ʐ��fa��S<__�q�l�M���_��SHx�uf�#���B��������(,K�Ss�pM�b�s֣�@���<G�b��Ne��>(��I�5�
\4d倘��-h)�U�<�� �\�zCf�� ;��\�w�{T�+e����S+:��@Q�R�2�����+���Q'<����C��N0b����G�E�~+Ȭ=�� R��,���9��J��xKv��^��n�P,�F,UC��:��B�]�gm!�iiCҶik�=B��?DؠU��8hcD1	����CS��/9��x
s ��(^5ɉ� �<q`�}q60�>*1h0�3}=�������_��l7�ӵ8�S��&���SH4��,-5�o��Xa�����l$1&=��P� &cC�U�y���8^W�*آ���������������f�T=<z���)�����G2|�]��
�=��MC�j�Y^�#"[�|V�R��Գ_�yp���7��F���xX��^5ĥ@$G�L�-�G,ϾA.ⱕ[��OnX�#k:�		���+�X@ظ�=/�k��Y�'��F-]���J5h���X3(��w�}��!}I#3��REA?anP�t�D�Gc��I5�G�БT��!��KV�r^7�J+R��VH1�.�)^�`�L��!��H����c�0��V)6Q�t:�E�rY�3'�e�oSsttD>��/���n ���@ �!��z�D�Į��\���o�=��u&2Qi����i�?ln���Q�l�|�9A�:�jff
s�Y��Hb��?�t�F����&�s�|�� �J��#�(Ǵ5q[�Ph�l�U�*��QagТ�N૤'Q�/d2;$�*t�2�T���o�|�n`6����D�	�=�=)��?��n�����j��ǃ����Z��~�$((���v�ǉ=??� ��+���P�PF0[�B	|�6j·��o���.m��Q���P }�e�����_z�6a/pA�����_�����F����/��_���тn�q��l`²d�� ��_���D��iQ���v����TzV�+�'%��zB1"�CY��>^(G`�ti��|ͮ<d�'Z1����t'��V#�� )q�8�'S(�5:qs�����Ցk?D����BA9-��F���@6������#�q'v��
l�s�π;ـ����Iu�CN�t�H�+��[ �1Kѽ)����Tl�W�:z�ŋ\�=ؖ
<V29���N@j��=�ڪ"E�1�T�W���7Ag��Y+)��iw�L�����$�]���~��ÝG��(�k���j<������W:mUt���=��z�φ�#��c����3�!2eׇ,�H�XH��r���|��m�}ol�r/Y����0�;���m�oѪ�˗/��{����4=��&���]"��B��$1�-�Z�*��*C��"j"�-ƅ�d�QK��g���µ���U~TV��@:�X��oː��&��ݼ�y�dOO(*ɦ �Y��;Ǥ�̹tbk�̂O�K}ͳj�nSM�wÈ:" ������As̞��|�5 �J�5��G��p�
s��^��?���W˕9���e5ԙ�˴��f�p���hSd�;F-P�i�=c��Lx����������ZF��Yh����uҥ�Z�G`v�<�ԓv�_I��\��u \r�Z7>�ɭT���������0�)`����n�R�e���N��um�u��|�"����J�ui����`_KΘ���O(eY`/V+�Oy���Q�S�c���~eB痡!Q��	��ԺS9�͊�9��Lq�����	��K'�r5��bVy�CP��S�C���T6����
���Y�0�7�SA����"��nC$�X��� k��63�v�!��z��v�nς��D���7���us��^x`�~
M���K��rX;xW������G"�Sˡ ��G��Ē6S����x=������Ş����^.h�*�F0�~���zU� VS5N��)
�v��N��	���	9�q5l_�+rV��~zK����ڴg�2S�NØ	�k�	�������իW8P�1	��k�$�ba���a	�N�t��p|FyN!��J����	�g���N�cF�
�����mrN�03t7�N+Y����q`�PǪ�E,� � ��`�� ȴ~'�{�)svM�-�+
-�m´Dځ;w����~�g��><�Ǭ��z���H��+��A@�=~�H����.HE�2�t�t��:�=d���ϋ'��3�k�D���tKp=�����rOŬ�,KL�%J+֑0�χ{��p��й��]^p�q"p2�y)d8�"Q��>��Q'��L��c���9����h�B��5Q��`U9I6}��O`�Zj�ѲlׄzC�Ir�si���v~{}#&����l5_у�)i����bw����dZz��}}鄓JYqr~��D�������E+轲 �h�`�,���5�>ᾑ��uP�Ç����n�L��[�!����-mrΤg�Y'�yU�!��֍G��d������9g��{��h�!�`�gA�G�7����9f�����-�jYZRf���jy�F��{R���^��$��m�T�p��_�~]I$�}��l{suus}}땞Ϩ{-�!��Yې��:�OډF��Nɞk���fD���Y�.x@(L��X(a�@�ŋo?��R�P�,�m������6@��Vt��<d�~˹�����y�>���G2v)�1�0�	��M5��N�U
J�F��؟lb�2*�?5�����b�I�����U6l�5���h���z� :��H�	 �}r1 ����Ӭ!�HvX
$p� �&������V�DC
��[;�|� <	D�m�������g2< �M�y���HeJ,�l��3���dR��E�_)�3įԹdA����4"�6��G?���"o��>}���=�v
��u(�|T�e�aqAX���)�Bhk1����R_8��8�6��su!�������q�+˄E��
�?�@˃�b�_/�Qd`nC�I�_��������ք�.�~�`dd�H�����1gI�� +��hS_���j=�w��3��������������[�CRrL.��!�$>�n.z�땫����2g�S�;��.�^�o�I(
Ds����-#�EN+��'�l�Uu{���ӁbI֋���ڮ��}9��xw|z||$�w��cm�q���s4��D�jF�v���'��� e-�B�c����$����Bl8��Y�y�h��]뼑R�>���:DF��pY{�R^��I٢��=b�sV���4��0��峪�Nr��������	)���K�/�̪����J��a;�73�"���(	�L���ղ��30���e���^��������F,(�l���x��&�QƼ~Y���dD��Ev-8b\�RR���|�����{[ۣ��B���)��6�Do���m���)�j!h�)�����)����-]�?GízM>ޜn���m�z�&��T�i�r,A�0���"ٖ�[�p���h4\/W9G(!�<�.1���)��g�-p��5����A1X5�x�7�u�,˱���~��#�q�+v�B#������D�
����o���_A:]�F��nyo$n��%�:*�[���"�6��i���l�^��+_�l��]7Q0Ǯ�V������rs÷��ņ��i���<X�1���NQ���������׮��F9�i�o�Ix0@O�����,��f����� ;V:��D�8v07�+��B��9,x?��5��'EmY�ڵ"��;!�dyI��u�,�Ǌ;2P^VU�+E��o�t�
<L.�C�/��AYj"֑]$��F��ߺ�+QX_j���VS4����VV � ���)EJ�K+�"Lu�P���(Lk���!�?�.���A!��G;#z�S~_d&��v�6�+mvYE�������*��J��X�"G�����Nk{G2W,8%0�����`G�ԙ����f�;9t����W/7!���T��[��&���������B+idq�'!�.oC�Ad�����v<��ѱi����W�X��M��l`J9ɤ���\{X�	y�RC�0c��G*�����H�X�N=�F2�g�=`��wP�G�FzE�˥RYU�ӢZ3��~zL��o�0:�ݻ�(�@���hY丁4��X�A��T2���~T&�ɢ���KW�(�|!8{:<N]7F�b�ccOC�����M	�;w����<���Z�vr�)�EH�
����P0�=�M�ZnS۲��N��^�+�#��#� �<Ţ�Μ�t"�y�A�d�&3Ep�V/S��)��Q��`1�gP�i�=����!j���~�( "�d9,&3�P����E7҉C��'/�v���ԅ�����x��t�?��C'hD�
�V	��{��a�2󈉖p����8��3y!7���z��+I�����Er���SJ�?�����;���k(�����&Me���:3�ݻw�l&��Ӏ��hP&�[9M�C�g"E��h�T���(�*�S�#!��j�À�~�!�h+�c��e�C
oj�SDR�k��4O�g:� #�h2e\� �#a��pj�hz������#��GC�����q��mrF����6F���� 돉%F�\�7�DhLZ��=oRn� Y��=�k��l�k6:Q�\[3Ǭ�G$�	�m����p�D�%,�]��tt[�&�=B���h����\�c���9����P)r4��  ��IDATҙ-2����<�q�Pj@TH:M���f�м�5�S��X[:P}�D�pu]Ϙ� E����lŻ�ǈ5DKl���Q��T�x�
�n�PG�1����v*���!�o���s�$Acv:�g�%�k?��������^m�R�L�+3�g:�����[1�u
���c�lf�'��E86��G�{c ���3g ��X�)�Gs	L�)EcmJ)*�pQ��}��8'�� A��0��������Q_g����L;���Bkg'�[�q	FE�$(i`���9<��{�.s� 6� ��8j���Q��T�#k�X:��p��LB�(�EH��1$P0����i���5�&�P��?��?�[>��3�x^8ġ+��f �t]K1Ju�[�ۢ��@Xv��9ܞu݀R��z��M�[(
<�K�^C�O �`�[�=#�����'���_�5]�t�;�O�{�Ƶ
/(������Pz�(� =*%%D
�f�͠��vK�s�*/p��s+� 3���_DB� um�/���Y�����c��OC��̄S
f���%r)�{���Xu�^�)7�
+�E�������J���!R���h��PV��7�	�u��z���ʟ�k��47I�^�(�}��C��{駡�t2���]�|�r6�CM}+�o�%��[�_�dUi��'!988 9alx��ѽ�i�]�P�Gwk�lN�%
�PGIUx�vu���BN�� ��a\����R�l���5R�	�-��MQ������@q��U�������:��D����Au�s2@O��y�����+���i`U������P��d��}�Cm]d��ˣ�M�T��gv�,��8�7륶���\��%���W�"�����V��QG
�oO�^z��{�A��r�w��6ζ$��Jղ=�R��:߶G�1
+�|�wH�s>�<a5�+�U�W^#a�1?a^��J�3`�W�@���W��.�ñ&� #~d��o���8�nea�=������9�5�����I��g��J)?͵�o�����Fę��*x8��]��Z)4ݹI�V�2i�:�H���M&cڊ���tuJj�7����R��(}9��#�� ���v�g��{'��T��XR�UEA�&n��CA���ڄ�M�HJ��mBM���[��]��@�14i��(�YӬG�;���J�I���|������TK7w�!�Q��$h~3���O�lL.�neZ����
:�E�db�bN&y#	5ϓ���'?~�o�@Z��T9�,E2���D����ۜK8x@����dM`��2M]�$c\����D�VT#��d�)��׍|�L8bAa4�M�
X�9Ѫ)`+�ea�	�wp��H6�v}S�����U�5s��4n�?5Qs|��/�M,.����c����ds0a#��%�g�4���xAq9��F�pi��jQa:��cz;�;Vd�#�����.���!�	vv���G��O����m�v\�̶T�G�R�)g�G/W�#�.de�:p��O���$�M��d��c����S�t�ُ>����۷^KV�ɢ� ���Qr�SŸ>�,8#�6uv
 �g(���z�H_��v��Ȥ�)DB�|�M8w�C��IiZxd�=Ƿ6@l��T�h��?�[�ܹc@�G���w����fy}s�Z�I�dy���]џ;�ӭ�qQ�mm����1��	
��|�e�
����┕���g���Ccx	�i�H	ӽ!O�B��2�x-F�kΣ�՞�蝮�/�����|/郣#nռ��{�q�, �Yp�kE�,���$�8hj��JTW)�֎�İ����\M��9�����W�7�W�AWl����E�F<�5_.ٰ��ޡ<q��LaL���,����G䊈�ZdB`c��y�����a���ЋD*�C�Y�i�"/݆T���sp�c���t����놌V)A�93��|~�T��N�1�V��x�J��EJ9՛�UTΙVGv-B�3r$ic�7�N٦�4!N^dC�r�Lx��իN���N�
�gd�V@LCõ;XY�$XT }J�*0��\�~]������மN�Χ�7ΩD/5`��&r��C�$��?�@��3��Rpc]בJ�O�?-ng�'��nhŀ/^P�G�qo�9F/.�����DtdgD��& �㉻̚�V>����v��Ȭ�\��Bf}Y'�|d��2�U�)���n�c�ї  �����C��ɏJ\�z��	�Q�)���>�x���|2|�!Η�kp�Ϋr�^�l;&JkI*Vm�}N��b"��C�:$��7#9l�h�%f��S���5 _( @��4��1�2��(�砬0,���5W-���V��v�+r@I�}p�GW6O&K=�����?�k�C��\����xJU�<�*vbг޴;A��}-�1��\��h�3��$�%�F�m��mlAW�zaKl�����җ� s< ���#:������o�����/���I����7��U�.2��<�f>�۝"�0��1��3@Y��l����ӑyѨ1��y�3Sb�Y��ka�jk+Z�L����a�S�����"�-WK��y�g.ݒ�;y:�X6��Xj�/pޥ�������/��� A�b���` �*���+R���	-�թ\f�Z��F�c#�y��[A�0�fa*%h�l8���� S��+se#�E�Uz�����E�Y�6���
hE1W-p��Τ������p�(����t\� �H~�r��̝%<p�d�N��b[�՘��`��uք�+&�r��9J"պ��C�������<�I G�{[�K���\-ytx�����Vsn:�rr�澛����Y�=y�d�"�L�G���+S����������ѣG[ۣ��ww׸6�����2	�G"���{�Mf�]/qf�4�zX
�gS�j�3K>�b7`
�p��h<�t�0I*��U���	�(�-�>��Q�7o��ȣi?"�I�Xx.Io���������Q6v)F�)�|#�܃b�6m����d+���&77� (Z:z4Q��Y�EfEp&�rr%�J�q�+�y)�c�ÛҒ�M&�\��n���`u	�y�~���-���j�r���_!%�&�:���:k���V�os������뱕��b�{�$+�@�,�
���i������N�T}/��T�ɴ�ֹ�(tʩ��ğ��4T�FX1:~0Yw[�B��2�<H�dR������d�<�:g0�Q0����&cu3�L'�w�(�D0������W0�Tb��&k0�)��F�I8�mV�E?���L �|��J�Ԇ8|������O���utt/\W�ٍ,�YN��rց��~I����pt+����ˆh�BQS��H揙har+�EJ��:�J����*���{�1T�ݸJ^����Xv�;R������ |"҂�S�&��K�	��4�6�m���-�!%��ū^ID@�8;����O�߿OW�0��5	���0�@����V,p*�[������3��:@te�H'TV�OMf�v���t�T�m_�ɓ�����U��ӊ�-vY�L���Ge�X>R��e�#~�k?�7���Gܳ�6�ԅ͝hz��T/f}b�6�U�zs�(N!����])�-�D��C���a6(�Y'rt���0I=di����ہ=��!�V�c���tua�,�i{Ip��_��Ll���N�_��)A��s�˄����qh�Ch<8��I��#�
��7J��G�+ZAK��YhP�i �yR!:��@��;�`N �y��-�x����|I(	��R?���{d�#�]��Ç��Ȝ����@���6��T8�<5��ڸ@��7�S`�QD����j�;���&�S*L<8�:�- �Sd^�8%����D�F���{�ez6�4m�(Ͽ��[+��Ao�$�:�b�9��j�N� ��|P���EMaW�`.���&�Y�f�yF�z	V\���qh���]�낍����_����<�D�)3[��g���-���kx���/h0e�v�;�%.%����'��L.i���q~��䃈|��짧�o^��y�Ֆ�\8#���icZQyS�M��(}�L�+ضI��=��	�:6m
���)���x:G_�5�������,11�s
��$�M�sa�O!���
��b�k3n��u������c�=փ|�rS ����АХQ*�5:�z�4*Wgs�h �����;��?���㗴�p�mp)�^�~����w���/;��f$}"�����+3R����t�\�E�,�����;�L8�(����|�>A�wk0���պn�gT���Q�s��5Ê��|s�����~��
%JΌ�E@:(F���R˃��*d8$��fų>�Ly���;����奏�Q���ߒ�^rR
eH����&��"�O�Z����N^�8NL���]��*�t}};��7N2ed��O�v��)��tLNNN`Cj}�}�	��>�닏O�n�U�w=�%^8�N)�rKn��>�z �.�,�6�X\�%%���7#,���cT��[HUd��<��L����)���kXg���NϾ���c�#�\O�2�=6�D� |���F�q�$��4=}�<�w�N~��%�5ћ��pW �ރ������@}�o��ݻw�ࠬ�7f!z���c�żP�2��i����O?���/���"��1~�	��ϔ{�U���7��[f�C��4r΀��3�i�]�HzXO��>�bF$��p�h��,s)B���63��4��!խ�z%��
Qi���g�� ���f^E�~2�<K��|^{!���m�dd♰s0�"i-�y�~;	��wo�>:�����E2c=0g�j�)u�J��?�o����!��H�A���p
��G?��fp�'�o�)���exd�.|�]3(�=WH�s&;��:YC�YB	M��O7�WX�ds��4H!вp�{���y��!���L���fd� �ԃ9�,���-�l@!B��wئ�:0���]���u����T����Ŗf�6��_��5P�-��.e)�N���Vs�kqE��D�쫬8���l+�.�{�"5,��\��c��c¾�Ni\T`d�� \l���܈������իm��u��<��z�����I�f�pً��]ӂo���<�%�_��s���ۤ?�E��t$=�h4t:Fo.u��EK�Zbn�I���� ������,�Tɑ7��������!����䀅+�7��R� r�.�u+�����[����̫C� ��@$I���$T,��}�N�p�4M��+|\�g?	�O��%�j�q���1,���I�����;H)AI/8�L퓴,���t�ӊ[���βM����S)C�I�M�U3:{'4tq����%���ͼ�ܺ�'�׉�O��1�$L��9�J���:���F˼�k�;h�ؿ�a��K@�k�m�B�}�!�C���jS�h�<y��GѢ={������޼9�1V��q��PKh�4�tF�G�� D�}�;�Z��ё�N�f��/,�mHY�\�ff�^ݔ�q�YZ9Si"��9tM�M��O��{���.�5v��T�ڐ�j·��_u0�aa���PE�2^]��/N%sR'�Rq��.i��:O#,��J��N!�FƉ��z���
v�A��^�o ��"�=4�y���U��N�{'�~�-�6"�Q����Q���b�Mm���i-W�nA�F�PB���&!&�=�@�	��on�0k2)+2@����+
��[c<5�A�9"�]b���F�3��Ϯ��[2�aō��$�U$��H�qc�7�5�w �1�{[�#���
@4	L��՞94������vw�Q<7�N��.eZ+-�������5����c��䅶Y�K��f�a*$q� '�4R�/�'Q�4�	�����ZÚ���v�.Mŕk&�.��f�,�t�w���+�(Y��U)�;�2	�I4�𦭻n@7B��朂���]�Nk���t݂�WyN��,SN�40����T6�L� a�}�
�Z����+��<�\I� ?��4�@:�իW^�eOOO�_Io����)�Th���y�ތf�R<4�b
e�
ȅ�~yzr���F.Hd镡H����Hd(��<�����3k�D���֘�|�Mp�A6e���*�|�����y���6�g<{�� ^�r�_6i\IG�FV��NC�w-|x�~�m=��pu��zw|��G%�Nm���ث�C�Us��bh��	���T��͛w��2���j����zY��W�O;;{�/�Y�|�	)�?��OGGG�~d.�sf'��Ҝ�vz���n6T�������kTL���"E��nos����O��%�_���*NL])��A�*O�`/(N$h�!�_�.��K
�#3�}�7��!'` V��u���M\qt*-�ꤋh��q ���*�sLv�O�x����� Bu��1��i���̙��)D<;;���o`/���t<x��g���NO.�`��/��B�	e	8�x!�i6�$H�Z5[[Я��lo3�.�k��m{p�N\G_0sb��m���7���V���듳���wP��!���k�F�q����u�sz�ZJ�b}	�ȭW`]���]7-��A2�v �0.$�e�$��K>d��0���+�	c&y���X����t4����\1&@x[#k�T6ӹ�oFĖ�o���2~b"�Z��%`�6K���.R��o�'Hx��A����r�G-���1@l�����I/8�zE!;�2i�L�%`������?i��+���M�D�ɇqA�q�(��S�r�-�_Q�uM� pF9��`�	�:��ni;���FiI���GƊ3[1��J:��(�������Z���A���E��٤�R'���:�� ��� 뚡A�i�8�Z�Rj@a���s���!�N��F�XYl���jY��0����'�wC'��2�|���?�u@�mw�g�3��ҳ�=d�jk�TK������!���/�B���ke=�`%u�:�b���e�Y6'��lP�td��<�b'�����l׊���[��Z�Y2DC �قj2�zp����b1�Wq6T���N@����v(��$̈�"3�����g�]��-믾�s9�T#��tC0J���
!��������A��\0^Iy��o�"��J<�oUk��a���zm��3��C8F��8��z#�;%��쩄�<�p�X���w:*�Oޛ�a	{�&����>��n��P�Q��&��zE3��$�j:Eq��)l�R�L��\x�#�����b�]E_�U�� ��"�G��l�@֭֏�� �Z�.�*K�_OշFA�"qM�x�a;�N�rICjS&��ď�����~���&��Ki�GC4�IX�R�<1"/Q���CF{/8�h�����lH������k8����Q��*����-��tG�a%u���Vȼ6�z����<'�6F-�>��3ߟ�(��v���)޶�.sގ�I00^�9�*/�pd��`��~����ԅO��n�0��\/���9eC�l��:���DF�	b)�${�p�N����'~��	�0��X��q4*I��W�b"S#6� �m>�'��@�:�/*a����f�E��?Ev��"8I t�L�I�н#R�H�nSj,�_tA�3�������6G����7��w�˪�X��T����Zn������첾��`�O�)�C2�zrr��ݻ+�r6x���I�D�K����=r��n�f�:E�:A42�V� �h����g�.�'��H�a�	��ڢ�\^cl~�V�̜� g�~�/mt�R?A�4Z��"�v�z��#7�,!$>4̙e$�����6W47�r�MK���]Q��*:@( _��
1�,r��<tB�O��U���"H�s`��
E��r��޾}K���'b�o�5�#�>
� bЊREp���΋n��Ç�T�C�l��0n�V�"=,��N�Z,`t����(�3���,��8�8>8���<���i' A'�v�0�՜d^*�j_=
v��y �,!�E�;���
a"0[�yT49�r���"�:�T2�I���)�g/���$D6f���
�y͖�kɈ�k���d�0���F��f�f�q/���+7)��V�����ogWW���3L������V���TV��u����.�+ IR,���yơ�uR�4 m�f=x����AO��j7�p��,SF�Tb&�B��b��nd.��:�U/�b�n���Q�A*tl�l�&׀$!�ʜ��!�l2MC�E��^6"mـ�ଙ(�"�G���_*R����$��I�*��u�,�SD!6fY����o�R��i_螷&SJ����N	j΂���W��ݯ�Kb�2�%��H��۳�{|�dF���j�.h]�(8ɉ�db���'����LGYY.�T0u���8�}x0�9 �TjCq�f,B�z<�2/2V(��<��|��GϞ=�f����8A��0^���	�	�dT"�x<�������|���l�V��q��`����AoV�B��@�eM.���n_�zE�J7�U����˗/���}'/I>6���**�ď��h��,Z��l!�6>!�]aI�h��GO�����M�|�/^:�+���L)ݝN3+d����;�1���AՆ�#�����F�`�/�uPi��߿��{2>���~�u�B*C���mB���m*:T(�����?��s:8�A��&�(���(���DE�����R�t�FP�V&tcr-F6�@���¿;��D��q0����!���S��Q,E��go/�ſ����I�o�jo�6� �K�m�$�-�}��������&���7ax�}�p�M�a�|o��y�Eoz��qX�Z�M���@"��'(&������X.D��[��B7¶ƥd��K��-�	wftR!_����U�ȬO:@0ä�z�Ȋ�cM|����Xy�J&��U���c�]��{A���������t��yw���䒞c��;����-Cd��n���35�j�G�!'4�s�JCݐ����s�T5����k���3�Ƥ�)
�)��<���t�G����9�{p��I��{�B���c��W�jei280�a3�qsc���/.���&��W�n����N��~\o�W��Fo/��a= ������o}B'�L;Y�+6U�����t2D&/��9�����m�Ŷ#�6(��!��r�!V���,˛(�S��Y:�l��א��\�����!��b��?�L;:�\���C	
��rZ~/e5	V(�p�a,����?¨�u(������/o�L�dڋ��S�^]��r���H�J~`�|<.����Nw��L&;�ݠӯnފ2����簿��˰f׊[�eG��A�L�)ՑBF����u�D|�a��_͂���xR�M�51G�	KH��>s5xM����f��+{"���D�ħ Z�(#�ޜ)\�u�P,������\V�:.nHW/,����z-�9s���=���j�С�6HV�%"s'')��J*��-O�}/M�H����/?<��a[�[���n$	�ta��� k� 9����:�q���t��P��%���cLj\V��mW/W�E��8|���x��u��t<���\��݄�)�NF��
AF��7@��3]���������r|��Z���.V�.���כ�Y��wr@S�IJF�r�4��G�A�9�eQ���k�}�[��_�xh�t����e�.���i�\��$uǐ�������t�F�z�J�������f�ٚb$��h�*K�(�~#�@"�o�~�ϱZ5HӬt^{��^w�Ҳ�Q����=�Iae] #�Ÿ��Btrs<�O
��O�����?���(ãW�ҧ&����O|�bcb������մ2�b(U�@{IɊ������t>�v�5�uiY��q����	Hf�3���n�k^�K�n�PN>_sߥ�����*SL"�/�,�ԏ/�(,�l$X�Y�V�H��8�.�PD�\��ݚ%���K!V˻6�����ye\��ѓ'���ȗM礚��,�!)�t)m�s�5I�E'���&烼@������"��A���x�
�El�"�S�V9��ɦ��d������&��e��M��K�'���� x.�
\g�V-��S����⊄����3�.!���N h��ߗ�u}}s#��T�>�H:̴��V������ao�GY��j�w������	r�)&g\fH��}�������'���6]���d�/O�/��+gq����Y�':SI+A4��$l$}B�������{��M�X�1�N�
w���.s�$�G�cq}�w��s��\[�������d4�cdG1'�5����ʫ���r�Ӊ)G��W�R#Y��P�u:���H�x��t��3�ړ-�����H�`�����z)�攧&e+F�l.usN�����pT�p��utt��Fz�a�_��������h��Mv���B��:	<H)Y��`�����8n�X-T	I̊��C>:\M��I�]�H�\���i���f��2�dq�]>��rȲ�&s�{sO��]Bܵ��O%�F���Uΐu� �Y[H��4��kR-��poi�U�]񧯾�Yn�n��d��ѣ���?�=9~��[Wf����-)ln�^ԯ~x�^�f����OoH���..��߾}��2�W7׳o^���.�zݬ��f���(��vTVR���0C(O:�m�_��F��E�2�ܙ��A���jEǐ���c�����黃���:ؐ�A:�����p�������7o_��a�������U,"	�b�)�J�2OV/l��!��t��|�bL�Nu���%m_1�����~lӭɨ�Fy��͊��D�0`�.��p�4s��?�|I���A��g3ڹ)��,���AI�zqy��/~yu�Ȳ��U�:>;nB��Ty��~�+hoY�3���M\�j�'���D���1���̷��N/ίyP#���3�����4 �FFE!3��hb�,3}@j�0�i{{>%-�pנo��45�?���@� ��$���>���>��������\'N�4p��<(za�=�| l�dD?z���OOO�1Jh�-��<�b��5)y�*w���>����%��蚓�|'''��8����-A���ro�p@1���q?��'?���������x���_~����v���:�Ys����	Q�7�h��ሉ��Ê�2隘&ǲ!]���LL����U�r�p6�Ms{}~�������6��1���K3(Jq~��׫u�^R��DG����&$[&��A2t�Y,W��$q[�/&+��H�	Yu����3ڻ���|����%�x<��� �l�a���6��c���F"�3��L:�"PR�5�u><����?�O{�%� ��AƧ�-��9��`��R��f�:�1&Le�صRNEa����C�NdB�4M�V^�Th��B�}9��y�M����I�*2�k
��ޝC�9���xRO�D�!�f���rV����^�|I[��ɓ��m�Z��ױ[��v\C����zXUo^���'��>#�����#���fmq�j����$s$ZW8�UA�����<���+>\��T>B�Z�r����@��	u�/�L��bBƧSj#K*>R(ߋ��������gM�Td�)�*�@�I:�������w�R����#)ް�'c���勓$!�� �[�U����"֋��ތ�uéC��]����r~�"nyѓ�\�<y�E�tԯOO�N#��� ��;���۽{���R�ޕ�"k�j�ۑ�I&ZF{��s+è�5P@�Q�s�e��Y�R�Že������k��tv�L漕��Ѭ �z���M��C�]���T/_��E��;.b�Գ岶�$���i��`��
y7.ǜY+����.U�W����˧(��@�<���������11y�]�]K��|�"�t���}e����t]���i�:Gp®�Ŝ��0+��8�	�����E�CN�u�8�Re�D�<�S��q�}^�h��0�"K��E�< �	�g!��ٔ��9�T�n����;�Gj��&�Y ]B�a����\���5(���Oj�K��oAI��M��@K��|��㏣��>x� �J��_���+�I߽;l��%������"CY�m��	��>/�*Õ3��-��U���C�{e���cP�5d:��eV����OP��zc�W83�ojy�N�y�e�UCon=�M�d�Vy=seGF��GBeF��ݯ�>����.6De�WӴ2d �����_15�s2,K�J �a#��
�鱌-�Z�"�~�;\%6d�iV��R(ꘔ�\2��d�Sa���AڻA+Y��!V �H��@�~��Q5�n)��#N~�ݻw�B5C��*�
�79#I�|!(��m�v����l���H�8�O�`��ŧzK�p�;K=��O��f���e�w-�>=$�Pp����C�:R0$M��JgQ(���[�|�G��c�+gf���@o>;;�"�ad��#ƂHH�k%a@��t�Dj�u�in(�@�)ח\��Y�I���BA�vp`{%E��2r�Ms7��Pc���2Y	�� �H+���@
�?�+�ؽ�	O:*��S\0���`�fY�:��`�}o��.Ȉy��㹝�G^�[�|U��t{��Zc���sY/����/��z�S9���	ş�s��5����Z#�^u��PV���lH�N��K�������ೣ��3�܇!�薀CD6�:��	$�=Pse'��L�ڋ
0��a���c��D=	�kc���:�ʥ��EM\�mV@�<��;;#��N)2�΅ p��C���=_s%�7w)J��^�[�b��vvyR��t��v�{ M*|h�G2���p��݂$N�����F���CC.�>�Q^��?|V��	^�)G�.b~yؙ�-�ʹ����4��5$��|�s�^���XR�;�l��q�s'�_��s�&��t�9WK��Ӕ����?[S[
�3:s�vR�X-��p��0B��S�M�Y�<aq⠚�t��Ú�ӕ)�5R+��0�-nf��$,�%�Y����f���b�.�\{�_�P�:��4�7��xv��wߑ'�R1:���f�(1�-w�Iy�����\��=�U-g$7�Uo�~.�v���Õ)-�����}��C�= lM��0�CY��E���v���.�L%�����5V�Y�&`�U7��=����� K���L����n��v���(�e�)��۷o٧������>$z�a��)Z_|���;;<�[���������2��%�:O�O-�''���mÉ�6b�OT,*|rx��A�W������K�5c����Y,�q
m�X�0ι@8���y$�k�O��7(o��E�����:�Aҟ���{����������>���v�FBK�f4% ��F�W1�ش?��Qu^f0�t���V<����y��D��I�E�e&[n�.��n1�ʞA�C�M�����՛_��Ϟ=������ߟ�E-����L��M��Q䛱]+���٦u���L^:�N�W� ܻ�^�"�$!�ڃ�X�[��-��i;1x�j�M�Y�B��$���d	���,��ׯ��
�9���M���f�6�>����|v�d�5I�eb]��+̬��]md��\a�谹��yfE�s���n9�Q��YG�#A��+t&$�R�9�k��OEb!��^��������9��	�O���oI^b@SZ)g�M�z�T���]�6�^��o��d}��?T������ (I8H��mzef����n�L������J�c�VP��d�u�e��5�`�T�#&�)�~�mjA��������)/�@uE����yT��)�ߧ"Df+\7K���W��E���R r0Z�����>��X���e�*�7�2:Lt�Zi���/>�)i��?�c��)3b?zt�vy�5A�>�F.	&���rj�!�v\]4�aS<�C�-ޱ�c�Q��)�V�M�J?X˵�!hw�m��9��Wl���N�	g~3�«"�	蔇���z	Y"�Ag���&��d&�x"��a���^0%V�'���t*��&�@i�f1�>u��v2U/G�m ����69	��ȪɄM T�{�3������F�RB;�/ލF,�f~u=�����%�:ѭ
K��ߐ犡H/�KM�s3���!a:�������6��~���M�|2�ɪ-7G�[�Q���}��zi1 �ms����y~C�.��T���-��t�k:���p�`�ŔiWnV��:�K��V����U�(���HlvXǧ��u)i(��1n3Dҹ��[�+>|�����=��\��8/wP�V����3���f,X�{��N���^�4�`��eoD���i{u�mD ��93�3�g��q�1��̸L���=㐆=��g�-/h� �i1o�d�h��7Ŋ��AhSX�F�����N"piq]�Q��+r�@֮<z+έw<^���sd�8�*g��h�6t�<��Ě ��z��s���ɿ�ihKaJ7)�����+�Y�_�Oh.�lmC�0��Fv-�(�v���R9��=$3�Mi�`�vkg�=�T��^�Op&�r�P�?%� ޱ�I[�
k	��d:B�2��
����\�D�����-��oQ!�h �fb����z��n3=����<+)Qg�9�
ئ�3���E*'�o�B*��%��81lVB��NFJ�I�!C�`��5���\Q�K+�@i��T�
�����Z�YtE23�	�.�b�g|���g�j1N6�!���)��ߐk���o�֓L�t{�}�j6cV�ZQg�?�l����A��9��2���/�G	Jz�Ȅ x{z�N����_�V8�apx#�o����b1�uJu����.$�PNG��7	b�o!�{C�,K���B�]
� ��0��#h�ʧR�6�0h+>�UǺTjČ��I���D΂:ʥ����eN��onq�-B0�(u����q�f��-��{~α]dU����ޮ�Z  �&�cT�$[%S�Ȋ�A��c��E�Z�x�/��yO�	�$!��H��{������_�L��c�>�Km��/ްh�ͻӓ�ӳ��'�H2��9rEb#5�ٍV��`�<ؑ������ңݴ`#B���a�n%����V�u��r:�,f-�a�c$�p=�qa�����"�ґ�*׹�hR+uBh.������.tm7kfr���#��]-��6Y����UYz�'�J��>|(�Z>W�W�o�y���-[��_����}���H�I�V�.H
����kF���5VH�dk���er� Y���9o�@@]�S!^SjQ��;΅GH�т��2��-��c���|5o-��ۃ�D���5�����E�orK�r	��3�մ���sZ����s��D!�Х������I*D�K��8���W�驥��u���(ls�5f��o���3D��6��U���׫���?y�������XɎ
i>[f����Hi5W��A�,������=�?::Z͗o޼�ݲ6�iNƿ�X�-�� ���lh$���¤��Wjd���o�0!�t�,,tć��i�N�Fa�sm�wZ.���H�0 ����O�=��/~qx�4(>����cz��]n��6!ldS���P���o�JgO�Z�߂�P�5��J>8'�RS%'��Qi���u@_��=��p�?��z5/�����߽x�)��J�k�#/��a�͖%ˎ+�}���|s+k@@E �E��E=��I�z�~�?��L&�|��M�H��.b(�ԐY9�oLg���k��)HlCXY�͛'��۷�˗{,�^V�G	 �l��,˪U�,�b[mv��x6�T��k&	'2[�죜��'m*ctʺ������t2C=n�ū��U=����Tn���-Ql��N���''��IL]׍�ˑ�Y��`~�h
{��Z���WE*c�:$�����>�\�f� 
�h��p�y�"k&�x^0�4K����4r�ZAE�`B�ˍi��U^�v~�n�T8�n������*��<Rf�U�vS��#��}1*S����)*g�u#GMG��F��o5�m	��B��*����m��E��_r���y4�C+cu�6��RIҳH�:��5 �	�ѝ�����Aj�h�b�U�`�3�1��@�J��'���� uK?:���]x����k����jY`��p�����<�m�EWSC�|�A�9�XѦ�X(�U��AN�aHyެDUuS�Q��7��v�Ϋ����?�v�3��۾q��k���؜DU�ګ�> �}��w���>� �E�!2�1�jj�����g�7ʦl0Kw�5�1�xL�!��<T���<�澷�\r��QhA!�YL�����M�>Rd�P��:==�"}�^S��]e��Xv=:���׏
�mv�v���`AJV���Иv��2fH��y�4jY����F���Z2�"bz�����22_�����@�R��sm�S-	�����\ΕNb��ζDR8�1��Ѧ/19�[=��P?� q���bD��~x���gϞI�/��@����b"�c�a��KiRQ��z����z�QA��y���_3�K)-��'''r��O��&V�ѣGl�"�P�ݻw� �ΒK�5sM��jY��ږ1�A3|1�<��0���[�7�hU�"�#�v���=��~����C�`��Iʈ���Cϩ��[��3��S��C�_�i�}b�	��v�6�
�̍",����8c���iܼ~{�ѿ�J���"�G��%�Je�9f)�#r�Y| 5z�Ǥ��b���� ʶ��Q�ӫΝ(�#����s)X)R���b�:�����=���C��2�u����;?�C�df�p���\�q[i�����h1)��V�rS�&p�2�W�	ùTt�3�C�67���,��Rrm��.�����e��RYF�o�{8G�nV��Ki?���H[@�$w�����,���3�����Nv�*�J��2T�#.�H��h��c�`u�"���R��ٰ������
��Qt�A_M!�N�j|�u��O�_�`4LPf�Ю`������sͽ�!�J���~�9t1���U��{(E�Ȗ
y�R��0	�p�ԫ̍f����p{�I��^YQ�l�խ��3K�l�!D�4�9!Ԟ�<wm�F%\���r�I7%��J w��=	�mbD��(?>��#9�Le���^���� �J�(�0�{E���6g{�y��P��w��
��`�R�S����� ����!95�n��zy(������G����D��q�$g׾�r�&b=�z�ڰo�7�s��5A�JyO�&������h�Oͱ��Ҳ�[[;�|-�T�ï f�VѦX0q̍`�����xd\����F�e���/�c��]��#Wk�����]&3�2�_��Ӫdt`���M����vaS�Q^�og�\��y1"�)0Z�����jmSQ�+|�����I�r�X�A��k�c��p	��C�ķ�&�J��hqo��7��~�Jgv�Z�lq��ʷ��W�	~��g_��/%�`����'�<��i�a�<�!��ڮ<2$F>��Wt�CcT崶C����0�h�	�u�����D���������3̺^i3g��.���@q|
k�Qͣ^�È��cQ���8�W�\A�N��vk��j�����M�a�`Į�κ�\rh��{��뉎�FS�6kr�~���_?�����::o����W�mD�ɳS[��L�.T���s�2Cz�8��� Pb�ɘ�F���ho<�o�M2e�Brx��!z����`���M���1��w�{���:����W92̞���Db�H�E�����Y�"�ӵ����q[
�ֶ�(����CS{���I�р������r�y�zZ������1���xE�٪<�<�\Lf�A�-�z�mo�W�,3��R������~n���f�(hac�
e��p�q9v����E�TD%S�&�no�_�����!�A��*��+��I�+��k���[��_��(l|b��]��VjZ��C#��[��|C���U��gdo��l�/um�Z��4%rF�)�T����MfS�ixX���hG�:�3ˡ�F��*�jSR���
�:&PUAA��-u�EL)�o�v&#]&(���4��)�,ʹ++��PT�aP��qa+Ff.�!f:k��7�V>Z57�2O�C�sp�[@��SaPHq�%{K���+�KQ5?�4���w�u�Y�_���<��A����y��"絛�x.Ճ��`:
���F�K��"��H�1�N��G����P�s��s���T�9��uY1pV��]-��5�FD�Z��)�P���~ m�x@z2�U>\o�ME�2>��83��`�%�����U�v5�ӧ��'�n��n�故��Z��%��R	�\!�OH�|���ݻw��w�A��<�����6\v���'�k���ϲB[�$�Hq	�:�3h�k�'h��K�/�Z�Đ/Ped���E��^	����r	��MW<yv|z.�t��!y���k�C�RSMj��P�+�>�s�m��U:ZT��8@��ē'/.��r��љ��y��zR�uuy�W�=� �i��8������Z'��?����>d�Dӈ�T;�|����XR�����3�77<x�l��e��/��ƫ�Zs[Ϗ?9=9g�H�/ vE6���:��;���"���F�$w��c����j���E cs������3�d��ê�N�R�h�<;@�"��E��.���?�4��+�7�u�$&_�i\r�؅V#�X���h�L�Mno{=n��6��a[�����g�(Z!�E#7_,i8+��SZ�%6�	�"_$�U�9�TpQ�%C���`���r������?:9g��++ݻvDW%"�+����5NԈ�M�Jw��>�ȹ�$���R�A��؞�;���4�Y�}��D��q6��YT�e�|����;��l��r{� ��]�,`��+���!H��u���K��� 1��|�]�ӲdF�e�X��d"
!��|�T�V���#Cv,�c謣�K�q�1����������f��-� ����ah��DGKL��*��)Q4�����Zf�jU9&��lI�.ia�Gܚ�ы����[FM�Q��K�6�9T1�D�#�V0Ǡ�[�q8��Ŝd�B������.3j��z�=v-�2h���@������g{�fC�g�5�hU�r��4zs
G9�]�w����_��  9���=u>ƸYrXNNN� 묾M�v��|��Z�(0c1�.p��M-XR��F�H�5ӡxd�aDʂ6���o;z�K2O$F����` ԅb�e������Y�&If�O��\�<f��V|~�����f�y���WJʇe~�g���P~wd���'�8R��E��<j�[�xb�soog]/w��ٹ��5�N>�� k�*�A[VK������~���;3zM�VZ5��*��U��O@oe(��"??��8���u�T�G?�8g��t�O�|U/!�Y�ש2�^YE��Y65���LpJ)����7I��۳����` �b�x����;R��ù�<'�Π�\�� s����oa��S ,Iӗ9tu�V�F�cԙ��F�k�z�5��J�Ok�c������W����*YX���d�_�<���@��@TP�UӶgc�Q:^���d��҂	���<e���Ϻ�뿗�Ա�)�S�j-�Y���3U%�!���9Yw�(�&�<瓩�GȕH�Z�)��)�"�b�D��;�{�ݻ���[�m��=�j:�cQ�R�֫��)ǔg��vA���Tzdf �����(�Kk����ގk�Q5�׭�����o޸-?��g?�#���/��K}�<kA�Y�R��N�΢�ڹ�Y7_�s�Ո�ZCD�&Y��sڵN��L�;L[o��_� ϳ�BШ���0<u�^Kz��"ښ^��?����}��+�;�Z���NS����Kwy~�	Hɭ.�I��6C��3)�<Y��D�"������+Z�W�[@���Cl���)�JĒ 9� �W��S!
�P�gV��g������z*����;'���,�|熦����ђbv|#�B�5������ �9�$,-P�}���d�����b.Z����|�&[�7}.���8��7p�YL�kw6.�0���ş���q�-�b�d=����?.{�T�`��-��\�Wɔ��)�t$�C:����:���l��2�j-�`��S�tL!��;>;O�����e<�g'�F;E��\�<O�(�&\- &��N����}l��T��zܸ��g'��?܆б���2F#�)��jڳ+v<S��]\�2�/2�OD�沫�wѰ�
��qb�ww�Sڱ(#��p��:3��R7ׇ�W�\9=�������z��2�Yrߝd�=��s�cC��ğ�A֜`�*a$7	�i�#G�a,�d�U	GKA��X�����v��_Ы��ZTF��f�i��ia��b:���a�΂PR8�q�R�^w jj//����)��=�}|�!�)6XW4x���{7*\i89��>�-X̶DKX��f�_�B�[L��:t�`�ì������!�Y�w�6�+~�U��&�֤L ��U7�r�D!	�%�l�5��E��U�_K'�rgk:W{�۲�_~�e��G��#C���ͳ�9Ȝ �r��	�+{"]'/��f����|���!�(ҭZ���C�1ӡ��^U��Q!�[�\8���R��@��P�Z�f�5+-�ն�u�M8��+U������z�ֺ�y`D%����,'��ܸ�"Ȟ^!��~Vօ����!/%�X���EP��D~t�׹�f��0�>==EP1�
"At� �(D'��e�~���W�h$���yOtyy	+��W�c��UR�c�Ü�{����d -�����K�ve�X�<<b�(y�"B� D<}���3[Q(]�y��!���S�(`���F��SN�.���moЧb0C�u��z֯0�G���Z�"��S��ڇi�1<A�
̔��-�)�7H�s>.�����]^�&Ԉ�3���zt���Zc�����JU���`C�Z米D�q��֤"6�DʙJd���R���Sf���AlQ	e�3��*fG��S"�wo;R�8ty���ij+��Z�0�͜f? y��	jk��S���O����F*wq��f��X�Ig�y�Q��}cӵ��{ĺy]�yon��a��J��1{�	�}�d��"�u!�h���L�ж�Ӣ��i�i>rJ�Li\��,�ܡ��[1Y%6�]�����@`�%�铲*р�ts7ٷ���2���Mm<X�Ln��������<��^�t���_> ��?H�]�;����F]MZ�V��o�w�[(EĜ��� i�b�8O�4�Q�ݡv�l�N+��v�#aVu�I�J���쫾6v����ޔ�!UuWe���׽�	W�a!ݾ,����X��T��)c&���R�y�v���������Kڴ�}����bo~!5�T>>E�H����d�^f%��c�4[2����MJ<a
p^�]}q���|dL�p_��%�PDF�xV2	�g�����p�e�-�M����ݺu+�"�v����������h�8����zZ���-���r[�S�
"��䃿��GD������s�S� 
u�#�%#������,������1�h�1uD�+W$WӍ*:�2 XȮ�U�F��Xu˒_�WSoиe�d:�4l[VzJ��rHSŘo����WN�D*��W�^�~�իW+��~�*fjU�N!�*Q�^��cΒ�ܽv�Reӊ���uxy~���Yс؂���UlT#n@����"[H�<�z����~��O>y�P�j7� ��u������j��
$�hѸte��R�,�-�V��d �]o��|j
7%%���`Ժ4���d:�;ֽcq(X��W��|O�w�[b���W����L���+���Y^�!N�(8;�'�D,�Ά��m@v �S���Sr�N���&���o�!�����Jq����NUF��?�豋�ŕ�[��o\���EՁ�Fw�(�1��S���Ra�qk�k�����F�ҦpL��KLC�[A��������h�/�v�"ttt���s9�(�����M���<�艺�
�Pf^yݺ~C����͉N������b�z�3Ia����[�����$�nPF�䫻��(�9�R��%n�g���o���ѫ�䤈q�5W�4�ln`�a��	$Mi��vG9p|G�����ľ���/R�������`��g���U�D�3q� ;���?��͛7����w��D���'�"�'g�����ڡ�˴Ϡ�p�G��Y"��F�t�XI5|h���Bq��u@�������#1��>�r�
L|� ;=>0eRmB��'�ffDz����%�px=׮]�\���`�)���O{!b	7`y�`����lT�C�bd��	/�I��	��wm2���ֺi�Ih��xN�4�.���Z��$D�$.lfmD+���ˢc7 ���p#���	�1TgdY8��M=83���p9.íM�v��K�K���(-��w� �v��$ŕ(K���'��e�4�Q���R��{��k�
d>��敱~�z&�e)�ׯD=1�6u-MU
�1�*����J�ea�;��-\�֤י�Eɞ	�#6Sq`MK����:U�ж�Z�u˯2���G��Wv𠴠���q�~:�� ӕ^�z���F���b�Q�	��Mw�q��/18���#�$ǇunQY:C��Q&Y����A��%�@ �^=�q׹�]�h�=j�7�8�܈��AЦ�>��.Ē��.�s�M�K�N*�$�u�������x��8�(��w��,�u�>�[7���鬍c�n�$��;l�r�l�v�b& �4붹�U���eˬ�k�f���
F]w���)��n/W�ȏ�^�렌!�:�L6��U/����D.����¨��a��Y���4[[�R���>+G�|%�X�&U��A�L$8�鬨�>��[�uW0��|nYsƐ��r� ��T����KZ��Aid�=g����QDk�B�Wƒ@Qv,a1�P�@��cf8)���xX�^���[\%��y=�yTM�̬��K�f`e�-*5�#,p3�2����zv~���i&�"��
��:E�0�Qo�iό��$HͶ�//r�;KH�J�����OSmأ�g���ݩ�)Kp� h�����퇜"��L�"��	���L�C1������:�(ؔ��U�4���G�o�|�D3,.��!����X�����J�u\������hJZ�:��0�+����4�)֯,��|\��tZې��)�gV���!zb�	�_����Ӻ�]fH�קG�[��.��˴��'2�e	w��~�7ƪ�A��)��b��ƽr�fܿ}uf�d��]ΣM<HO:�5c�܊�C-����TM���r��;!��蜅�krK�2V�D�8�n��j�P,��̣9�z0�����Gᇄ�E���>`�f6�Q�~r�g�\=r(
������\����RL.��/Fj0�	�<��������Ԏr	�Sc�
�QR�D��_%�q_�����*�f$���\X����G�%�-E[Zou��
+L,�i������� 'Z9X�&ZS0Uk�r�jʟ��
�?힨|����ml[7�l��"Ÿ����PB���J'w��yg�T�A%\��y�������۷�߿��Ԁ�d&#���ZW8fZa6�un$�	�y��n���m�������pJ
ZPY���B�lڵ��r�ׯ_�;aq^��˗�;�u�쁐ɜQ�k̹�WC
)�E����_3��;�c��d4e6P�r$A���4F���3���Ja～ Zs��J]5,��aӿ�L��R����>��������n�u�/.�Ġ�����=���/_�����|����p)�ϙ8��{s�T��<U}�D�d���2��r����zQ5��r5�-���D�9���|���?���T�;��7�xڴ���:�W�US��)�ʪ66�5|�˥8�� 
���;�ѹ�e6�F����:'�#G�q_E�_�).���>���;ƀ�M�bd�� �e�c:x�>�Òñ��<r/ �ͪr���f0�����L��!^��lgW>���(��vfxmأu4�L���4�/�J�l�Nfc�t����D@w��m�������!Dvȃs������Q�.�'g�P%�¤3p��q�.���Vz)Y0 B�7Â���es��H��v��&����Gf�9�"u�:��(�I6�k��85�u�.�����x2�����޼y3St�b9��	��(�|�ً/�>}64��@�Vܦ.Peڦ¸S'J3�����[o�S�!���PM�T����<�x�(��CV� �u�<�X0��|$�_�����ɓ/����������-��������''g��s�h|{�mu�qШ�0l��tt��A��}�Ϟ� Cc�oۄ�dG4��{���d����|�6��r1������@e���U���A,��P�eT� fEof�����͛7��珿|��|������5lnJ�%�giL,����ᡖ�	>�q��"��gͽ����� *����'''YjQB:-Y�V��l���*��tT�d��Uq�,���b/9d���p���7��6��k�&��K���OO�K����pxz�Űj����}tq�3�JN'�|-����}�����Ȗ�8��k����ۣ�?�Y�Ɖ�}m׸�Q�@	o  W��8�����M��������
��9�p�	:�)d�f^ڌ��x6�k�{�n�����Y�Z�v=��%J���@���y`����_9�5�/e��)�XM� !#�9�x��d �Z��d��0���iY3٫u�"�Z�[�Q�n��u�g�%���Z�S܉�V�B���Ș�E�t ��s�Z_���PW�;|S���AD�8}[���M�[�� C�i�U�p��vE={��+4��J�a�q��E|Ht�i���$QA�̍*.�+��*�F+Ql���ʵ�l-�EĀēsy�W��|����{;���cX��sP~͏^՗(׉+'�*(�>�U���\�,�px�..�1/N��֫X�*q�kޢ�������`��ћ>�;-0�<��m��X2�Q��i�n�5�Q�%�/dg;�Js��8@�0Z�,�0!(���E|1�|�ǴB��9����e͟%���T>
����f�����(HR����-��o�3�R�q�y���ъN#��k<@��\�Q�I\�^���Pѻ��JL��tRq�������8��g�i�8>4��C8{�J�3�<��5ԆZXrw]�j�2��`H�l��ԭ��ê�3���ނ��iwϒٴ���ӗ�Sy�rY3OA���*S`b9*eM��H���O�?==��9ElRg��sϘ��wy1�B>8��pR�]��r&����n=z�H!�˱D��L;��H�n�N$H�A��5QP�b��k˿��liK�����ք�LiԔ̕�e>�����Pk-���~�7� I�fF v�,{K%إR��l�`�Wۣ�i�y����yt�V��y~y�(u7p�"M2]U��fC8�_�'$E��fG�����5�q1I[,�|:��rd�0[��,5�	��@KL!ou$�"S��kN8٘�<� 
i	�a 2�g�u���>o7`�&0�h���?y����;;7nܸs�69.��R-���
"84�h-������.���du6��;��T��ཊeҔ�v�,KW���ʓ�J�If�%�F��ً�'�c���ޜzZ�	�7I��&B��Rεz�	�G����p.�i�-'�w���_�[�F�Y>8��$t�</� D��P�}
�{�Sg��q?8�M�a"\�H����=�� �"t��[n���Ľc�O��e� �ͽ{����ȝݦ�>	�z�DpMz�)�1^u��^1��A��4��G2S����z�\�A��Fc�v�mo5a�C�(�L?:Tz�Q{�����p��
�I�_�N{A���bZ����q�-%�]"�@0���%HW����S\�r�D�nJHI��Y\���7����(Z������of�T����9=﷕{��|J*�p���CR��o�2�#Y�	���#�#1MY�<ɔ�٦�F�Fa���۲ԟ?|��>}�
4��,����K�+�����Z����J+m�:��)ͭ��
����������s���nX�Ή: }��/)���_�:���U��PX`� ��4��W �\s6WTN=	|��0�����\����,9NJV���k���pq����#@��^��r�vp�j�bU�2�o�׋W�Ut؋�jՠ�ü���s�p�H/5�=��U%VR��ڔ���D�*�K�c9*h�X	@db]!lp��!C��DQ]��ϟ�g� �`�r���R�t�u
k%���A7�1�h�獵�
��\Qƨ�V���#�a��.Kq|z�G��42k(�t����Y���� �e�{�}W��m���5��O���ի7oޔ?�E���%b�����O>���ѩzvB��,���.�P,3�O4 �	u�|���P޳wp�tr&7/>j�8Wօ�>�@{�7�L�����)�ԾKe9h�1Σ��ӧO��j��|����w�������������,'N֜���c4��{�O���Nk���)V7Ax�)������'Od������C� �V,�P�B���5GO,mU�f,O;���H��g�Q{��k׀Ǒ�x >6�幨Jy�[�n��|����Arr�����>�tpp����h!<�2���	ʅ�8�o�Md�g*� �\��Ç�Be��|B澱�t�j;������0��k�W[�Djvo���sH+��+�*��X#��V[|~}
�{��O���S����ƣ-Y۽=����b��t�������^���6^ pB��5 >�2��z2�ȽT�s�զ">��$��/�eo�\*��Z�[�66�sls�n(3
���w\ë$$i��l�D��>� ��.vu�.G5R��0%6�uӓ�/�1��[mZ��̹��՚̓��Ͷ�_>}5��RT�Yۣ�3A��̟�bV��lDJ��Ө��>��m�F�u�cP����8�=����B�`���w�ζA./ϭ��u��qPB�-�ǩ����$�w�\ӯ�T�W9�-��L�ͬ<�'�Ud	j_{�59#�����z��7��o�Fކr�UFg3$^��/)��u D�Mq4CTV�u��arY��ﭡ
���N�lm��v:2M�h�b0TE#^�����_����t�� �a��g,��5�&#Ͳ(CYaXv�bT��/b֍h�P�a���������[ט��Ơ�UyQ������!�qVt}�!�#�#���^T�L��})��(����~y�h\-�:V����{���E�j:�4��"߬s�+�!`hSXi����{����B5J����7��!م�+�t�X�Y�E���'�5q�"#k�
i-z<�*�sV�n��X`�w�������#O�F��Y_Ro8j��Ӹ=�\I1��)����ŏ>����e��m���_X��;�Ρ�w���l,7�wU�F�fV~��5��W���+W�޻u��]y�������f���Ct�4�� ��K���?iF@�S0H�X�k>�YN�/ҫ�9]�uUgF�,�qN�a<�|`�,)�8KĴ�"3ي{�KL�@�b#�'�ht��^\�TS�NN5m�-�����&��fo�ę+�h{6��2{�Gu3289�1Y�a�:rF�I��rhVE,�d2��e�W� �sqP���RO��VM��Tl��3�@��~E��u��sϠ�oZA��5(�	��Z/�����d��'rc�&:�1�02^WJ��IcG<q�1�UT��G�����o����ZX�6+�R��9�G���-�K�#����t�r'�&�Lm6pC�5�٢7>t݆?��A�Y�h~�]y/��f��|DŽ�!��al�h����h��e5
V×e.�"�@��nQ6�\F�tF^c����v}�X7�\������͵��I�|��JTn��414~L�0��(6WbA�k$�à�<%�'9���W��'����ͅ�[$ڻhÎ��TF
C���[Ig�Y'����0��%������酜��k+qaX5�ȯ]�&�Y�H�+�e0eC흃x�8��?�G�6[~P������#=y�z�2H̳5I'E>K�Vٰ�V�2SUF���ec�U���;;��E�:�Iw���&3�,�ٙϗ
����Y&_�-JY�,�I<&�ś�ypj�Z��\QD˥�?��vG�Q.%7!Q���6t� 53��������w
�<>~%n���6�c���Q�u��E��MN������4��z�("�u�-yNN����E�-�
���qъb^��̵��T�U�ˑ"y��\����|����rC☯�%���ݝ�^3�����/��(җY�RaC3��f�K�ԄDy!dm��x6�c$�.�Ɉ��ڦ�� �$Ǯؠ��=J@@3�7�/�d�|�h���j�~�tU�����w��@"��аs�E�����]��q,ƭ__�ve��cyjYKV��[H"��YV�D�1e�#�^~ʡ<2�!(�7�����1��m
3g�ok�ZD��oQ6śa�=�#�p!�P���j{.~�F�����>d(�δ�A�{z:;��p'kY"B&//�� k�Ԋu��u�Z�*��k
�����l��X@А��h�������9_l�]3�T~�:������m�,V�������3�MǨ�5)����VR��c�%����7Br F��P�_./�<ͅ�;�I4[4�`� θZeU�#;�sz��s�T&��p/=���N�y=�����W�z���~�Ν[r��98@����������ӓNA{��lYI,���7n�-��&�p`��7L:�4EY-/�)d����x��7o���◿�w޻wO�%	�Z��s��#Z� �&Yb)��Ⓥ.���(@v�����a�m"S��.w%g��?���!�a�ʠq�2R��s�)慎��1�!)�=%AY��Y��~]4ө����]��vw�QU]�z{2޹v����y�E�d��X����?}r��]Y[	NG�ɵ7�VǓɕ�WţĶ�^�x|��MQ*���_|!
����P�f;�T��8��v�q1mz�Ν��]�#�&��u�C��,�&�'�jj�Sb��q
+��K�����|~q��B �f(�M�۬�1y$�z���VѬ��5SѾ|��Ȣ<c�M���q���ߜ���t���:{���޸�z5-�1i�&�P�;{�𯲢*�H8���h��1����'�;m� QB�g��t,�������z�M�P��J?'�_�a�R1�Գ�D�Q��XD�k�o�G��Pl���;B�Q��Id��i~u�p�`���y�GA�h�Rk0�����^�#��j���6���,U���t^��@���;�h�O�y���N��h�i%~�q��W��m�F�C�Og#-TgH��=�!��7EmF������=1�HF�p�����'��$�'s:����z<��ɡ�俭��R<��2���K0)�E��x6��E�K�Ih�:��a��E��`T���(#�$�����jmF˖�����G�"��.u�o:#�>�R[tƎ��h��
��b�j[^��祋��cY����r!a����ٖ,�(+��w����裏n߽����/RP����wƳ��MAT�x�У���p��՗�g�y8n�
����A �<�2%A(3�I�`�@||0(3d�;�CV����o(G�R�<�8}��m��w����VH���	U��`�T�.��Y2���:h�\����t��`�|��� V`U�zc�P5��t �`�)�	��qp/�ݺ�9*t��+#�t�Qڌ�̤c�wŢ%uP1�;�(�a��7/����]>�`�+��{��bbH�YE"X&��Q;~N��H4*>���(�������'��d�[?Q�i�<!ҥɪ��S�$5�����C���JX�mSJݧ�u%�Y����/t��P� �w��ا�M�5�>
�K�^P�H��֑�:d	��koc$61w�JڤJ�U��@��F=���9n�Dt
N�t7,���K�\�oo3�B�o�qh���7�\j��f�cbf䋏࢕[��zf�}�����S��W`6=>a��߅�P{B�f�'���G�
��*�����i;-��w���x_�i�td���P�*#6uQ�{a�9�X..��da{�ׯ_e�Z�
�Õ����bM��j�Y�Iy0J�<ѽ�@=wiT9�7�m�ތHZi�����h|%3Dm9`��ۯ�7UL j�΄�ǳ����؉Ja�ކ?���@]D#���R���e��QOӾ����GN�	��:d3`Wr1�#,��D9�Prp�J�?�&�c0.�hl,�s1c��:������|ތlto����g��#��ޟ+3ػ*���dn�K�2D��lclӮs��%��x:#"��@�~*��8�}^;�z+�GB���>Js��R�1�'�a6�Z����� 1�h	`$�l�5w�F��2L¸�H�Aɝ���)c+�A�d	ކ�C�����(���M:܌�0�M���bc7taS��V��F���x��Jer3���eOnH����k��F��Q�_o߹y��}���Cf����1|�2o,���URʤ+�uT�+��
��ߩRj��A�>�uϘ@��b�d�+�`�?]^K�7ES�ƗF`�
3��X2$�X�zm,J�x{�kr��U�'���O)=^b2�J �j���$�朂�9����[�?����R���?��,����?�}��r���~��ÇwEN�N塔g�2�q����G�:��w%8������ݮt=[�)�y[N9��
��nJ�r;�^jipҘ��*��hl3���bs4S�p��a\.�)!�|gk���ϩ�Ȭ�i�tr�
Ϝ�H�MP������ܘ�x� @����4l�T�U����r,����ʝùS�0�e�.U-j�&`�e>�4$ 6�����zUuAG
��R�HłO�3)��Q>Äj߽�s�t��o�\�M���V�L��M����S�\sy6)�,'d�0�k���S�*l��U��R��ۘF��?�3��e����%��/^<~������G��ц�'�R��cn���;C#��T.���|磏?y��1'�ȃ<{��ᗏ�q�Iem�����0��z�T���`/�$�M�G'���.�ݧZ&V~��|��'r}௯\%�l��X��Ϗ~�#Y�>��Ns%�`0kn�O��8ٻD�2��<�J���ʉ��\�j��+�u�d�3]ߪݸqC�F/r���� �"� 麠�׍l��]}pueU�=y~ҧO�ʒ^h_f��'���Fw��+7�l��T��'��X�̩Xc/6�����$B"&���.u�����	l�G���<�hT.�
���B���i~N-�D練ʶV$���A���,6�nV���# h�,@W��v��,����ZΠ|?+�x �4��
-��#�R+�
3�r�G'�D�D�����ʔ:�����/S-l�l��xf�l�,S�魡G�(i+�$�[(�y�Z���4�;!��66b�M���Y]�!�_+����?�ͧ���=��DC��0)9EI�3v�eγ�y���ϐ�#�����m�����1m�٩��Kb�W���Qڱ]Qa2�9�P4q�h��k{{��ݕڣkq���d�g~j2e���h胤�|./���w����f
��zL�����6��3��[�z�E��({y���۷�v:Jid�C�ݼyS���9������ʹ(�
<��*�1����3���T򈯏�?`,�
��UX���?h��#�0-}�-���<���(/$j*�@�5�^)���dz�����ޓ_�l���q��&O9D2&�d"+�X�_%���۠�u�Z� HLcSI�5�$;;3=���P�䖩3QO&c��oK�P B�����;�i�-��!�)ǠR�9jŇ����9�ΐ�*1=��Y?�K�z\Uׁ����E����5�6-o�zu7]��H܇I��x:�%���� ?��k�A�-c6w��ѵ2�
!ejZ���JM#P�� ��S�R-Z������|{�ER��7��>eZ����
�T��S���3_�x�.��=i�Q�_�;�Y��;��Tٓ�ݲ�T���T����Y.��C�1�I��}
����^�}���]n=i.����%����O��tvz!;�!q���c�U�ٚy
&��a;,b�T��v��G��N��r�m�Y}��A��	�o��y?����޹��/�kp��Q�=�s��-K�`X��B7�3����y��K�n�3�PAfJ��i$h��V���#���D�c(��*
+ЊS�=�aSm�7R#��[���"�<	���Ƚo(�$:HDc|
��W�N[ū2d��3kC˔Y�6X%f���-m�hR���j-
#D܌����S��da)��Be�\hJ+�V1�e� h�}��ˮIhP(.����nnM��%�D��_�xv|���WP7uGJ�MH��+�<��MU�a�Qk�̑qS`k0J��ǣi�5��5���̸)]%��*=��*X��'��.��b��N�>�����K���E	#j��!3f:��G�Դ�h}���wR�{�ԗ$��u���0t<�*56���"���
h/k	!1�H_$Q�}�$(7)�E�|zr*Z��bg8Ym��t�&��"b2�n���;�S���ޕ�7�_0+��%�w��_����o�p�v�|��b>���R�\,V���Id�\ ��_�����7�\�]���4�|o^�#˖�1��	��e��`�#ug���b-�sR��)�AK}�X��x���د�u�����ꦫ��Zw�۩�
c�n�8�x���ծ7hbBbO�Mf��-���^�c�%(PI�=���C�r�By��٣G��7/�O%*��z�:��7^�Y�1[����y6zc4��ӫE��r�u:�I̽m\���+�����o��Z��]�|��7�{�;�n�k_S�%����>k���w��|�Y<������/�u�j^a~aYP&6����H������7�z�#���O/�����z�����Y������W�Z��=���j������7�!�)n��BeF�^h���9\�=���uG����#�d��(Q�Q�Kh&QB���#'M�\��A�%�8�-��DG�#��#��^sb�Ț�zpenhP �f��π�F�[[ξ�F��"���CE!�q�|���Y0�|��ZʗN���:N.��0$s�ĨX��zFmmS!�I��*%��IG"T&I��&'G$�ٳrܦ tDl�zh����
8gy��@E��*J��،ꥷA1���z)����Y9�����"�^�rxp�G[ ޣ|�<���ɫ���������t2�%�NF�#�8�ˤ:���ܹ��o~�������?��C�y/�=�v��,_*ǐE�W�.���c_z~qI�#�i�S�N�奘%�(�x���rY��^�7���|���ӟ�����k"Ͻ2B�iY5���8bN$����	�_�|��I3ݩKn��`�MR�e5��N��<y��-���|լ[	��VW�����!YIr�Q%�%綌	�%�ڙ�V���}�1ae��O���_�_���zkw��m�n;�8�O�|��'���s(V����t<��f��`��8��udѮ\�"�$�ytr��]�|!O#�(�|�������g���<:~�䩜�������D�"2� ��>).}��ŋW���нzLm�B�,ौG���T,���O*��:��\qQ0�Z%��B9�C������w�ygk� T]���������;����eG���B4�<��'��&W�]���vE��;e��!f6P|:���#��R.Bd�N
�m#^���DI�X޳\Ħ��3f ���������U[����j�`�́�SQZ��D��it����>�?�t�)���uʼ�!S�r,:�����:kՆL�#�cVs��Jm�R���@׷Q��s	�8L�L�,uP\|Xgj�ZLV���lZ��d<���t4Z�"頭�mO�o�����]�a�3u�#� D������cDm��V���A{�!����ba�7�J}��l[��.��IxV�]o���^�O�l ���n̏�v�Vq;�6���|���;	:�B��i���g0C����ܺu��z���5Q�L��D����y"9�צ����g5���)Ť�2Y�Mz'� 6�9"�ZY�Km!Yi�h����Gr�/^|VZ�v��4�4K)�3˨��n���gR���r댉)0�_%>ҵ+<T��7�3�������J1��j��z"<;������w��l:�0ZfړĞ���+ ���ΰ�M��Q�cn�Z�3hY�N3��&��n��U�	�c3ǻuT����,�/��Iݨ������<2�	�*��<I��=��0h�}I�gB����t��sp��0%�B7.�+WF��ԔG��S���)����%3;�=�M������s^��.��w{Ey��� ����;��T�ľ\i�8W�|OlEԼ{N�ϼ�[�W%��Y �VE/����4@zۀ�/Rs��."�[.uM��Iꙝ'�+���y�L��}��իW�"r̓1 �����`u�7�P��`�c���*yE��<�s�H�h�`�K�OG���x��gC���nn�+6�hX���p����~B]���rȘ���T��^
k�2����ߌF%cW�:��J�̝�'
c	|b�b	��x�2Y�,�I&E:���|@̕w:ke{{�X����\��趕x�:��,g��W��c�e���^X������)Ոl������3�N0��n���M��g��r��U��=�#��WJ�ř��J��4	T�tf��x������A}e�y!X��|.��
��I1�4B"��Cǧ�E4�װ+)�BK�B��2��q%�y��a��V�Wi�k�ϵ�E(CРA�k]�t\����_����va��XBY�k׮�؁6o�mLvP3������&��F���f[������(Bd!�'o?���E�Ư9�k�~�/.�3��^+�I���ط������æ�h���2�1��)�GGG�eM�9�?��[d{��b�6�2�QQL�>f{�"a���V�GCɄ�OP7�˷5i\�XK����T�Z�Z�zg��Y���]�����(��[L�=aG�[��Ϊ�F_4��ƨ$Med���)vy��b��6�O5n�2�C�0��8�1�U]�R��6��V�2N������ҏ'�8��?�B+������DEQ�o�y���~[�y�o������N��"�����~�ce�ab�ɱ�����͛7�:��{����L��|�����o%c�tkAL/ڣ(���kr��'?[�֍>�e(�x�My�{��ݾ}{��+w��_��?�����Nk썁G*W���^:�t��d�1\���3ԙQ��:�����:y�;MC���՜��|�+p������d�h��_��JP&&�ƍ��冃����+�VA<��f쩶�%׺^�i��߹sS�O�@�)�V
)�<�����4"S�c�\�T�r��''"໻c�[�`~�H�����g/N�5���AI��N��x6!���]?�G}�(5�;wd[?X����Z.�Q���I�2h~M�3W�<����J/�z�H)Ps�4S�:�)./�ޥs$zUn�xO>º^b<�W�nZO��������Ӄ���^t�5	a�:�����h�/�h�{�߿/+ ��G}$���oM�ym����h���)ACF8�܉��G�G^{�G?����ݏ��H!�5O��\(�����4�t�B�c�!�4nq޳,������}�P!�)�V�Ud��˥�!C�j^�`|Q,�>�z�ۄe�$먴��[�_|�ŝ[�eaoFL�R}Q���Un����hԈ�<==���~��<��b�����&6b��ޅ�|��[��*ԧ`"CX��I�yH�M%����}0H�.k�*UB�nu��ܘھ�U�;�J6�o��vN�Ҙ���Ĕ�ÂGm^!Uq���|�;����y�����g?���F��#��K4}OwfhPV�Q=�R(�L�p2��<�� oO��ǣ-�L�¨�i��S��#R5��r�ܴ��~"� w�,z��w?{��T��NǦ;���*�j����,i�`I%�a��y�!H_�KĴ5s�r��s§��~���R�J�ҭ�H:������4!yn�QR �su$�d��ch��*�FE���l CHY�� ����EaӚ�.��s��Ȕ?4�i7���d\�0���7���opy�����ά3�����I�U���m��]��"���_�[Wt|j�,���90�n��[>a�JU�↕�^KyEٯW��.�k����0�4�2���0kJ8�����#�!�'��r����Et~t�����G��SԘIy
���re�c4Rh�?�Uie���+kxO���X�M��϶T���K��55ķi4�}�O!#�J`z%3�I1?Oy�Jm��6J�_]7=�JLx筶��Ԝ��[m�
���4K��͖CX�,,�~{�'�Y P�3��d�ep3�����}c�j�)R),3ޮ��1S����ۢb��0�ͪ*/r&��$2i�A�q�*�l�]�8�`�rN��<Z������5$vn�g��6�5tj=��o���hT��4�{,3E�[V�*�WY���{
�؋Ɔ�t���ݓ��s�Su�!��Q_CŬ�}̘��V)�D/����FYK2#���(l��f�5P���5�6���t�\c9�'�'._%�+�VYٔ��{b�5���J�P1��C���!�<-�f�����G�W�-�_� ��s�Y+qÆ�%b�X��3��O������M�,�Z��[��4�"�'��QW��"��梍���R1n���e�4h��%$�؃��+Iٔ�+W�{�Rt+��?%ߵ�4ÓY�R]Y�\�:��эKe�L�(��rE�l<����F	{�3~'�Hl�X،��T���L��I:�%f�;?���Ϟ�������MA�2��a��Le�I�y�x6_��.Qf��r��]^P�������6�DJ$�{���A{�/��Z4����%�(�������8#pT����ɳ�D�p�������R������6o�~�����\��HD*�%��[��
�Ͻ|�RT;�Z9�[n �$_�t�D�W]�"���8�ԤK>)s%�եno[-���	>�F�@�H�=\Qg����g��n� z֒b/�&QQ���w�������GdAZ뫕璓%of1�,Hm�@2&��=IY��R�i �<��a�o4�^�}GR����Y��ӓs_�����"��g�pdk$�UѦiE�8���Xɵ��tԵ�)Ve��G�Df�w�Vݑ�
&I�رK3ԗ����`SL`���oP2�p=����)�T�S�QN�m���"/G�c^���f����1gbE~y��0��y�
SK�~Y�,��a�LGu3�OT�2$��s�\���=����<c�/..�=C�d�����rĵ�u�{)�,�6C�[��G���f����lo��vԥa�G������#�����[ʖ�,����kw�%8a��4g������S�g�w�U�*�����r6�^���Jb�����Z����-��;������޽;rϚ�<kl���������������� �$
���,�<�`ܝ��3�c���jtM�����w�&Q�mm���������oݺA%�\�@h3�Y���/b���k�Y7��|��"-�nݑ������JA��9�v)n�ӧO�y<x�\]��O>�D�'S�R��ғȭ�����\��_�������[ځ>���������_����܌\_��=1�"c����D:���e��Ϗ䚲��-���8ݧ��ߖ����U=�����o�
p���}��w����<?~,?������%O�_�RV�ƍr�"��tO�>ut��Uљ�^�qSV��O�}�v��D�9�����V�Y�Gh,�\��-�sy�웈�|�>I��=�g��ᣇr',�NǓ��9܈�]���f�P���D<}�\��1d����ջw��\�KMc�	u����d5~��Vg����sZ34�\�q��͛ar�V�\=p�Uܖ�<�{�������׾��|���?}_�E6]�!{��ycю~BO�Ө�|0��Ղ�(H���$�9ةF�O�j����'4\k�NT�d����Ǭ	!�W�(���]&��ܹۦ^b�l4���}=aޗx��Hܺݺ�����8CQ�˥8se��-9&��6oڣ����/>�����V%���g�5UVk�IݬSQV���6�۳�2/��]��o��M�y�5�Z��-��C���������:��^;M'����7�����D�܀��'�Ӣ���>�>�z����"7��,��G��LG@�GX��������v&AM�bèB���ř�Z�:�]�պ��_�:zqt��M��e�-�K�Dg�Q"M�8aZjC����Y;�%�h�x�y��M�n�f��G��b�Q�1Y��
���2�u'��b�"
Kr�/I�R%�u`�ՓzjR�oo�u����@Bx��U�p���51�W͊���8���:پL�M+%beUE� v:�a3�HGg�P�Fr�zq�^ɘ%���GL��-����}Q -�=Y_�[)�W����Q]�u�YUw��(Ԫ�1�d�A�Q�$�|�V���R���'�9�"d.Z�n�+�5��A�4�F�^� �.�R1�oM�����A���?̫|�E)�]�H���H�u�Hc��Z̶��)�N�	���h��O���S���L��^?�q��Q?}�:��1X��}��8���u:��;����*�g��.ⴢOSq>����|�(����v���i����la#�.5V�	���<Q���%�~�727��ގ�&����B
	H`�oUT7��*���i�F.U���-��ᎠI9�@N�-�� 9p��l �뭋��;׶�����n�`�}��ƹ9l�� %>H�a��3���h��e^��`޿��h5:7Ϯz�����o�����K��m֨O���t����S�jw,��m�>��B�)��G�SDt���;�|M�DT��8W*{�k�pO�|5�h�yEl��~���JU��8�f��FBS���3��T���/��9M����k!>
���XJGR���-�5Oc*�!˹yhYB�6��\(����r���\���Sa �(Hܵ�K��U��_�(��u"�E]�N|@��iL�H���<-�	���kH(�tE��F��Z���چj���O���Ŕ�{J�ܼ�.��*xy�N,�BL��څ���W������
p�jt O��Q%�y9]䜘ԫMVyè�(%�2�ɸ:�n܆�9�X�H뵙f��3Xn�++��L�q";���K�i�fj^�����/ � ��)�\'zs$�Kx��H��h����g���\\ ��iM�������K1MBt�����!H'�y�x�p���N+�SFښ=����/B���mf���H$�F:��U���O�e�E^��k%w���N"�;4��	�I�,�Ub��~�/���7�~�]A2Y��AԱxJ���u"T�]����@�����1�\j/xb�0O��tR$��`d�x䚤8!��0����I��km�~Ҡ=�X�q"6�G�I��|-�I�����Çs��S𜑊�;?@��Ћʬ����RifV5��ԭX��8Q0ߍYW�jp�c*�d���,�mqo��<�6��^���|���D�wk(���FX�6$��n�Il=w��`�uV����N���N�DH�\��2 ��\��چ����8`�����,�&* }�)�\.i5|����ܨ�9:�2Bj!;N
W�"�̘����V�3����p�I��X�6�5����˥~���~��O��G�������t�������۷�a�X�SZ"ē���o}�[�����_}��(�i�m\cTk��	����B�Jƙ8J���<�"�Kn������~�G��!�ItgЀV
�K��A����{5Ls����LxTY(T�\�K� J`Z�X��{~��w4��>�u�|���c��)k"�䙭������6��1;��u��\JNa���Ԋ?����(��M��>��s�q~�:M:J��ؒ|뭷Dcܾ{_�.4����=9�T2�`��ea�Jٻw����2*�v�s�Ĵ�+�u)W������Lϳ�5���LI�-9P���t���6-]�WNpbi��dih�7�����{O�<P�49y����8G�˭'\!l�a
N>C���'�?��o~#�
v����=Yj�w�}����I������s ǫM��ɗ���]��R��"%��W���,�]�N2�7���?W:ѫ$ ���DP��ɕy�7tI�v�q���  �x��C��M�j/�I����&g�e0<]^�R%��4���o>��S���W��SD�����O��$$ͣ}9�L��l��^�F\�S��ìܕ�G	6�&
�r"����9���I�����N�� e�e�vk�/��;�L&#�V9�h�X^�{6Ӈc�Ђ�ŉ:s\�`z� ����[�U#*1�@Z��$�����TU��v�i��\��ǻ�l�#_7j�,"���7�!Xnk8����M*'&Ҍ����������=�w_���z�S�BN.&��q�0�G��n��:��p�;k�K�o�d�"��,GC׽3@��e�i�Wi���}��z
c�,�W�=YiEc�,(*pӌ¬�N�W�`�q Nv�4)�~��:� �3�5�����z`[p�6{[�����nqx煁���R���~B2�`���[����H�I&�ͼ
�����R�DQd�t��7��\���S%�s_�x�m�=N�A�h xm:xYY	�0S1��8u��|�,Os��Q�@]�<�}�'䘒���g|U8}3��H'	�{�VU���w��B|�E�����eI8:�Ϣ]}AE{`Z�����/�[&h�4p#zfm�v=:�Gu�5� �W*�r{(m�fZ�i�b��hN̏����UY�Ymp��L�U�Fc9�y5j!��7ɫ�h������� ��.��(���J��9L�-��L<��%"��Cs�aA1Sb�\!jU[�6���S';�i�@�@�g��8��'
9B�+�`5�<ƭƶ��UͭEf�EMl���l�VC54-m�A��W�[�VZ)lć��O��.=E?��ޡp�
�� ���q荛�P0��x���s	Z��̺zo�_tuL����ٌ�s�]�S�����J���t���|��N�����qٲMYoq��|�kj�a0O�,�u]��Z5����8�6�l��E*,����`8p�	���:!O���k��5��:"�Ezš/\�C���;�q!������jKc�u�I�]��`i��h�T3%��ǀ��΂O�����J��t�y9���x|���q�Q��[��ٕ���~{��xJɗ�Z��B~��=Y�Mf1dIEr��>�2O����c��x����]�)��6���s���OJf5Fg0O��E��3M̎f��,{zĊ�	�WE_�J���Zk�~i��_�w�]�����Iߨ���w����ѓ�/&c$��<�����Yk%���H�y���u��O�k��M���@zzK~�|�����Ǘͺ>::���cg(��Xt:N*7F����,@#�#�2.��w�q5�������b�<Qc#�um7�M���M�<K��(a�Ra L�P����1��(afPbE����3ˬĕ+�١��J6>�w�1�x0�77��\т\C��^�:�-Aj�1��'J�Wn�ʕ+��33��_zj�5|}�j��x^(`��p�ڐ���uCaFמf�d݂��u�H���8���{����\l�=�1G2�dr�bU����]�Z�-=2��>��C�H/6�lÐ ]�aÖ[�꾷�k&Y��9g��rD|+�l�Z�:jPY����Z�b��<�J�u��t�A:�p͇��Y=;��7s
��t��S�a7a���ә�� w���7#^�ʉw[��O �Al�t&�y,x���KD�%�̤\
�"��1�a��l����L�A�ź�ı�58�nrk\,��b�W�����:�	�w{�ƺ�R��C�h/0�[��NOO&���7%�W��pf�/ʪe.,�&����t#���X2����zYg��nI*=�m���Y��
�
�;?�r ۹f#�0�P�����o �9`�'�kN^/�I�h��b�n@` f�߫�jsg<�]>���p�#���:�i'9��=��I(H�HOw5kf2>�~���*���3��?z����.�!���oD�6��u�DA4&���JN*YfO�B�T�dR��?�������{�o���;%�KB���+��t��̀�^��X.�g6��sC�>a(!���lr�<�P�>|���0��fFo;�}��ڈ3`����.��΃�;�����G���/�����7 ���$m��G�`d�E{���d����"_ȫ��ԹI6��w�ܡ{8<<�JW/O))z�*�[GMQfг�={�I%,,��u�Q���`�vN��[�6.ۗQ�H�Jo{+Z��iJ*��w~v��J�
G9����^a��5�RY�v��F"�H,����<}M�t$6�� I��Hrpp@�\���������?ȳ ��B�O��ָ4��!q��a�o6�H�����޼y��ū/���D��HU��g>[��E��A�l���\�*@A��8&���I�� 渗�!W2~iE�����b�?܆�R��"{�6y���j�A����to<h�ί޾��`��b:yp����~����v>iW7�w�� ����^M(t��5��t -ou}��E�-�K:��ҡ5��M�Cq9a���3�T�:}��bf����w�ޅ_��Fł�������OisA�A���uY	jf9f��'ٸ���}pwc{�7oI~nn�Io�S�����<VnU�i'�2��!��3Jc��@�@�j�tE,���5N�D(7���� y<_�Y�@�U���~�K-5�Zk	j�V��E-�V	_��F�2�˪���N4	E;��=,+dV]KiAt����yP<���v�?�B2I��Q���-���Z-��8��4�����R�"���pBBF���"�k�/i֓{�{���naX�m�+t2�A�dbXqbS���1T�i'e�jy����g�`���	't�#� V���m�eZ���ڈ�j�����I0�� m��/�`�x�17qڃ
�<�F�
�.'��ue����1���u��]���m{%l��b��9��N�6t
�Ffߵ�P�i{Ұ|gB����|��(k��	cKζ�	�$I��6A&Ł2�E��!�(��'��;pu��O	9���|6�{�6?3*�f�<�u/�W$�$�.N�h̟���p����4u�/WD���+�+DZ⥜�9��0��{M�Oן�X¶�6ę^Rl�
3�H;%x�S�v`�Pc�2��Ngi�z_�S�l;���������x�H>ӆ����M3��X����^K�q�j�T�E�H�E�q��fri�]W� ����c���zr�Q�0^!�f�T�+K"x%(��2b����q�C�2��&��PWG@����P�N�",K-�|.�`NDY�Uq��N��	��aЬ�ޗE&�yX��PS��Q_]�_��-���t���i^�O]�9�<x����b.%AS��%2z��IQ���@�������]�p]�`��G#��Z��>��dҒe%��u�j��p:`�+L$��e��T����P�W�x%1?���Oq��Z�&´@>�z���]1�I�!\@\2t��L��"]]b��D�dLP-y�k��/���#��Ǒ�I�C�G�� ��K�����K{��Q^�.�Y���q�i'! �"W�kD_f��Ԇ�9�:�|\+�vX�8�`����0x�ੑ���C5>��*��С9��B:��6ȃG�t~v��{���0q�`g�ʚ� O��,�ɂ'y���$6+� ��������rI�M�Wy-5Q$Fo w������K|�#@��8�{���,Q �%ː�A:�R
�%�@�RFQE��e�4�J)��J1lk0ni/��ܧ���d�Q�r%?2@�Ң�.�(����d֡��rX�^#���m��`�9�3 �0K�yH�ݻ��M`��p9az �#gZW%�7*kp���V���@�WJR�%2;b����-Y$A��C�Հz���ͫC��B��B�0�Ny�#��~H0�`	��fpj�.G#�`�#a�cзXd!oȋs�¬D�
ӆ/E�'Y�&���j�PNz���8��4�/O�yNh=�4�j�� !YED$��բEs��<X
���w�/�f �̣���"��7���A<z��jAQ@T�&��ͼPVrӥ��6TS�l��D�D����[�5�=�	�$�0�����+��A��u��i�ѧ������0�?5�;�-�\�Oh�ٻ��豟��<r���yj��,����JY}s��5J1	E{}R�Xf�Nq����C6)NFW�S� �j�*����4g|�O,�Bg�4�9�"l1pj���+K#	-g�"S����q8� \l^A�A�A�:h*:>�`@2���ߣZiw��F0�	�/2%������{48Ϯ�&�$�D�&��끳hJEj���>��[�3%#n���rQ����k(U�#��n*0���&FV�#��-@�>˄�R��ڝ�t�X[`�?�S�ӝ�{�uF�.]����?�cN���]@���:˱Tn%���Vk!��E�3BW�ݙM�@*A��3J\6�@�U"i_Φ�Ǒ�&��V�g?��fw�Ƌ���S�A�L�'�d3o�آ&�`�|�<��bS%O����Y�V�B5�,E��썍>��I�-j�THc��#��8����$��g�g�7衮�%V�$�&�x�b{��Ǒ �?��g��L\����q�^b� yA7�	����s��m�0Wqj���!]�v$��v�/��q�ۆ�q�4���Q9p�+�(����J�RDI+ttD�K��,ߠ���uyNW��PD��Z�豃-	ON50~Eҵ�6��s��˚���񕠢�UCǣ-�w�~���b���a�;��~�B�K�MΤgf�K�.Ɲ�4�=���r�vP��cpi�W��Y��J�G��\h�&D�",2�b�0�=�40�ȣG���}@J����u�����e��R�1d^�*�2)gZ����K-8J�}�����5Lwó'�	~g�ξڴ}��c��X�cľY��ݲ# ��L�
u@޾}�s�M19i	���&�VE�X����xn���5o�
��2D�(���N���Kޅ�Uui�
���L���Ef�$Q������.�:C,AiK*���|UҶ.�%��Y�؋�_���/J<u�20�/ݐǰ�O���#�E�hN�O8_��t��"(�z�B�RF�9�>��"|�Eo{c�gfb�Ib��rUg<���9XM������l�㮘 �@k�g�9W�����1���XWg�oZ�A�͔��\���v����e����+R�)�a1"�%�^-8��yb	�j�`��fCСJF4�z¬��l���BY�,kഓ�\%VY��κY%�5]qF�1^��5�G��E6��8�>5-Y@���/���$OQ@SCb������l�y$��L�qGȑ(��ڎ�KW���&/�?��
���1'BA��r����ߙ��fޮ�_8Q����mW���\[n�$u�%I�rB5�(��JXl�����F2	q��Y�`�[߄$ ��O�~o��ɞ����2
���Ɨ�A�-۾q=��zk5�����N�,B�T6�hs���"� y����L1I痮é�r��vv=��d'�l{|�I�~{��2C1�)�W�����������t.È� ��%u�Pc
4|*�IM��V$YENG���M27
��|�U�l7�[e�+ÉY��hJ�1wS+�E�+8�a�:����i�e]�z�;|�|��V�w�aʸ])��{(�~�,�U�!�|�Vi�	9G�N{��/��<�dM�,G7k����4��I�'�Sr�Q�G"�)kf���(˖o��<���ŭ���|�=}!G[�x�'y�鞞\2�)d�LQa�Kt�Gt��g��F�T��/*��}���tf<ݎk��y.KQ�USE�Z�rN!uiUV{��A�Vs蟽�x:_��6�᪪�|��!���V�B����}M2:x� Ѹii��XK�����9}�noo�V��Z汲L޸ɜ�iޣe0d���룓���0�����+�lJM}�B>��D*�m�e|Z$�T�+B�5m�h1��
f*iZ_-��z) ��tZ^ON����R�&K�O��L�.E��j�`��{��!��/�߼�Χ쯬(PL�ټc�C�:+H-6�8�9��+(\5	�.'��tѢ54dJΨ�fɭ<��K�A^.�Ր�OI� �"�
6,S��(4�9��V�%���O�%2�(����١���)���?wwn�d���y�[�;yvT� ��JO�%���d@�Z ��<���1	�l>�m�v��Ndx� +��=�Ӌ�U-	 ��'<s:A�ܒ�Z������i��	2#u�:����g�e�\*O,��6�]�gm���eY��!�E�L�Lk�+�����X.��^�b��۩g��L(V�P��h�]Dp��F��7A������/� d1�������{�Z鰖�5�Ʈ�B�n���:~{��l�+2�A��XP'��*�_?��Z�3G��V즔U��(%�ōN�0,���Q�2��a���.i�U� ��i���Z�����l���)��	fI��q]m1�z1���>|8b�8m٪���ђ�mnnW�$�����4���Kඤ,0KJBھ��0�<G鄠��2A.U�v����x�	�y�,%hb������\��������Ϟ�E��E*���t2YU<m��Bʴ�a�5���Cf���������hY���<``��:�G���gqrF~��7O�j�֞L��T�k˄t�̄��ۃ��|��m�X�p�Ke�i�9:K}-N,�?����9�_i�"�g������)M[���V9�r6pc����>.\�,@<�,a��,�J~Ѫ�V�4�a����ɗJ�u�ԑy�IJ���˶h���ʅ��rU����R��p6}"�y�d��&i�^ξ�Tt6-�T,d�:����ZL�;b;
R<��Q<���Hy6�'Ӱ����7v�t����ΨJ���=zm��?�A���]($2��@r
?d]��̋s3d7�!�G�.�6��M`�S�!�0�6�჻?z򃯿��-c4�%�uZ&O���>��;Rn%���c��tM����������v8P�9�ʆMF��75�P?��	����~�+�U�ׯ�%��Ĵ�uMF��O>����ʓ����?'	���rN��j���Í>�C�t�+f�E�nD��A���b�|�5ٸf�&5�^�e: e���Jٜ�����޽��������{��|�}���t�O�>=::�M���w}zF�zN�p>�N���߹3]LI3�>��������={6�0���J����sZ�U�^E�@����#���Ŵ��U媦��#�@
8L���늬������$;�q��{�>�3Q,EV�m�F����?�����Oo�)�Xno��W��>c�*��뫊�y�/|�������������?m~��nz�h��1L9�?f��14��dI�^�zEq���?�<y|r�䀳��ں_d˩[��tR�M�������[o<��z<L����o�<`견$�H���03���YN�u�&�퓋��<�����bNj�����z�hV��d�L���YJ�)Qu+�-߂��r�>���X-f�^<O�A� ͖c���)U��V�U�����K�i?#�4��%'J��*{y��-�rE߼���r
�k�M��h�� P�B�'�I�VsEԉ(Uj�3�Σ����k�[��.Ws�$�	�(��H������(�����$�=/����?$E1�޽w��e���"bS��|���0��
��#��Zƙ�nƃ^3`���AH(؈�,� ���nx[a�e���H���+�c�r����J�&�,����s@^-�c2/��I���	=���W�t�&�x��^�y��a�"��d��@6rqI�`��Ȭ��Pp_T8y��B�ؑ5��4�fnI=v�0�tN��N׳UI~*	�V��
�"�Vo�ꘅ���Ɂ��u;Z����a�pV��g8+ �ry�r!Y�^�1d��}5]6�z9Y:�ƽۮg�ً�K����NwB�&����<х��������3X�?��Ql2�Nf�͖KI��B銜W<.�U,, �a-#'�shnds^��z��U�).����j�i��_��A_4X�Y}��3+/;mP�jh�e9]��!��P��`���D��
�������q�`�2�x_	���.�¾3���!���} /�`��\��c���2����>R�4O�"$�F4�N�m-�e��"�BЧ�,�vG�äC�	Sx&d���a�9W�Z��6(�К{��Nq[�J��il�F�d4h<15�{�[��_{y��� ���MF�^��ǁ߀�Ȗ7e��H��g�jI����hK��"y0������#�֋�ON	��+J�#׵��$.˘ЕA�9��Rc�	uaą�;�h�H��ۿ;�k�&�YfÙ�O?���z~xxHQ���m2�p7�ʧ8��Q^���	?�l"��r�¡���gb�:(5�1)@����bط|�CCT!/x���9C���d�x}67���uy=C����z8�Li���2�Q�A��g?* ٦V��#�����ا�)�#��i�L$pK8,����"�<9ZA�/A;�!�Y����M��f f��*�'����><�{��������GZ������ސ�IT5�R�B���H��.ө�^�YəV|��:��c�������Ѕ�(����c�W4�߿������#�:�R�^@[r�����:J�SF�Q�]��'?����׿^I�$-��6c7��FB�Nb�r��l�S��m�cX�Ւ���JW#��<΄i���w2N�u���Z����-]
�}��^�ː|���-<8���Y��hAF\_F�6��٬&  ��{�(�C7:�_��[it�^Fu�f"�P�`%�7L%
�A��8�}�|��0��:��"�爪��4�j6�(Hߚ����9mڢ!<{{{�/��P03���_P钪��6
�o��+�
O�XI�[P�,@�xә���T����&�;g�����TW��Ԩ��~��1���_#ƅ=�8�a��"ѿL�8��ԖV�D����+qy��I��-��9�z�	Δ������ss�wn�d�.���|��7������Jq��K�))ϲ#�.�
����͛7�,,]�����?������\�M�G.�s5�R�6� ��aa�i�ˊ�MDt��*N)E�I�E^y`�#Жɀ����U�)���#��ǡ��������ׯ�fN��R�����s�D��v��	��d�D��운µ���RJJ܋�#�-i.l�y�?��73�2r' ��S���j/�dֱMmRI�V\�*��J����_V��[<��u��Vs*q}�o �Ř�\Ir������_��k�����T��&�P� �BH�FH� Q�J#Ka^s|�界 �s�}�t��L�G�y���9$�l����7�^�����k�[��z�X�kɼ�)X�� ��K:�w�r5�\^]�}��Wϟ�4v�w�ҡ[py��a�>���ty�ػI�p���{��ѥ�r�s�-sQ�M,ez*BcA`e�P�d� yR ��Í������f�U�N���(�7n�1�\�p��	�(�����}�r˼�9z�>x�1}�?��p�M$��wE�E����{�G7�჏�������G�WF�lb� ��	'�Ƞ<}�����K������w�Qv��	OXN��
��˺��ۑ�������+&�0���� ���j�5��)�22N�Ǚ�6ԥR!W�F���<Ө��@�o�&Μ�@&録��ԏ-���Ɣ%�M�'RHg:@�Uξ�Cu" K������)�>������g3\9@�x?��hx�^8 Y�=UȰ����PY��t"Hf0�	c��I,AhХ�â-ep�Q��gp��P�_�s%
���.y�Xy{S�qM�N�V[	S�0�J`ͳC�����:� j_X��$ ܜ�����#�����!1W�IF��D��T�]ɡ��w2%*u���Rr��I�\��t m�Jy��'��D�iL��U��Va�&K�x��{ox��З}�]�u:�ڈ+7ҏU�����;d*J���'���T|�M�����f��+���>��; N�rR�NB���w�gMb�*��{ɳ�7�_�̥ur*bpk/��<�sH;�֦�ч�
H���R$LeҺ4�|�.� �g��Sn,L\ū�iNc���m@�* :®�:���������{u`wb�c�9c�ɠ���o����%���U!�`bm�JB$�ۼ&�l��:�k��Sh��׌(V�	'�n
�i_O�ԥκN�aP���f`�ɸ�3�z<�^�>'���~��
��d�+��3�\E�݅J�:�^�2�"0�St�T��2�h�f��w���À�&cK���ey�tW��6rs�w��#��_w�x��۷����<+���N�*�ꧻ���2���������J�Z�][M">�J/cD�Ce,!�"u�Մ������G�&0�])·�}���4����e�Vt�&��p�4�.�-v�K$���%�$r"IX|L��Y����ΪƎ�d�!���W	E$/eZb �Ih{���'���zNk��TH��d�41Iɺb3��;�<�_�H���ڀ��\��v�õ�@-���K#8*�Z [�Q�Ig2c� :d�:� ��9�]f��&�3%I���_Sx	�>z�<�ʆ����{����w_9IU�W���v.���)��7�S�J����&��
�+�f�,]Ve3�v��^�J�r��������$��|�^�x� ����Ϊ��?���?=z��/��+%>#!Uw-vJ��b���y����~�O��O�����x�����k�͂Ovy9�]0(��~��G.n�����?��?!'鷿�-Ȱ��mπ�C���
���B	 l+�\�����%W�u%�D]�6M��h�����eV6_.W�,&IL���J�@',sd�z8�����A��i<2�yH#-ݸ)L�G�{#y�������۷���-�~8�JG�f�amP��)2�����"�����K\�A#�HS���կ_��T�D�c�2zm�ϴ�a6��R��8v���T�qؑ�>zdp\Ǝu-�DwK�q������xs�񤐇��q���E$������� ٺ����?x�w}=j�%��]+����IJ�a�dI
=	FH:��mŔ�LSà�\JG�7�K�H���b_-'ʫ2dy����ة�w(NT���@Q�u�4+%/v���]ڔ�����g	��/�X�w,�d^r�	���:>��Ri���lm�DKN�"��v�|���P|�ɏ Ͻ����q0�M&�A�����AEgq�}�!�h�9h�D�<�!���\�(���,�E�����.ں\B0Xo����z�Y�uڠ��W0�9��>��b�Ď�5��f�E��K�)q���ɼ��CHgI�֙j�:B�Z�H�,!�K�)7�GؐXb@4aW`�c|�]�U�"}������*�2)+����q�6��Fę��H��
+8U�q�P#8ԮYw���vE��JDpڹi���o���X9�,iy{�C�Έ��[�^AN�[$$�l�� |�io �)�g�?zDZ�͛7tSS��E9����'&����=�orr]|��j�_U\���o߾MFv>[�uEv.Ȉҭ��뷇gtK����br��x>��~�]�xq���|�����>��RBt�mr��7?�����7�^9O�$�b���&��t�%nw�5����8;(ҍ1Z��1c�9�wFnr�֧|в6�ǯ_���	]�.W�;�7��z�s6O~�$��/�Kr:x%n�!��'���������w�]��$IaSX36�B?��+9��nݢ����9=;&�x��9=��;�9�1~!/�Q����)d�F:�!�(S���h�SZ��XC�q�6���,�tj��t���l�ք,�����W��i*�	ૅ���,p3���]�)6��N6��L��YS�|���	��>HRޭG�7f\�m���j���¶�� M�s��RoC/5��6�[��=Ju�6?;��oC��7�`&���F�x�ۑw��3�D0+I��TQMXux��(�%��@��a_~��qx�|N+���wӦX7P�`�Zà)�ӦF�i��3�a쭓���/�%Q�Q��!���^5�%��	�㩪�r!Vҟư�,����D�,�v�(���� ~�J��i��PE�WOg��fBB��x���>i�ܰE:�/ꓚ������I3�b0�4�J^�R��
=!v�n��2�\g`8�2#k�[ü�������:['y��I�+x˭��>�O�b�J1e�MWggg���L�Z�٘��5G��D�a��ciD�<���S��|f��m�+ș���YdʌO���|�::����e���������w�Ă&e����׹�?����D�^]��:���	 '�"��4@�<�vK��6�1[�ͼ7��e2�1���lKo;E�HM�R�̛�V	Np7��=��<]�TDxC�,�g5K8v�s�3��,��2qgWPq�>��F�؊��T�b# i�ZƸFG��Bn�S�ÌD%��b���"��v\���Na2'�e�KBn��>�[���8+M��ՠ�(@���&����6�>�l�,��x	�%-�lJ,ն��[�0K&�t
�d�?g�¡|ztt����=�d��䣽I��L�i;sf��4[蔘� 9�c	�79%�2���!�`Ʌ�.�p�6"+N�x��k�S��-8���	S�3sn�S�r^����2t�N9R�k���{Dxs*�grR_�92����`;G[�2�D�*�ֳ*w녊+H.���k#���je)���K��Lάj�a��E�p�����ˋ�!��u1n�&��R+c��i5��:�vS�i$G�E6�<3�$xܧ���=зB�z��w9�0`ygxB�#Vq� �Ў�V��v���H�C�:��+�j�y��a�Y���%R�dV�$�#��S
N���s��ɔ2æ<x�<�B��������5�נZ��pA��L���3���BEPJ������ѣ����e�����oW�y1:��W8�h�����buj*vĐ5�O�|�_m�r<�[j=8�b�8-�AnU��a��>63
��#j�|e�24	֤��w�b�eA���'���ԠӺ�Z�8�on��QχC�ZA��& � M�B�\Z;d�X	֛{���t�re�6'W2l+�v-��^�(��y�l��)�H���.2egtF�ͥ�A$|dm�7�x*�����-Nk�q 2]�� �ۊ>qPぱo�7�H�(�H���3C�#�l%֢��ܸ���9h�s�w�e<˴Ca��2��V^c�b��ᨀ���l��x�VG��fB����6f����=<<�J���~F��駟>�},,Z�{�����5�Y�1�!Cq�OI�i�n߾������)c�L��#���7������64$d9t��i�X���G���h.��IP�]?�U?�Y��Ķ��̓trUI��Lh�0��e�R�K<|qq&�UJ�;Q0�&D��/�j�)j ��]�!�f���JN$v]`���-fv�4}v4�h5��s	���D���\n�����Uh��Y��3A���`��p����9�³!o��!�^!L��V!�a���!�'�_e��t�Wh^9����9�arͅ�ٌ?媥��<��5$�hUm�0Ѡ�K>�2մZD�*�|H�H5����G����}#P��ٔT���J�M� ,Z�Xd���L��Ӌ�ݽ{�s��~~���Y��jB3��D׼��],$�>Kf����}�`!uǺ��r:@�x�C�#���Ϟ=����9���5�f�A	=@������q,,W�� �_r�Y��y5pv�X2���2�1c��h8r��.]"�>N�'Bvy�����G/_�_AB�������o޼9x�0���?�d4�w2\ey�bd���ށv�믿����(�XZB���<�ɓ'����c��٬���^�g���/i�J���]������ܾu%p����o��ce��T)
0+i݇���&s w"�$�*�=�:�uh ;��:u�ه o+$��3�Op*&�k�:��±)r�$f��k�5�?`���9��F�8m%�u]8���<x�n�n�lJ���k ��F��%K�Ca�ރ݇Zƙ�s���ux!xI:�4�f>r�@���}�D���&�%��;F��F�,r7��a�J�b�f��T j{��e@\�=-��&D�wH�l�Q/L��͟��Y~�����ML�Z��iuގi��NÁ�%O�V��#����뾲��������v7B^�}�Z���2QA�]���\YF��^�dL��$XV2���Ҡ��'��M6�;x�g���`hh���C��Z���B��9�J��Q~G�	@F�8�1�� �X	M�F���I��z�&I@���Rdkc�/�T1���Fg��Z=��um��ɨWt��i���	��ԣ͔��uH%m�2aI�Ƞ-�мN��Da�8;�!h���qE�N���S]6T�{����B��T!�������[�3z:��U��?���H��1 6
ֽ�RAH�W8��DP�E�K��\��[)VH��&�W@jI�椏��T�(&���C0pJ���{�����ml�lkh�'s&��RC�i>�m�MDt��!um�&1]]�H�����c�}����`�;�pLӈ.v]��@-�h��K���AX���UUBA�n��x��á���߅��*����N��T5Z���{�;�����bB�Y����)���r��"̟(AlR&<�<M��Ox�5�#� �5�f��:�՝�Y��]��!q̣Ŷ��R��d�6��9I�V�L��P8�.��]��_TD�9GH|̤���=�DE�ִ�
S8"�����o޹Sre,���]����(��z�6�m�(����|��L����,��f�|��d��t�џ�G��\�������g�W��r��ٖ�? ���.��ս�P\:�t�@�p�*��K�UXY�^��H�0R���1����	�����T����Exqy-����N��|g�-����j�I@�@�N���$i�����}��w�A$*ju�����Ln5�-�'��6Y�.�l)"�>��߿�ӟ������s(v�Bh0qҪ�8�oP-��� <��L�
@��j��"5��O�@��#��؁���s��x�@�p/�H3��j��\� �I�z~~N���1��,�E��׬���J�����F�ʄ �p�{cC�6�8a������A�C���A��Cg:�}�6�z�X�^?����6��.�8m4W2�2�୽=�^����G�4�U�R���28[�)�^6�j�,k�� >����!��s0wu�\�z��7�L��Uy~vv�|�X�+�KS,MQ�?N��7����c��|w��(4�o�����E�7o<������o�����WL��%ޚuZ����$:b����7, %��|w�m�}��0՚,o"���������EPnlʍ�;}�=�G�w��hb�Q-&9,�޽��DP���5ra��'�|BK����<�Hn���D+|?L�%�D�A�||�J�Q:I�'��lt����lK���r�}M�>��nO���7."�ΎO_�^���Gy�IKcU/y��1��q�nA��t�U���}��A�<����^锌xۢ��1�i��@'5�\KZm�Ï?������ON����������YA	�8�>I:`�DX@L�i��Ag�:;�_Lg6�
�$�A �_�7v��<y��~�S���d����d��&}��������p������쒾n���\$i��z��*y������F��d՝�p���놂�dNG>�-�F�I������e���L�_������jVe���e�_}��G?� �B˳��=;�+���ܽ�X�/	q[B`�Y��q��2[�z�a<��`c��9��ӓE]�>��ߢ�lnoa>����ۣ�ٜV-���!q�.??=�}${��k\#�`{�D�,m
�=o,��r.���=<��I��fK@5a�T��wb_f%FMN��F����T�5���,<��͛��v��(�~pp��͹�r�JN�����ݻ�3��鷿{���ֈ��w���蔧@4����������kKڶ۷n�1:3���6�K���d3�$l<���·~H�������Rq��Z����7�n�^[ٌ�l�ZE&�x|NN/&d쇒���c�ǳ���#DJ��|Y7���)։Б��~N�rx.zh�#�����S%���Wە��K������q�r�'f칕�bF�"六���T=�����[:��W�O�H<}w�w��.
�J�6�ð6�D�B��z�1cg��h_H�g���TW:
��x�D'f��@�6=�U�!�X��n�� W�Ea�h�����2hЯ[��l���4��|�:��rI��7�N�3*������S��e%�e����PA&��H1gF�L���ɣa���i��ɾ��(S�e� �c/T��@M.�H�t�K��/3F|$;�۴�Nymt�W���]���>�4m)|�s�^�#0L��]���A��Z+�@$�|���O 5�4��w1���׸F�f��:���4E�Z�Ȁ�D8������z^�h�_Wqf4�H9I�IG�K%,!�$q�9D����@M<�%�,=$��	����d��p����T[6�,�	절�D��A����V���[p�L{�c6Wsƶ�9'Zٶp�̌e�Z%��f��b����REw/�E�0�3J�R4�K4�y��Y���ǃ���F!<�,�r�NR%粓c�:�B ��'$�r<TK��C�b�����b|\Ir�`�Q���b���#��N��:Lmg[�D`���8���zvU}���!h�@��`��y����vO>�lA"Ǆ�%Os6��"�-A������,�Z'/Hm!Wi�!��l�$���,�TFF�H��	b`�A/�߰���e���Э�ۦS���Z���0)3 ��S��㣴\��B��Ǐ����g�)z���'ޘ��C�.��>��m�5�R�Xp���]l�=DzN{�G#���W}������9Xr�H�I%Co��"�o�9-��~?C��Uڭb�uK��d��\L{�8�HJd�Kol������F���UY���؄��3��M��É%]2����os倫5��tֳS���G�p�j͎vۡ��Z/�r�6^�z�/!�\�2Z����I{��4�L�a�i�i�q~��+|���|e���:����%�mam�-Tv(Z-�!��ȕ�lR�ȩZ�#9_Q:q�
��5�b�9�s�k����tY���AB�"7Z+,E���F��i�vX2��[����O�OϞ=�&7�����rZ� |��̋�����u������6�v�o��S�j;|X�d#٭g(� S�?�8`� E2�L��EK>�1���f��0ѦE�[@�������D.,��s :`S�X��WPM���͛7]S�Dƕb"4���e���EH�)�wM=�F�/E�n[^��d��z0�n����+�9q*�M�%����I�#%9��P�����[����;�e��&n߹��ɓ��}�g��+��5��$!�N�ہ�����t�����),�� � MF��ߏΘS>���j��^$�2(�lw@S���c�Ҿ����Z�Z��ӧ �|���ʋz�s���l`a}.Oc{;4�ԭc8������~�����}��?��?J收o0`f^,>m���	Y1���)��Z<�%X������h:Q�P+�X.I�%H��J�YK_3I�V�jO��¾"���L�i�~����گ��qX���8�Har���,AQ��j�F[��������?���Ic0�m5�����/_Ӓz�)�|"�oc�{$� 1��'�-��H:�t��m�!e��&�?T"���W_�g��hW(�n1�3YʘQz���!����)o�L�<;����I]����U��h�bДelF�*3x����[�3	���}d|��$QdG�y�|1f�r��x�\�A\A!)���w|#DwKF������?����y�xqq��*�o�`G�SYV�
�v:ξ��.����7��cz���K���E���o�F�Ӊ0�K�Ni(.X. �R�Ӛ��zR,��\%�}�퇭�nR6H��q��	�9�rc����O�S�DD:�PG�6.�G.�=x���5�$})Y�D�F7nI�~ۓ�F@�1fSu�����Mf>~}J�����l�c)�-#ڋ�]@�����ɪ�b*9,t �O/xd�݃��˿�������������/����h�1~EP^պ³ �� �+3�3� yk��´2�t�gg�6��#I�GX�^���Kla~���-��uSQ̅�ĴD��
RaɗИΩ�.�0P_� �/�΃�(@�ǞX�퀙r����M��ă�Mr>�@!�Ay�̒�-�Նb�����F.�8u�����HGc�6��V�ז�Dq|'|�]�ܬ�#ձ���axf�H�_|�
ǿm׃�3a�m�F�0���%",�0��������Dth��2d��Xl�W�>ޑ,M:ئT�i�:�=�֙���ѷl��eJ��;�P܌e�����N����\"����_W�Y^���jj�)��,�_�l���G��ץ�黝����2�������/Z"m��:ɛ��Ub����-����\0��F��1��\��9<GFX��le�$���)�G���n'ϓǳ����xĽ��M�f�5���`�a�xe����pW�D��"ٮ[f������̅�@������cN��QP3
6Sx�I2_]�[r�a�\|��R�8��/����I���ZϷ��jә��rx��Y��ǉ��f�<���%�R�_�k��H,8K�+F7�n�Q�@GW���<�O��<�bYZ����Ԗ�I]3KQ£��r�D�MN�q|
���g*eR�"p�'\���Try��~q������%��.0�����C��BKMڎ�hՌ}#�ސ�P�~]-�'���^�<S+!����/�٦�xRSU&���B�D⑧��%��v�ףXq�\�P���6f:�h�UHz�g'��,��b�r�ĺ(̖�`1_�����E�&���	���L�y� �o�+�R���q�Ǎw��1e"��3�N��e��K�h� ����$7�[M��2y�S�)J�$��J�pZ���<֑�T��%�졆�Mv�Fڋ�{Y���U�A�<\FjUuh�i���g�~�����.���2Wk�B��b��5�5���mi��@5'�h	�߿���7o�\���B�[�&Nґ���l�1�8i�q�Í�<xd�$(S�B(y�L�N�^/haI�KTV�r���$/��1˺e���al&�W�)��/���5�_N�uz�ݑ.��6Y�t>_pӉ����[�ӵ�8 �I30���)�*��#�lwqK�q�9+���A��0����p�F:�V#�<�4�`�/x����"`�����#4�[���1@N��̡�� | ��� Nր#`@�m��
��� ���k��emLo!���=L��YZ����
L�8G�$�$��!"e�Y4�r�ܭ��L�"/8� }�Wú������o�����oc���귕��6��b*�G�
���� I�2f��6�76�<�{�;Л��	�u�T�$l�W�gG���y�"EkrZY#�3�H�\��lAB�hM�:AxZ8O�l�!L�.^�z���������_�xq1��y.���fۛ�t�����`���O��>����Z�E(r��n@l�j�l��w�k`�[����a� ���I����ٜ��Ѡ��y5��7w������l���/D�^�wD�o)����ݓ.�A�����}��9	-w�&�jg��H���۰5� ��zs���x�Wii)�m�H�Y�\0�b(sz��6�f����ɱ��| ��"�U�\V��������[��"�JNɥ�k+J�ؔ�I⢁�Eq"S6^�4n���@��E�@�2[`�tl�1��L��9�>�<?�sg����'���Ͽ�M9�I��V�!Ad!Q(��x�� ���|�O�'�\T=�ޜک"�S�v����n|�X+�"�'W�_}�%=����d/H��q���z��?|���}���NyG���5O�>=99"�˛���t!��R�'��e�l�8�H!��4��kW��w���Z��2��Ð!I�����"� ���U����o����?���+����-�SY,�O���)��nꀜ���R����I��ܜ�ʜ}̪����!@�_�\�d1_~��A��?��}6 ���s������b^�z�����HO�H:{�:!ekE�xv4�§@�xI�(�%�����xEMD��jY%#VR��Z���b�}rf5Z���5��ry�����b�K���8?~�]�����[�vaL<���;�������������
0�]�w4�_���f�4�\y�jߒP��`��G�C2v��5̪��_~9�>��ß����W�W�����_���"+:��D�ސ�ez��tY2�}ck��z\��Gz#����9�d��<R�|�'��b�
�TC��	A�"�[ � 3��W�W��-mV��I��H���l��R8���rQ�z���~�d�"arR�߼��#P}9?�U��9��+5����'I�]V�ʂ�r�}Ē8�k8z�R�$9,�*����E�"P��
)�g� !:h�-q>w84>U��1�����o����֤�A�F'�B����#�� � S	�U����Qp'l��i�ҡ�O{�&��Ђ�+-x�2�7��&��CSFR5�'*"1�����e�:jɼD�y'g)�Nd~o�j�,�P֔u.�?�����F^�T)@0��>b�mO$Y7O�I隔#�L��w�2���뷝i��Yˢb�7S
��1�J�cK�KZ<��$��"A$l����Rh(�B !H'޹k�F����B̫U="�E_Pj��g�~�),����H�Q��,k�?�a֋�DF�%V��-��Um�*�9)�fH����9�^_v��e6zֲ{�[��!�1�`f��f�������r�'�J�|KAڷ�gK�j� ��d�Ԁ��t�a����U����Qm.6�o��� ?�O�w"j���촌Ob2����^1 7��~�[��Sa�5��V���C�	.�߫ݿ��q&󄶹�NISO.&p PS�E��w
-�
�������l�k��_ ی��IT����fR�d9"��m�uJZ.�-5^�&έFB�>�^��on��d\@� �F!�&���k`��[��k�`H���x���N�=�=swO6@�4չ�Ҿ�#�џ�je�e�J���7
��-���hv�6͢�@�l-�c�n��/�ż���$� ��à�,����$ږ��ڝ�eQ?�pʙ �Ā4���.E.0Y%��{�br�p�k�'&	h���K~J$*!g��.��;;#(IR���ڡ����W�Q�]�i���\#���^o�ŋ�Rx]^�4�T�t��v�B�4��K�!��ߴ
2&w[��!��a�Y�ry醰q�A \�$�$�"���f!q�7-!�� �Ip���8!Ԟ��T��R8�^��O(�gx@d�{:,;Q�n"|H�1�^��ӿ�$r��p����d�"�N�y? �Bw$����Ǵ"�An%mv�U�{�y��< GAI��05(��7Yi �E���@��Cڝޏf+��"M$7 �Es1����g�i��1d@HZ ���DF��cmx@�7����GE����Vt��(����㐧3�ɣ��RC��c�h�y�4*b���qG��E��6�>� �?��*�A+�a��^�7�/���ӊ���ž�8i��Q�I��q���봲Y�R�����W������ʘ�#r�!������*P��R]���)�BH�W�\v,�i�TG�a�0�,�"���]KM�FG��2�����a���;w��o���t� �'��H�8��b-X�1ՇN[&S0<��x��o:�t����w�{�PÙz�0L0I�E�CgOޡT(>�G�c��&�:-����)e{2�ƆC��<Ud�H�$Wu2����pV7D���h6H��";	�Ƽ
:���I�P��w5��!Y]��Q	�]stt��������H�O'״�8S%s�^��&����	2�u2��tۜ�`�<�$o߾W��2����tG�P��,V���o�P���{LhF��۹�v�����+�6�gX.0x���I��\�ys�'����?���U�����>�=�ƁC�s�m�tŃB�jz=��`%�)�;!�����i=1�Z��I�\�JZ�Rl-���88R_t�o߾]�]�zfڝ�p�c(�G���I�m�u���=x('�y���o����xpp��w�����|㚬*�כ�����!��j��R��"#�eg��| �h��m�{[��M��ʢ��؍=
�I��Q�S/�I�x��bR��|��9��9�?z�9��?��|�����A
-7I���K>��˼��2����{�}���gϞ�9|IOzy}�HQ���It�u_E}�D����su�p��ҜG��&��G?"���ɓW�^�u�޹��'����3���g��lSʚe5�R�8T�$���Ew�b�L!މ�:�}$[�H��X0 9
�A8�,�W�.�<�u6$��z)0�j�R��ˢx�Y�A�G�1.h1���[G��Ne���(�����Pׄn���.xk��n����5Y�E���
e���x
(+�N������(qe��:�E�X�I�� A��ƦF P��kb4�y�9�6Nʊ��ں�Z�4 ��ӳ� �WL
u:^�]�^F�����8��G�i��%i�B�m!v��f�rQ*�wM��65�:�4�W��+f��"���;E���.��ޙ�M���f%Y9+����y^��]G"�uߛ� -���A|\j��z(�)=�߳l�z��#!>��6I����;�d�`!�0������#��\��ѴK��ߠ�Cq ���B���EY	j�J�[d.IZLNω�?�,%bh=��^\�5#5��pc�z:E۶�Q�<V����
^��j%4��;*QJ�F��Mg`q�A���k�NC��7��ø��`�:R8;<�5}��Yu�K��-M�셤C��\;]�-Ѱ�^A��Ks�:e�>���>�j�
�}�ܺ�w~~��+�f�,�(�bqvy:�$�ƾ+�y�픟=�4�(��V�J�@�t���Չ�,�:5��,�̻Z��s��iE���u�  ��IDAT��Yb�L)��y�r� L��]�,3�\g�M_hP�jA(�!����E�"Q���]��@����ػ���44yo�ħ乧UH|~=!��Ū�-�H��$��A���p��2]fb�=��yrDA��,�H��wsw����^�|��1.)�-�������S��M�.2?����׫U	��T���0`:O*g��^&B���~Uڡ�GDh����3��'�,�|י*Kac!m_� ��"W��D���'���;�d�%-^	�l,7]�U�
�3�>03�j4bQA�l�d�~�,��(��N��+�F�����&=~�Mr���%�N[�S�]�I��Q��	<�~��,����n�F�dW���ѩ�<|<��]-�,�ӝ���_:�\�\-��x8�����;�E���>_�D~827���7�����']��ΐ����ePϴD����2�E�6�9���{�nm���1��tv
�>H7,�ַh���� �G����C�35B�91�1�+$I��j�}!cc��`�I�}�z�J"�r-(s��k��ٜ�Q��f�i?�WH吀=z��޽{�����h����b熬�Ũ?n�2MR.��@a/@hK���<�2�<��jm���v'�vJ� S�8����'��M�>�RY����9�]��EYX���gJ�d�y�,�G���Њ�ӊ�+Q�!KC��z:�ggg��Lw U%�����<:��%rR�Kvm�g(�~�Q�\��7��tz�6noo�����k�F$��\�8K���}���d�X����`#�Rl8����&-1_��$c@����yv��j�C��g�4/ƛ;i޿���[ݑ�p��X1�1e@���mGP����eh;�X`@睎�Ug+��I^M�����k��^�O'WM�wqq~sw�/�:�t�66��od%�Y�_�I/��S�����#�ɍ��y���j��[��i�+������4�':��	/^�e>2���_D	��<�:5�T)�r�q�)@�)�"2��ޚ�9�Q-�nzY�~��%V�s@�e��3|�A�2xI�թ���cc�4U� ��x^2��$|��X���L�,;����s!#յ�����wS����I�\_�_�{���>�/���͋W���|��H��Q��Oq�裏v67�
!/c�9`��ѕ��.fSFXoll�$l���ǇZ���R0M-R��y��B�d���/(���'�x��0�|�	����Yu�����dhy�mnl�W�_/�r��T���ȿX�
��$��:m��OG}a>��@����3�R01m֠`�N����3Rד+����,v�Ϗ�Þ�R��I<X��^Y�rF{7o�G<���>��?�Q���hX^�Nc�Z�3�<����%p��p�� 
9�����I
�|���������n���o����y���/�G~��ݍ��|�C�MB٦
o�+ӓbH4B*˶���Q����m��7C`M�V鐳 �%9pՊ� �+(s<ч�wrr�����<,�<�&c�[�XNJ��Zd���Xۆ<r���	z�&}��q�d|����[����T�?��������SzJ.��R�S�����4���fp���U�L�}�����iYv��� ��V�a�q�Za�!C����R43[�e�3�$)Ǽ��]"?���Vt��h�d��d���ZWW���NKe�8C&tv"f��0�S�)6��ЩO&����g�	5]�`y>�����}�VYz$��d/�)�z�g~T�x�]�N�xM��xZ�k3�%ݼ��Y�B�Fˁt3������̏�	�׮D�mH]��
��I�!	�*�M�����^YCgV[T;.�=���#'�n�h��qM݄���5sI�XR@Jf����p�T���h'T���-&�./�8�<��Ǳ���)F/��MQ16�Ne�r֌��Y�ȠY��is�5ZE������fX��-�se�,�V�95e�JJ��&��.�q��3�^��GU]i%,~��Y�n�փ��PR7e���O<&J��%B-�b4�,����Ȱ� �Dd�	G��{�W�
z����a�Nn�\��G�d��:d�d)SY:���r��ek�{Զ�z�v�^"�3�f����I�`��yW4��47��T��+R�TT��[u�Q�&�|���V[�T;V��{��\8A�UG��B�-P��0�&�-�{-hqBn�)㬘���k�d�H��6�Y��'��2VE'	�,gP���&j��T͑���4u���ݿy��XTJ��LD
鳽=rfv�R���xM~dz�,  8^r+̺ZErw�*f��sCo��`�o-�ws����^�gx��E?�͏7�H}�͓mF]�WtW`}�jO����̵D���wڦ���%ז��8�F>K!��m_8��V�3lX?!��K̝�I�r`�K�"A������{qKW�|�?]�e�֭�Yo��ǹ���r.���'��M�N�5�ʑHG�7��b�Y��O�XF�{ס�Źƅ��Fk'�ȉt#VG�m0( 6��1�-��ȭƊKdt�hgS�r�iU5q(��A��D"��_���6A��k��Vޜ�"2i*��Q���ZƬ�3M�5a�C.Wۢ;�����Hcn%v3�dY��:��J�4�AE�R����y����l<T
o���[C�,��w�R]��a6~JQ@����l��\<;>�6o�Iyv���Aހ��!IP{��:�-i��e٫�.�لӑsnt�1H�떥(�$Jj��N�]��L0K&l����p�HwR�q:2��*�	��HL�ʠGN-]M~�J1 &���F��)|������,��Y#d��0z5����+h�F�p��h�@B��<v5�'�~����vҫ�p/�2���O77��o�����,��u%���aj
Npj�Z,q�葱5p�I��*	����8hC�8��i�5r��J,HaCtqN��Nr�V���ŹL�B��K���DK:��0Ҟ��n��_-X�`����yJأT��� �����E�y�2�NNrE�@�GQ~�"�b��y�1)Xg��xsG
<�9&�p4��S��g
�&:�� ^�����P�Vxu�8Y�1eB���s&�u�T���J�Ӎ���XD��u~��d���I�Nn������+}YZ�7���'<88�}9>>�u m�(�M~��Ӱ�M�K���B�q,1�(H���)�)��<&���`�i+��E@暯�z<�1�OX�����f{q�9� �u�	�]󵋙Y��A�N��j׈��gݒ&�P*��IO[��KWJ�A8�� ��d�����4��\phI�)t(�6;����^z8G��"��A+�����Ϫ�~����<��e��K[�D��`H:m5_Ȍ�^1�0�3�GD�ח_~���T��&�T'���fm-/l�S>>���ЬJ걿��|�>#�ँO���N+Po��Hx&�5��H,d���,���ְ?�3��P��Ӏ	O�TY"���ӫ�]�@�70Kf���J��1�1`]�V5��7��/�oޢG{��	���3�o�;y��Ǐq~�ު��l,�:ݻV>�֡e�Md�
���jm��"�Vw
�hV�u%�t��&��>yM{�o�n�����d8�$̙���O�5�aMxR�c��7n���}p�Q��ۤ:ΛX��]�yש�B�`Dp�9�uy�|���	�د~�+~���c��6A��[\
)S��~Xy���qf;�9��v��Mo�e��XQ�!sby���b�z.y�8y���E���6����-��=�'� fz�l:m�	�%<��t�s�����*0Mؽ��X�D��1�Q��[eK�8W�u�6>�4i�;�9�v3:+�[E;"�*��RHѦ
"i��B1S�X�lE�q��m��ή_\��d|i����e�6S�:J�`=�&�g�(�wR�ϟ�����-!��gC��
����qҝA�,�a��Ԧ�n[m��d�s!��
ǳ��Xj���ڒ��?ko�$Yv���s�Xs��j��F���!�� �H��l063����y�Lo�2���HP(��Hh �@wWWך{fd�w;r������MX[uUfč{����矛kg�u���5ݚ��:�X�����&^��/�f�rWx�NS`W��Nln�ْ$�f� ����)�d���Z���
-�8�I('�Ӻ���H��ixc_n����*A�I��I���cb��o����sw�EZ��S�ƚ�ܦ7��#ɴ)/K��9E����P��:��7i�ڛp<��*���?�΀C�WD�e?��.e���~�P>�-l�O3Sx��x�*�52nM�i�����Z��vW�Zͮ��C�K�	JX1����dB1?R�y�,�;�3�4K77�;�����ի'O������+�'���H�����&�����뤽���,{���&WdP���?|���!N6?&�
�8�C(��y'�^
m,2SH(A9�	&��w/�Yku�,0��M�n �Hu�s ��xP��E~y��MW���x C���BkwߤфĤ���p!S���n�]���ܽ{��Rn���K����Ū�ѕX�����艐rGQ.'d�!l�u�3R�[�ʥFb^�I�d#��(�N0�$!{��G�U�X"���,uv��P��eoo���#'W��ȧ�N��/��ݣ-�(ۛR�~�sR���MR�L�s<�����]a4Mr�'��(gd���|s�?��������>k<G�-f��2u�ekCez��v�ep�L�����M.!�f8ޢ�X	'DU��I�q�Fml����[^:ﰒt+eU.sr��r%*��:w�RZi'W��J窫��08�	Z�ȮQ K�)��� )�8�2r$�dGj#w�Nsw#���ߥ�y
#��覗�#��N��)0��^_c��J����l����K�Y�$>����^[�+��� ۈ�� �)��>E ��...J�_]�n�Rd Q�JxOV�%-6�.�І:aB�Bs�6��"1�,�ȅ��4�j�+�;��7��3��9N3- ¹��PA*:�ר�4:�Z�k���@Z-('��_��F�<Vb�DNt�2��+��
F�U.�%�e�j7��v	���i��u�#�	�t�!JA�M<��Ri[1����8i�Jf��qW���VY�4 ��6aY�H�N|��ݺEwۯVS� 9�����G�*�v����~�&{�I�]:[T�钴q��b�$U���ݑ���	O�!=V���Fنק'�zH�2���F:�<_n0��;W��'Bz��S��啱N��,�:e%�����M'I�q��DK]�0�>Ů��)�kc�����lg;��N��%�1e>�j���әl�j�Z�B�3�'�t���G#:�������[E��Tm�,��ˋ��'����J
U��3�~�]~�+�)�<(��y���h`�K{?���8b*�cK3$�EC^a�N�ӣmB�����Za.�9{��B�U����?_�"F�͘l����,��
7�/�)89_t{L&E�˰G�^^�������Mr��������F�'�m���[�A��#K�1��ϯ
�V\�d9��]I�k�]�/(��jz�9�5��ɔ��˫Q��ǿ�\_���:�������4���t_I@�?��tq�דT{�F��Ko��ZTg��y,��E�e�m],�I�6+��.D+L� 8��Tz\`S����c��H��"RN��ipzvvyu5�\�����:�Ϟ=��C����\p��ϑ����ɴ� HR)�$���޾��o}�ӏ���|c��BZ�����6�`
��G�9��I������ᓏ~��-�~����׾��r9?:9��O�����z՝�����Ob��{��v'���EG� -2Hd4!��`���9�@P���ÚT���g<1r�M�ꖧ׆6i�b�����x������V܉��ٺ��	�����j{s�z���$��P�岾��[w�Dǅ0�������c,Q2��1�&@��Y��lX�}�t�w���L�>����O�N��?R�t�����j��t	:��1R������u�o����'ik�A$!�����\L+��e4[�<+�l���k��"���������)�>����走:p��$B@�Xf�Z�Z���5�8�r�v��`��ՀT���F,*+������}Ӳ�L�k;M��kY���{��;m:c1
��pJ��oDc'X=��S�X]� ::���ec�Fo1�o��A�hg�ɐ��[M�Q���-C�nU�D	s@�+�#^n:�\�Ǜ�EC��T z��p�K
��[
 �Ia=��$M,��(ݖ�Υ���U<cw3�)���/���:2�&L�G&#Z���!��0�2�U�c�V�˱y��Җ�^��`￉�/:�����8 �s�����a�A��K�o�Cy�(�L���B���$7�[>f|��@�r�ʌG�0y%�]��ȑ?Z��+�=�ɢ'cL�K�0�&�dA�L_FͲ\6��e2nF&��Er�L��+��X(�tdG�1���Z�|ʯ��`�1<g�P�D�dC���D���+X�ܲ�V��� uo�s�\g����$խ��He�D?h�Ʀ�L���(��n���-�4�m�E�I�4J�a7i�fJ������:��e��Mt&:�Ö���)^�is�9��tA	L7���:=k*-j#�
a�ONN�� �gJK�v^�5��w����[o����z��y�iQ�������&��4W���K���ݹ����f�Y'7�LTD#��t 7�\,2y����b�wZ62(��3�r����T�ʈ��8�����2�P���c )߬	���i�Z�ׂ
��.�Q�������n���u���;�����n{����h/h��t���MvG�*�浢8���=�E�=&��4�
t�NU��iwM�a0�#٭S��:N�:@|t?���@a��+�b�g��,w��~��矿z�
��Yߠ#G�����@JeGj���r�� ~�����yghUX��5瞧#z��r7P�3[}���C�2��6,��u��'Sέ�0��^;-��	�"2�5��S�؉� ���)T�L�阍H8� 1 �5�\��$f��8 L��	Hi�B����9_,������|�\<W/����	�w��*hܳf� ����^�J:��+z^i}X�'p؎�Pi
�"`_�b����İ��Y�{�r�������{���7az^�~}||!��9]�l����>f9%7��2�^4FT�q�ܺ��j9)E�5 i����
f�1��s��z�[	��#�����F@��,CQb+���������D���7���
	5�&�І4��l��:ٿ�gD��#��3i�#/�
�N9@Xi���qN�]�E>f-?^�1$-���^���=��W��C�i�4����d��Ț҃N��Z��u�.�AxyFnT�O��D8�)�+Kc�I�Ύr�D��d
L
�?��|���y�)�����ի#Ҋ��L���Ζ�y�O�nT�LvZJIy�"z�W�O��j��G5
�X,(v���z�
6�d�'N�t�	�.�<��zϠ��N� 8,>t.rM��Az��-�lhM���I��40_6j�G��X@jһ:5D ���d�ҍ���(��ȕ��f���Q_����.h�V��-t�[��ٮ�R?���(����쮺ϔw#� y=[Q�}�p���G5/x`wh+���2�U��#PH��1Hf
������':n1*�bЗX��j�0#麥��~�@S*�S������Ɉ
`��T�a�V����2?���p�䋤� �4���6�Qhc|��]��A���č���T�PP��~dd��(��`Ȝ�h����^2N..!�t����O?����d��WϞ=�q�t�s8>��t2i�kJ��{��{����?�m���)]���������P��/�l����O6;����_\�=߿��L��Ǐ����'O�G�׾�5h`CK���������%��7�D��� Y�J�Cl�-#��s2m|f0��!RQ���8>8<|��ѭ�M>q�����[�1��'��D��C�kab�jӋ�E�Mr�g��V���m��&���*뗸ă�,fE�yrRf6GY����ۻ�颕�?< ����/3��S���[Jos��B����&�+��
�/���b$<�!�UI��.I�ŚM����)��):��'pcG��c�	�o�~��ע����7t8��q��\'�f���s�_sڙgޠ��!o0�x�����ZY7(ٜ��``����ʝc%���A�&,I���.�:/��v��N�����8��.i�xL&���S��x��#�%�D'Z@	rl#+�,�^C`wm���p+�8G$테���d��N$ڊ F�M���{�&�X@�0.��𝊚�Sa��K*k ��VG)���C�穂
�#?�W�Ԓ$Q�Hj�3���{4����e�a������N8ܚN��=lwC��хX�������lx;����6�U�Nx)Y>�}V�|]��x`E�2鑗�U_�),�`Θl�LIi�ޗ�l\Pd�>�����&��AldЎ`�'�F�����::W6"C&JN4�g�K�Q� ~Sͩv�⚖�x� ���`[�7Q��J�)�}���4l�n�\	�
KI�{䴘�h�ъG�7�%����L�ҜZS����K�,l=me�����[x��Z)�7����k	M�;��4U��8��Y�zy�QDq>7�>�w��D&Ok�(��73W���&�)��So����7"?��h�l�HѢ���8��VU)RJ�F�e@2�IDR#+g ��/C$�ƌ)7;eɅ�0�R�v�DOW?C��t�5A�T'2��dz}z1ؽ���6��.OO�oP�چ����)�c�����7�����==����.s�]��$Oq_���=�e5 ���K`���^A?��4�H :d� ����&�<ˡHsӌ(��}��;��G"�J4RN	a�g��\�K΄�I�
��$���A��?Q�u�[�����NϾ���E;$��������
� �w�)���ב3B�z���=�d-3
8��Ϳ�����������/omop*�#i�C�]�a�.��SGǚqrZ�I� �in���-E%�=�`����Õ�\`z~r�rEd*�NX��	]GZ��L�=���Q�\��gs��+��y�j���1:�eh{ߩ��e�0 RCX�?��4e�{$~�`n�J�Ec��ahB` Q7ZX\=�'A]D�Օ��@��E3�ԡ��¶w�}q2��%/�D���&��3Ե�Z�K�#�ޏg��<f4%h�.U|*S�k���1��q ���vM���E�H@�{�e$#�u���DYrZ� �I;�^���Yu7Q^��^������Ϭ|G/_�R!�-�t������.�tȂ��R:��)a1C�����A��`����HG�VX!�"io߾�(SL����O�p����U�k�3���\F)�VvJ`��re�z6}u����~�l��L悶}aϩVR���DpyY{����y9qio��۾�5.ol�q\�&�g��կ_��.������~*��i�/}�j>���<=�~�+�,N��&Н�#b�Ms�X���Gݎc�ϋz%CQ�<��1�H�kAkNןL8�0�����/j���x��s���0����������InI\y�D82�}�Y-=S�a�N�d��U��v�P���K�!�ɽ����k����Wx;>����;��C�^[ř$d��s!
���S[���iO�Xs�AF�	0����εt<�j��-�Ʃmy� ���جT;1�?���߃�)&Y��xh�ܲtڦ��<�F<��;99&#xg�f��<�+����"w[[x�$��0u���tb	4D������х���cuzt|u~1�\߽{���ߺu��� C۲�ˋ<�������r݂�ӱ�PVG|� 
���'�Ю�1�!Ku��:�Rd�E8An����D0f�|��������C�j�;X�S�����YL�����Ǵ�!� ������W�{{t�omo�ww:���?��yϑ#����ϖ��#L����A?�>8�e��������������������]U���-4&C�Ur�f��8=�ٿ�����ksg�G;=,^��&�7��f�#�eݖ�)t��@D7�L4�4��5,k6�ꍠ=I�X�Qk�h��Q�p���� �Ŝ6�!Yރ�[t��׻�����wy�<��?޿���[%�9��4�JWHjn�Hή��Q<Wc:��p�R1[.�"gr~i��t����Tr�E�Z�p��QI��������ј��>���r�o�Ty�֐�e�����l����&�Az�����L�-W�U_���r��9f#�|�����/�\��D ����D�3�{V��6�	����.�D�н�V�6��$z����???g�nћ+��������nVs�o�%�D�(L�/��@*�$>����|�v�E3�(�:���2�4�az2����"�Vabf�W^�h�$�R�py��M��L����ϸ�U�w�+�'hQ�v��b:i�(�I�
#�JX/hzP��7���BN�[3�����t>��h_�G����ɌxW�w�]���nZR7�,W�G��ЬK��҃U�,*�M�9����o��Z�'$�Ҟ��s��Ht��o����f��֍���HA��	2�1�Ck�pJKx��x�D᷵�Ȗ���!�p���=�M޵n�'B��	б���6C�I���i����S$ ���^�lȧ��nI��	:p�U���ƚ=���c ���DMX��3�'/�,	i���2C`�_&-:ܳ���~��	y<�L�C��i��]RL�S��~��b�VȴIG�m����u$%�e
��˂/��G�y�S�b���P��mv
v���ja�<u�O4��Wk?l@	��,1�(��Ӗj}��������j���)��l[������ԡ�L��*�����X[(��{���w嵁?��<�V㍍��
�x��=�v{�#�F>�x<A	�;�`�V�3bŞ�3	c$I�4#��Ϟ={��1���K���wT�JiZ)	�έ%�~�ەiP�5"U�H.���,j+r��w�_phD�
@d0aԦ����<C���'���ﮍZ�	����c��+��M��bH��ӧ��ݫ*x�����&��k� �ΰ�?��#���S&Ep�ao�T8�	w�0�"Ǆn$9y]i>H:�f�D�Xϖ3,�%����h�h��"u�ݠD5����F?S�6t#��%h�T��I�C�a��2ì�3'8�xv�P���y��&n?2Y~�h-G.�_�O'��-b���I<�ؙ4!�J�z�D���(FIlo3W��4�
u~r1�Z��FĖh�u���}�A���t�*R?�5�3�R���	--��
���'�b9"�T*s���?xZ�T�{��t��D5�(|l��\3��ܺ�u���t�1��~��_����!���>���"� �[z�ʹ��N��)��;���"��Z`.VK��Su�b@�|{ćB�\�t-(̒`C��!,�~��)�k`o@�c�<zU�M.sW̴Uګ�;��R��~J�"�d�0p�D0�A0���h��ғ���
ceB��g�����;n�O�C��|1K�#�O��ŠmIBY�������Ny��:�VX��!�F��Z �R�#����� +	�k� 9��d4��3=��C>C��ֈ�8�W�Y�$�~.�Ζ��&�W�� M)���𞑞.�90�����@f��H��������6����qj-?�h�P�o|��������/e�����Z+�t�]�k>7Q�E��9k��G�ͼ��!�Lvrt���y��׌�X�3��2TG�!��Р�9x GGGH���$]J����'O��?��SL�v�LG��3&�����-s�np?,��@�ͺ^�np�	˹��Cz����ޜ}��{W�O-���mD�e��\��?�sm��w^H�[i?r�7pR�Va�Yj�ҥ��
>�R�1��ɬI��q2�{G|�F ����V���iR����ɥ����<H�9�>*�u	��|�e=䞐j����V��Tǘ!�Dm���W��}�p����ݗ�9Ku�{�VvW|��n��*m��8=}z:�a��<�5`Z����۷o�[�"��|����\]O>��������l�XXa\!U����]�;�{� �?}J�����?"a��"�ߣsM_M�����ߤ{��^2�?�������fd�om���~��w�%��o��oV���[�xzD�U��<x�+�w�1nz~p=}�����T1e^���tt��e�����c/�[C+��v0��~/-��(Y�1o	�M�d�8r�t?��dJ��2	G����t��2��;!H��5�0	�V�˰��� �@�c�Jש�G�^�OzV0��3"���dq*t�fт2�a���x�%�-�\��	�'�}J�7�@�T�_1��M��#hN��k�J��&��6�X�����^X�b@����P����}�'�Qc��jڜ����vǼ��I�Ɛ���*��,�#.��A��1��*���L7��i���5��|�&��#����]O�k�֓�Ź�'A�H!��@��=p�� �������Τ��ӹ���j~AA���.�۹rs�Jl�� ��$��}�s��g&!mꔂ+�  ��J�)�%��X�F:�4m{�d)_�8#�Rʦn�L���ZZK��4�9�+`�6,���<��FG#�X�9K�mD;�u�C7�R��VqW��d!c2;�w�g:^I=��L��\�����|S�����,����{=��P�}�k��,(M�p�ж+a@#5��5i�Y4���[?aWG`AWKA�w���F Y1ѐE7FX��T����C�n�8�i)�����onm�Q��&��EvJS�
�����[sʬ�-�e����j�R�֜Y������.���G#���w�7x��{���(cT���v��PD׭�$Smu�}���S�"-ҕ��&�𪦉�|!$�:��lݹs�~EN	� :ɒ9Z���@��r�����c��ɳ��)�/@�	@L�g�ټ���G��JpB�'_�V����N��-�	HSg�<(�:@ɬ��x?���9$�β--��ftƇ1:���cd�#V;eX�T���Z-�@�	Ӝz����8a�b��U�$ì��'n0��س{~a�[M���2�����#���������E��2���Ϲ¬�� .���B�����=�^P�d�`Q�(�d�
�V\��3GI
	G/�4��~��2�nJ����C�k��2Q0�*�u�J�6G*����c<%͉������C:M��0�.��� ����ܦM�������)r�����/=�ˡx͐u�ő���]�Ӎ�(j����{��������i��4�W孭mRuU6u[3"�6��eC��=I����{^B�W�^%<iZ(�vL��e���5ѓ��x�w�ŷ�e��(���dM�ώ�O�@ Re}��C��2�d/M��� �I75�,H?�qk51��h�QdX�&H���6�i1�d�)����/��H����Ȣxcch��x��z&�"?`)�m�A�R^3�u#x4q���;�aj5k��ߒ�G�7�	��V���{���7�j�Ӻ��:�{��DF(s���meP�n�9��I� �JC̥F|�Ɓ*��e	�9��9[�K-FP\`r�����9��'��<rW�mz
�v��V��t(���@�8��A�%�g	���]E�F�|�R��\�m��a����u�Xn�H���N�0��bQ/����^��&bc��WӪq��a���Z?_��{?�����%E��b��L2,��&'��P��ӟ��d�=/x/���H	���T2�kNT�y�Z��Q���l�tB1=�rN�b�Ӳy�
s�on�Ѣ��趱�K�\Y�J?������ZV���x���ы�â7�^��F����ӧO^�xA���|6��B ���"�{Y>%����T@���=S�o�� n�Ε��<�yMM�����Ç1��k/�irS�+���(�2�eu`~G�T[%i���e�������5�����4�.nt��)�t4��S,��� OR�/�l�`,UG�|x�܆��-��0���1�$�?;;�Bz��{��1kJ/��z*3�{;	�^�wdt�(�2�:Kr
[8��f�rAzuqN�~zF˕Б�f�����<��ޘ϶�^��〩ӭ����E�cM��reQ*�k���X@��,�r�#��������wY��1��b>�����|~~��?�я~$�M���$K<x@2�����Ϟ~βD��j�3�跿�����ˋ����#���o������?y�9��/���ٳg{woӝO�ώ���8������������8��r	y��_����7'�|��&ڛeo{����ť��vz~.!�'�O���g��x�r�`�+��έ�=rz����E �A揾B��2	/�-���݄�%�[�5�N l$��3��(�.!SN������,� �"�p�o�����.Q���R���qAv"��MVћK�lY<Tn���uk�5^�/���a���	N�t�H#Gppp0�\�����YB/�*����6�>B�@�N�]�/�h���ҙ#u>��EfYvzp���a�Bz��b�j��[G�{����㤍m��1�b�jJ�Р��Ɛ�[4�L�.s�m�.�.f/^]]] Z�J�i�Ekm"4ρ������2��@��eŚHh��nHn��F>�Ml!N�7��!�R��L���A|�n�S�M�����-2'`��� �
�V�5,����:��]t���{���/~�Z�g_��}א��|��N^~������B~~yq]�Vk��%AF\V-{��,��՚�(+a�>�|Y"\�9`�S �H��]���z���D�1K�� ɞL��Y$F�&�Jd�)�a���X�n�೪Ywn���bs���O�e�R�"uN���o��d}~E����E����ͣ�M�iL�6�+/�˒��۞i����&ݜ����f��c2���딕S/1m����P2��JϷI��P�U"c	h��Izu#Y�̥2d5�	gd`���`J��j�5;�"�H�Kҟ�U)�0���%E�o&�${3ǩ�̈́)��Ѭ��t�+t&:�&M�p����w��-��*Ʀ��N*�캥�-R���j}�K�B�Za���N6͊f�,��vJ�%�)���*�u^�	2;Aa>�8�ߕ:��uR��ȆEr�A�4ePR{K��N��k�&������	����"���%�T�ԥk���/-���^QL�'�~�!�f�S�J�<c\�mZ���������%�D��'�N�/�K�Ni����~l�UB�(z!����@V1(J����D4�Y�ַoW_���JsB�B�cӥ�Xu�j��D*�dk���<Ro�m�o�7��u2G\��%�<��J� �|ș�����r�0Xo������hq8:J.�ѯ@�!����W�����r����Z:F�Y��AVЗѐShF
����y��`�ģi\������6u�L���$A��~J�A�9I�@ʂs�P�$l�tZ+�
����vvv�C�m̑B
������ߦu�o����dQm��w2��f��R*��a�MR��"�#I��Ai[_�k��%}�x���]�[��|��9I)z�_�I���Z�G�$��B����sj�,܉S:9��C�%<BXkJ�O�+�E�c��)�aP�^-��6�F�g�@)IS�I=l��`�V:�����)�_`7@���l�\vs`�_用q�l��_�~��Ν;��aF�G� �jO'Y# �TwB_甀���Kdxh{.B)c,t'�r�)�k%��O=~��w�_a��{�G�������b�\�Xu8��6R��J�Ǡ��RL ߁ծ�8c7�y�P�a��=Ń���>%@�Yj8yfD`�0�ź�!��+�` ~�&tKim8G\��)ɶ3�-�$Pi�-������ӵ�	����kf^� S��J���cU�1n���8���l�Y�D(�/�`~MW��8D���񢼼��(�-v�� z�|k��e�K�y�b����_����ΰ\]� �Ă��>��֊�sKZ�������hEZy�m<���~�[@�?I/��a�b����\:��*���3��������s�&W���0��F��X�>�._�^+@d�^�έ:M�����+i}�k�j���1}>�Plf��H�6
_�ph=�!]s���Z��[8w
k-#��D��5Ӑ�U�2F+1� ���7JC���V�W������ ۴��n��ɴ��I%'MsC�-\���rV��y�����2`@g��诲�K�����GW �T������VA.�d�.Y.�٭�]i[�4-Θ��F^�aP�B`��d�*�S�8��?Y5|�6��{���˧O����;F�f!i�o}�[��\n��ɧ�z�~����O^����c8ܢ�������������w��Q�;���� c��|�A>��^�����?~��'�Ϋ���?���޷�{Rb��#L����~��)Jt� �YXJ3���=i�����������+����}����}�s3<�J�t���~Ew�9?��g�l p�-:ڴve��Й��j?�F�':wK��ґ磮@�zX��қ��#aG�b5ؠЖ���+پ9��J^���*�l�Ev]�7�LS���U`���:P��4�5 >6�FH�����\�]�x�駬�NOp�ɀPPϳ�8W暥CD�[n�(8C��9���d(AJgZ����d=@)���UZ��=f��ҧ66��{��弄�����1ֹ錦l���m�":�B	�e�G,{����� Hܰ���PB6��(j�N�J��!� 7HB����7�^����������>Ű�G���б��X�Z��΢�����.���2���X*�&d���l�h���B�#�����΋�+Stm�"�(�5<p�:��c����[֜��Ɓ�.��o�2P�����V���@�r�s[Eʅ4B�k�q]�1��y���͖j��}^`�S,oXC��Fe"���6@���n�[_M��iY�I/�-���%�v?t+�=�����+�kde��,4�T\I��4/�1g�yJR��"��.�CͰ���ru|{|v>o���[���f�.�p���L�W�Q�5��N~�:��&ҹp{����|�����yfo���� O�G��2s�^o�͘E��h��*��iW�I���!��c��dD�� �v
Xf[�x�.����?��A��	D��@k�ñ��i����+ALPd��,a�� &��ܜ���.W�U��ˤ1o�*P��	� )����IC��?<~u��6�ܽ���E\��9�9W��Ū�؊�����m�z�*-.�F�_�pi�x4Q{� W ]�C�&qmG?�Q�2c�ŷ��	)�
���d�6�Ώ�Θ���Y��j6㙅�\s0,V2��/e"60���y��~��7Gc��In�
��9�?���{=v6BZ\��ӆYx���ܕ4���j�m^9Ϻ%��l3�\)�Y|�d'W�t	C�+�蹪q�g������<$U[���\0��/2�Y��&�2�{5!��w��^�5�	�WQ�zXZ
H���S���=m��z1�./�;��ùj{gd�j�3�YU��\�{HJ+OICx.x�@F2y��s�"� ���	�zRg��|E���!L�B	d��L��zI�F�"Cᔥ�;��O�3я�iZ��D������UY3[��-�e�`��H�^� ��i��-�ԈO�]�L�1���c�{���6O/��w�TM��sYͦ���+�o������R�:X���|4�吰����b�C���ϝd\>�Q�x�h���\ckx�8M6��P�~ttz�����3�jN[��с��߻s��?,�>��,�Q���3.e.h���r줙�
q�V��劅_�tz�$���*�wb׭�0����΢�=�wd��F<F]#5OoC!�����B�#nm!}�&)y�&��������'�^�x)�A�>K�yi�� x�C��E�È��5�a����Ւ��<��i��.F��P5��7���-r�76��/^���,�:$�h}�x2������|��-5;C��i{�I�y�j^7,��D��V�6�����]I��� "�L^������6���*���S�@�I��bI
��y}��,�t�șn�����5'�VA����4W���|�<m�g�z��L.�nM���m�|���Ɯ=_���)r>6#���ڌy�E�AEn�*uX���&�p����N�����F0�*aD)"�����u2-{�����M�g�5��*���x�z2�S@z������z�7ˊ#%6M�i�Ě���b���~�4	�0G�����۷��"7g6��|�~�
����l����@ݒ�j�,C��5�/Ͳ��&���zQ��5S���I�Η5OS ������Nk`�JR���G�����_V��6�����La'��	/��������Eb�����
vc8f>����xR�ܥ^�I5�����	����������b1�x�v?�����y�s��IT(t�&i��b*�XR.���`0�/��W	bf:GmCC��B���,��TjoS:������ô�֗�D�$��"혋3�fs��,|D�4���q��H�VB"���I^�rQ֕�̐��cJ�oUϙ
�%�zg������"y���w����2T�_A���<�B�VjZ5�$�,�mpеZ^�]qՀ�m]��V"�X	�)�z�IV^����rF��1��!9ƪ�
8w=a|g�[}����M��Y���i�G��3ºn���V��&]�'���^����L|]Hm.;p	}jEna�ƻ:�y��CFW���
Ce�[����dW�T�G��x�9[.
��_�6�fw�qf�c�]zq>��Ѱ�r:r�J���[;[���/>s
c��~��b
��EF����B�669�D��J�xdY
$�Ze�E���
rog�e�c>m�gSZ
�_~��o����l9�Px��#�p5�6�����y~t���������_}��������c��$�[���������B0���{p{������'�Q��K� ;Bo��6���|�L/_�t?������k��_ ���������?��w��,[�tϟ?uz��(�e�\5i!qf#��sF!��l��g����Sd�h���>�����g��J7s%/xz��`-0]��D�:<ɍ��VNb�//z=��0�7UW�o%���M�C�F�
�;��r�di�ԧgy���3�"Y�!K<���8�5��`ks�E1/�k��:���4\�f����\�oe���)��'���H��Y�
ց�+mtۡ{�YG !ߛ��t>�C��j�XJ��zr�R:�F�9�!H54�B=[�!���<�̻������bЛͮ?�����YY�R�+x�b�)���7�|����Ӎ��f�<��V�G������+�d��t�;F$��B*	H{�JGJ+��#�����Xr�n{=�\8�`��r2{�������S�i�
s���S~cẗ�t���d�Na�E��p�.Mj�K@��` ��F��� c���
uHf�A�|~�J�VxC� )i�!�Z�GGb%mI�;�Ŋ<���N9)�[��YC*�kY�ʐC���J��,�İ���p�d\$?� Bn;��41����BF�$�@<+�B�	�1KIt^Wx62xD*^�x<pŰn��@���wϟon狣�~�c�]���4�٢�k�W\��i�V!��ް�!
њS���C�q3��N� RK��G'h+:7V�@��_�u�Af�94Ȯ:���y@���$4�,��P�M#K�f�@^+23��y@�"RN%Q�ɈH�����V2�� �P�,8��i��[I����J��Y�<C#Ϛd-P�iL=;�a�ja����w��Qk�`�/��fw2%�	ˬ3Гo���-�&��S�8���}:m�%'�)��@/6U!��-�'�[�����
9]m麁x�;h��i�@�'\��u��x�!w�P3
�w��o��\2h����d JLw��r��s�to��)���9�&��k��j�Zl2Ǖ�'W�:��+�nf	�J[�S�38�%���T��Ŷ�:8)�!t�D�v���	Z�=�F�J�5$��IQ�&K1R���JQ06ũa��y�)7|PPdPFB�cxwڀ�7Ң���� �v�B��4B�In4�{���#�@'�J2����4�\ D���$���ma� ����'�Dd(`��8x^�� 3h��=:����1���������k ������������ӧ�n���i�(����Y2
�\��_��5�������1�kP,*��	�ٸ�7�'�h.//���16��8�3v��Y�Me��~(6�r���4
�ȕ�+����^���l�,�{��� Ɇ#� ���)�C���z;�\�H�x�V� � \�T( �/����3����6ς�'���"�����䄑&�dh��\��D^�*�((���\�'�5���t����Cm
/Px����779'���Ν;���8 TPo��N�EA����fpd,Uj�}a���)���bV#��AAUɀ�4�z��fGQ`n���7�YC��0RC���+Z�\zGE�4q&ۘ��l ��Y�A� � ��S�rk2Oǖ���gƵ2�q(�@#��tB[����X�[��Zb�e���἖2&π�8&�S߽����oMu�Wb��2�om2��ּ�
��4l.�����I�9i[
@��N��Vh�m�'M�Sj`L�2�_�\NV>~����ɹ�:�x"d6�n1��4 ?���"��׬�j�-'%BDi������}5����8�Ӊ\�...Pl�>�{�]�_A<C�>ʘb��͝Py(��f�@e9�v�p8/C�9�2a��X+7*��J�)�v��jp�n�>�Ÿ[������'�|R+w��ƨ<��o�M�ݳ6�\�|�B	)?C57��һ����ч~���U�!���ȅ"�_�ʇ�lZ+7�⇄��G��r������=���a�@s�^i#+��"D�,U4��؎�3�^J�5�N�	�iBß�܍�C��GG'��Hiwpe��f����˙Z���R�� �lP��{jD���f�d�:�G��H�l!1'�P��}R,_��{_��W\�Ф��3������D�{w��]�>ṀJ1d���[��s6L�t�#�ja���o��3ъ[�q	�OS�$��K�7������ďIop ���_H�m��ոm����wV#o=2.)b7���̵ˡ��QO�I!���ٳg}�������H�LV�.E������G?"7��˗��L�=�\ko.d�>(�͓���ʟ�9N.V@�5��Ƌ�V��L�a��>�����~�\Α.���!`A(J���A���=?��f���EgL�
1<�Th���hr*mĪ�xym3�1�P��\���<��|A隥�1�"�g��+��b���c�Y�߈�AII�'��.��͢+���H.*XteҊd��~�mzR�	8����a��C�K�m�p&d(b�}�l1'�B���Y�tXL�Y`��_�|-� �Ӂ o�>(�؈�S9����=N���Õ"z^��E�����+�gn�����b�B"�K9��p}��������G��yzE����+�>t�,$�P=6�_�'{�*x٢Q*�٪b�:�yQ˝����J�a �e�1�'�Za���q��"��8M;8��&k�X�.:���-���~�����tx�`/H$J��K�j{{��#��d'h5���Ł�V&a��#���t�����Ç�<U�g	2�;\&=0�{*Ѿ0f��C�:d-�e,���%gX'�U��>8M��p#��U�׮�B����:����+w�Y������s7�?�N�Nƛ��umw�f���$���T;�;\�gv���ĮysZl�{�����������5� ʂ�N���=~�����y_o�o�*�q��o|� =\��v�ɠR���yKF]ߘ�;�%�o-�7iM��B�If��$����	:K�p(�b��n6:��+g&C���]�Qs�An?w��6W��L�mt⛓�bQ< i���BqA��il�|aZ�#����l�)��2�m�Z�V�\�E�䅩iy�A济cƛ%r^��"3@��$��|��Y��Ҽ�RqB�u"C�F6<)�4Vm@ڎ�z0����%�F'b���$�85ጘ,+
��έ����:fS��u�� Qk�e1�:��r��Wp=�7ǆeRX3��T�N<D68��-yJ�fx�ӕ��Tu{5��%b�����,;�{�;c2��$Ђ��n��4}���h���l�4�;gIV�1�'s�u�x8�Vϟ]��%}�r�L���+^5+�Д!6)p�)}2��<�����(����� tS�i���		�~�G�yc
�h����>�yP�Ț3CSY��r�!��JL���Ƶf�t� �9�L�ơ.�2-x���X?��%����s�uT��Ir�$�Id�p�%�U}|z��t0�
y�`s<\̮��f8�_��;����σ���YK
=�5�4��=:&��^\-�w�z}���9=�a��>��Y�\mlmJj�Pװ�������Ͷr�ɳ�E��n8�	��,R�S�&�x�'�[�>�M���3�Q(�<Wl��8\N�>�r��gSV	o�P��t�ȃD���
Sh0sC7�K΢��^�#�$!���
�xB���ڔ�!�O�������JS��g�wn��=�S�_���E��{�.]����>����ׁ<`��)��3F��@�(�1.��"x�l�߯���gۀ�2�� u�2��̞3/�h4(�Z�рF�E��[�/[3c�,�2"i��VTpyh@��

�*H:����)���ȩ)T���%I��W�8�)����Ra�o�0Xurjto�7�R�T0hH�5
�dU��u�l�zd�'��������镏̒m��5���G�P�X�^z"R>�o�f�g�8��1��+sL혘F��C�'7f��pͿ��W��`���c���r
B�\&?�cL.ί6��A�V���'�>ۜ���'-"�\Yz����O?P��/&g��_�WfA���!ØFrR�X�#�N�ޝN��	E�l�
~��C (����$�\W�a@��j�i�|�Xqk�tY�P�,��e�-#�K�I{���U�t1p����@���Z�I|��!��ݯ���o{�9��o���;��_��9��S��B�DI@�b��>W�ⷍm㰋�)
�_LBĨ9
����w�����-;�i<J�9CP*g^����W�L�<�;�2�/e��\.�ˋ���$ȡ�M��fi�><vG�'1�X�+	fc�O�4Biޡ��2łt@!������d6��|��r~�<�F������dZL�	����<EZ�m6C�w||�W��[��x�ьZhz\�\���TKB���˽,�������Wx3x�8k�Z�&�I)�+�j�e��f4��jgs�oM��|v|vztt�����#�F�,)-���%:+����[,��'��Ul--�Ƃ,�,Y�"/*�4��)����fkU�kf�wF��t��,;vk�4CA?�W"0�?"��l�Ç���n��h�y��&re���~B��gg5�,8���W����p��ģQ�A�}����y�\�����e�%��{W�2�0'{�	��|"��@�'O�~A*v�6�4-�V̫������r��$9�IJA��%�')�Պ���g�������������Ý��bk�}�쒭���=���.g��VBE�B�ILY��W�A2�]T���ݝ!��rş��J�P���eJ��Z)�+�H���Y� �Al��RX	`�s�s�lI���|B�%Vm2��>s���8M�ʨ� ��߯.�`���7���e���˻�����߹w�4��ߦ[��L��Y�- �>c�9�d�"�F1@N��UF8�Qsl��|x�|I�m� IM�i`���?�@%3�Jcrv�Gb:�ЅFر�M�7���n�ЯKAzO�G���|�L����8w��85���	�&-q�|z��Q�!��Fa6c��\�v���x��w���&�:��+�a��q?���QA�v�Ԋ�����[ۛ�[sm��p�Q�G\�,�Ԇ��X�TX"�L����k�5���UzQ�_,�e�i�ֆCi��ǵr��b�����^bJ�.�S����������Y�(�Ӕp�y�&P4i�N�Z��tYG,��A�K�]Y8�L����m[��)k��hqf�t������yE7
�v� A���EF�Tg�l�4gU��TVE%�a�ɚbS��E�HO˔YΏb�dd}ɖԊ��g_�������B<��;�.�G K�p_��p�?�Mm^sOp��j@�#� ��J	�E�`g������Ar�C��8���A�ƭ�)
N�I���(��s���<��qt|+�P�� >�*����]T ^��&f&�6¯�8���~���$S-.)W@������G�;�fߴ�Z7#��1����~������`G,&s�"�7}E̛��ًy�\xH���uay4UW��l/w	�k&>����2JxP[�J'CTWNy�CȝDaM�<�:;8~c��{@�oqǟ�c��&�����
��<Z�X�ւ�%Yb�Ń�].�
)�F	O1�{�.cgZf7�Bࡄ�i8����O���b�Y�ٹ���V�A�����(����b.G�)j*N��F�z�ќف`���l
8�d���P���#� ����8����Y��>ez�[����9R8�`��U�PA�`��a��`�D!#����ZAꐘC%��v?d�z�'}��˗���J�UJ	9,�n�$�v��q&��`��3!"����x���l���C���-�M�~� y64<��$�K&A��h�_��I#���7cP�$�8O�D!�#������4s�N�%Ut��;H�4�E�Y� ��eXh!."Vs��s3�R�31c�$Q���!�˅�2іp���)�w��a5v��躼���C���EZ�_}���ݓ�Ut�.@����-#���M�K2\��wKU�J�\+Ny�Z�E�r0If!9r8�������ݾ�Cq#}�<&s�(H�5��98�5W��W�}E11�Gg�� ����~
�*�k��Cߨ{��kYDC����ji%5��*ÔyM0[�h�
 �Ri�3ՆZ�2骓|P�E����J��G"���'B�:��<|fȿz}5��506Ċx�p@3�*����@�������|f�L�\���,|���)��g}�	��L�8Y�$k�L�k�x�bD'���P�)����7bV��SF#��cz�o߆�����ɓ'tG��lعM�^(�}��a��bU���"+�(��{%�!lD泼����`�f�c����LՄj��R���]pf#E��ikh�w�}���}-�l�'�(�d�ԇ~HgP�= 	� [L���5��p��Tq��EӇ�¾_M�1�?�	l��4I�����t��2n^J�q��Oљ�s��b:C��|�FX�ή.i��t��guY��!�O��3��O�"��nq���p�-_֨�M?�����x5����^�ln�s�`����=8-%d ڂ�y8�A(��"n��4l.�kC�ѹ ���x�5��Ao�;�^�ܭZ�{<��PqW� 9-K���X+�^����1]��;$�ي�ts{��qe��'���'?�裏ښ	�3I!AQKB���X4��]���oۡ��t:������ ��ܼ�i�L,��b����<��u���������".����W�8==}}|B�ǟ|��_4±G���u���F%s�X��{8<�1�,�v�h�'�TI�E����T�����*Ze�ʏd��Px����M���@���$Y��f7�v�N���@fR��	�����/��P��Ig���O��o|��U����ѣG��`.(�=�8��O��"Z���Ɖo�XZ�VY�$�3� N�B|L܌X��M�7����@DYq��67��+$��r���t
M�u�K�+-����{�+�R��\v^��f��QDj�f�����.�7@4�M�Wfah�7�:���L�ܖ���eJc��0�V�� �w��p���iѨ�c�U�I�鴦&��wr��R�X�IT])��g�4U��(�N[���v}�Š0Ȭ3G����-��Kk�\�]���!�(��:i�gN��ՒSo�<�L�ḵ�`x��7;��dB�e�8?Q�TS��l������N��Q�hҙ-���j����7�&lK��Lt{�erߕ���}f��<��IR$b�u��}����C���fO8��"B��ʤD5���+�*©�*@�Z�?�*>����r:"��@���@"=˔����9���]�G(��f4����:�`0')\:n��8d�� ��e8T+��^@
R�y��d�p��ɼW\%.�}��p�	e?��dţ�3aF +i,ȳT\L;Ŏ�nzM'��j5{>����_��p|r�X���;/^����x�I]-���V���Z'(�sɯ��k8L�T"8��  W�cԫi�����In}
�՗g�A�_Ud�	�\	A��î��kR�&�nh�#�4�G��q�	��P�����GH�dT"o:�Hn>�p�!}�F�ϚٖM��g��W�Y�U	{q\|:���<�ׯ�U��H1ĦS���Ԡ���D��yH��\�Aě[��[[I�;o�|�����%�i���f�k�+���(ObBba82R@JO��PVM�F�,3��G�m�̬	�Ed�L�
�h����M"o��O��вym�Huƴ�M	Ú J���#�E������]�l���idN�'=i>(-��p��۪1G$�8�8:�Z� �P�B~y.(< >$�JR�s��݃��n�&�H�������&�F�xp ��/e���p�׭�5U�0@(P�ز �Q���$":�{�k`0�;�(&�{@z�'��7�)/BY��vjsJ�n ���^Ϧ	����(r=�8���f搶C�&}-�p�6!<|�,+�0����3�$!�XXI��,p���Y6fPgIn�$��xg��׵�	h8n���v1[^r钒6�4�ֈ�i?]��Cb~�l����zi���vPF4�o5�P�E�X��n�~�a����a�I�����}���ͧb�*W7���0K��-Y5&�eIS�=-��,s�r<�#ưǪn��Yr���ɱOBMf����'�r��L�03�D^���8��A����\g�`�q)���@:��y�@��b������0�͢D�-���hӜ,0g�#"t<==�t�6����&֪q���n�Mt��T�3�ԕ�G^�"�޽�������o�\���rp{�������Wҷ�kR�1\a">8�1��?L����-�A3�}�8��BMy��߽��������?{t��O~�>��ٳg�e��t!�ʐ���z3�����)�[pMͳ�2ٕ`����H(x��P\P�����'����I��!��Z�N��OϾ�������t�`�>���CT�,TYb�E]B�>���O�R���k�^�J�C��+<���:4J�`�Ii�۷oC��uz~FW���z뭷��d;AH��R�G>wݝ�6c�N.���I*�D�'��:bgLt|5[���?�������gQ2��Xۚ]�(�K��|N6��n����4�!�Mf�������p��z�"���ڷ�~0�� ��j�8xP���M�%�7���.:�(ڷ�"m�Z��(�qb���a�CjQUV0hYW���U�F<X5l\�ώ�<y�����5��r���YaP�C�[[+�#����t"]�Kn�H�B�.����Ǐ�x�����իW�h9YA*�(b��J�_��1_@����ϘsN�-��=��,䘔u~uI�ǔ�Y6��臻�H�H�Ir���pď�2ᓳ������[{_y���G'����g;"����3a�"��}��&R�y���V���,c\�Y,������Dq����F܉"̾��i���ԻE���V�E��e,��@����,pڡ�?`NBۡ$

1n����\�n�_�	�}����i����X5��O���O����@ʀ�����
�b��˫���^/�^�*�UӒ�%�+�ۼ���M��i�f��Y9 �t��Ƙ-
���L�0��R͌wVA�{��&�O�՞���N��o���_W�yk\�K �
�3�S�L�8`�&� *��/��
�%�#W��$/>L���"���6ĵ�\�l��\��P�bG'��/�S��w�+�d]jvhA�e��м5�Q7`:��K���[�;��uS�L��Cj��.���o��T����
�"y���]���RE�Y>����A��:n��T"=�+I���ǆl%5ˋ�B���v��xh)K��:.��3��w�
!���L{OR��r��{�l�ˢ�D��l�,5�hCt;��T^v6,�doK�T����k�/v��p�Λ6D��i]6���ag�
��^(�Y��׈�F�Ä\ȃc'�G������_W}n�1 3`�p�际O���59@+�}����Va&����>�(��,�7�`����i� ��F ��w�&!����o�:����g�v��Yٝ����e�l��+�&$|�J�|$��S�<�;�jt�'yS��id�g:c �鷶x(�ĺ���x��~B�!������=�m�j^faMj�]m��7�;���B�m�"�
+�;�<�LeZ�� ;Rt�\"d�\X��4! �L�� j^�ڰ�N�.1b�򵌄�i�ķ��{�h'ypv	]����NE��%'=�sf�'4��a�f����vsY�M��pbb�bZ�Re�����m���S�u��y��0�%���3�)c����`P� �څ^�ŉC�[/��X�T�0����׹�a���)u�:̃3������
w�;�"�r4�tT����d�'�3^ɠ�\[�p���C�YZp:�X%�=88 ';n,zÔ{� ���q
6WB@�b+c�7�Y�3D/(	1�-쾁y��\<�O����!7�4��'j���eF�w�EQ��NHM��CS��,H�N&���Xm����,�7CB.#u=~��*xa�p������TTQ�\Nzr=��r4N^�,�$�F��S���t�e���p�,�UE\���gc�H��+Ӣ��uKHL;N�STl����:C�!� c�ٍɬ �=|No�M����!��wD�Z&��N{� ���X4׉{�6擇I��&��U�r኎ ������2����"����K)�|������.����x,����uww����1��fB�
4��LD��<*(E�%0S\�Cl�)��`�`�DKȉ��Y����؜A�\wZV�N�D%��b��V����A֢ٚ%���Ǜ�ǉ����0�v��ٴC��c��j"�Ê�|c蘮���~��Z��":�=!��<�Z+��.2k`|"����
���YH3��[�'8���U�ܚ(�������=�������9
l�"��M��%���t+���Fv��B�\��Ҝe����&��:�u��+@����1�t���!#5��b�?I���?�ޫ˲+9���k�We U �66�p���F#�+�������GZ%v�j�L[��( �3+�����v�=դ8M���3o�{�>ۄ��:fW�6�V��U������p�P�MOA��������=C�"��5��Nֈ�Q����+��hA:��m�V[����b΍�dp�M���}Z�n�=��K������/�l��2��8��E��reŘ讇r1��W�!~3�H����/��~�O����>�]��p�<	pz4d�!�L�GF���@)C���@�$36�K��X����	����.m�7��6��d}��G������������4H2�����y��d��w�t�����͎��t���O����o��?��IK��رW���@N=^�K;��!��dYR�;y���!������l�ƥ�Lx�3K.7�L��Y��pdH���y��i�:}\r��l����x3����7�T@����Z�`e�V:F%���8���q��+�c{�p�E4�r�UbY,�������f�J�4M`e�5s���/��f/��q䯍Z�)h1�����CV�j��ɓ/�Ϳ���2��@z�>�|���+x�f���)@aRS�5K�_��6Z�B����ȴ(�t�oSt~����%�Qc�ֵ��lT����5-64{��n�\��6T�\��Ф=�m���춝��`�� ��D�@�7��.�}h�(:��ȲLV�����FX��� ӌ:gm[�"���``��ޜ�C�P]H(3�1�����A;O��������~�����58��<ѬdL��M설�Wh�-�0�a4���p�!�����2(w@ �M�%�G�\�j��c)\��O;���8�ɚ��ih�lt�(ݾ�m�a���ܺA�ǉ��4�0tr�d�*7���_`�8�"�����o{����e���Q߰�j�&s��A�<n�6=yv����F�T������ڮcI7��O�3!cY?�;iX2�L���,{�/�X#n�'�@`A���Ɖ��-�_���\�~���"mM�̠LC���5,��7���X,޽B�ҵM5�=)�M?�T�����;w�,fb t�n_�>�(L����n=��ig��PB��2g����0w~6*�z��^/
E�E�ݪ�������zM�{GQ�y'���I��{��$�e�,K��6��9��ɯ�&���9@˘H͔.��i�)� |rE�q{x8C�=O�����b��KV{Ԙ�������꘷�;�\Dhdh�[)7v��(��i�r��Vv��2�Uִ�jM��|��˓�#�dy�Y���ڿ�>�#�ЙL0�T����	�I*;wM�#�-�3����9�8���Q&uId}�mS7-��I?�ш�q�]�6F3U�	�~�e����x��
���g�ىcR!3�.�b`y�h�4���L��iݷ�Т��������O�Ԋb¡KM��H�)���A���7����1��F�;�A9�R�Q�� �CzLo���9_��pN�xa`�H釻w�P�E�|���}��X�������E�9D��(0BZ;���G�$�KNDAPZĦi7��DX);5����c�4Gi0>��8�(�F@�0$���q0�� Y>��3:�$qN��A,K^�6�B�X��2R��~�3Z��̼C�~&<=�i�(0��2~.�%H��.�^,�+]�T�Z��z�w$:��iAP�4��jT)->�
P٨e�<����6���2>��9�f7�`*�}􁤳��|4�W����	�X��,�^��!���~�Gu��^ǫ���BP��E
]g^]h4��<3�e��G��#Z�$'v�]�*������:Q(f��>D&�w�y�dL�xD��v�xJeP8-z��z��v'u��8>9����}:n?�я>��'md%ބ�خ��G�-�2q�z�
/��U��!�)}v�Y8���d���$���O���x+�$$Xh�C7x�����m$��0�E�
��ƞ�r�IA�V�&-1�ϖ~��tzuu���[��Uw"f[sED���t/5�<�!�O��6�����l>U�ߙ��a5	e�ױoi�����KøZ�����$<��!3���\\>��{qEX�B��n$E�ڹݮ_�x�U\S2�pߕ7���c�ȩ�̥tvzg6��R�Ul����t�O�qf��r�G?�N:J�d�T셧"�ڐl�8���)���xsejT�@��S��'�FR��0�sJͣ����zt�?��(2׶��u�]��]�$���w� ���`�Ψ:8:<�/j�>���|p�w�8<>���S�PC�¼���T��4_���i��b���[�đxSu����9�l�TՔe�^��ȉ?���͵���&J\�U瘄�WAr)c:o�5Sl86gS�V�$�\\X�]��"��#�c�������������������~���_���,��|V�<�����x`Vx��5���-"ÍQ�E��Ш�Nh�"Q{Ӯخj؁����j���A9͝= �	�KaG�=?�6��7��Zrh�����>}z}q�6ОIQd�yU�l�X��'ji�nS��OO�l��v�+߻���}�Ng ��bH��fh���T����QRт�>�j�V`t�^����0�DH�IՀp?C:��3��ɬ==e���٣��;G��R�E玾��v��`;�&�/ Cƀa�XPK�p��$�/��X;贩kgX����E^�cN�V~x���=��(�� Ȏ ��s�{M��)��!��>�j�V�6���,t`�SN[�Z4�
��eЬ��mc�F]���HJ�6�rT���Zbu���lG�%	�łk��(�W��D*����n���Kp�{�H*#��f��&��M1J�y�J<W�4y����ϛ+$��".�
A�����B�T=k�D8g��p
J��J��������y�,�l@�bH������w�Z��Qd&����J�Q���-����5�L��� Sd�ִ?}ʰ�ѳڒ��U� E����{i"s$/�kX��qe��t�CϳW��к�7�LMG
�!g��cNl��ug_Z��!@��D3�z�ckJe�>&�V���},��� TY��L!9�w�F񢢥���|�B�����/�ɠ��&�$.�X�)D��e�k1 �Jэ?��g��B���L�w`�:����;�lL�
m�d�A�-���=E������*�C�m�,k���B�$�>�@:�:q�RZ�vp���ԐH@�VJ� �5�������;����w��0\�%% �P�0�^��s߫2`{�3HX�#aN*EdT�N(ɢV�a!,��	�4N.��'!� �!��r��͟��ge�~�[���"�ĸ�>��B�'1���A_��q��)ζ�]�|���ݣ[\�2������ʙ�9/�. ��Q'�=IKL=8j��9Bx���%�,�Ҝ4L�͏Њ+��u��	Q��Y��w�7p5:O����k�w�c����Ha�&�tO��4�=��'		q�IBW����SQ�r�|R�,N�q�c�:5Hk��hx�����$��1����\+��Y�A:1W02֨�n'�k���^ܘUH?�����ggg�M+k���(Ӭ �^D*M��4]�}�1�g=K�о���"��E�5��Oc`Ɯ$4��cI���1�7�q�4Fb�P�J=q�F��G<	}p`��+�J��)�d��j�4�$��,$&$��Rc8�?"�>AR�$��Я�����M�3d�uBxGP�����e�����-j{������p���ԫ]�=��r�]���9������:�Ɇ��8��i�"�8�s��#k��x/X#��I�)]��Ow���d�",�-v;>fr���R��xrr�⒘|��D�2}��!}���u��@Yp�S��x܋�(�k�U2�J!��
Z�  �.�i�
ާ(�\C �>@����+l,lP��V�3��' ��m�3#���W.<���vX:%uɔ'�4'>�|m~�Ls��w3!d`��\���.�1�1�Y�]��lA����N;���e��q�o��ؑ�Zi�<&�?-���^l���CD�$���z����������_~�%�~(H<gaʡ]��1�۾�<�~�lxR/&�J|`4��\�ʦC8&x���p"�R��m��LiO�C@�j�[p�yT��1�j��s%�}sͩn�(5��N;�a�Ѐ�v����/�%E�w;f�ߚ��9"�]x>S?���_�x�+�e0�ڽ��o*��=�J�;�s����dݐ}�a��|��g�z�.�-��|�I����p\͝���\d�;�xV.@�z�]c��;$U�����|�B������x]�޼��ml�\ne���J���L���/~�y�e�s���a1�7���;�R��l1�:}���]�4Q#�xj/�у��9�8�(m�-��i`h��Dָ���e�q�7�%��E�Ť7MJ�!%cDk�K���Ǐ�P^��o���cT`tJ
2�Ա��B���o�
 �:E����c�WEj����������C�_��_�R��=RQ�Hy޷�~/����� c��k�qc��ruC��­��[���鉉G�,q�K��z����*dR��[��k]�vy,^F�N�ʄ���]���؊�/J�
Y�D�Te���L�0$�/��<��$�
6�3t��.mu�ĥΟ�Rq�దO�����B�$�+���$?�s��fϮe��*xN�!��e�p�(�.]�(`��fkSy\�)�?��^����t���9jTP6@����,�4����=��� �b:�T@<`9Ȅ��i���SCMyM���4/ck����AH���>۪pyi��N�X�>��gϿ��?�ï��G�y�����9q�ԔÞ����%�&FU�3ca[�K�e԰:N��H����6!8�%�8h��^aߑ#�At��!D�B)r����=��J�2�=�_H��Ef�w~��.�R��Kfw���JB2F�Yu����.����/º
�m��,6�60#Q�M�Y�8=E� �+q�6�Ak��fgn9�J������zA��.<y���xfo%ܛ���5-u�ΧE�!=݀�
k����z��=����!0�r����^ �v��B3�zm6�QbM3��lDC+�a�����f֛��Eu2�	��+$ Ɯ+�K�lM��p5Z�F��^�-, ��M�q�C��4����כ�d��g#R�B;����t�<�c�W/���b��|�Im��0��������?�-уU��:^��#� ��*L�M���	�g��?�i�v(%M�h���m�x�ajc��[��ĞhY�y�x�V�%R`�Z�x��tZ�V����:�!�$��n�
���	������a�~\Mv���w���� � \6��T�D{��S�M,%���G{����+Ai��<��lR���7*���Mӵ[��Q�:�"6;fg�Eg�'3�d4&�p��ry��t��f��a�Ҟ�ʊ�M8X�Y^�̋L��9ͣ+�߼�Yd7�/NW��п$�h�J*w�Ď�ZP<2`�N!�	Lay9�ikf�\�hTĔ �0�3�$/�J�������>NZ�!T4�N�x\���Ѵ���y�$JW�ݨdX��U����RtT�,�A�2��<�@:hJ_0��]6�J�w�;ƀt�=���M�����	�w�9^��w�o��c�L�bB�߁LQD�>U�Ki�KL��QǱgV�n��G��y���8	���`{��+(��p�V;]H!ߝ�lSԽ�B�d�SwŞp飄��M�%w,1�/O�)����/���L<u�����w�;�C��y2�v�e��N2��C~��$�*�/GZ����C:����
�rb�� @�� ]���6�1�w�}�nJWx�����c~��Qh�
��+UR, X��QzXr��Tқ�\�d�[�c&��6=��`�eF��
Fm�	������ȑv���3��&�<. ��4��b6`T�.!�ٯ�~���IS������|��@�2�|:�@��{���}���s�JG�������W<Dn�+*n�^�'y�Ĉ$��d)ٮi*�E�W7�2�	�D�v[��Ɗ�����K������$h\|6�6���F0]h��OR�%Ba>��=�V�b ��i'��})V���h�X,�qy�l�f&��C��hCSe�nĮ�	@�\����Ƃ�C3wY_��%̻�<����%դzu���û������w^��x��'�\�1��93��`�4��F�3$�J�gD�I�1��nG󀓵4M�b?�\t�wp*���/�����#�
�,}������]�`�_�Ê`d�d�=x}�����]���U9�N�\<�Zi�dw0��?cMM�Zj����l<)|ַ��vq=�lV�r�-nNFS�f���O�|�].�7�l"�˶���޷f�b�uZ�#�>�;�����h��)4��׷���Z�2O�on�>��~���)���o�$YSkG��j{|\�f'��9����/�*c�`�Eyc�����ʵ��Wn蚬H[�3D�h����&�{^S�ɬ�,�FU��.�G�]q}���/��K���L��YM�K��l�L����Z�`'n(��	��n�4(��!��e���'<�,��-�`o���"����	P�!A|�o�qHA�&
�e&\��B��]�H���`NmRy~�!	����xI⟎hJw۞�C.�@�����λgg�zy�٣�˫W�.�?{L �ϟ�$y��)���tzxs���?���LЫ��㓹�b����c�ve�9V��{f@0���Я�4���v�,��/�YЙ��&+f>�
�|����w�L~���Mp"+����w;Y���]�~���)�%���IQ:�TN���i5=�@;J�H�e��g�D&Fs9=��Q5�#���;��$�.T඾�x}'P��L�7�	��kƳ���s����$DqI�8g���˪�HP��3�u!\j�.�Erұn%�H�ь��+�z�W7t4�5�W�6m�Wb"�Z�6��}�~�z���F���`��� ��>��!o� b������VK�t��Δ��bs9i��=�Q,���qo�so(s����zC:���ϰ� �feJ�b� �K�8�@^o�;s�>
^�7���F�;�@Y ��/t!��K'���H�}�4|,h!o��u}�ʶ� M<��,��f�KQ �g���Zb��h�M��Y��]�ŝx>bZš��Ԕ~�a�C�����
�<d��cB���3�i+�-�YA0��D�To���:"�|Y��o�$I=�����N�F���TA��ߪ��Z��G����.t�5�P�����$\%���R�������Б���chۉ똗ʧ����r���������O5Z~�5�_�n�bX��z�S�0
�K����ie"�7ҦB��Z�ӂ,&˜�f�J��2�� �)do(MCX#h�s�̴��P�����^��f�Pf��d1�\�HcذH��J/e�D�cΙRd��0��n�S�	���y}�c�,�>�[̒����Q���B��1N��qFJ�a@��}��Яd��w�l�� Z�C#�6iup8-�M�;}^(���Z�N�z��Ɗ�? �� O��:�4�c�c[��d�9+������Q��͖z�~5���X�j�\y�l�ٓ�Z[�6--8��Brx­Vl名���K�u��[H�'�}�v|��Ը.A^Uu�!K��I���v�W����Rx� � ���
z�Y�!A8X�
m�ea��>? �Ú"{_&V�{����'ht�*��a�b��@5ǶYa9�����#�d?��O����7k�9���p� XLU��8xe�P����Y����3��Ǐ��ή�n�<y�'_��E�ݍ4O�'�H��CJ���%F�yMAK9��F�/�E��amc�L�U��k���+[�aP�5p�̥1; �h��L�1<1hSĭ�!��=~��LM��&���r�,$����]�5j]c� K������*"��D8�=P�������}� mi�x�d��e�m�ul�#3�ہ� �3��������6��\�>��1����ׯ_�`@<�J���q��M06:��;��q(�E2=@�G��..��I�"d��%3S%��:k���?99甅)�y��W^��((�=9f	�	�L���������	�K%atJo�͉��|+5���2���
:�-���~ �F,�T��)=y�f��u	���Cd!d���T�'˯W�p�*֓���'��T��
pQ�6"�ĂzTa�d����d,�)��B�P3ڏ��LM<�f��Kv}}��rI��e����(�ȍ@��ȏ=C�Ҥ���� ���,�n/^�0>��P:�+�k.`DCI�\���=��@OEez�J������_�t�,��Y������1�I>	�"IK�9O<Iv;g�j��U}{�좝6���=�E�O&C.C����S����z�@���\�� "m�g���3�U�
J��ҝ)Oa� ��c~��� �7+��O�<��E�dD�خ�E#�54쾡zL�e���y7�
�
�Ǔ��n�'�*�M%$W����1�(�H%|����y��4�;�̭F���V�5a)+˔�>�aϥ�V�kJ&��N$��R۩�����iHq@=�5-<?����~��w���E�ꫯ�|��n��`�J,�O�]s1��\��FgP�Z~������ߌgc)S�����/����b�q��{NR�������ɗt�/�|��������Y�g'�ˠ����elXv�}�}���b����yp�2�Ϛ���e#�</�������.���� �h�Y�8�����Ev�f��eqsK;(K��\p��9:���v�Y;���%�.�s��+��v/fL�#��Fa��x�����K�ݎue�����*MauǮ�a��wd�0Q �	�
?Č��c�s�=��Ӊ��L��0t��9HZ
�z���^~¹FL*f:F	��M�q�c�_n��a��e3���ŝ��K�����-23�L_X#�ݠA�A��s.xO�o}"b����������x���!w��2b �H�:����&4��#'�<�,�)� ��ks��S�*7K;O4/��w��`���	ຳX*&<py��E���ـ-�8�kCG�Xi���7�"��[�J\y�j,$e7����Nz�c>(�*5j�9�2����C����w^�cj晄7{������N{f�L����HK�~!/�kg��>c#XBah	��S����z�8��I�,��(�ie���6�0C�r̡���ާ̪WT���1�����sJ"f�������a��A�N�Jm��o�	,��+���0t	��٠�ƌK�[����S��"�6*�Ml�� D?*uB�%N^��v\M[�se�4М���:�N���	�(Ӑ�J�����r#��N�d�ݪ�$ߞ}ȝt�̈́o8���9�w�¡�����9�	k,*��������蜈�OH��(�0�dB:�d�L�K��W^p��AQ2�T*]
�qa�R0R^7-ij�,��t�Ɉ���!�&�[�Q�R��y��g/lV$�9<79x����)c�<Yd@=t\5�r��x1<��}��]퀌Ä)>��5��Si|8<��f�������߅���������tT���[/U�X{�����o�S�0ڶ E���}5"yX���}+�E��JN�$����1�R�� g�d2B�SG
�`�Y����S�c�9�����RЦs ����c������{~Gs@��kw�\�����O�x�3MR�D�9f�W���'_�F��ݻ{vD{\�HH �d�w��j��׽oM���GB��]/Ṝ�<��"d:"��uq�U�=��������g}U��i����� e#M�#��k��p�[��|̒S�MM����g�6�\t���2M�F� k�'|#CH��(w�$r9@R���01�`���;Z%��3�,��Ç�wP22�?��c�����dp"yA�����L�L���n$Rꀽ�&�d쮶�DR�\.H�H��}	)�m��p+'���*�nId:!Z0�b����;`�&�&&>t����i�x�-#m�ED����fO<��D�O��g^m1�p�ŝ���cാ�,m#�	���9�Xt5�!"��	� y5!@��k�Z��N���F��-	@q58E�Rw�BD{k�Ȟ7Y�mU��'���Sˢ���+�%���|/�o5�46gi0:M<B�b6[�9r��%��'�1�Դ�B�h�A���Y�8��E�8P�i�5��DcftB� �_(����Js�0�� 0LM@J}����_��?b�4�u��)���X ��gy���9A��MI�7놫��N,_3����%x��حI��\���]�����p>���\-�m{����R	��ЮX#��ba����*`�Dc�
�����)2.$M��- �Nr�_>����↞��Fi��~b3#�DK�4�R<%�2����e���p
���q bK���w�%�N����D�M�j��4��j6����F={�	;/���\'�h�&�� ��"�QII��I�c �,��᠋���:egXMt��X��w�W/V|/^__�y��$�v�p��dY�FJҾ�wE/ݺ�(s@ȵ�0?����"ջ�}K��'f�J�ܾO�G�$]kK�������h�rn���U�:��{���ѣ�w�^�~��vˡ(ҡ�;*mM�k��02��R�4����D���?��`�I5Ƣ�d�Fr;�Av���֒P-����0X5�B)�✓Z����o��i��ӭ�y�Le`����򗿤�<x�������7o�� ��$" ny)�������-���fR��n7���,eqh*h�}��(�����ٳgN�q	?�v�~��\,�i�ċ���C�'kDgȞwZj����o�d�b�ݼ|zA�;����D�f�L�����իWA�c4{�~�)���͢�Lj4����?4ך?��98>�\TeZ�d�'�cG>�<W�a�w^]�D)ӆ©?�l:�&}ۤ�����6k��6�����q$�����E�Y���t	Mި(i����p�B�`.4��f�k��Z��\!��Tc.��YB�ӑ�ysuyy�	�Y,�4��@⮷�,/��p
�	��4�o�}{��"�I
����Z�C��]�xS �bސy�P�C1��|�[�R'�C�i)�&$�.�a��7��%��P�ӽ���/�|$〠�S�f�L��B�q�N[�.�u'�Iưk���SR�Y�[r61N�Hs��})w�ԫ��z���4��>Sv"�H�5�u�K��I�BpH|z[r[%��R�n�N03���֍afV\�q�!�6�$�B��+�)}~:������a���mK-��R�;���(�$���=�2B�n]h��\�zϊ���P����k�o�fz�./Jϻ�f�IK;�&��jH�s�^٤��\�`�C�qN�� �賃s�g��Q!<a��=�������g$���`Ԓ�˾5��܅V�a�����Y-����}���K����JއM��Wl���9Kb����BJ�r}��Fm��� �h.���rN�޲)��`���&�B��e�� eWT̠s!W�_��h ў(�1!��+j��i�6(�w/��K
Ջ&蕢>S�^a������I���4\ig��C��d"&��r��V�R��r|v�+H�+�k��KD���B(�C[�gm^ٯ��
>��e�z4I��c+/������UQםMW�J��1��}2��R�����w70V@�p$�%� ZɆ��;�s}}��c���4��(��ٳ%O�������(hW����[�"�����7c��j����>���p��=z���������z�X�T��V#QF����b�\	9�N���o?�d�t69@�!��jޭ-�����8[���w�⭑娐���Or�`;V�r���N�P����S�e�0D��^�k+wo*Pt%8�Va[0Tb�S�^y&���A�g�Y�s��Y�U6�@�w�?��7i�и:�8M���A��{��qh)/�Φf��/^"�g|4a�:�b"� C�k�-�X��E%[�a҃,<�����	�N{F�TM�#�F�Z&;:�e�26�N�nS�p$y+��.sb�$"0�B> '�)p$���<����Ǐ������?�1��Ȏ����&a�/���?'C]�sBX6�>	"0<�x� 	�3�|���2[�>v�W�^�(	����?�i��8 %U�JF�@�s&H ���|<�x�p ���NA�wJ�/q0LmC?��[f{�g�%������������
mB���9�y�bU��N8�-E	'O�h�x��Ez�ZG�P?�|ҿ�Rb��8r?�K&��R3+���f�K�}�31d�p��&D1	�2ɾ������4�yOƕD:\�|y����j��pq�HF�Kܰ�NS�r)7��ze��W�V(S�]���)�C޵�-$j��N���v������?���|�;�f����si��P��K	g�L��m�ݾ[ZI��J�N
ͣ�"ǒ66ݎ6 V�Z`̝r,�TDkT�f��OM�s��B��-�6�L6`�����T��S�OoSoߥ��a�&	���CtZ��[�7�I�e�\^ӮFs<s�*m��j��8`?tZa�6dfv ��d<�ү�;:ht�;�S�d�qA��Y�8�_lna��m���{;.��Y5RyW�SH���i��Ϣ���a98�2Z5��J_��rj�˩��0�� �$�Лr�� �t��4�3J�e����>�FY�	[D�K��ʹR�;#4l�A����$-���G10s$���RS�v�`$�C��7�8mT~ z�˸ �M_�f�f��l�-q�-���u_��Iք�e�����������dQ�Ơ_�]IY����q���A�R��,O�MS.*d3�����;�4z��;�'7��W�E��Fp�����I����X�����
���ko�0$���⠈J���^HE����Km�'̮�����%#-	��'O���������S�R��!W>���Dv�a4et�;�VB40�BO�i�D�i�'�oo@0��}xѼD�/��ӂ��&@�f�x���­1?:�(�f��X��/)��`������'S���D	�Z��HK��K^?/%��Ԇ�������>��3���-��@�!�ْ	��5��"<X5��`�q�*� �
ZR�l���a�l�X�C�bR)3�,CFĜ}���n
��^����_al�!��[#Wr3���������?#8$��â�<2A��4� ���"�WW��W�6~��血l���6��� 2)�Z|߯9�|d a1_��+�d-?s<#�(�����,�b�?�b�^�?�
n_g�� E7{���>㶼�`��{���|azA�a*�Z�5�z+��u{�����l��ڴ��	�
�h��IG��B�=/���L/���X'�d�3~%X{Q빺A��ejr�Y�y�m����s�}9i����!�q|q���o�����}y����Qk)vgz��[��a��Q7J#e�����_�������a@�f_�����r��	hW�#�S�;��E���y�A�H�<J��l�D	ћ��+� ��+���?�����0+1��ז�X�F���zq S�-�)����ܨoZ{d�ǤN��&lP8�#�y�&�_�Q#Ԉ8�)�:���{������Ȭ_�W,�k���~�W�hIĥX6�m�l�^����� �+ѓf�9P!F!׹s����)�y͑Η>'��F�\1��9���A2����-8�Gk�@����b�۠?؋��	z&\_/����%���UZ��S�]�ӟ|�6������SkHgk[V�EͶ{s=�qP;?��d��ҕ��k@��9w��.6d����m�7W�U�E� �$7��o2�y��\�0�))B����v#��[�ѵ�w�!^�D� �[hM=�n�r��'i�L�m��۩�d﹫�]�n$�$��DI��c"B����������=?�NS
OΫ�PF��g�=�"9]�E��RO&�V3!s�!3�����,G�#+�?���G*���Uo���{��Wo���q�"��9A{M�`鸿Vt��DV��Ȫ����L�bO*���y�Ȇ��'����J��¼K�(��\q�G�� k`��_.& s��*�|��MFl�,�ʐB�8��,����٘�]��;`܀��U1M>�k&�L+7@J� ��a�5���� >�cHo�grWr�ّr|�w�_ě�3��Hqv�� ����*_��?s}}�b�N���v�r<�+����9�� ��$a{�T��܊jM�"�B�_iu��C��PQ���Ǐ�ЉwM�K�p��Я4$�亥��޽��A�E������w�D�'g�	�%H_1~��E"Sy�-��}��G �\���ܣ��~>��!�[)�B�UN�\5pk�=�����A�߿;\��~I��M�ɳM�1�Y��F����݀�ؒm@>�����K}�7\�^0¥�SA>��%,�8N[�*}A��IY��)�ֹ"ˇ!E!��p�$���r���þ��Bi`�s��K7��,1Y�GP�w*e���$nG�[⛫����7����wk)��O?�����;4j�z.q	]�MF�lJ'���������(|/�IL�EiF����0�^�WϿ�SP/�Eh/_��.V���W�Lӱ�"R� ERd_��� 3V''�ܼ0���g�xME����o^е����A�(�����a2!�!���ZSd)��G����=��d<;���./�\b��H\G8~~�Dv��&�m�j�Ee\Q�}x;�+d=��Q+�[>�2*NO���._0�O �QR=�!��%���.�oFk�?/ju/�ޮ��g�Ig��8�8ѐ̹p��G3�-�P����@�
�jA$y��Y�H��t�=���K[	隰�~���c��N���# �P악��in;�8�%:z�l�vlPKna�Z;����|��	}��7��M����e�m:M��������`��?�w�jgggh�
3��H������/�$��Bs!�a��u���G̓�O�����H�p�o�`��4T���vu\zuq��i�؊9P����{�]5D�]���$ܰ�۷iJ:��`���B��3��&ˊ����Kf������S�>�$�-^/�g=�@eZ�G�~�ZƖ��"�Ώ晏���?�\�Y����]�D@�^���F�D,�_����y1��T����v�&3#�ϊ���/��]����ւf��9�¸J��]���#�c��o��/..Z��1�;�P� ��n9���� '̮.�G�>vr~2y�D,����-����HQ:XQ�`$��S����[֒ca��rT��E�ק�J~Gࢥ6$�n29���ˡ$�B� ���*��c�� V�kT���_|׊ՂR�@k�.�mI��}�s��0ۦ��̯���FМ>�h16�F���b���-�҃1�Q����M���W�����4�yr$���v�ev$Cv��W�h��ŗ�޿zs���H�'0u�@�p���0��3��K
6rV>/Rk&�?�T�!��/���ᴗ�԰V���#�`�ؑ X6脹�H|�4�;�\�+��WsIx{h��M;�W�
y�<J� �h`�ơ��]�xF�R�-��;�%!�C�
�0Gc6�,�c2��V��W�p�'u-�9��l�<���%��U��泃quL�@��n{x��P��Yj�!+-c�����7�,b�y�t�hy��E͐X��)�D-��K�%�Κ�sWpb)�U���>�y�]�]<*�0S���z}ف��f�9�@��7A��e3e.��Y�	2"(h�k��)�	�eA��55fy��^�M�iC	�$�:�߶qaV�=m�i�E�շ��Z���%�0��)�k���?�r����Uf�V�df�)��_>��s?�x��'��D�w[�p���~�0}NC�x٣9�%�Լ�i���R|��L�b��FC(�v���8�1�!�l��`�O�k񌍹�E���Jm4�2��y\D/t����4�-X#̱!'��R[g'%H�t����2� `��� M`�Є&����K���&_�Y�I�����,����R������ľ�9D�T	�l�f�mf��qX2E�N���=���
��Ҵu�Ϊ1$R:t�ɵ$�XU)�Nx��&���F�9��fXzo���*l�����e#S0�	X��G�jN�
�-�ßKΦ�3��
D^Y��i��Y	�9l�Z[��4��[Q���UAz��j���v�b�;&�mq���O��w��?	�'��ѱ��%[�'U�~F��>�`�M)�n����l��hX1Q>W�C��*�؈P@t��ۂa���&/�˹J0&��s��
�A�74�E4T|ۉ��F�?2y�'�)|�k�\���`P�a��C�A> 挀���\�0��}��gDu�Z��|Bz�ѣ�¯��i��k�L�=;���&X�ESI����YF�}Ea�>|���7������McZ���u�t�s�����0(#]��tYZ�4^ʘh��,�����d_�ɡq��}a.iz����;�b1�p�a�G�O������L���
_��N��Sz�r��A�Q�Y�h}i�!M��g�։�Z�'6&x찉3ڏD���{��h]��SD2yo�o��
�'D�,�B�狀mI�R&�!fc/�;�LiaїH<Jd��[���l>�'��Ï~��<}z�K�9��N�YnTC�L��,8�|5��*�0?u��Bw�� ��>O*���|�]�AA���a����ވ2�c;�Q��Z� ����u�$��4FqG+	-f�+�6=�9�S�����RU:��29��P3���Ϙ�cef�S6S�A��Rt/���3�C�#���'��U�%˥{��ѯ�O?��^B�%�"�R6l��ua\�.QV�W��*p�nq~���]I=f�2"���\8%W�v�}�xUS_�b��
��[M�x[vۄ�$��k�����ѸA�ߢ]N�m�в�۩q��8��nX����B,�@�������;����,s����i�f �%Q���Âґ6��0]�@��iV(�r*ltM91���
���|�7�ꁭ(� �z���{4�G�ryp�c��jƼ�lО$t�d��$��K�X�d��*��2*F�����d>�=�z���AF[�����l���9% *�^�S�� �\^*������>Ӵ]߰fv���r%M��H[(gb#غ�􀾽�I�� �	f]�����am�Y
K�� �V$���g�^�z�����1gC�݁e��f�L�\�^A�m����`�����u+�^�U�bc<����N�7����)��ef�&��ɔ5N���������PM������1*-�Q�H�P-K���	ږ�L%��CϞѥ2#��	K8Ҏ�V5��i��о��(a�`�������]�G7;e�5+=j��*�=Q�s{��U��x�!���O'V(�RːMA8I�����g�sA��]�'�����_{��N4�b��RN���%���vB��}��Xnv��Q�:���!LJn�#�^\_2����2�48��y��˿)W���YdfȊ~������}ƥ l?`������ xN���r<��wY\H���LY2���$V!)@��n7�@Ds�9�ZI�4�ի�L��Tc3&���w�?S䩦��oj��3S�6<�
������'��� ����f%�u)��]D�]���Ed:�9�d��1���� ��h9��]��g�e�`�1)(u޸��(^�!K�������>��4W�8m=x-s����R:,��ɒv��>�থ��e�~�'`�b[ۦ��);�r[��6�eBi�L!�pa���u�3�
�*����+���i�r,�,�MK�-À=�ng�XI���E���R!��B��i'��K�L�jS�(�W*C����Z�d+M����������T����b���rb�V�'秓^W���v8v�͡lK�I���%	V��@�$y�_�ա)ڙ�&z(Ecճ
������`��]J�,	x�܎#���w���ǯ�\���l�)7�ݛ��<;��(/2����Shons���Υ�#�p�9��%�������<����p��&�w�}p�X��HÜLv��wmh�޵>�|\�����^b���jD��i7 �i��>Ls����YJ#�|� �e�U#���<��	�(ǰR�X ��U��S$ B���䂆�/��K
-7fs�Yig�1�K7Rbr�U�aIOǒL+vb��#�������^ۻz���q���U^� CY���`)�t�ʤ��q5.	�l]So�]�bWeUp҉4�N�/^|Zr؜�|j��V�*�p5r�,�oQ9ɩ�]i��h8@�ȩ�'��)U�q��P�����z��jąG��h\��@��.6����8����ɂ�~@m��I@!��pj#�/Ip|�q��M,� -/.���#���so�)��՜����b��F4�=�M�̵O}�s-���\�v�K��4Wt<⛰V1-�01��a$� �\x�y!�
�b�@Z�����),*^�>��Aʄ��daW���I�rZ'MR2�q��s��`�q��_>`�N�� ?5
{i�"?_i�	�G�BB~E�PVH��HS��%�P���5q8-Ҏsi×��� NI��j�HΚ�k#Gܹ���C�ͮ&wt4��BoAI�pp�O�`�kr�+�������m-�B2��"fl`���ܾ�vg�n5]�P�~>+hJ����Ϗ��g���e�^�������ǿ��I����l�*�|T�㪘V�.8v������v%��w�*
�Z��6/�d}��g_>y�ճ�e�r�kZW�Ͼ�C� m�Ts��"�	4̈Ͳ}`��:h�j��tMz�YȢY祖�C����{V
��
�%sW�7�5l JVN�7���n��5۵TB+�lj�c8A��]�h\�oo��QS���M�������W'������������Y� ������I�<Bq�kf4b/��L�D8{A����Ӫ:RL{�==Y��=*���T`FB�J��\)Az�!߄	ͻ��MI���X)��,�vKi�5�ۅD\��WT��x���Ʉn����eM ��$���_O�<�|�XHrZߊ��@��FEB�\P@�K�ߐ�B9*������>�w��d�o�n�&���N���r�]Կ��ۆFu~��tF��z=OV����'er^�A��m�@騈
�=)]��t��f�(��{���L���.@K�9XAtnSm>}y�%�V�{�J�S�&�h>�j��O})��J^!�4�p%&P��fS��ݻw�����9�8��Y��h�V���;�eJ�NU�vc��^�l��\Q�E
�.��;t�#�>X��)��x������������Q��\�ޠ}UN[| �>���h7ϕX���7��W/_���5W�N(%��c�q���p�����������'�zW"�VT�׾��@ ҍ^�|A[���]m�ڠ��F��#��B|���V�H5�$�
���)���� ��,J��%�Ͻ��ik@,`iZC�qrŉK���̱�?��B`�K�#�:�p4 =
��ܶDg�hX%�~�����,P8�f��{�O�s�C�ʫ#i��ν~~	4�΢�oh��]�uS���J��2x��KA�d��	-rc��7>$Q���PӦ�}����/����ߍ���Մ#j��3,���x���1!%G��[,�ҁg�k�(pSyrnD�a�+�g�h+`>^b��ɒ�U�1ʞ>�ވT�.v�V���j�V�"`�wl�I���B����a����G&�2%2�$�x�ջ�����ޝ�)d�>�N���r�	�(|�$ц^qr~�l/^Z�)c��1*y0�Uh'��;N	�p.�;��j��3&ZbW�D���d�7�vqX?��ݠ]�16�y+s������:5m�a�Zv�k��٬~��V����(h�T�l>Øc�mO̳���aJk�5�oرl@:��}��`�1X[�p^�E�~�3��G����v"%�y�fD���D�c����F� 4�bs�
%�(�+��S=u� 9�cI@��^gìkA������K ��իW_}�U5��ό�#D��IA�����5J.!�X���ʢ?	�T,Fiz�>��y�ٞ�OMr�%)z�&�t��lt��NY\d���9�O9-�ר%�fӬV�|^�+��f΅Mi�}ٖ�c,m7z�O?�T6��ѣGVaq"?�%�P���5^���d�L����iP��/���Ԍ�J1y�VL�R&���E���`@��BB�[�D��'����HR�׸���f>�͡?����� ]�� ��OJ+�	�6���w�iDe_/�m���`vd�/��KnH*�	'V���8��;1x�L�00&@.6�,Mc�F��'��*p�q�U@"�2,��Ʋܝ�Xu_�3��2�/���!{�[�ޣ{��I�����9Cۤ{���)w�����ӧO�֗�.Y�
Оh��80ֽV�уÃ �Y�~J�U�P9�����i;}���d�D�	)�f�|�?í*���I�3�(��г ����R
�Q�%�:}��i�5��5�{Re�d_
eӫ�oJ�Q�{��]D�{%������k�b��(i�4r��!:؈��Л�H!�J �Q{��iq�\/�@�[�HQ�OO��y�� �+�6�RH#�m͍��p�+������R.Ц�!�����U��RI{�Q���E�/N�>�&=�Դ��@�4H��l����Y!S�G�P�`��C��N�gy�ϧ3<,_�L�hl���d��Q[�u �e�M�J�_cM���MH@0p��$�m�J2�S�x)LO���R�v��sh�v4��xl�ZT7$tpOoڞB�Y��=c?��-���$�7�������_�����T4y!a���{���VlX��i���\1e���_ܐG�nݩD :;P�=A& 	K֤�7S��C�̜@7hL�i'h	b�!�ù^��W�4akAL���C�Ls&e$�킘}�_R��r�4N��2@p%���ɝ�Ù4�ři����N��L��k��i~,}����&Yh}�ye��;X��[u�x%_J0�~OB�ƀ<�s4���{���y���ff,|`�Z5@.�S�����هh!x� ����B�t�Db�Hro���5Q�0��� ͵�e����$�.bc���@p1	̨Ƴ3Z,���'�s�R=ѯ~ŕqzv�,� e�@0��F8�� p��p�i�OL)����A_J�.h����#����ޣG�?><8 �;�v#��umC�h���$��۶.����{{K��U��ONN���nX5�]-;��$����n;:y2��}��~y�ې�qO옋��8K@���-�O����C�9�#�c$`0�@u��'������n�C��{��6�@2�F��M����]�=�Q�)k��e��-#�V[�H��x6[���J~�����us�=y��
�&�܁���~�!�8Z�������^�6
�j����D�M���M��b��^��g �F?�çw��	� c�T�b�����S�l�kƅ�&#��y�N޴�R3� �d^�i��<Ԩ����|F�=Ӛ6(G?�D��4��ر�B�m�!<a�����6��t�y��v���,���jձ���z42;
AU�+���������G��͑�O�&�gQ����g#�)�r��I��ktz.e�۵QJi��~��{�9d�=���9%LR�ˡ�q���2wH?�p	?ɹ�K�砐*�������53Z���\�V��k?K�l���,�Q ,l��@}��X�5��$i�d�����(jZi���ׂ�T��ؤc�ez��¹�3�!V���
��_�$��:�Ț	��]9W�f�IBN���`z��6|���Q�-{e��;y9��r��gԤ�k�/W��w��dL��>�'t w�,)��2T�W�{.u[HTRfH�x,N~��)���ݖiAr1�����]:2�p�\�����s�r��u	�g���s+.ru����a��ͥ��e�r$O� ��L��m�ܘ��4�i�*$�%��hw
�1��}���`|������5ބ�X���(_e
n�MT��%/I$�Bh�3� �h�����0Z�<w���� D�c���)����Qu�jp*�AgJF�p`�u�fM#/��vqsx.._���TQ�2L�!�7z�S�CB�L�l�$��+.���������-a��R)���3��f����l�>dy1β%	�ӹ��g4��5M2�E���f�M]q���.�xɿj��f\Ned�� ��nM6��p)!d4���]�4yEg��8��N!��X$�*�N$���B�3�v#M~&۠����p��B\8��V!�[�οz���2.�����w��"��.��(���	���_�<�|�}��!�&DJ��J-2=�����$��C�<g��u��Ӫ��N�懳��`J"��س%�-�ź��;�w�{��/�c�Ft�K�f���9==����͕Ę��3X�-��UW�gBvR[7dG�Eֵ=�~��ф��̋N >=#ѐ� �9���SZ	N���T���va	�^k�\��i9L6"�S�N�Č��W��9�	�m;�.�f��knHG��x<��E�4UNb'�i�ڮ�i;P�����x����W�M[��?��w��~1:&���O������E`�x���%T
8��M��[�Ae˸Y���\A�����$3�Ð�����d�p�3C��j7�z�M�炧+��b�������F�l"d��1�����)q]Oۇ,H1�Y8��lͮm�}��x��|�������Ib��������"q���j���助4�T/9�&xE�)�A��v��Џ� m�ٌ��o.��c���3>Ӵ-��q\��[\���"<�8�p��!2��L!n���N�"F�He�M�^�H�#������|!�)�9�!z`J���s��|:=��Fd�{���K���f[��n�+�^��_���UByJV���Il&#:������cj�ɏ��݇hx���&�-C����;w���"���rl�#�����e��O���&M��p����@�"����yD4h�wϹ�-h���ދ���������yQ�`�:{�Z(6�����O��<�ZBf$H��7�z�BH�褌D p`E"�-����1%~��v#ч	"�,E�����H��"�������r�Z�Zq����3�Yջ-�=������>���?������e��$�m��IX�P�<$Y)/+	�.e����W�(��	ߍ�"K���@�R+��su1&�ЈΙ��q(PB��{�v4l.B_q��H3KfMד9�Tܐ�$��H�w6�qp��$��$��fͥd�����#�?L�,0��?����^0|���8l��}B��7-;�~��$hɮ��!�"\7����vH�u7e�l2��Ӫ���M �oӇ1+����)x	������r6�}���>>`�_�dZ"�b+A*jE-���lnh&��+2��B��J��f�T��!��SbM`>��Mz������नf�mG�O�
H0��M+��6��IY��K.9��@�M���s�xK�Rsȕ�H:TyY�
;�דn$%�#9y%�Gd���Ps�]�bB���e�Ѹ�LG�t���$+�j2*F[���B��,�gR-�>��)��:�?=
ҥ5��[e@!�d$�ڐ��@����
�Ѫ����L�␯�]CF����"�:3S�n6���[Ҵ_����؝)�D��-�7�u.���qWfz�vH5��ꟶfPU$�?������]�s�ȶi��9�M�^��D-�����}2�LɎ�� y#;$'�a ��4�b�V�5�H#�����a�[��N��M�c�A��W /ɢ�[ސ:l���kL/�z��v�M]�4�� I��zw��PZ	L>���]~���_>}�G�G̋r0?�{�V�l�u�@�z��v��RJ[��R&L��c;�D�
�^�}�!��Mݲ�� J�L9���/�K@���ɩ���6L��7Y�owd,����nϖ\'�\�^����W���cCS�M�:��Cz*��f���g@��2�;8vm�z�ګ%�����~�Z~�駝8����$��L�̴�8�x�q!��CN{p���Vū՛b��Q�Lp �Z���]_��.������V̫�\�Qz����2	`t��G��i��={�<z:�!����wxq��K�ۓC �q��/ow����]�{HMfd��eq���o״��+�F�٬..^���5�I�$W��]U��z�g��@�d G��b������!h��N������d�A�)׭�v&1� >'��(��~�!�bTE��j�*�ZZ	��4���,72�].<�S��ӂsw�eD�DpH�X�kmi�si�Ǩ�Z�\5��}���W��=��V����w��)�(�D�?��ɛ��Rn!P��\F	��k�v*�MMAZ�dR�֐;�y5��钣� c��G��~�4V�^!1\ջ�x4��C�����t�Nj���-
i�պF��O/c�9x��aj��ud�>�<�����,�d,�1�I��`�Ф��Tl��F��t�؍���<���O��ŵ�����K� ����sr,�q_ 6����yfӢ���kj�M�I]B�uC��R�37��zB:ʱ��F}�I*�� �ث�jI έ�x.9U�>w2rM��tWpَ�������3ͻ]�lR�rx�C�Fr%�|;	՛�A�"�g�W�0��0�1��2����^BSK* hq�2�s��Sp*?`��`ڍ�n�iy���3b�;-�͕d!� �F�4�q��q�Zx%�d�`sTP�<]��H�)�a�L"v�0�SΤ7+�D ��S��������gÈZ�+����h�|I�3<�.J��[eWd�e��Da�����i���௒V���@;�b�#�]��i	���$S��f�q��+()�̉�ݤ��%�(LXL�S7�^�x�k6g��h4�W��e�X@�>%F*|Hn�ؽ���}��!���!�Ř��Y�����Q��岩��l��v��[��@9ISE�?���+���{��c��U#��'R9,���9;�	� �����,��zؿ�/F(��x�Ν�1�_.��L����S���=����a������dTn��v<&��z�񩶂'�������НP `M"
��v��J�F�N���.-ٳ�����߃}@���r|<˄�j2I�&�c�0������@L91;`��y"��?�5�B:�����3p��d�ZP�1�/~�J}�;�)�cEV�՛3�@�h�h�4���:�a��$j��N�X��R�B��i0���������7���կr���G%������х5F�3�ᜓɴ%�_��-��G?����:<��P�t����&Ȍ�F��ڞ�ci<�'EL�e�2O��測S���`>�5�4B�@� 
����O� p�B8 1��/;tr�P��ul�^�Bi`(˵BZCl2���8����f���4��)�5�%�^�+�	�"�'ggtM��"$�馐��ǂj���� ��\�������}������Z5j�c&�X��S�m��Ŭ��j�=DT��J����`��g"G�JH����� �
��~�ɺޢ��(POwt�h��b-'��Ʋ	��yb���O��z��v>/��(w]4H���ׯ�X�\��{ٍ	� H:�>z��r�c�#8��R�S�H��T��'&O)9`�	��Oj3�`���ZC l��!�%I��	L��FC��%'��E���X���EI
"��q!M�z�a� )ϹL��!���`�{�h��}��Ya֚-,Z�]ӖL���
J;c��dz�)\����&ڀ-d��I)]tHxH�'�d	�K�@� z�^)���8�ߦ�1�5	�,�ձ ��*�U xa���e�� rX:	V���� ,
��@�mb�vG������o�iNPn�l�Ĥ�����{�����Ӡ�sI##!�)�m�R[p�Z�a���>�H{�&ɮ�L��5"2r����U � ��HJ2=��汭�W�f���F-�g��-� 1X
(����b����;�q��ф���̈������?o�@v��bK�ԃ��9ع��=��D���:�,�\�!74� e*(�4Bj�lzP���wP]>N��-�S'Gn�6*�G�J��J��:�ٲ�%"5���E�Ѕ�Y��s(�ȋƐg��Y�P��P�Q���v"�D�~��G����[7�}�]��{�E�pَ�h�}~��.i����xݾ}���g��=����@�ަfӳ��F��
S�(lٛ�r��{�坏��F�X����:�ň���#O�܏ܘx;�ɳ�`Ի���w��7��������=\�>�5�9��F�G�!�1iJ�l�m������5t-�'ĩ�ͣ�v�4.�af�N^�p�"�9��1Y�O�vضFQ�yk0�7M�b�2w�G��p5B�����7&.�lS�h�<N�G���p��v�#�>Y��B^jba��tJ��f����`3���ԢZe�qg�r�i�;nCܕ��F�g��W��c����*Y��yQ��G NJ�`h��o/n��C�� ~�l·uؒc̪4��ީ�i�"O4����6I�C�2`�� ��x}Ӊ���_=9�8P�k���ם��6̄�@�`n$��r�_��'��`z���׼�"d����t>��,�u�wM� �-�4�z-�B5�ۘV��Pң�*�S�z���ߕ�DO(�%�~�O�J�"��4��Mk�-��L�i�@��3d����|����.�1��,����$XB�dl&���u�) ��Ts �<8��,�fF�����:ػ���EO@Gp��cQwuyIrW7���腎���f�y�*�S��#��F(�"~O���M��e�Z���:5��^3�:ބS�b;dd��Qn)�l-Q�͂�t;��j%��y����OS������{;�^ù�Z���9*�)�r����{��jDA�����Gy@�Sc�Jܚ�M��lğ"����W^]avLvJ~+�c��:��狲ˠ�qפR�l:��J��dXl�ì��΅'.������_9��q(<��ϟ����-��޽{�������U7�jlJ���\���]���/���9hɽ[ٿ�"����dOM���<�iwv����Ut�Km�X�(!�hj��l�=��Q�_�t� n��r��x~�B9t�ᗿ�ͤޙ���/f�8WݺZm`,u ���N)A�c��0
��x;���['S_�}mm�8�Ҹe��¶���	�Ϧ*�kG�t���:_,/."��j��m��4�e7_mOĪF�~��p�:/w� � ��~݈W$>z*lʩ�]N�m�ݦ�7��a�^�s�c�a@�6#/�k�و�Ν;����#Ӳ��3�:�������V��YoS��� ��v�Yor�\�[�k z��T�rj�8�7���<���^iww��T���n�Z^b�R���k��M�q��n��U�<x�O�3��k�J��xS��^9\.����oÚ*�A�>}�R��w��_�*��j�V�H��;��{������͛�f��	=����9B]߁t�\�r�'fHp���zբxu��ў,!��:D��|��]à�������"�Cѵ+f7�3��{��-��~�kE�9�CV6z��n��-�ȝ�j��(�N5��b��i�A�H����kA�G0Wa�u����쌈��!���ׯ��̝��V�<�`Ly�z�����/�6����&�h��](�0��!'.`�������P���)a�kflod@�hĐ����@1�ne޶�̇%1 ���d��%�X��|��zcSq��-����R�6�0* ���)o@?����T4���RY��AD�(TKW�$Y3@$:��,��g��F�UX��0�pț�^����z�
~��Jp"�@�)��
(S�:�~0n>�V�
[�Af6�Ut��x��Ғ�$��8b�s�yy��)�����1o�t�[{�;M�(u�(-9n}�屼���+�'�[R�{=�����8i�D�"����п�}� 2��놾��f�ӭ��
Q���_e�(a��g�Qȷ6E�R
��	�ǰ�!�z�����􌟟_�����;-
K��c3���aB����b�v�3�H��("���Ҕe�ɷ_��R�E�<"��@w�q��[�6i��|�����5��&l%�r�  ��f�f��X,��g�JB5y�"�&��r���TCdy�Z�C-RRZQ��5�~�x���5!��U[�k�QL�]��Bz���)Jb��QH[�6O:lc��_to����)Pd��(!�\L�[E���w�� �$���^j�>�8V̙�d`%w*!~t5#�;/�0yI{�f��1 �.���O�����r`'�9�b�!V������ro��1�1��g2�zr=�R�z�	)?q�B�<0�}�.7�H�&���$,X��`��JeF ��7�n?o��~�I�h��p�W�^]\�%^�B���s���.��Ŗ�,��d���uk���iU�1R�b
c$��Ř�5�fJ��"e0��}����K�aC�l��,f,�]<�8��rT]��b�l��TM̌B9��F�t-��`s��ej"�X��#΍�⩇��%>;�<��2K�e���G#�y�2kL�m�Ak3g�F��9� uuc�s���0�<�|��cj���)���u�KV 
��H:�ۛ������&��1B�/����j�`<��%�Sx��h����Q�J�e�R� 9,*����v��H��N��dNr���O�B쐚x��E5�"��i<>�k�lq�}+��U-Kt��	�E@ +MU)��|E�u��MN<I*�=��R2>�ܔ{�-�	��fJ=�F��"���H�L��...9�Ё��B���Ƅ0�xh�
�z��Ι�d�/� ��4-���2.������Ve٫Ҏ\T����sv�46[^.����������R"&~�݉�yH��^L�+4�
4(r��xz�f�ya�� ��.�`	�h,?��זi�,�@l͐�� �A�����b�J����-L՞,�r��0ޙl��G0�0�rH;5��>_lt��'��~����_�A��`�6,���O\!-��LhIv�j����\�Ĕ�H��bo+O|��{�2����h���0����f0LAfM�9HC�Tx��F��-q;~��_���?Diw�h��D+B�QF������EKj����9�C��S`�����w��e����Տ>��R|k�o:�pbW�N��L��"��x�S	��b.��I 8���9��6P}]0��$�r����l/��RL,˿�1'G�lBe�")!|L���(���;�o��Ն���_9�.�"��S ���Ѹ+��Ш'��^��?e.'�Y	��h.P�-[���lL1�����/�ܹ3�ٓHX%S�k�����.wrr�Tr͵�JM�J��0S��D$�m��>D�A���GQ�68|�L���^�~��(oc������D�(��^5AR1'4��^���|��Tl&X�x�6͂���2�~T�I9^m ��G��;����틔fZ�]��ߏw�5�������r����f��\�~}��X�<�G��±�����i7J�&�.����D柽�v6y�������z�K�qp9�~��W��h�,h3���L�}�v��'ͪ����!3>�Ȭ6��t�^����R�I�Wd��������5�~��V�A��=������a�$󊊍UPe��T�o`���;=}M�	������	��ȉ����ӧO�7ol��I���e���K�}v&_�+|r�򓇱}w���,�;#���HJ�F������ա*���2��e"T��-��u˟nݺ%%�xy���΢o���\V�M��|����4����<�O�J��y�@�����j�բa�^;���ے�)w�!��߸T�/Y�cС���" ��F,��~�����. ����3U<8�rUqܧ�DY�����zsp��w�Xx@�cǸV��* $/ɦ�PV��+`T7���d�BΡ�	���Gd���6�d��&�C��` �U��`�Pn����3"#��y�AvA���4.Q���zh���^9�*�<�#��2VLJ��q%H�#NV�B���=�슮��&�ܩ'5KF���������J������N�P.3���3�����d�DS8�'S\	���#V�$��D�1.Gt��k	>�!o��,��[���ђv�(��	~'�6u���ݣ��)���w_n���qYJ�C��f�'�y�!��.C�RH+C�r�6�Tf���쯉�c�3Q�h��2]N��uo�Ha�,P��bN�;�D�&q�E(�:�>�� ��\s��F-��1T2�X7"��)� �#��̐��L�-����
e�?+lT��h���L�@2�İBn�ŋ�GG����_�����w���֦����Fw�Pn�'e����Åu2AEyW���z����B�c��a��7��=!80Fg����C�u����h�SW�q��1q�� �S1�qPC�t�L����2#���v	��<T�F1���i�ԘJ��-�'*d�Q^�R�Y_�%{T&8�W��u;
�_�T�0�i*'�2S<S٠H&��������[��+��n{��B`n����D�PB�F,��Je~4ʩ.Sb���ǖp��HByX<����I�{��l@��(o���;�$��vo�H�BEE�;��Pք2���ϛ�mHU��.N��mS��_��ŇY�7�y�콑�/�ǳ0�?pY�M�w}��"�:]m"R��`tc�!_�i��D,����;7���
����+��2��T�˴��:�aMHS�آ��s�uv�tB���<�ٓ�%�yh�.���!=�?)]2Q�r���϶��:0E�	I�P��=�P�S����t0Uς}i.���Pg>l����Je`\���8t�3����K Q�|��pT��ͷ������[�U��P�VB0��Y�)���XZ���)����~h{U�A��ix��F��*q\���}R�RYe`�JM���iO&� ^!�%�́fjZL��B��\�RȒ�Q^B3����]��˹�a ��ݽF��(�Ѱ��5"�c��ȋ2s���)o���HC�T%5�gD6��$+�
b�z���u}��/�;@��H�Q�ͥ\-�5��j�0/��j����F-kD��*�.�u���'_��!��F�F�XJ;s���,Ɉҧ�<y���?&~^�&�;�q�ǌq+���r�A�$�ב�<��m'X�W�L1j�hv��L�f+�+�]Q���a�c�=x�����4 W�XU,���5 .
�sï��=J����U�[
�w���	�62�]��׮��?�v��r��'O���>]~����|_�-���<MS֡U�A�G"����J1�����]����PDhgir�b��=��n�@<���Z+��s�=�ˮ.����T޽� O�2�<w{{rL�#����L����ȟf�b)���_�z}�)k��!��k�+27��C$�=��5x�ƍ�ã/���ޒg������3�yU-�*�>�o[�_Į��MR	��B��:1Ч�q���S7U}S>B��M|�Btn^M'�.���#)��<_0ثqH\
������0ʤ{X2���U������S�+Jڵ�V��kGC�7����<��Y�M�I��:9x}��XR1�o��]�D���(��k��{�OB�۷o�J�_,./����*7�R�'�m�^�)��b������bn�p�
9\���ׯܹs�id������y
�F$�"ƞTHك=JI?�̶�ubG�Js�#�W���HdkZ���w$^�����Ϟ<yB�Q�����$w9F[W��d�5΄�����}�R��P��FT�e��/_�+:88���[�u�f�p�#9����<,�K.BBüLݗ���1$p�;:�S�m��;��7� �$S��XWX�ZnO�&7,'W۫�z�XӚ(i|�"�Rq��oBd6o� �j����7o�$#W�*���DB��Y�G��V��z��<�w��}y����t@�0��-��<�z	{tJ��=9�� u�&�~��M����y��K?r�p���h?����J��g�B��o��B+E�,WM�I�Z�ׄAB&q;�gX/.����Ϋ�s9g�^dU
�@$|\�4�\ܝ��2�l ����O�%7��n�D>0�T6slC��u�?7���w��+x��k�nv��L�ր��:}�&f�l���j�Ը
s�����#�S�H��O�z¢H�����Y��0:U�X�c�鼖��y"O�c&/G�`bO���ѡ����6�Ǟ��Dx�n�+/���N�I��I{��a����z�w8�!�̡������Yo���!}%+ӧ��t�
�d� nM5�m*"Oߓ�@lZ���D�p5��i�f��Bi�fD�?���Q���	���2���:���w9��u�[����$�p8tc��)$x�,��E����M�d
b\Ӭ���씫WZ�u�.��xz�i�{�n!��JǊ��%a�ؑ��H����8̔�OUX�a����g��0�#d�^�룿��h��f6*Ptw��!���5!n��<\%���3�dQt>���^R���wB��6�
F����G��3޿��h0�8D{�6�M�0q28w
mG[��i�3�����o~���b�Yv�ɝ���P�����#�$��01��0�o������z��_�m��B@�����Y��|��q�;������LS���M��A�;�L2��������L�1"����!��V�8<<��1H���A�+x��w��'��z���z=��B�8�ֹ���t����Y+�J�������K�T��O��+�`1����/�H0���î��)����	���<z^�������6��/����IO>����>��iVxfK�l�s�Mi�oRc�Az}{R�;(�i��!�p��N�7�~�IӺX��f�������e��v�M2\�����}Š��o$Ev"�N5�\��|Y�l�~д���RA7MgTlП�I�Q	l۹%va!��f%n��|��O����ܳ�)άr�v������vu���6�B�{�nD�m�T���QF��@0B$ľi�='�������Q#��� �[&h��M�e�x)�o�e������J��
>m�E��ۯ{fc@�Ɔ���]%E;|T��;5�ʈ��VZ�	ڢ���j�&u	�60'H��:���X.��\Xi?�X��ZeX5�{�,x����{B�Z���H�*v��iM��s�8�	�S��鬗��:؋0Z����йa4���0���pOa�r��qe
�ȍ/��dnX��X��j�kG~�D�v���SгD�a���p�(^SnOl�Q�Z��m�r��-J�w�
�t�4�g:x��;V��`X������T�&UTi$��n0Ģ�P)��ɷ�Ԯpun�)$h���/I���%Z7��ܑ�B2$N�y�X&�Ԁ!�өZ�}��p�j�.B,E3x�ʝ�8�����/;'0��j/	�[d7𴒧˥$0�́�.l�_�g� 7<rD�
�Ւۻ~�:�B�ѣD�A,�/����u�^�9Ǎ)O�z��#.<����a���Q��S�Gn;��:턪�pvp��H�N�6�c�vZ�@�.,�#�څӠ�7nܠ��_}@'WU~�Ͽ��V�LB�H�j\��mm��Ge�D]�۷�М�2J���_����,;a�rN�0&�睫��֐��fSS'�u>�a}��@*�W�_�6
ȧ��
A5���#F�B(�w|RW�Χ�g�}��ݛ���ftz�x�zKE�f�S��o�k�8�������_+k��:X�[\M5���I�Ĵ�E��I�&�"�%Kq����.$j=<8R	l�|4�W` ��ƨ��� p��zɗ���p􂡳ӌ��U>T�=�z�*8�S������1`XA�W  ��IDAT{/|�a���@vGB�k�k�P�]�6;��Qb.�԰6ա�MÙ˼��klD���S�ԫW�`eT�d���	�<t�|���y����P���@v�gVAf;S��8��r7��f���\g��ܡw70��b8]^��^]�:P��yg�-��	������<��}����&S�����X�bnS������ν���,�K� ^�:���y
�+yR�Y�C<����F�4Q�A>���S��ɵc'_#�I��P� �j���[׹e\d&���țu��Tw�-��H��\Ьt�ȿ4��Q�Nx�0
�"�;2����%(f1iwwB6�t���E��� ��"��є��l�2�mso˄YN	5�MKmRg��$��P'Cp��zlԲ��)g��V�aoW�}��K�YK�0,~�&|�OtK�&�5�a�9���omT4��a�2����M\NEt��!OT�+8�� ��5�Ѳ�%Zm֥��n �d�+P�5�/�;���m��-BZ�`�A���5 :Z�ƣ��)�Ш�nbQ�牦�.W��6��w�ugŹ�yI�+a�l����"��rS����="�T�����.1!K��Ni}�i,u�!W��C�Ws$�oL��j�z�6������pCa�-�S�J�~��Vt7�) �Wn������(���F7�'72����������8�!�S�c3����d�{\���J�Ҭ�S T	<�4P�i�7���� (�BsF�?�������Ԉ�YX��;nz�O�w�.��}U�����ɧ�(�\g�n���׈���Ġ��@��8�g�(��$����a���s+�4�O�Ŭ��(c�	Yӧ�Te=�L���ӊ�V����#���(�|� �y<���C�kyF�x�t��5/�X�}����k!�FgO�m)��+z��EUʮ�2J���M�vf,KP]{�e0T�?/"�1\��qH9��R��̸�[���7p��-.JBcm@ׄW�=�M6�)ܸ�
6�&�[�_>b�(lrs66[�T�s.��U޿X�<51􉢍M�,K��&���{�.�4�b���9޸N�����y�,�w!������x��ʷ�"�.���~WZ�N��#���(b��*S�b��]v������ET�>��ͳN+�+���~�2}m�*g�jX�ӔB�°F.nө�9�u͍�#sw��=U����ۂ���r��PZ�S����ގ��#��y`pAU� �q#aٔM��o?l˝�4X �0��{���/��Ͱ֥�t&aK���Z�<_�<a���!�� FQE���5qI«�A��2�7�|�,!0E��Z�^�idm���(3+A
Ъ�b�X��Du����ZW��J�!���b���r�b۷ؙ��F��:���^�;��X��"n@+�a�ӖI om.����*#f�����L���HH0�^A��Uڻh;%�p�`�N�E��t�*5Hd��Yk8'?lVkyX�{����]EL�DnȻ���U�����A�y�.�h��R;���u���oh���kE"�DkO��7Ж�jtM��x�v��[��x�`C�#�k��M�:�e��҇�CU�H��k#��9���ؤ�+J�u>#C�/��ZDk1�D�[��j�z#r%;m ����N98})�� ��n-��d�F���`�4x"YE�1�.�@ *ɠ�+����v�}.�^^�،�t Ҕ �(r���_�͋�yQ�l(��r1|��7J�S*�gU�]9��&�Z�vQ�9�NXq����&GU$���yW+�bP��e>���s�2���f3�dm����˻7O���0 �9T2�I؟�/�jh��O�'ʄM_��5+'�i�g�Cw���v�>[��/���+��4��Бc��V�r�0���Bg"�rvvFq���Ӹ����%}��o��H�z��H@�(2�`h��w�3v��Xv-+�����M��'�y���{��w�w�܉�h�E#3ڬ1�c���z07Yx33�Np|3�����(�Ê�*�R�RG�wMW���Tu*k2��Yv@�M��|�|^�\�:^]�|���EΪ\s�X^6���p��r�	!�eȇ�f o�F_,��2�0����&���4�<�b���k׮qno�q�,�Zd7���=��X���-�ɧ��2?X��8�fӭ��O�Y��ޣa*U��!�c�1 $i*_�<�%�x~~���N�n��O�s���T��*��	����xZ	���������\����1���d@i71�ʊ��$�`���Fg��w���[�ݸq�����@j3o.�����<y�M�=X��l�D��nݢbϐhc�|�SyA"YE`�iYf-�8�E���l��X�ǥ�9y��X�9�jq)~�ά��x���g�E��i���,..���������![I�rT�׀�����3����*٩w�\k챏u>���&�%Yw�<M'{.�ׯ]9>�_˙Y_�Uy��������+03t# y�Թ�%41w�c������Ѩ 6� ꃁV�A~�W�E&3���?������1�/����{Q:�U/�<cd�B/������G�.fR�k{��,��ѳ�I�!6���>e�b���"�n��� ��QV�(r��/��%�ę-���d��6�����0�2_�e"J#fq��Y&��A�QWS��n���S
B�>�
�y
��A���~��X�U.�Z�:y��f�z|��U���}�H	(V?�&c�@����ʥ(�vF}��b$d-���猯*��Eu�Ռ�:y�|�Z��Q�D�TY,EE�Y���ZkE%��BY��i�k5�'z��~Yo�^b�D�D*��<�J�o�`E��h��Y,�3�ƽp4�& ��PQ`w������=d�I���K�Ms��ذ"�RF]q�q:x���b���j�l"L����2)���=��n�FLA�#*z����a-��PK)\�?�'m��,ײ���?������+W��wR�Skw���`��m��)pq0���z��he������g�}F>�܆!�6��E��h(t��gО"Pw�|^�ߋ�$'eK��S��*��� �C��(�:��hn3d�P�������	~V�P^��@Z�O�z��A�����?�H����[Ϫ���O�
E��읏�D�M�� ���K��F�K SJ��HUe�k۬C۩o��؋K�~t~��	���{w���������>���~T��-F(l��.D0���`M�]+J^c��VcC��.��˭k;"��ȶ�x���]s(C퇔̈́`�YA�@R�tѿ���C�Ƌ	�����b��$�"�*D_y��K0D�w�p���}rcd�զ�0�9�C�������D &+9j�U�O�֧��l�����6��zcB��i���� Ɍ���̼�Ю����a�x��X ��J��r��L�&���>����_���'�A�[-Ô=lb����/�X]\h_��Q#ڦ���.�n�Lk^���s@rIu+�zZO�z;�s���zA�D^��S���Q�M�I4�m�+��Ь�%�w���0u��:ԅ��G
?ȘU�~��	T�F�SJCҢ\���+�p����N�:fsX�*y�j��)���Ӳ(r�	�Mg�m,���!#&���x�3ve)��,r�	��e5R�XsQd)�b���cX1TD<�zHhް��E���� BE������Fm����5kƱA-=�\�����ƥ
�*���хNo�G�*�DI��>�iҔ��gv�TMa���/x�����@)�S�/����+�L"p���X~\�pa�1R�Q#M����Jwx #�G,��nI�*�OA�\�T"Z�\���uy��*��N��ǜjV`s[�P+KI�-��kI�8��R��4�`1(�|zz
�<�T�KM��¢h����F����n��q�O��CFZ�>��
���R�}|b/ׇ�	� OJV{҈j��-��X�"�'Z&����+ o��OvR�D���..N_�����~�!D�������իW�9�m�T���A8����P�FuG)'Ϙ����'�=wIfg�:؋Ǎ�בO.H������Ue�I�=�����/^�2޻w����_}��Ϣ3���d�"UM[ÑJE*��O>��������F	�����H6�U�X13n��O#�D�,�Ҽ��PavM�Pn�E �+��o��Vl�l�IO��xM�%���G?�#9�>�+�o����B{�������&;d�&��{B�!p��06-Te.�h��C���
��V(�m�V�I��f��K�N�\��Q���(Ȑӣ������.�=�JJ��\�WNcNڭ���J�Ç���%�����S���@1O�9�C�4x�؍�`�j��z��J�^�����de� O#���
��2K)2%����YL��sۀҞ�>��y��i���ї��g�T��ד�h
II�`W��U�ϒ��щͿ��2f�o^�ڛ���Rc��Hu�~�
�tά���YG�ؕ�����F�SV�����4ra�1Slf� <S@6�C��l��M?��@��~r�ۭ��g��Z�j0c^�:�r��<��[z٣�#�7�j�X�+,K���7������Mwf�BD7�CGT2�ђ�<�9&ט�7��h��y�9��ʹ` ǇU4Sq�ܸ�Q׉�3|���t��.{Ӯ�H�/���������XCl+�|ܒz��Tl��l������':�����=�3�yBc��P WYn�����iQzNT!~�d�b"{���`gL�bO�����e[� ױ��*k~��2��heq�Yh��Cc�x~	��V�+�sZ���A#"�����8ݿ���y&��q&��C���rAA�씄��*��==��%�Jg��/��Yn?�����L.�6l��
W1!�����ĩ�|� �|ь|��=
O���`�4�U<DE7�)�P��#�4qe��(��XƨvJ9�ZKc/���\��m���t۴��W�T��q/�nA���1�4r^#�qt�+:P��>��a��ի�:a�%��Lʳ�$D2��6�X���b�z9��ݻw<x���Դ�ӧ��`���z}�0�~�E��Sׯ_?>QT��)~�K�h9�*�t@�MIQ���,*T.(&�i2�,�/?Ƚɿ��� ���������]5 ����h�y���6î̪ Y������.U!�EYn�����-��,yL�!U/}JF�����=�,����qZ��f��,w ���©��.��UԂlt��/�@X�ꝼu���e�N�yW�c�T�a��p��\�S����򫯾�G����={6ٙ��=��I��X꽠��Ղ��"ʘ��݋F7��x�&�-z�Z��胱���r+廨�)3����|�.�`�7w�^M�����@���wbs�訸J�
d��m����h�y^�-6�45�t�w���;_Lk��.�Z药���[��>v|�;A��f��׃,��.e�e-��H����c̞���e���"R1]/�x�駟�ı�v����Wd��Lx�X̠��t	Ъ�X����_�^��T/z��(@%����N�oM���������1���>_*��Yo�B����rD�35�t�z@����H>"���#�@���"B�5��*s�ԕ'�S=m�i��N����45�5d��Y��Mh�*lV�(���>aJ���c���吢�H筈���T��Z�Y�0*T[�˘���T��P�6J'{9��� C>��Qn�/c�g�S#���v�fj8�J��,7:��
}�)syo{m��^p��fe:��Q��jq�꼈��8�:�w�4�u�)BT�7sLXV�G�@E����*�6C���l(�$�`�PM_\I����I��
Bg%X�m���Xʯ�f��콂|(?�b!��Љ����=HP=����S��e��p: �ɐ��Y�Ȍ𒺌���UϦ�q��8��N����G�jNdRT��+�����!�lZ��MU7�%Xѵ]'ˋ�T�
ȃҀ�D �$�t��4�0G�U~s~��x�q���g��`e[��l�]py���:� O�e�����YF�,lҭk��s0�!�/u(�dφ�Gvɑ�=|��<���oQ���Z�<lk�f l��b)[&����i���<��e=۴�/�/�z�Z-~��ݺq��ū��z2��>Y��hyd�SF�U�|�[�]/w��C��[GTk9Q'�"$�(���	�`��nR���J=�r�L��35���6���*,�j�iY��aYu���� 4^|��{�<{���#�iq�u���Ҝ�� xZ���D�ef��u�G�F���g�g��j�e��5լ�Ly����%�d*�+��q:���_t�œ�wvv�3���D�/U��E&���>�?��P���γx~�TDQ2C��\e��_���?�p��a�!%Z��N��L�c}:�E�.�0r���F��}�1�!Z��CJ�|��7��,0���ƕ�63��Yk��Z�E��e��V&Q��qW�P�KAk�y�ڞnS�C�~���?�T����˗��p�G�٩�����O�Dޏ��voOl�lQӬ� ;�s��%P(�H#&ep0�'%d�R*��z��\��HMM";+�!�4k�+��X�/.N��H_.�ߙ�Ke�@������*R�k	�傢��G��rMn�I=�H�@�X$H��(8R7O(F�)����R?��q�L�P���
���	��:�.x	B":��*y��A�s�z��d���f�
�*f�p��/�{�]׫�� x�Qr{1�`�P�Å��T�
�(�����lVy����_��  )�E	����|������W������͓�o߅�Z���k�7ϋ!1�?�=2��+��)�P�[g��AF��9�S1D������ׯ�8��8�爱��z����Jk��B��#���gً*�w����~��!��P�E+�)E�z4g�NpA/��Dήَj�1��%ղ�|�#r�h��^�t�z�47�?iVk2�*Yt�<�s�E�}V��`	0��"�4�p.��[TV�j�À��兲Q+NPS���%��ͭ�t�_G�3��ӱB<����)x�����M3�-�1���N������s �r��5~U�����ݒ��w[�&��q>Bh2E�H7*u^P����'����>S��L	�Iw�u���8�����좪ǔ��,�sX�	�R���g���3��0Ϙ#Ko����+����|w���yBV#)3ۋr�Mu�3��t�t�ҌȵejE�*!���T�~��X����Fb2���[6�#�6ԫN��Jo����^��|Ga��X5Q���uL���A�8nѐ�W'׎����c	{:��[������q&�|����ܹs���n���kQ7��R�i?���/^�ϰ��S~#%o��%{�\ML�ӧO5������kMܾ}��?��������ɓ'����k��_|��g��ɸ��`P�8qt��r9�\�N_�f	��*�h�a��h�~Cm�s�eE*d&Y���G��H�I�,&h>�9r�,���&?�䓳ˋ�f-�	����B5�!c�X-��V�@���g�\��ENϝ�.KJ��s����L�)1'ܧRud�F�m+͛��v=�$��F>%?{1��������}�{���&[&b��&���b��eH����$�X #� ��\ϼ3���qR�J���ޫ�(x��J����l�y����{�{:A�
�~;`Lzr�	]��ׯi�)���D0��]��YK�O��2l�� Xת�3��Q�f�W�,�ѯ&�Ġ���ԍ�O���+�=1���<�$x���L�Ft�R���,˖�Pw�D�sB[��s�A�m��}���
`�G��O��1&�@E���)�!���*�f�*����+�v��oX�RK�#��$s��MP�̘�;`�����f� �Q����jl�&T/z���@$GʿG��h9҄ �Paf��y���Ge�߾��ܿ����a�ڸ�7Yjrt<ݙ�i� T�����̻ݽ�;���g��������_���P��Fc=��E�O�� $W,*2#/䀟��*��/�g�Y~���bMW\�f4�&'��b�5k$�P�w;�7�$$l�F���H��L�3�NJ�hyn:՜���XL�����	��b�UZ�$�w�|5�<v����}-��x*�Ĕ$*�� =B�Qd�%���#�NN���+-&�`�Y�W�0���Y�`�Տ �c����jS4���t�y�X(����v�0����\��J�*CunزЋrE�oTi�U�2¨l�7�iN�M$eJcd';�e.No p��)�JԢ��JYl��˫1���yמ���|�a�sC\+N'�����|4��[������#i�OE�%�2��u��Ã=.���jD�*������,M�Sbt� ��PX�S�D�	kj@ؠ��I�@�C���3�˒��r�i	@����s�sҟw./�\�l��Y��x3wjmg�q�Ґ�v�>CK�}w�Ac�fU�F��S#�bA�7��y5Ld0�~�K\�釱%�O)6XIK V[N��������ŹfW����k��AXf�n�I�`%}=��,�gA��#��9p�}*��y2������%��L�7�]PJy��n�`�i��
��;�:Q�H��ȉ�ۈ2��bH���������F�^��.�ŉw"b������}�91Ş��C2G��6�V\V�N�j�9�EmC���������O?x���n\�B=~G��Z�ы��Eά\}����0"Q.
�[���ߓ��C�����-�g�����^C�����.>�%xx�mt}V���L�?.�4����,gP{�ONN$l �IMF��Y#O}0N���ߪ������ʪp�ZT\�iHW�:�`f�5$������kp��$���䶣%^%��-y�X
�0�J0��1?�4�L~���G(��D颟J*.F&����>��02\��[�-���4�y^QE4"r| ��R�����E�T]҂q�7nr]�6�/�#��M�.�%[&`]��VR�ш�mH��E�gϞ1J�c��B&��P3{��6�xB�B��
�y�é������5o@ê�uxVv	��a�sd{����5���Sw��8���=b�`6l�B�B���1F9)R�k��;�v0�wɿ>wO�!1��,�<-�I1ڲ��u܅ɴr�Dn-�Q��|��f��,�=�5�p�5m��\��V�������W���czӀ��/�%ިpp ��R@l�<u�F���.>��<�R�g1&F��O���%f�(�|4��c>�ؒ��K�����+ׄX�w��g�a4 N�	��s���G�ǁ}�kmњ3ݎD�0f������jT��X�2"��:߅�/F�nSh���	�R�2k*�ST��>���T����p�fU�A߇in����2�^�VJ��`�Kcx��KJ���&��چ�?�BGU)V���F�u���k��gu$Xݔ{*�~�ƍ+W��}��� �������V��2���_��S�~��[o}�������E5,���-.��9�"�?�g��\�~]"Vn�X	X'��lV���u�[��w�}�/��/��=~�8�YnR���?���~��7/�x�ɭF�%*����2���Ռ����Zğ�I�\;=����KY�{����<}�����`_\,��Կ�U����o�����N-m|��J-��h�ln3�e��Jf�*�ܫ2��ju�z�v���N$�W^��z:!d؏�to�bҰV�Ow�Ν>�@�����慵��ˢ]Vr��1�N�2#��s��&L��We�¢�Q�u/4O�޾Dp쮐���ϗq�;��Y����Pڈ^�����'1rL��H�ȡ�㯾���Ç����Q�.q��F�H;cF���A��S`)�P���L]Ol�c?J��FGGg����=v�]�҉���oQkN:�.[�RR��A�%^����a4�>�l�	^h�\_�&n��t�����kx�^��s]PA�)m%n��*�������4��r�-A|z{="x�e��(���X�&`� �R���lu���2<��T ��m��/(����^������~&'���[z��}8utȁ����)��bEۡq:N�ήz�g�0��B�L]>1��=�\"��rA̪!�<tp6]+A���X�3�~��7�ļ\\6i��@g@�m�r ��d��P;圦�4vw�f�4T�p����7��_�T��u8��|d���R�81h4:/���ht�.��2W��$d�Y�CC�\�K�x܈�0�wP�#*���IV��-γ�����g�rrvq�b� �R��f0F����� L��_\T�<H�m¹��>�u}�T);{3�q���c���a���Q�s�<�R&��
k|��$�?ף�@������ڟZ^���<�j�z�+36{�/���,;�M��Y��_��E��Rƚ��H@EC�J`���v���|��;�T.���V�uu�Y��έ�-���2]�ì��U%O�$�b��zFIUs�׊�q�Y���}�����7�f�Uw��L�ud��e��yķӧLl唷�Dk^)�%q���+���"	��f��c8Ǎۤ�7˺R�@��~h�vx����;����r($|8=U �<����b"޲�5�$Z#�����;��s����w�Zm{B)u����#��*�XO�O��P�ż�L'})ڭ�_��x�uYO�JK	xQ]Of�w�۱u�/�$	x�v%�u�H��7���t���=Z�P�o�+Ts�����_�AJ-+:}�>Z�^k]�j�R?���\��ť�g��/Ξ55)�+شD�̞�_�'�Th��G�� �� �MZ��;��6��P9��\Ν�Ȓ�Y'���D�,��x-�YVuc�:��zKS���p�vë�gg���_���O*o�p./u�70�e�[�I�U�'��o[Z���0w���5C5c��ɓ��ј���	U�������bD�8SF��7��i�5�	U���_]��2`�S%�8����㕅q�#��J��W����l�J�R'�{�i�� �a��������>�h�i�����_��6]JR�ru����)V���eY`�`Y��]�k/�Y�N��X�������� ���د��*�����R�"��V���]�}6<Η7<���3zr�؉X���)�
&=�͸2��d������!r���\�P<!z�����ә����``C����0��������/_�d�F���n��_cѺ��E�2�~���M˘_�kG����.�~�ޭ��兆�%��^a(��u�����L��*ʝ��`v�=jf�
Z';�ݓ��UڦW�\z�@91��L2,g;a�v|��ѣ��y?h�`U��G�����/~��\EQ E�6�*��'�;m}j%��D3�Q�H!OЉ�[gI%zY^-pu1�V5 �z�v���K�M�x~z�Zv_�H~�.V�����O��j�'+�V��jCLl,��H|ɛ:���^q�{��\%|���`%%nVbrM�}�F��F��Tz����!yW{�CL���:c`���6�Z!)X� Ƥ�`4��=h��j[~A��������oD�<&�ª	¦^�R$�t��������8�=�
m��b�j:]uŀB��2S�����ؔ���[���5j�J���˨C��n��Q�NN\)Yd9.ST�U�e��j����Y_R�i]yЪ��(Z̸n����Q��"+�c/���#��(P�}1/,K�&RS*�<A�E�UD�V��8��oݹq�ڵ㫊�����^Dd��O����ΫW���w� �����;wo�|u?3Ч��;L'3
6�b/^��u:8��QZh.~A�||E@�h棣#ڠɴ���������vr]�����{���/��'�|���: '{��x�}����9��0:��ry���$���}�r�d1�۷o������tž��+���� ��	�\-��U�(�:��n#Z��ND�� ��+G�ns yfK�w�Ɋ����¤;�јy��];���O����v�y��3�v3L������Ԭ�����L �����������}��ݻ�$P�4��Z6�/�Iy|9�=:��.��'��p&�^N�s��1[�\Q/���p��%�ͶY>��ͪ�Pn)���!rQs��̒C�k����.e�D~�a�>|(�$�կ~�.m�����{�G��̬��Ꮧ�4��.�����\
��ݫqՔ����j��jMe>/5����AVOk䅹2���7�����CBi��Z���S�Ԙ�
��k�A!l�~7"VGw�O"Q����K��j�c���)�+7:<���u��ѹ��9��>;��'E���:�e��=��K[X*��	�eu���������6/��R�z����gM���;>:�r|�+|�⢰�.��[.vf{z /�E�NrQ���6�U�3� ��i�w��_�g�w	��y�p�4��zl���ڗ���b.����+\y�L'�cf#2�'wx����Ǐ���,Ö�.A^HV^*}DJv�1d��ݓh�Dmv%��C;�f�'�0#�JH�J�h��W6�g�'�#��E/s���L���F�`9����Ί���dׯ__���#�����h�+�'�Ob�$Z�PS��f�6 �$�Kl��1f�;D �SZ!�X?f���|p`\rp)X���ʍ2Ƴ�����`N��/��E��Q�����QWʷ�]�-Z<B^x� U~/����3y�h�`M�d֓����$������x�9�!��V�k�T��q��q`JVP���ԑ�*F���5U�>��O�&�M|6��,MqBd���Ɗ%Q<MZ�`�=ÏN�@M�֟�_#�4���=�)��f
s�0%���UbA�0`�h~;եB����%fG6E ]��F��0�-��$� <iK����7��Ɉʊ��>��ca��b"gQ�D7z��{x{u���N]����>�{���ߗǿv���i�O���Fq;am;-�[��M�^�[���������MZ6��\��`t��4l��xN�]cU�36��w�?}�Lڝ��0�g�n�p�J�05喹:r/���fg��ߜk��~,�f����͊�gF����re9���@���e�������SG�ʭu�R���U>�����'?�!�~�ĭ��.���q$��]��M|뿻w�/�/��C����lگ0|k�C��-k�s�����+�d<���*��`�� �q����1����">@q���Q�W���LB����ܩT�C?�Md�$V_L�N3��Q
h4���>)9��bӢ�����Q���b�^&�k�߹w�\����=�*G2`h:R@���'r�vC��vZ&˨��%�e��\��
��_ik��� �����������VQ��I�'���-+��4vC�o$�!]�K)Ӡ�1�3��\�<K��Df���rO�8�v�.{��3�"eQIGaS��+j�ir��{{'w������d�Z�t<��$b�Q(*}��Ss~��Ѩ"0uI�.x���[o�5ߝ�'������U+PN�]�Foᷟ����"B�,����(��W�W��~����e��\T6�]Q\�N����W=g_bT�U�5�9lG����"U�Jn�2�لk��/.��ʹ�W䓥c��0l���v� ������ϔ�ڵw4��n��%RQ\�
�	��<>�Hw�D{��1�'��;�)��zFAE�RM�1��F"&���ӢM+���"y�|^j9������u��@I��b�5��h�b��D�Ti�\3�P��o2<k�%�NX�o��ֲ����;C�kH���d���FH#y���i��GMo�˟��K��|q�:������S/w+��HL�&M�C�6}HkEkEƅ!ۖ�����X��F�Dȃcܼ�3�fj01D1�8�(�����{�ꑎA�?��p�H�K��2緋^��|�c��.
�Sc%W`�o�nhh�K=c�_��N���"�%���{�Z��G_T"�[�n]��,SI�q���w�}W��g?��?���%z�S�	9@W�R���h��^�Z�x6y��0�H��`���!^o��69X�������_|�Tয়~:��<|�P�T���g�yʬ���(ל�L]-%�m@�Fx�y�z>\�iU3K�(���%mbi����7o~��7�^��`3��iT:��@��<Q>r��?����ݻw�yeI���"���&����s��e��w�Y�Ww_�KekxϮ�[cI���e!�^]Mx��h���N#9 e�<�ĩ�=���m^��r��Ȟ�\smHMR����?���3��%�Ḧ	��E�x�\����hl�$���SW�3a
��!���έp��b�{��ǐ��I���䧨W�7���~�"\��7�שr���4mӁ!y�ohTׯԸh]�����ʌ�����%H8�>�l�$�yocb�+���#љ�����	+�dd�/��-J�o@iF���]�FIە��U6:�&t�6�Yk��ٳ���ۿ�r8��3$�����o<::�@8+��;�d�r�*�m�:6�|�f�B�N�t��r��r�x�M�W%�m1S{`0X�(+"����bQ���Y���h���F.����
rju�NڜT�2����<ܺy�S3н�pɓ*~/g#�~��Q�e�t�b�ĝ�@�����Jm{t0u����Z[w,��M�r,�;V���]�D�j��A�h5]9�^.�ے����W���l_G}ɞIȡ�|�wQ����׬�JcQz�\��������[���((Y�,fs�i��"U�|�Z���,�P�"+��� f;{U�(�^�֛��}�4f��)SsSJ�3�M@"��0��VT�&6��\��/Nwܾ��26�b�ͲG�o�\佞���&��G�IZ.��.ɓ�zvz��UE��_dF4��n_����X��Ζe��J���-��Q�fh6� �%զC�#r����N���*�ޡ�,�,o�C6�5�J�j���3��v>=��Ӫ��|��by����0l��Wr�bdp�NG� ?X�Z�����D��DdM�fJ�W�c̬L�T�xDY�zCQ~����z�7��Ix�|����?�D(;���G�����z9�D�w�٭���ܮ{zt�2kH�9�u��p�X�Aȁ;�||2�":1$Kk`l#�F� [��K/�0lD���,jhö�A�Y�'���]4��x^\�=���G��D?.V��r�EiNP�M���D�`+oy�����m���B�����w�t(�~Dl(�;�����������W�\�$+Kw��}وg/4���էQV�Fʀ�n���L|��`b��|<��BY��n��ֹ|璉�"�e*�D�;��O��^�_�0�)e�5O��bD���N��o<>�e�Hl�������>��͓~��LV�4R��8:�wS��-���-��Rt�x�?���9��.���y�2��}�ԭ��I[I��US�z:�&�$˥]�6�X���+�H��~��ԭ��4pvv���3��#P��Z���v��{^-7�Ŕ����jL(`�Y�{�F�[�]�n�j�$����z�����&��U���2��ۧ|�2�d�F�_[�������{7�]��́�><A�З<h��фɥ^����|FPO0J�~�:�{0�:jn���������&�>xr�3wƂO�`�����"4^bm������A�C9A�!y~<Z�q�@���[��'i�(�N³hl�����\��ʛ@�U��iȽ���~��w[pA�S���&ҋ���]y�n-V|�4��E�ʧV�:�1� �R���Kt
w��Ҽ����Ώ~�ǈ�UƮ_ە�ڛ� ���(q1�ӟ>y�����?��?�6���'?�cَզ��Zwb���}����o}��WO�y��8o�4�q��p6�>K�F�U��H�QAO�dy�M^����#�C$�����o�Π.P��O�ȯOщ&nd�\h��"����q�ZыV)�N�,��ҌsH
r���
���;��;���෿��'���y�ΐ��iYj��R��ys1��8�����S]dH�R~��1���Cg����iY.��'X�q�;�E4�څ��ű(���x1B������_�l�X��/�ܝ�������?���X�_1�Q�.4�g����u�%�T�;!1����܏��@�hUG�#M[�>�р/6�h�Ղ7�����7�Sh7@^j�PMwd�����p���:E�J���"�t��[�Cu�bԆ��>���D�+M��g�j���`Ha_y�Od
S�7�Ҷ�P��&r`�s����'줓M8�WtBk#txHp�S@0���J�� �<���0֯�x	���n$�Y�:�Q��y1`Z�޶�^g��gtq�Q���>����sYhY�?�P�co��o��o$��%��X���sRP��0���	��m�+��X"9V����}�]L4.�������G}�mx��!|�\�|�]EW|���b�F��;����<�ɇ4K*�7��q�w9��'�&[#G�����^].�����'?��/~��q�tZ��w~5���l.u�f�1��8t������5�r�_�w��Xl;Έ�{
a���l�׃����5�O%/�n�yY��{潸��x�
���!w�AӦm��6p�05�[�x�Q��8��Q�+�_�����{��uWf������,?�-�3t<�T���FG���/���Γq�&�T����F�Y�
3^|��x�3��[>>[�x'�J�teE��<]>v���ƨ�m��0*���X��&_�:�+�a�O8�~6Q�Ufm�05͊���Q��73z�Z�QQl����t��d#�������p������:���Y"Q�
 H�]�q"y]��8�5
������U�,��������ԓ]!��7n�A�����!r��?;� �s?�N;;SR���p�V^�|����{AU�ܗ�LM/7��<x=�i���E������ˇ_<�R3T��Zqg*�u~|�Ja��tz��,Q��f���hA�,�3�A��g��z�ڵ6 ����e5��
�\5�y���,w�F@��#�X�T�
�,@z����7���)�#{{�;��\w��CI��x�U�CL�����TI5:� J6�)XD+J6���t�vʃG�[�޺{��$�ie��b4%?3����A���R���u��e`�{������8��,/���Nd#��`cd{k��,��{����RM"A�<�͛7���dt��K�`�ދq��m�����ϟ˧$��o��D�"��m{ �	c��r��T�.�u�U�;�nZ���#�|d\�f#�
��hϟ���ε�`����n�l�랓C��ye}Z%4yE�g4�zQqʡ��;�r�[�V�o�ӛ�61]:x�Z)S���c���|�g�����-Qm����A��2e3Uv�c�����k�z��t�5�V$�gE��N|a�`0RɅ�X��#�jn_�#�":�ߋ�ӻ-'!hbh����Ǐ_��~)o�MT����
��a��J9|'�g�&�o ����?�K/"�X���@�VS�gONe��>A�C)z$G'�TW�b*�j�Ŕǔ��#��݄KM"�j$:�	�� G��D�J��x������0`S����t����N��n�V<��#1Z�� M� �o�}�G��5�ٙ�ԁ���|A~�Cy�㞁k>b]q����7w6���qw���ɳ�m�÷.���d��72����y��~bP4%�l���	{'�)��E�)2b��:Q�)1	q,�e��>���n�	�h�yf���C���+3X�)qU�ja=�� �-6N~f�u���H^�3Y�G>�2nl�+y4����*����R>�C=k�u({��2�@���iI�h�b<!�VY�\	GJ����]�����5��VƶC�)�UaC�����1u�?:!]�~ �����WL�r�'����V8�Xn��4�s���P��atCIWd�U̓�z����Dq͍��22>u��:�|�[G���_n��Ji�0�I� �C8R���F��}�C%���I��M�Tg#hzt6�+mV5�pT��7o�1w�o����_�����?����[����g�}vtE������������_Xl�"�)�KpH��Z�v��Ω����n�$�)���=I}i��@J<u,�F��J-R�x��Z���;��g���G��o��
�����f:^棏~��ɋE�ވ�U�bJ�B�Cu|���H�Q���ba�ƚ�ٓ��p%x��T�]rt����R*�t��� )U'g�]=�聱���'*�̀մ�yV��7q�{0,�$�F��6�^9��I *�����W��qIy*�x�����j��#Αگ,nM�[���y�H�q�+�������*2�����t�Y�d�u&g��NU�
��P�A ���%�-�)[K���������g�H��/�,���j���Ps�y������_D�)P��nݛy�{����nő�������/�Q�5�Osd�o��Z�Ja=����>���/�~�kx�isO�=|@�[f��A�����8�1�����/�]�	�3��z^T�/֮��Ȉ*o(7�8���@��ڵ�w���.�9��kf�8b�&�G|s�)�U�9'�0�E�s�΃Ĳ���=���z����V���T��Z	����.� B��E-�xvM��!V��_i�4�w���#_C׫�#qh����Q�y!�G�1Q���m����=���LøU������s��\ޏ~������N�=�Z�$+܄V<l��F�A�j�0%�Ǽ0e5�<.'���������mD#��N|��P�:d�/ԡ;�m\r<�͑ϲ�<6�-k=amex4��K��p�q�m1��X1�����*{��o~��W�먊I��〻����ow5:���
!R��;gV��@(%1����1*S�r�����j?8�\�3r���rE�L ��!�2��s�4���}�7hZ���
��4���ȇ]��K�?#�uLh��{�����3Pj�$� |�<���/L�������Q^p5�-݄#ⷾ�M<%9���nߒ����|0��#벡/�mLLY�-mVh�¶�kU������o�V���w����kѴ��o�����w��n�/	g�X1zn�6��NA��N�O/�
J��+g,_!Q� E�,v��r���~����xƥ�aWt���&�M�Pa�κn<w��9��F�W�q���,=�g
v�K��G�!i�Ŋ�QI�c��	�Rj6Pҩ�%j(�Z�C/��6 t�@�X�b�fO��r�`�[���z-��:��}_�|~~\��ԆR|��[����>s4a���v���ԁ�%jF(���	����0�)�a|�i�Z��gT@�/�SG�'
�?ln$�t!������PJB��6^~�����8O���.�$�k=��|)����ދ���~CY?��j���cIy�B�����#����2�����6]�y�D�8���="�U�A�o�˙<��,̿�����;;]��Rs�4��繡�tHrO�Дg\.,P��Ak�ѩ &�E�������*Jbr�!AC.j+�7�w��Y�Mߴ(S�aK�iG��w�12��	|�u�.����!am�a-O�e,�1�	��b�^o8�V�����, �R��F���L����b&�MA�B��2k )�t7ۤk7U�\m@������QM1zyr������q������S#�a��# ��&��"{�h���<D��������U�����!D�Sd�D�A�^qD�s*�o���_&�*q��ޠ��
4�ID:�A��ѱ�g�:=$�s3���df�Z�M9E�R�O���*y^)�g����%ġ���[����"�	rY���B������u8����u��˦�N�����ݻ�Q��Β \�η'P�)Q����iٰM�w���!J�S��b)��Np{�Uhe��G��^扺$p�8h0w�N|��sx��u8����Yо�c��_ �����w�ٔ�EG:^'iT�s�a,**"�8�!Q�n�p t��98�Ah�V&�`4���uIφ@�NK���%����������dr�qW��;��o߾-�$��:�C�x?t�iﴭ�$M=�X
�>c�Y��L>r�2����.�$u��W����]v�#_{�5u���GO7�)9�pb����^�RĜ���GFV�ଷѸOG������pI�L���2���x
6,�o��$�8�%㈫�P6���g�=�����[nZ�<H���+=�m9���%��x'�Gy�ϧ�s��ڵm�i\�/��(�\�s��d[����g�������� X�u^�z���F̓�y�����QR7��w��~�������>���x����oN�;��u�gy��<V}�&J��s(W
)�P}	;��$wcfP�s��]N�{�#S�u��6Dqt��z`�"����t�d��_z֔P)R�Qu;-XCⶵ��'��Ӷ�3�ϗ�no��DV�`��?��?_���ǧ`�@�'��K{�����6�R�X��<G�ٌ���K�v#������6n&��� .>�+c�'R=)3�f|ր�%��6�Q4� vJ�\g\��$M�n�y�=����ة<��8�fp֟���6����7&�	o�#�3z��d\60��2����7��Y��>��nv��"sSdD/�!VZýi���W����S�:��f���}v�)i�2��q��duއ�E)��$��f�F�,
��?��T-��t����x����}�.m[&��v�F
�P�v�i���@�:�A��ŒG*TS+��4�bmb��(Ø)�Z�uҁxI�5�B���r�T��X,�j�Wu)0Ж�������C4���E�ErA�%�L����CGv$�v�v���߹-���/��u�!9���r������pd����K��eL��NҠ.�H�����a����j�{�^U$�Hцc��]�vh}zgw�)O�����/�P^���(E�A�2I�{
��ӥ��W� �.W�S�t�}	�=���/�0=ǔ"w�h��wi��N�  �Y��]�sj��W
���j*mm>X[#_}��!�2,JF����R��R�<CH�Ɏ0�%�+g��8�����C"��Gp�&�>Lt.���ȳR����$�%1}�z�@ʈ)���ω��8ϳiC̀���^�3V��s&���Q�\�F�{����Q�yL|R�!�dG[�W���D�J�y����@�i�ʰ���.���z��e��e&Z��V�D�Grڂ�R�Wf�FP�@��<��X�����G�������ݵs�A��Ҳ�"����{����'�yn��֫�d4[.�M���������6���~ZLsx
�]-Wgg��9?�TFbgq}��bo#��,������A�c��0��͊�������H��ٳg��'cz��-E��ܹC1��3+���PV���S���j��NG���:X��`�����u$�]��|<
����bN!a :(VA�ˍꆹ�����%R@Ʒno�}����`rDBv�
%��i���!�|��\��k�z�^�:��r�F�����w�Q�&�i�5O �:U$�/|��Ie��_)7��l�2����&qI@V[7��{�;������84r\:�����1�+�ź�����Q��%���F***��M��X��:3���lZ�8㢀��͓ �y���IL�fjFƍ#�bi
4�Nl+��<0��c]������E)�o�W�~���h.�q�����+�&\�	��P"}����	頇Z���1>H�Ǟ��7���ܤ&"����7��46�V���zV�֨Tm�X	HE0�e+����ur�?��ף�e�d:ɹ�쏰~���Adq@�ub����)]�7�9OJ����B_�:-h���޺��N��f�f�i��[���&y֊-3�զ~�����#�q�}�D+r�X�ti�E~���e��
L�x��ȶ���=T&�x���^H��m=2�S�?
�c�cz��Fl{�1���Ea:Pl���0��F'�|z4rY{�GwÄ`����8f}�t,�"؎y�w�JC�(�ZM4�;]�` ��P��{T��Z����|����n���/V��X�q�!@&��<4�'_�z��)��|n�\���~ʉ�s �2R��g0>�F�a���b�h��֨�s.{����L$�cl�	�1�6X�'���JV�i,��J=��:V&FAt�R70���Y���Ҋ�Y!�3Ī@ֆ������x�ǵ�]lO�W*�Pn�mD��m\��{G����܋�nAy!���GzԱ��-����:Si�&eYcUSb�����#,�#��N\1����&��4��8��sy��p����|��a�<Y�|�̎v6�eK����H��]�_�W1tQŞD<� ���b_&�sO�$VQ,)ׁ�*Z�J��H�z��$��O�#����]�Kaԭ`$�����l��7þ�� ���j��X����c�r�k���N��W\5�����n�����/��~<K4)+��ʍ=}�񠥧��iZ�w/�F�Z��\��P�TS���P᫬*~V���)Q�]�F����$w�O���2ya��<�&�N�I^M<yl�P5� �9�"�r��|�<�5�����j����q��~#_��F�{��4b�ji:W�@z�_B�-�E֖���NZcV�!�#�R�V燈GƠ4�Ӿ��v��B�!��:��E�G$\6�S �LR�c��;�g=2����O���@�?��Rd/T�a�F͎k����Zk!�jx�]��:����ecB��p��B����D�h�`������NQ�K�wŷ�h�d�u�����+Y7e(�PI��9�;Y��v���f<}��x� �'6���U��O���l���3�Z��ȧ����K/�*7��hݠaR79�g!x;4OY�X��k�iw0U\d\+����QU��l�t�@����qk ��K�ȯݹ{rr�^�ށ�q�3e�5�s׻0�5�؃�z�H|c��
� r��l�q���8̫b��8�'/��7��0UPc3�裏l�5�ox�T;K�$�����D�Ό~@�S�9y������S�vqM�X�f��8��G�q�r��h:��e�L����ʈ���t��ҋ�d1OOD���s1YEcjF�`.YF����~��$嗲J�����r�:s���vJ'
 �
�[ò��H#��.Q�y\=��dJ��Z�h4�G�S�ѩ��F=�����hp/�'͙ـ��}��>��4BM%���o[� �D�c?;�堍�LWn�
Tt�93/�/�]&��/,c��;��g;��B����)!3�r >�&��g��e�����FI3hx�<�n:�a#��V�۪x.ρ��E��a?o�F�������7b7mR��lQ���s��� �z�̐9i���"��.\^]�=�Y�:8�g�~���R1�����ͧ�~�����?�����>���ok�b�k4R�r+��H�f���ұ<��ٹ����T�P�ӻN�F�%���W_�9�X�C?sз:�aL!�\������Z���0$��uZ�w]/�!����>����?�PV�Sx��&r�Yޛ2���s���/Wkyq�@�֊�c@c�Db&��c����hz�����E6S�ҵ�B�X���头�kD���zy}y
����p����
�+@�p��j���@�t�'|M0��M�3��")��]���F��x Ղ9�ֳ_�ľrKM�^�@]MG��t��ĳ���L�q�y��pM��*��	�����f�z:��U�5���Q�FM��ݔO~e7���޵>���<�ɠ�q��t�3r�Z��̖���bhhk qd''#1�IEe�Zv�HB�8�s8�ΟiA˸V�=�Qۯ7k�m��Z
�C�d��j3-���G'��SlҴ����r�����}�Ap[��ZL��#��@"�<���P�齝��?;G�/��(�a��s�V#b)���孃\������f2�ޑ�j��O�e�T��^�T�3���T��S�Z�Γ�i�r�����v=e����9Tl�&�Bؙ�����]aYS�b���w�M&�F׍���g2Zۄ��1�`�w�����#NT����Ҏ�:�V�u�*5���V��� �w��19����j�q����ׇ�~�ֽ��ݻ7J�^����c��Lw�Xњ�W�1r��ƙ�T�d�q� Ȓձ�&bj�TL��T`��3dz��X�Ľ@-ރ���_{�m��4��n�j�0r�/v��Y�t�,�Y��Y�Ԛ��i�TL+�5��)�
�ℊ���y�wwwi�ĵ�K#��t���z�C�tU��,�N��Q�Q����n��D�� 	1�\3Ȫ�8�!���>�6.VG�DU�� �+1H���(�Q3Q*�\$��i,���_���lU�L�����|ww_P�S��Hr6��X�(�HК�v���?ME�&���V�J7�'�VUS7�
@E����s�a��s�q�ޫ����b2޻up�D2^��f�KEJ	�)��U*�Iv[�3��V$[��oڿu��;��*�m��gϞi ���nzNw�!(���tp��UTȑ�h�����4[|�\\ul��f�\�ЭL��AԠx&�(�?1�Qz,������-�y���Rl�Fr,�b� �,����f%��)k1����Xe��Sݵ��0� ĊX��-Q�r�-�&�J%BUBF�1���EY�f�ܹ#K��mrͤ��B˿��T2��vB�%fg�R�_]�%w2��J��-�c%^N�����5:�cӉ��A�E�r��Z���)�T���w�{�������+���8���a����<�B�B���t�Zl��WEκ��N�ӬS���A����Ū����R�Do[�8L��ξc�x9�ȇ2<]�b��l,��z���|�3�����o`��󥅊)���zY��#��u��ŝ�N|�V���3�S��}���4s��/��B\(�^�CyR9�r�G�J���k]�?e�����FQ�1{-�M��"ol���B��ԟ�B��ߵ�������Щ�2}�bҸ)b@�>d����"]�	���f'�_�^�m��c���N�>���n<����{�h��w?��ǟ?���6q��j3"�*g��aXMn�q�:yogO�W��{J��m,��L1=�ytf�P�T���2�]�I����~�(��˦o�啬�8�E*v�o�`,Xִ�^������U�	�s�\�M�Vy��Dq}h�#����c�*�K뼸i%)�x�FNO�����$5��4J�>���C�g3q-o�n�B�L$D�W�l��c���PH��N�xS�р�CrGǋx
vg�"�$�(z^Cм.I���������Hu*W��$2��t .�9�䯽���^c�|�j��9��K8��Jb�F����<�[Y�h���uԪ6@��s�-�/�9/�X�1nw���M>��w�SP�-ʲ�y���x�Q��{�"���GϞ^�)fF�_� �|!�轐�=�nt�a���ͦ
�$�۳�s��HP�绌<x���Z�E6� �{yu~zz���D��H�3M�kpL������F�A���h�+�M��Җ�DRӋ��o+��_����������˗�r�M�H��**�jL�X��^x+�����_��5��hy��s�P���u#�^v$���?K��Z^�խ��X!�8�M�,��wrd"����lw6?���ubJ���4��Kͱf�x�q�����A���4l���6�&5q..����V���)M���EG%␯���`V:���TY�Xgr%^�G�V"���Yu� �K�\\�㓓�����yS�T�L�����WiIlg6��O~�"��\/���9�ן�ɟ�v�|���G��j�e�5��3�1#��k�l�u�=sr~�{n��kL{�����Ю!{���y��ִ�8t��� %�+]|0��-:J��΅�(��Md
S���V�!�4$�bO�{8��3�<�Eb�	3����0wɂ(<�`�4��C�,�VC������<-0(<p�Hf�L��M�����R���O�
�}�����F�ׂ��81� іh�I������A7�Wz�E1IL?����e�"�E���$��a>�q��#��b��12~��X��֧�
y��˅���lr�p��zma��h�;�ѧ�)��;��+Eo�x;S�KM.ۨ�t�l��"���D�J1�
r�c����&��+�� 4��m��t3�R�"�ӈ�;��H�㞒t�h0+�{}y!�w����g���˗_}���#`�׏?f��8p��d]o�3�&3��JL�fj�Z]^����#H�|WM �wie��">���J\zub�@&Z�@;�u�����z�7&�RBu�2n%<�M�^,�Rm�*k�(�	j���x�(���Y2�ƥs�z�۴U�̪MecT�bMM*N{׎�ހ�*6�k�C�4��,�>�ݸ7��^�O<g���~��ua9#
�}�ZɢAIo�������4�Y�$HVr�ˌ���7�z��ҵ}0Ҭ����ɬď&�H"W�ႄ�7@�I�οzOAP���>��Dǿ��x���p}V%�L'3Lb����j(&��:a&Z�j��%ڔ$t_�͌��I�7�K���AsDȌƇ%ώ-Y��d�LA�3T禠���+N1S�Ŏ����{츻�@�T �W"�l���uݯ����
��A:�]���f���>�J�!����҂Q;������e��k�W �8���Jt4ۜ�v@7FL@Y��7�0�a0U��z��%���Kw���#��+�P��M,�*M8�/��s�2��|�֖	@�8�>��(��m�P\�"���>�usu�X��bgX��qI3�lng��cm	�ͫ�@�1�U8�ᘇ��Zqo���iߺ���A��sǋ���
�ϋ뵖M*�A�}�y��%�
kK��x���d&�	����^rg�`��4�?�%�޳������y2�V�C�uI5�����"�G�K����$����t8x��SGGG�������7����c��xܵ�{.�kv0{!��P��jZ�lF�W�}�W��KE��j�{��ޗ:�,��l��+ӝ��txጥ3wv'��Mͣasg�.���w���k8�]�~�x��s�"�e��sƳ�ecB�b�=��v�{|Y���<�y
�����˲�\~�H�q��t��l��d�D����X�����U�%kv��ݺ �Ȫ�^�<���{��8#�-�&�Na�Te�/�h}^nOt`��7�i�0�CT�6�eA-Ǿg'�L�z̸#������t9�C�����d�&��ht�v;}�W��^uRN�z��7���1AL���[��`8N� �	����jO0B�x���ҩ '��82��8U䧝Z���&��G�҉*ώQK�9#��G��T2��$~�
0;⚉Ci���>��g�f�-ҩ�{"�e�Nq�±�/��w��1���o��z������"0'J�������Q�x��u�@�\o�<��)!EJ.C�3�1�F\3�F3��sft�cjc�O�S� �S�l�!�]h�u�i�y.�͢���^��q!L���E�}�N!�]����Q$�6<�Zy���SIVvE�}[o���M?a��D�
�
��,�zڽ�֟�.�X���Xu`uS���v�ab�d'���H�lf�s?0�=���ӊhd��Ů���)���C� p=����" D�U�GWWWl'�C_�c%kծ�"�:sF�/;4�q�
�������i����>�'	C#Rè���:�at!0�}��qNB�Q6\�`)3j��B�����O�Sy
���"K��"?�L�y���Ow�p���\�~���τ
��E�ɽW��E7˅<����*�7��W7�D�A�ԻN�;�+"q�lW�驮N�r}��e���$b_���'O��Xճ�K��?��?��__\��?��\䣏>��,'�O>�կ~����T���AP�eLVv���ʷ�X�/��� �Ar��ܘVVvE�75�����|��7�L���bq)��}`&"� qz|��y�EZY��1��4nf4K������+���s�j��J"w�b�U���������A��x��/+t*\/�>xٍ����Տ���{xG>xq~�i�"@��A���g"I�"ܱ)dU.K��˛kH��<>B�f��싋+�E�d �J�,����3B+��&/�3Έu��"-���5��dͶU(�]�v��{���J8�ʡ��I���r�l��J�k5z��ggg�4�H�F�FY�ѤP��h5��l4���G�bHu�z\���L���D"�ǁ�$�п�O�l|ˮ�d>�(c$��<�ޔNQr�%#o��I��`�����s�ɫFWY�0�P�E�gY���W�H�蓾	&�s�P��u(��R�A�T��ļXyo-�r��J�1�{3W�>I����`o.&�����D����M�f�N��j���z8���s"�(7�H�Y�t��X*�",,�Cbj���v��]�ѥ�����X�J2�i�a��M�aG����4��(򍤱�{*�e�<El]r���{Y�����$iT؛�sS��4Û��V��*C�=\{�5�}��+����)�*��j6��A��(B�Z�	��g���:��η�ѫ�=�r,���X?���^K��A$���U��Q���v�i�_� ���%-�Z~;��N� �d�aCoU�OZ�nZ���m�<B�4��� nD̰0�Tg] f��bԸ�Wҗ=F*�&������B�ɳMQgH|�T��IAI+�����7-E�چ0c�f���\M�����#���c<DY��6�;ܐD���m�p�.�#V@�ަ�j��):�8���R���n�j����%���2�y�<���f�s�y5�7�;_u=�b�&C�
R#C����J<���Ʊ����ک�w��c�_y���ѰfHLb�{:ŵ��)�tQO���E�a����<h=Ee�-~!�0��X���5�U��n�Ͳ\�|6h����"���֥<1�t���7�c�=�$K�����*��q��&�f�ăf�ﱈ��?���^�V�?(�^�0ŀ��H��f�	]>=�m]��W7+���,��څ.r�2��`�W%�;!� iX��&�M����2�>�n}H-�$3eIRN���<����N��`���E(g�Z���Uf��y������ѓ'~��[o�'ِ��hyw1*�I)0=`��T�Aۄe�F�|��6�9�	k���O,�1��`�8c����Q��H� <鲈������a��4���!���5�DӸ�AW&��-����'֋|\&Y�DG)�&
I���Y`�m���)齇b�Z|��굉��{{9%A<0�8�YU�.��}�23w|����$W�r	2y��]�e~��?����r�/���׿���D��'	��+aF��c��6�d�[ܡ���6X<h��%>&�B3����A�K����L���v��S7-:�EYqұ%T�_J��Jp}f~t�����H9�� >e<��Q[Ʒ�gO�I� �7��јVh��b�����|�Fg��y����^'�&��|1��F� p��O�E�n�v�Q-؝qH�{C�0�xK�TL�īOG��x�\��������`���c��Ž�&�7�x������E��	����F�t:E��|��K~�˩ͦӕԼj��CR�ʏ��ܬdl%ܞ̦I�Dn���X�̲��}�U~��w �ٯ���";f��q���&��l��돤�<������Vo��3�1�E���>Z7����Z�_4ܦ�̠R�ޏ baO|��Ⴅ�,;��ȷ��dP�C�0I���\�^�8�(�F��~��{\�5'���c2���mJ1 ���&P42i�b�$�yY�p*G&��G�ER%eXt[>�	6������ղ����
`YL�=̤�6���g�b1c78�P�6�S��(��A��X�!q�i��f���� Z��e̱e����c>݁�BnE	�xk{�J�G�Ħ[/��^���ja|��|9 Ū���o�F�T��^��)� �������h=�?��4��#0���v�}�����O���9*J� Ȳ<�������`b�<y�(�`p�b%9!��G$��dBJ~8�{G~��o~�y�������H�[���S�R���eu��@[�W�hZ*�Tq�W��
��N�C�ttr���K�ֈAy��wO^��:�S�;�#?|�ч���D��?����:`��jݶ��LY"DK:݀�a|���F�D.E�����Q�o����R�ؗ'�d�����/�&���zn2����ǾiGl߰�R���d3r�Byȅ�z�.��J��x��WaC��BK��'"\��	�ъ���AV��A�5q3�l�D���������Ewg�����x����B�S��$WFuߟ��������V+�v���l<�/�q/����3%���7�4����ŋ�c*F&��3��z񩑅�s�o�"y�GgqQ�	�H�{�{ �1.��up�9,�Yn9đ�̶���bXCߓg}m&��~�z����E�-��T����AeE���XR���)��S�2+��3'JWn��B�2VKM���l������{�:A�]�v0�(ػ޷�C�p@�v��p$1O�͕Ę�}��a��K�͉���hńN�����	]�^,�񗽶�r9��݅$,I6���bg���\�>�3;�v-�D����Ztl�&ͦL��NL�����k^M�w�oh��0�/0�m��6���Z�V'LA�F�8�,C�R1Za�Db�e���D|k�J������Z����-$I�z]=��]!�,֤� ��u��u�h�rOl�*W:X�g�����K��  U�����^�IRY�H��K�,i�������y�V�����Ԏ��8wN�#����� ��\�7�p�����]6K�0ߝǞ��pߒz�5���G1dy �C������}VU�B=��ț���Ģ�S�!�Q���a ��{��Ϫ�H���`����a��\$z��؄;���0��o�[#�p���إ/��$�s�a΢�ͽ��v��~X{X��7�ӌ����kh���Q�+~o@"�W�3f���=|�Y�X��F]KfU���s���MM�AO7(
�7Ʒ��:� ��E�����H�zћ_~�%�5��paEkk׶��9��X��e�W������N�C3x����X����l����B4c�L� �a��ZwR研ZV�o��a��̻`L���U�bJ[G��u��y'b�(� }s��=p�H0�\'��YWOH��9�D�0�S�}I�f�g~���x.�A@��`:Q�U`�ۯ��>���
v7�lT�8��ꕬp.����a�_�{j<���d�9���1����;����o}��Z�cF1&1��B��c�2Ͷ#VO<y�?˰���!��g頇o����������(|3E�)9��{W=[31�T��1�p�kQ�,�`"s�x���sH��R7[pk+ၪ��[o���� �
�<�����;~�et-AE�]��
A�?K�w`OeoP�����*�%ͧV;�#EU���T��[e�W�A9��zR,�B��1� <�u�|I�!�8*��y�c3�Fm��#�3�,7N	�<�3�lt����"� ,M��;�t�[�(V�}d�դ��=�3S�D���_��;w��fd�%$�SK���c���N�N�}U5�&X�^�z4L��|�x���YMe�@�Y�؄������u���&A���(\Q�#ܹ���r��3�}xKԲ,3 ������Y�!Z�\�tf2b���T������U�k���o	�9�3ᩃe��rC�$���W�%����F-��JQH��,�g��j)E��	�[ּ�1��|U�v~�EMǣ�����~���,m�Ď�tb����s�b~�+c�RB�?��'��t�x�[����)�����ǆ�-�g¿4�73����Yޗ{ΊT��pFJ�뫙fI����|����?��?�_.(�b�d���rc>��sr\�~<T���B�o-��)d��Gv�(.Į|�bp���f���ȗ��ؑ�p�8ٴ�m�v04]]a�z:Bۓ�{�P�=�9�d3�*��wz;ȼ�i�{ɶZ2��;�Hcj��a��c� �X!i|�T�6p�=����A]�FK��;�mpfx�q�����OF	����3�jd�vp�e�V:	�%b<2��!B	���d�M�tЌ��Ը ��S��M��?]�M������UFQ�]��|��ݻm���������)���ՠ��7J-GD*`V{�}�����'���m���;===99��_���-��|�\�\ܰF�����JN(��V�i�z�f�O������|�H�#Ρ<�t������Y^{���2j�����6�m4`�V�� �0�2��!l������yQ��^�5`�7�B���1�\]3ז)w�)�����.�7v]8���t g������1��yӸN���b���￙:Æ�g���<mt�]�K�!��+0E�� ˻���My��	J}��T(t�"�����wd���A+����e�h�"����#����fE2^s�J�j8��F�BV���=\/�4O:�gؔ1������*� �P�����ʭ�C���h�kS¨��EB�����{x�{�cO)Hw�f���N��<�t���V��	�[�n�o2s�9˔NN98�������O~��9]�O_�ӝ�A�~����ͧ#��[N�(qi���EИ��C�4��]Re�P����KE����I������bd�w�3n\ ��daȟ�w�B��[�$/ڣ�������0�߿����#P�����I1Q�j�������l�@��i�eRx!&��J�W��bU��J�֟P��i����WYY��O�e.�L��FaH�y?-�7�u~~�"暮��'��L�.����9�<�8�p :����M�n�b<�	�n�SJ�_���$k�|D���mL�8:~)!��Ǐ���XCD<:��;ߨ�g�>1}�>J��$ً�Us6:�y)'K���(��m��=��n���Bi�$��.n1��M]�%������Z�6؃��0;2~�) �G��tjr7����h@��Dz��@�3���!Hi*M�@w��i0���Yd��6��$�[�9)�\�^�k:6`k_*�al�X-q�������|��Ql#���(��sr�ڣ)JP�<b���v.ހ�0$�S�\�\��s�x5��$j�:ht7�f}���Uo�@E�oY�SǄHc�JHj ��`ćM̚!뢃���KtYO��n��{sƙ;b�{���¶,�7�q���&aY�Y��*��n�̉v@Mm�;/?�ۢ��w=���r��h�I�6L~����0��z6+�yR9��zñ���sZ�$�	������fl"�k/�"�&�E1���:�#h#37��
y����[��3�a��D�V���	�lQ$bW�#����Qt-���wO�O/�}������֭��S��E>��KU@��P�r�=��L4��#�
��y�!{
uѶ�(�E�N���y�#����D�}��7��WB�XT��(խΙm�{4��P�5��Nv~���P�P�.�rc��^�S#�%&��s�X-ђ�s�V�����n��`3���1b��+/0�FP�Y�j���x2��>j4#�3�^�^߬��E}��>T'�Bƫ�H�HJ������[Oo�p,h�<eJ�ص�������@ҏ�6�%����}g������:%�	�)~����_)�_��|.�/4���nS�P�l�C�G����	���,��WѬr:�&���x@N
�%��/�z҉J	��o������V:�ƣ��BBw��Ag�^E~��~D�$��T�j���0��Anu� o��?N.c%�}����bfL��g0��cд�c�ůs��X���k?7�<�f��3Q��\�ES/sKJ�4V��䃗`q���,��yC�-�����K*�ҽ{�����MrL��x����P�5R�sO���1aʐ���E�T�A���yPz�Xw:�s��o\�+�]C�C���:�q���ҰfnR-�/y��ք�T�������y ���9��h����aŉ�lW�'��ݻ}��㖩g^A�ړ��t���W�R+�&�onb�>M�����1��S�f^��7��L��z�S��U�s�p���JX��'�e���5>�b��ΛHs`z�~�].{$>=R��1*/	����������S���j��n���Ѿz�H,=˟C�H����䣥��jNvU�p��+�z�z�eYߍ
��~`(�[b��F��ﶳ�#�?����Օ|^B
�#�G,k"
�ҳ�$}(cL�%��Ή�yjW`6i6��c�y��x�'����EY�*Wde9O/.M���ԠO,t��f\9GV�SW�S� ��I�v��G��Nz�m�@�6��i֕��;�hc�Ϣ{�L�j��%rV� <t�!��n��s�53|!1B8#�|�T�j�|����+�`���8�Y׷����L���;wn�M��V+�ͺq?�c��>n(<8����Um���:%)������Ә�U���������ce4���f�P/1b7�"A4��լ]���Y�ɼq��\���_G��H�J,~���r�ݝ=T!�)��׈��u�����ۘ�t}���^�_�Q�����nY7���ӓ�B!�u��4��dT����"d�FN�<��'O�vߏ�Ι��(~��g���"iǧ�7WW������:M�����!��憵� �dD@[�ZZ�����D��8�.7g���Iq��V�q<�:m���A���SE܋T+�>G����!��]���%�J�y�>'�`9�:�'���҈#x�}OLlz(����_��3 �{���H����8�)�c�'�h.G�_��_�ӟ�ɚ�br̏Uutt���(����N�D�lW�e��yy�O&��=z�M*Ez\^��5�Pa���y�œKS��,Ө������objꪚ1Ʊԫ��F��$� �\V"0eU/��z��q�bzI������Kn�nCǞڒ�ή�n0�/�s��ѲgØ���*�j���*�ki��JK���2�{��T~��o�������d�o��� F���ꫯ�z��;��o}���8_,�S����4���=��G��ב������g?��?�u��q���$�qCy�����	D���K���ǏE1�<�y&e�b4����%a���h�ф�(
S��ܬ��X��4�o`~�ř����[�ǆ�;e�����5��\I�È�yP��6e��w�a��
����T��M��u�7��Q�/�i�J�f�)�C�D~Vzh��t� J�\��{��_L�^-�����+v
p�n������C����Z]h��/E���^,1�t�/�8��0}�фTȟ��!���k�G��
���y�B���;*����$H�؏
N/�B��s�>��!��M�F;��
3j�԰�fu.��k�޽s='3L�|�~ �B����e.��a#ݫ�`�h��`�+T�8؆�YOVe�s�w���DC�	��J��!��<��߻`��Cv��#�_��^��	U�pKn5��ف��_�8|���I4h?4Z�W
#$8�hf�cTF%ˇ�7f��Z���^0(��O�w���<ꙹ:F�jۋVX[��O�]Bf��9ih�Ja�ġ���љ>��5��a��Sh�u�q!�C��2�LftH�����b"ac��i
�Mӄ����J[@�px�����4ʅ�9@���d��Ƴk�y���&�M�St$`�#�䐉>ډ𰉟L�UP�C�iB���71�ź�0(�&�b�q�2�#+��_��;��7�u��J=c~�$X��|��v���!�6TA!�C�;�V	�<�p�Ն��� WC6����d��Q�X%��	`	�'�<u���S���<�|�D��d��Z�d�1N��}Z�g�oރ�顠:���Z'��������S�h5١<jQ͓�iGR��$nҴ@v�'S��_G�Gq�3r��҄,�^�nN��������� 0t�?d��jA��2n�����3\V�[�}�����A�9�iK�|I�R� ��v*�i����;Mg��=c����i)�FY�?T�� �<M83�C�4���ܰ/�jh��������3���F�,�%�'o 6��W<�ܴ<,��8�C��:�%��gp�#�ʹ�!R�����?D���N�!�'<�<�dO�?�6J2k������ҹ�)�Ր�>/�Lז���͈#�'�?U�칄����B(}�q�X��A&R�����#m�1~��^JT��)νqϥ�����%_X�%�oM�~Hn���C.����3K�.�n�n:�a�wũ���;d=yS��������%D�Wr$��f��,?3��h��A�9j���H��:����6��!!����V��Dp�F����+/�H��m�厢�'m��9D\aСQ��t7I��/��W����2���D�{rr������ ����ƱC����Hc��� ���6a��p�g���#�%��Eu�_��l���
w��[��� �R��ڨҜ5K�dTkAӺ}4���:���n�v��͐�,R�(!Ɔ��ۻ��4�:�Ac�r������Ⱥ�
~o���r���$��Gգ��emX�S C�ZY8�^������Z����t�Ҹ�5�F���'��������(�����!N��Ƀ�b;��!̜N6 l�wl�(��?�X\'fl3�@Ji��������,�޽3�	i�OB��E�\������S����hi��X�pq��	{r�8��^[X��7p͍*m�s����~���>y��>|(1�|Q�Q(7 �`����S)��˗/�3�Q�e�/*
Y���C���W���o�a��3��9�1M�&����o����̳]��t<���`�t>�Z+CUa�<y���ϟ?�;��1�F)ݍ��z������Tǿʖ,�������hlW� ���G)���j��8ˇNl�!8/��c�N>�:ׅ����e�X��j�۶��EG�4O��v��{����L��� �.w(��\\CKl�z��G%�Hq���w�}�2!܌�Hw*�����S��ݻwY>�ۘVNM�j�-ծ��$���1�w�ܹή��KT�G9�Z�Eyzz*�1�̀`!�jˁqz@Z�/T+�"���� ��'�#���$kHl
��cn�4뭷��������x�R������Q�30t'��:ů�(4���2��(����Ɨ��aKo�w�y�G?�џ���s�D�A��.o��?�Y�=�h	�a�zk��Q��_�ŉ�����p`:uL��U��E�����*���rY������5)z��Z�02�:U���X�f�\�tg�\ޗ:�L�ɲ=�+r�� �6��&�5s��9�V���#�mj�$b3�&+T-i��EЊq��Q7c�[���!6	m=�S69�r��('ə�=�;[7���	$I���@�ϯE����/���1�i���y�&�#[Yn���\�����Z�U��5U�;�L��� ���o`�.{��dByK���F3�Đ�X�r�RŌ�B�U�.������&ڷ��)F���,�.;n�NLj%�z��W�kC�! ����V�'��Z/3\��f�p���q}t
�{ݼp�=i��X-�b�P�gG|��� �%{f�6�AK(��f�p�i����y�^4 �٨��"���/+x�Cb��b=d���HƉp���q;BA�nw����J��z��z�0H��8G|+HU�N�ŏƲ���� �5��0.WM�s��APdj�Vڞ�BY�v�z|S�_�v@�:a����1�}@�6͵�r�����×.`����xr�sr�p�,ךB��	����Jt��9���;
����&f�����cdxb��'s-I��ĥ��Sbc��0���.��`��֩:�s`�'��q)�VM]CL�����{CT��+
G4����8��d��YhR(&��E���I�pֺM��EY>�n>�ʶn{1;s@	������DЩq�|/#=�d�.���w:)�A�����SB3��3H���l_-!�����ȇ�H����6�,�ͦ��< .�h�A:V�[̠H���a�Yx�U�6ؐ"'.�mU���&�Z��!M���4�S)b*(F5$�!�D�/5+]3~�<��[o�sY��p�d��Y�N'9*Z��o�:��ʖ-9pJ$o�N�����u�۬���B�:�O4	��._cYFy�F���#GR�'�k���݆�s�B;W5���^E��\s�:�>v�]M����tHB�c@-@��/�Q�X�|��i�e��j�c[+�>�hm(���ݬ��⚻C�d��5����0@�8o�b�zD��Y`�g�X8"(@։v�Y��#6��J�!�������@|���L�i�� P#ʄ�jS���	l��$�Ԣ�=\++����w2a(<���&
����L��:y�Jz��t��1�DL"S�buA����e�EOR����e=b�A,���.$q��;>:��#�FluJ	�74�7޳�^����~���o��$EĘ2/D��ۑ���s�5O�'�0�?���4n����׷�+�m���
�ـj��;�YaCi;����R�q���5�p�}��ro��g)n˦Z��L�c�
�D�h��V=����\� �����XZO�i}�Z?`|fƖ�� �"�;YV��t��]���g���Gi��S�'�t2��I�XܬeY�^\g# 6������ؚ$�^mZњr���i�Oo�ڗ�d2K����/�~���4�̦TD̠1�{�K�kGL	U�=�*Se�E/���_����-�\���	Yh1M��.	�u���U��B{�={��7�\_a�#ó�|��W2c� W�PeĴ��ZAg�^hL�Sk����4uV7;=��uŁ9}\��5��=_#���j�x(u!���$�)>��1'q<��.��a�7t��3�}���# 
��w�Hf��l[7��ͺ�։��2'��wѮ���������eU����j�����
��f�9�"Ҳ�"!r��x�%t��~�7%�`�ŋ'g�jӣ�92��.�*�@E�b�y�� 	�w�>��K�E�C?�J������4�[����)[f�$���Y�H;��b4�r1�c�Y�����fw�����ٳ/כJ<��˧�^2g��j-N D�!_:�J4^�i1��:6.�G?��w���|q|��v�p<��P4<�|���uu|tdM�Z/d��ʚ���u;{�w��}뭷�<zD��K,�p���8�.b*��<� �A@�ƟJ���ֶ��'���h;���h�7eU��H5^߼6�ˊ�2;Q����bɡ������a4F�Y�����益�c~s���ٳ�W<����l�#?ݹ`/��(��!j��)v�� é'#搁��c�M�E���D*����1�A�tY1���˪��P��=::�ꫯ~��O�O�����*�'�ۤ.�����3�PoW����8�vo���zbp�
ώ�eeĥ�j~�����b>�c��Z;uS��R$!�=�c�]�����u�ط�4�̝}�T�I�*�Y���y����ȉ��	yL��Ʊ/V�1���o��#n�����h!L�3�r�ȋ����1�A
3c=��I\�^� ��R�s����"�<�9Tx�҄�t��6���i��������A��h����c�Q��Tb��eAT�eJ�)y��!RT�JM.F��ڻ�ӟ����0����;w�?�ϟ?���/�dr���R�)a��sgW�8���z��x��\�q��H�X��~�/_��\3=�VY��1�&[6��R�.-gBū'��ә���ز{��ь)& ç�ɇ��� 8p������B�4����C���0,��UuxpK�������p�T?9�h7K��Gv��&����I
�2��:�Xn.e��)CO��a�
�R�������i�f�ܸX�D<B�*�x�j���*.P��9n�i�װ��V���]d�#b<��v�'+��e! Ѡ���Q���M̠f�i���5Ư�:�OI��q�	F�<E��l=)U4�`�ǪJ���O�l+�<��l'Ĕ�����_�`d��u���фo7��UX(;����C:�W�J��G���hr����ۘ�o�U��qw:����zR�R�2��aP��E�}^����&6a��}�t�;Z<@y�O����]l��dO��׿R�� �� ��tZiI�0G� �5|�%Eʤc#,�P�dX \\<*�߭ΰ�!�t����}�Y�я0"B���-ZI�+
��_:�r�`66�9C%�h#��2���w.Z���k�*H����Q"�I�؏�@���ZN���/�_��@1��U�n�RE/Z�6�.X#Nr�x����|~��g�-nz�s�A�����"�y�?b|0��t�0z�2.}��X���zi�6�X��v�%��4e�e?8Ek�<�B|%�{2S��Ⱥ��$���r�(�*�+�M�4C�H��Y�ۢ�CD ��G���*��Q�4���2��{�F=	��7]��CũS�T���'���'� ��/��y���~4�p��j�Qd��Ǚ�[���u��:�'����ȿ�"�U}�k��Ɨ��=�͊}Oz�9F%��{,�(㇦��e���i���z���i��#���:��*.�S
eH��܏�)	kŁ�ML��W��L��:�f�dz,5�|�l��r�.^A�L=җ�+�"��"4���C�D/0�ę<&&�i�)���S�"er��Q!��xȧ|J�D�c�J�Ob�/�����q�5�]i�*BSW�x���:i�ֈ�mZ'ZV�"���9����o�����5�6��,��>�D�ڠس`����[�br�:pu&i㠗z�VC1?+��GZ_�X��@(W���}qȦe����n0t�W]6�N���W�:����)�z��v4E�� T��`DJ�&
��ǳ�Be�5%����m�U����6պ�����|E8��"߃�x�hՖ.�Ӄ���#9&�8�����R���K���y�� k��$.�4�+s���L'a�����u�Q�\3�]%SF|k�`⇥��I�$�g�F"x�.a�� ����BK�t�so�BEB����6��ܭ<����7ޖ3H������3%�IQ�0�u�j5B�Kӝ�Yi}:�3^+�m1��s��&���੧�H�G�y�k�/�0�%�9�X՝�X����(��x7�+�G#�mþFܒ�C-�`�'MN�F1ϋ	H�7����ͳ��I���j��OQZho.��ʣ+_()���9=�gD���S'�3G��Ծ��%~���@b���?	���R�Sp��]w����󋣣#N{�6�GRN�	�3�|��)%�r���,���X���s%k;V��:m͛k�
H������`����?�+�9;?������0ۮi~�������/��/��,gn
3��h��R<\��)�;��X��}�ѣo�}��)Ղ���m=��i����ă��W�Դ(0(�C��S��ѩfQ����=��Vy��H�M�O�����x,�E��ٳg�<�4����q ���s���������^<?�)�8�����&>f� 5v��*��	�bϭ��p���#�PuB�i^�{�uY���A9:��Z���S��"�;K��ֽ���o�~O����I���><;=�C�2 �"��Q��*�.�!R$zB����:�>~��_��_�?(O�{den߾}����k���,^V�3б��Ы�c���6��O�
��X�eY���T��������jp�c��$�#��P�g����������r��E]s��;[j`�e �M��1��N]a��S�(ɱQ�]�oX�~2�n��I�%��T�����#Jh-�L��vqe�$r��E"��3��cC�X
�����	�c�UDQ�^.���Y�I䠬���"3�Y�!�>"E8���Q¹/r�d��<���H��D���ggt�G������Ρ�j���wrF�A$	�\~�)W�vZ���$;;6�P\-�k�&�'x�x]m���Ϟ���Q����˗/�>�x_�
7�AN\�^	�j�����?-n��2C��Q?@O���򟱟k\����Mc�ir�P[���a�|���5ld7-B�g5�K.�6�#��ŎI�50u�׌)��:�	P�������#7K�k��E���WI���y�[�L�
ޫ6������#���x�0GWB)?GȀ�&)&\ŠiڐhP��|�n��s��AF�"�О��õQ#��t�0i�JZ��s��f�P�B�Һ!V_p}��8��x�t��s�����a���qgw2�K�U_�PKG���4�C�F�@�,���y>)
.��@#g��cO�ijմkPʇ3]Ղ,�vnءܻ1����d~P?^��T�����P)����$$M�ۊ�;��l,τ�\�沗/�����|��y��Ey���mŚ�tyװ6�\$ݝD]LƜ40��Ш�C� 07qPr8>!OG	G��#&�7��NM�	��l��Lq�2	o��"�֝#����E	�7�b4���m��4�	��Mw6�=rt~}c�"5�f������Q`�lM��6����k��z�:V��V y�:� ����A�ɑ\���;g:$憑3w��Ĩ.D&��}�I��8�CN}��夀f����ȏp��5-�:v%p3�;c�m[�P1F�*x*��k�ja�C�"|F�+~�}`H}�@�v]� q�(j�5�z,����j��QH��j�s��LG0�"_���S�Ъ��[l�i�8+&E�Ի�b��=�\�q����\��w��`~�V&	Ħ޾} �H�c���c^P�6���`G�[�6��c��0պQ���:l�M��%!A�n1��@r�PJ!fC��{<�-Q	��j����|�X		{.��㩢Zz�݃s?V?���츱����>ML�S��i�Hι�D��c�zk��,G��u�P��D��J�M�,E���.[�	%�5e@�&Wo䔁����"�����>?9�=oCS!c�\	W����e0�Ҡ�:|��:8bŲ-�Nx&��S�_#�^�����2�nd��N�Z�~jow6�bf�ʵ�T1Q~z:P�#:��2%G~*�,	:-�����~g�w��J�	L~I��N�b/^��L4�f��3GŸ�8��tvG�}>��T�3��>�U:E[�&�ynVFҋH��U�z&2�؆y^�I�<� k�w���˧.�zUnVKm�)��D���cU�V��|��i���ԅ����V��}�D6}R��f�XF�ڌv`Sߠ���	:皃�#eW$��Z��,/��'i"&�y1��rݜ��&v�����r��g�uXw�+hM�(7�,׃��N��n�ٹG�AU����8G�|]����M%߳��F����6�nv�J{�w}�	4�����]�R���שN�n��S)0���N�MSE2�C�`�I������D�(L�yTf>�K +�c�%W*k�j��O]\^��Q�(�	״�MH4�G.�k��Xlq4]�V�Lf��u������C*�E:g���7&~��u�q4iM,'5���t��쏨�"ܣ8t~zq�m���QѦ��8)��֚M�N��˾�$_�M-����8$ڃbR�nL"AS!+15�t2/ƣ�tr�Ϗ��ܜ��\���c,��{�݆�j���11�2n4��D�����W7׏�>q(��ŁG
�ȱ�����tP�g,�b�g�Q�Ѳ�eUȿ����O~"�\��6Y{e�8����A�v�+0�ًP��:==����'�Pu�34$���D��ݻ���E�ZW�gr�b�on�:kx���.����Kd	�]�~���?������Ǐ�G�o3ʍh��������w����Й��z�Պ|d��*{��	O�ڌ몯ћ1
˩l��O؛�Jv\W�q��X�XE�Iɢ��2��р��Ҁ�_k�CC��ݰ$����N9����+"2��ݝ�[�f�<'b��^;3<��j���`�{�PSc��,pyl%s=�iO���,I�C�R%sF��:���ͺ��Q6�8�j�T�ٻ�<­`��>�~Ϭ�T�LA�G�ɣw��<�X%fUf�3:H%�ڻ������~��/������qc�dF�'�"z?���=����d<Nj��HCkt�1́
_�,���Us#�]oh�qKg�'f|�����Vc{�����?���/���?|��Ǐ��͎�o?z����[�;B5�o�Nl���C]A��*�&{t�xk�Ի�hr��nt|ۆ��u~��_�O_qhdiAX��������,,�p��c�1�ep�!�}�0��2��1��%׉P.5x�K�yh4VԦHS1�
rjg��Ԋg��1T�����jo�%��'�]�a�5��1����*PJ:V��Ў���=���t�\HX��kΥ)<޼�oH-�2�����H��_Ȱ��!�hr9,%��T}LC>p�m���p��t�A\����W������,�O��:9K{w��r<+��`�/._⯱^���z'��6Z�K%Lyֶ�8�(9�6l
�6���%��(I=Y�6ަ�B�$L��^b�a>Y5/<��gx~�����q���<;���zTK�UZ���M��AH��c��dL�Vm8ӯo�����A7}�w�`K���vB�a��z[E�g����hz�nk�ؗ]��ZNmx� ΢��IF~���D2,=���o�T�:��xt�+�iB2�[������nGH�E8�M�C�]����L���2-~
1G��^��q��/�J��vL~<�x��ÄN� Z�$������@�&Ɉ����ӈ�zE9Mi����P���/��x�bB*Vc
#&wxo��$�8��)0�.P$8a�����o��cZ�bF#�W9ߪ9��[�U�Ŋ��`��seY��$☲��������v��c�$�eŚy*	�s�9Tv��%��A�|��XZ<L���?�/%z�˚U��ɓ��fE��R�=[��7�i��"B��O�q�*���K�D������9��*v��Z�Ɨpڡ2?�
voƲ�Uei�j؇&�ja��>((Szp�Ώ������Êwio�ʭU�W����~2�H�����?�i�聡k�-CJJ
�R/pF���m�C��Q�c>�d㏉>㑉��'�4tlE���|���C_�K�r�m�Ⓞ�l�J�4�̂�I�]�<�i?�/L�j�S���FVٷ8�tBL���0a���{�sH%'�mh�]7ĬD@Ψ��P۠�®�g��l�l��OYK$G�/>��i��"O;%���M��.�YD�D���u��E�;8'�߹
����z��p��b��leWVj��ЪN���d%~J�?�>��2�Y�1A�lb����^}Yt��N�niO�f��D�` �I��̆��i_|�avZ:��Kx"�@��P�})��)�5�_&�R,Q�wG��ٙf�!�����'��]2�
<�!=62�c{�N�YA���7�\\,tqgY���cAތǐ]��s��o��>��u%W�b�N�_��
�`<��
Pq>/R{4�����O��*�,m*�N�O��|�#��9�-6.��Q����I���Z�I�����A�xK�I�
-�tӉ"7ϧ4n��r��w�^G�$��i�)OMp���tLˡ;a�$n�JJ��d�"FL�mmyҢ�^8���h:�`A����e�dmM��`�6M=DW�n-�
~6Zn8�M�|�X[V׉iP�vr����Q",������Q1df6R��O�v�Yg����f�Zb?l�}����T���E��E��A��=w�̱�E�2��r�!da� c�eQ&T/9u3�w����kkY�v��K<��'NB�@�.k,���L��D���c�+�>m��R8��˚��������͗1���am{���f�'6��r�&��h>�ȳ�$0�X�� �[a[ɰ�Z49��B�Ԧ��7���{G�KlJr��)B������	1\a���]��r%j[1�,	8��Ȅ�q�?~�x�M��={��/>'��(�(�ʶZ����T�]2�1Di�`Ir����w���ݻ�ɳ�U���9��}���g�}�� ��a�6lǏva�<[�f_���Sz��tk$\�5[^̓�+�&�bO,��1MCG���eg5*A� +�P���3����O���o�e�a2�2�5	��
���G�8�A�����Xύ��;.��h(Y�F��YxIQDB�/:̐j.laȯ�������	-ڭ[����9�ܣ>��Kw���l�F�0��~���t<���������� �4T����7�X�T�##)v� 	��,�e�&N�o�N؏#��R;0�6]�w�S\h�)��e�8�G�`e�k䬻������Cc:1�:� 	A?������v�8�c&�X����d��8�նդ/O}x0r�{@�ϋ,��,���0w>3X�Z�$�cZ!z�.0�&ل�z��Y JOB�@�q�Xa�bC�7����-chM���L�&��T���H���	��
��N;'Wյ��j�m���*s�h��%�B�'�������jI��hc�:|���o�u�27�iO�	1��@�46DȈ�V�NQL�+hkV�o���d4Uhu��'�@L�0gI���Mnd�iؚ>�bnI�S�K���w�`a� re�mL�0/���	
�3<��� p~9��p��u�4L�?3zMS\�I)K�i�U�ӣ ��P�����ϙ"��t����^u�n�Z��c0����Ѽ�)�j�WoÀ
����J
&//.�48��^u�[�Z�gԊ�oT�8����`Ycz(����G�0윉T��.���*��}�����#�����8=b�)�$�u��..�LGh�2�&Q�goAC�oģjB��c�j8�VT7��&�X�[C��z���!%!����"2��'�(:(V�t%����GWj�n�u�1��Y���5��9/8}��,��+��^8�G�֗��D̜�� -vI����[6�ͦG���I�u��R6��z@�|�TFb�'��ɸ�!S�Ζ�n_e�R���g���j��l�1:��ϟ���#�$֠P��I���x���uz ;�h�S�O���^�AfS@	����ˡ*�9�G0R%,)0@"ǩ�S��V�j��e88���'{�Be8�0�S!��n&��
,�;��x���z�2�%��6LB�#=����W�>�r7�A}8�W�(Þ\?����f�m�Ɠ���ܠ���V�.s��7�ś�Mb�K{����ΦpC\�i��5s���y�CT2���1K�B*<��p�u���g��ݐA�t��Bu7�>���;FY� �2�v�)�1�9���Zt׊���X� ��b����T��0�w[�dZ����*y}_�����S���I��a��;f��M��ZgG"��q�4��Bnk ]�g�ۀ�#i��gв�����gmE&���&͠�c�[OlFP����ɳ�y5~� D�ք,[݇�RrP/�������Pͱ]�X��3��X�t*ړ���@�m(N�k�u�|zD)9�)��_H�-��r���)�,!&C�n�!	�}�Ϫ�0�J�<�M�_8p88˷n���e! ��_ZN92�A���Zuz�~������y��=~)�pȭ�����{�p�y�|��W]�C���{�ܹ�c�Z� v�����|������~ʲmD<��bn�%sI����^��&�R��sG!�"�Dd%c�"9��v�s�l��	��0d3k=�g���D/���Qũ�Hg���Uj[GUi�?��ҙz������fݻwv���9��݄����I¤,����l1��q/����Г>�x�"c�Œ%�~�z����YB��\����Zܬ7=͎5Wt2V�m�_j�P�M)�V"R��������$�h~��v$�P48���Su�t����u���4�\�"��"��;��=���>5�fPJ$�U��:N�n�ܼ&�r�ݍ�Ѹ1��3kl�$�lv[-o��,��j���q=,�I��8v��~�r�i���v�	���:�W�
�ܢ�uvVrP��_/�pT���Z�j<��&3H�<��$�?;C�������������,&��)��ڻp�\ΗK��>	h"��ҋ�S�,�l�D��qq�0����y3��fUZ��.nn:��ԸP7mO���-�fGg�ٽy�*� ۬�)��X���� ܶ �NP¿VN�mpH���>�;�Ͳ���<�����F�Dfh�Wo^��g�V��\,�V����s��\�����횔����%\��+r�j�1yH���]^���Lꆚ����S8pƥ���6�WX�M���. *b�v�5��G�~��_A�c�2u�٭��|���~��_���qd���������;�ޢ�a�����������r��}tr�X�����f����z��9H�p�^Q�C�e4��	�
?i4?>�����_��'?y���y"p�Y�x���E���u��Q�2�0�N6��%�W���x\o��/�u�у[�y^f����Q�������jM�xSg6K�Ra*��|��Ն�@I�k�����g�gޔ$ii��&��X4�t���=�OU��㼜�������/�� �n�a
W�b�S?v $'�s1�8ٸj���.�z�}��~��Oݬ�:���?�($��0Ć.h�R��}�)�������pfC�����,�DI�U762����fO�%}��� ��^h�Mj	���P�vyG�欮.�lvʸm6+8˝�����<��i�ٲ�{����'�G%��������`�Ǚ9�4�6	#5:_-N5����Ï_��CUl����Q}y��c�T��r岧]h�`FY �����f�6[�gx��W_����4Ʃm�E�f!�!6�+w��73���%��9]�(W��%���G>�n���jV\�,����Raf��+c��hR�zO��S$��2�Y�8%h��/��c!爹�)����M��.W?|�-,V����h����Z(��&n���I��wE.�m�`�/���X�A",`Sy���zJ�<tq��)�a_Yo��C��b>!�ۯ="��Y
}�2���/w�<U���+��������o��j���rs�Z���C2�3ʘ��u4�ͦe����lஂL��^�6O&~��0SyP�h�<��� �S�`���<�߃`��L��\RA�r����QSOVxvj�r
����8�?
��(�VG�V9�q��ۈ����4 40���s��p���!���$i]�P�;��]����,��#�۰Z��$��j��	C�s�O
u��ј�q34�Ч^�ŀ���mE��IRn?�9�ߥ�L�CK����K�~���i�TZ���߃J���ŵM�$����[��B%�!yyk[���x�9(Ku�Q��FN���@?��2�����p ����Z�����]8�7�{שN�9��}�__��]^,�ɤ0��nە��vݿ�6�����l 9�vhK�ml�D���k��[�f�2�Y�xgmop���}QhP�@�ܤ1[[�, )��Y c�}RL��>-�X*�5���e��j�UB!��U��/�-~!f^�qh��>�4Կ�������秝�^J1ܹsGe+]�&�8��p kW��`:MCU ���0�NSTV1<�;oz�'�;#�� U�k�~[�z�Ӂ..w�XqqZu�$��	����{���\�h��2Q���vܮ���U�<��W�("bO$H85S_^�)S���J�r���Y�K��&�qM���5���z�ꭷ�:=����&��{��r>^?��b�$�_��DWi��Z��v���p+:I��LD#v����+��4���ӓ���G����_������ӴÈ)I�}g�QP�N��B5x�}����d�"HT�`+
#}�7�D	V��>����/..\hx��q3�sV��P:�8a��:����4�BDsC�i�u��`��r�1+��Z-oq���-ȃi��!������%$��H�����,m^+��n>���D�"�������T{y��8$M�*�3�M��ɒ'������_怓gON$f�9>��@�j�1J>^]]ݿ_h��X�{kn��x�TX-�����S��hA�2Y�;�~��R��Y�, ~i=ˉ2מ�$���l�X[aCQA[�����k	b���D��&~8�U�,_0���ҴM��s~�g�-Щ���!j���v��a�����%P�̅@�|BK&��I�c�k�c���؇!��Xv7DRcF�Fm)<�"��伵��8�=]��-�S�B�6$.f��)�����)��њGć��h��P;��l�̏�����NN<x���O���͠�rx��e��i��`�b?<y��?\]�u}�ɤ�b��Ί�f�
?�RbE��ry�^op���'��m�h?�v�^�na\�u�$��{ǆzcY���,hu� �ʥ
��o�Մ:=I9�����?ω8[	��s�Sމe"�M����qϟ?�Q����G��*��y����w�����.�Ϟ=�,����>`�_��`�Jw�싫+�Xw2��BP&7�K��i ��e?�9����W���Z�?wm/Ͷ~��	����,O}ݷ�gp�_|����)�X��,��+`5ת��{?���b�Au�Em._bS)���駟"��Q#�|�шՈ���_���O>�cB�DأfL~iN���~��O�O�g�ӌ�<��T�)��Z�aH��`X�i!X'q	j��4�I$�AJ���,�t>L���8��$��z��_�P�����8��D�5p��k����#���3&ݖ�Z������ԍ"&�C+[L�J	���Z�hg�*x���{��%��&?��WBB饽�c/�[*��J���ӊ�B��<����F�7��˰YX��Ϟ`)��L�J�򵼂������{��1�����-��r����dp�-a�7�+I�]9���"�é��.�x�-��a�3 �(�����`��HJu��I9,�taP�,b(�Tc��������OY�Ȑ����Q�ΜA��vP��1�)���^^V꓀��BB�>n:>�q1*�ow�U��QF���k;�􊬌I�xF�0��F;u�~B^����|���@B�*�
���O�Y�����G %%�?��?�j^�z�� ��ҸD�����ïP+��.`'c�VU�q�Xpms�\���|b�^�;�Et`"�'�����n���IΎ�T���3t���y���#x4"O+��ݹŭ	Q���C�!��P���斬��CH��dn)N?]$�5}��PMw��2�����d���^w	oE�n*��%�פ]g���	:���x��(�k�i�O����1hRp繢G%&$�Q�i	����4�G���m��lnW75��G|�@�Kb�h��٨(}'�A7���%<3�>����'�z��2bU��Z�ð����n/7HB/�
���CC�)��m���]i��x�}�o�]m���F 3����V_	1�,�;~u2$�8�lf��.,�?��L�2f!a:�r`"/1����:�9i2�R�,�	��G�tas�_o�>g�i֧�!�p��ݶo���rG����,�]�n)e�[;��Y��@�=�q��+�ʇvp|ۦM�P����F��Y�����IƗ�"&F��Bk���v�6a�.�N�K�S�펰6��L���˛W~��ʳ�����R�1������<�rUy��EV�+���־Y��:]hW��cДih������q�����FSb{?azJ�d3 ���P3�]����:�\ҹ�f�;=��vCSm��j�����a9heV	5r�\�8E"ڀ6�"vaLjXW|}P"���r��,��+��-&Ѭ������ė�L��3e��@�X/Zh�f&~ԩL���X��-���(B��	�ⶁ̑����!���Mo�[�̘?�o�\���X�d�Y����}�Yu(G���mt�:��N=�A]ɮ�כ-��d:5��l[u�֋ն�]ݳ=�(�G\��|k��1�F�h�|����7�=�>�Dװ�d�J}�Gh��������h���`��uSwnT`�'����� ��G�Ma����4��W��N�ƥ��ɦ�-NK�,����,G0X~�G�
��m��JEu�ůl�/�7\֪���5v��d�p��nF1��V����|~�pՂ��y;�,61���"7y#k��6:��J�X���N�#	�@�8l��zn���^�^m6-a{_�#m���z����ҹC�|#\P]Q:Pr}�H�R_�O��M��b�f�J�,�o3�.�cIQ2e��|���5TJIڄ��D.�6�(���t�Z���o��׿�5\ g7�j�B*ɑ��6�%F.ӈ�$�\=�D�oX']t��IU��s�,Y�\GJ喒|��+��׫D���n
M�i}���qa:����mk�eAw��`����b�t��t}���[(�Y�o�*��E�fORL����&S�9O��BQS�Й�b��|h9:7�z�ȑp�Zs3�K�l�1�v�͞Mq�]�$���͊2`���zN�c��___��@�D\�����NS��򑍠.�/n���jg��B
υ"��j�W��ra.��'��7z���9ަaj�S��Y�n�y�9o|�x�2�Z�S����gg�w5U�*��(Za���{�+k>}�(���O�hs����h1�3pD�g��vE�!����Rp˪�ƣV0��-6�����U�7:���z�80������S}�C�=>4�:&��L!��)�o_�ڈso:�L�XܛC9��|y��-ˠM���s�0�
e�m����t2���'���z��¡>=em�������'�ȣ���xF������;�',��1��b�����������u�\���y�7P`1��ce����3-�������\�G'��'�1�r�gܿ|�z�^���G��{�ȹ�J핁�2�n�'O�`�qK0�nl:��v�1�wva"G�3N���wGq/V��}�#w����͢��pة�v��}��-W_}��o~���KhBN2IG6��|]�ʳSN���/� �p�ղq�6Վ���t����T�S�/��_��*Pmw�-L�=/�ۿN�0�>���65�ga>VBr�v�v�����,)�m;ʊ���m��m�n��WW���R�ڬ޽��Ç��6�������Њ7o�j>��3,�U�n�-�Cy�>L���.�7��s����ϟ}���?�P)[$��1ꍋ�XU<�"&��F��>{����w�r�x��͋g���2���l���v�����ח�ϟm��*��F�d��@Onu/����ӆ�]��;==����_���
D�e>��UC;4�fK�a�\m�4�f�͚���;Dg�]T�} �p(���[QmX�G6�O.�Mo[*"БL�C���a�lfw��)i���;�s|<�	�{�T�L���ﾃo���nv�Cld���G$f��*2�Y�Q���(���`�*1��ÐR� ��
���˗XRl���ܦ����"��#	8�T��fuBmG�vӦB�6z���'��pNf1a0�k�^<~�[��?|�=脿�˿�%a�Kβ�_��O?�����y8I[��5=��S���^)/p���UA�ʟ��+�E��j<����n�u���W�?.)��GGt����B���x�^��l�]W�֣Ѳ���*dc�7b�4�͒9nU�L��=;����I8m�`�"�ZGPz��r�Z���ƛ�vq}��f��uuS�X|�PO$��ڹtۙ-�r��UE7�m��ҍ�^�ٴ�{�ҝ�	����c½�g�s��q9�҉vvT�,�lL=$�����ew)
-ϒ�G�uE�ZD/�IyLp��߅�OLT!ˮ��iʸ=C����G��7�!�Se�^�X|Nb1���7��Hz���}㡎�D<F�] ���^�Eu\t������4�t�!�a^j�_C����Z�{<�� c���w>\�u�Ĩ!2�����6#b��Yʷ+Z���y�Ei�ݶJ��p�V���.
�`GK�{�KL��.n�L~(�B��ꛦs�=��f �j��1� �~��wrr<��Z5��B=L�F��'ҏ���1�^��`�C�\,R�٫gQ�d��	de>��r��(n��$hT����fe���8B6�:v�8_{��.�����8��%ѾF�kϣ8��Ł]���<Pr#�n��Ec��6�X����t��oM�`9�S޻��e�	��PK�En��5�%�>�"}p��C����p�[�#� 6d_j8>є�)������jX作Č�N���77��ϫ>b���߆Q�3y� -2�Q_���؜{?ҝZ�;h:jW�Q;��a��@��`ۊ�w�V�)����r2�$6A�tD����),�(PMi�ɳ�-N=�Di)Ί�:���ժ&�2"j�]ݲ��~a�ĸPU���R�])D�K�\7�rp�w6�A�j%�f)S��m9��^��Pi֞9��Ά�о�B�:��
�{�P�r�R�G����>���Z4�z����ؕ	��󥁺%��A��F��n��6�B�E�n��P����^�6xWR�)F�
ŢZb��R�C���} y�O���d)@�[�L�x�B>+RB|
��p��X�W�J��ǂ_%�j�=����7��r�c��z͌�XP�ꖮ���}"vըڸ<���D92S#�lUGU��~N�^�o04�{5X��9����WC�3�,��?��Gx����_���'�'�{�0K�G�<�F6�p���h�
\��7�$��g��h�||�x,���?�Ih��4I<}�a) ���u���jI��:��T3�Z&��s5�����ݩ��v�76<��m���O�$R��=��mG#�����B��$~L�X�+���Er��l*���i�=�$~�������8�D��8��o����f+���5�>1S�̜�_l�[���jC5�$g��]$Z�$���џo�(�C� nА�i��h%��� H��h�yz�~޾}.�a{�GV^\�XpG&з��*a�8�%��� ��Ud�eIi�m9���<UBZ���a:vn]ɣ�nCX�I�^�V��N�;/y&��I���h�mg��Z
�Vr[�B��{��w����ư�#�t�6e��@vnVó)����#vIW8@��,�,�]��~��11��l�����o��o?�����w����Ś��~Ɯ�; �7�N�Rf�hR�z,	�%-$�&�,�;��K�Km��I�z��U�2�����ZX0�OEC.V�S������D���5b�Z�+Hf�O>�K���R 姨�-gڛG����M��u,�4:��Ç�~��93�5	�X<�}3�^�Ȯň ���<�1dV2�~��ĘpU�h(�|��ᖓ��oHo0���>񒋙���re�Dș\��[��*-k�#܋7�o�uc�_
��w �?��V�S�]��N9u�G�&��?
�"�j��	G	�+9����`�,����Y�;�S�mR��Rʵ����=Y���sCt��%�9w�����HQ�P�����թ(�Wf� x��tQ󻃴`�G��H�� 9a(��S
]h�i������sA��M��ۢ�v�ŋ�����/5��Jn���w���@r x��k�p�?�s&���!����t'PuV�Iҋ<�������_|��ET=���	�e��}��6�F�ni�2q���16�O��6r~���27���{�=jž3�!��a~��_��9K_��v��|6M`����$u1,��B�7	����Y��d���GD���$@Fb:H�ܘ+����e��g�~�]jm�����\�z����j�3��ڪt+�5����6va4b�u6g���O�9�� w�,��-�m�x_�Y�v1�ՁU���p�B����ߣ�����?�JR_48_�d���(��!#R�I�|r͂LS[A|M^�ݬ��h�k�A��������k�zsĸ�'�����Mۇ�O���03McZk�в���{�F�K��h�}���
���,3��ą����]�e��c�e泴 �Z;�}�y� �+�Ao�=}���6��z�X{Fj[��٧gB;����A4�{���.A��8�F+P:!y�h��s��/I� �蒔����.��Y��YU�α>�8����aTf�Ј����5m��W��Gh�a�;w�����㗯ވ/��+��`C�fp=�>y�����ӏ�c��%���V�GC$!��\��GC�������e����G'
*���뿴w����=G6p Ktr2�ݤT�G��Q���v���Tl+�O���~���<�����oə�Ja,+�٦ g1/لy2�:C�s���]t�U)�H�ΆP�ր�s"UkCN�up
]C�H9�i��e�N+�"Ljl6�e���L�4R�����Ql�������wV�]�6Sl�/��
��?>;��Sf����jkI-&I��qg��j�o
��"�폢�n����Ar#Ej�T�;a��rK>��񛰦rI��&
|d[WXuV ����)��XI�r!�ŭ��#�*B�.B����!�	QĻ�ģ;Ԉ��ؾ����Z%7��t`o,N������ߓկ�|���Q"�&������=B�p�W��m�?���o���͎���Ģ6��j����쓓��ޣ�u4��P,Hn�D_O��%]څ̚��}S��^C2�ͥ3gp��(]��;�	��e�XX����,֋ʞz�3����s�9u�u��{'Ϻ5��
v�����Ne	C���������H�KH�L�ѡ��H����&�4ь�o6�ʲqC�륰�P���y��e}������F��e�G|Qjɫ�@�m����_Wj�%oae;���3�����{x���auW�a�3h����;�V#�7����oE
��5;�e�}�:���ml=6�/5��V�^��e�]��ėi�EiX�ê�M�Gl6t{���_!-��w�y��_
�mh�����4C�q_й�r����V�x1��
����6�a8U����)��B��0�l��Y����n��Og1l�*�*����4�\}I��`Y���@ˍO(��;>>]^�>g��r�=��.�պ�{`�H�3���^�L7Aӭ������0�\A~��@٥��~�T�w+�e��պq9K]QW&i9�Nƌ�F.��~������)"�|M�8X�r�p��6;*��I�!ti��y���p!lf��'T��>�j���,ۃ=�
�'�V��)
�Ҟa3Bvg	��U>%�9��^:�;���b6#E��dv<��B�2��x$�1���nh�n���hkK���&o:G��e�3�����t��D�P��eL�En{1����o��	C`��_�N�=9�|a����me5Ȯ��1C��l��Ũ,�}�ûwo���n�1�Q�$ӑ<�@�)�-�Cgӷ��<B�����G�u{�M��b�c}������R5��þ������'�|���OL+���Ew�o+c��]�9)%�'��.��F&�f���W��=MBi`��@P9y�򥂗X���S!��G�����__�v`�sM�Һ�i������z��m�[o
R�qn�~ Q�����*�`���X���&�ni��>}���{`NO�,Å�G���w�K�s�N<zI(ɦ��/���<4T�a�r��`�w�wKhDj��3����?l�׫7W�Ϗ�*�$]�������6z�ӷ���;�__��)�F��N�blh,��S}yq�n����z���8���zi�;?3D&;�q���xn:��4FF#A�0_B�'�h�A��1;�c�;1��:��q�)�⣏>�������b�q5�W}��+�8��A��nv���3n�Պ����6�p±�l$�����~���#c�9��|�n~r|q�&o�2�E9��3l��Y�Z����cM���D���&(��L	�b�$f1�%&�Ê���/6�1������t;��-o�z!1�5<b/x_��/�W����T��I>�>y�Td�)��i�B8�UI�L����Bُ��f.��ID�����
���<y�V�!C �)m~�Y
i�&�z^��Ù��r)e��G����^�����jS��_Ckv��9==������������;��-�������ŋ�B)RoW,�Vm��9C��̧h�Jq�;�:�y})]g���,�`��&1�$62�QZ�ϕc��F�(�Т�3���Q���1����ZrC�sM�F%�'5W�WuW��ed1�Ӝ��U	VW
</x/���Q�O���M�^�W�����!*d<b,����&0�Ke��nV�r�Hu�U۵���x��oi�m1:��s�����!�)�.&�(��
�b��ad>���V��s�tHPS*���ZH1x�Q`�VJ�@�`��8G@�"�?b�O��4v�TRk�4O� %1f��@���[�6|��ÙO�n�@�E!;����<���b-z�;�����Q̧�ZPrƱ(���b'l����F=o|j�B��iGY.�B� �
��h���[�ڳ��/n8��� l&G�G��Gɧ���P<8�:��}
&�K�a^��|){޼���	]��z����c��з0D��2�Va��Ҽq��o5,����lR�{��}��c0��8��8qm>����d2��hm�%�"��Y*Z��9��u�	�01Pm���F�(O�B�SU5ө���:@�&56u6}Hz3$�K�5U)A����u�cƼd:ͅ'�+	�Q����y�	��y�7�K�alw��t���^�+�^m&��h�$×�
�BPZ����=;��Y�a,R_<���|��?���ￋ݇��{rBz8�4d����b�����s�aؓ�����\#�V�K%x��w�rnV�)H���<X^A�%���)��urr����`Oo��
d=����fhqX��`�EB���y <�	N�Xg�	��'&~�lv���4iΦ��N��E�&���3�����؞L+�3~��l��g �ړ��Ԉ�.�N9���s|60�|��G���'����<g�I,�ǃk㨢��YZ������S@H�X6+�_s���fi�H䌇�Gĥ�=,��a�Y+t4�i��l��r��M�Ӭy��Љ��|���HD�%��mcLa���*�'jD����E�D���<p��cp)���t�� :˾I����l���CksKna5T���H�:c9��sI�g$�
kH���]]Y~��j�����R':|�gEw1�a2P���R������߷�z�g?�ξF���גU��_�$��3�P��]��"�M�kbd���5��f��A8��$ �8 Ԅ���KmL�S�2.ź�HSJ=7���䯩o����ҋ���:?XY����V�xs"�����q�֜;�~�������k�o����9IgQ�{R��ͪ�}��)��&�8��Ҭ�싋���un����dn=��%B�qkk��G���H�>f�u�H,�������Gѥnσ�o ȷ5�ᘘG����	Fp,I���lih3��2'8�����[)Ir^Z�<ݳGi�&�9�������9i���N��<}����i +&�(��T�v3��.d�[�T�BG/�0kX5����YvO�.���tH&�����[P�)����l����kd�U`�G�mԳ���V�]��X���0<�;�\Ϻ���Ij��X��܊m���F0=�A���R��u6��<=9��/~��`Wڔx���0�ո�&1�Մ�>����e� N}���S^>*]��k�ƈ�d�[�1�����7����i;?s�g�b�1fO�J�����pa����{�j�q�f����3I�D�9j�44�]�hHN���JJ�yI��8�3j���i��,�i�m[�`��~��ɭ[��EZm��v��&jX8?�6��XC��o���g��c�g�
�9�¨M�l��J��Q�a)���g��lܣG��٧�.:~1��9�OrǦu�:H�7�Ý���<Υ->��1=�[�۟���eC�o�s<�Y�gE�Ӕ�gϞٝ�~�i�y,#��+�f&&��<�;2۷1B��Μ~Z�(%%�f�)�E����v�Н������f�T�~[H,�Ç��y7�O����a-����R�. ��Ķ���t�5߄y{�ܤT7 ��/�2�C^�f�>�j�J�]��l;��x���L�#�4T�ED���Zv�Z�O���H��_�z��a;�"�'�a�9%��B��(����ӎ�{�µ�;Y1}�,��f�-�k��Ƕ��=@�.Eu�O�Dt��P'���Ūy蚴ny�
H�j2L{J��A�^�zeϳ!�)���R�ڀ0�����hX2��i�� Q������W˯Ȼ=*>���05��
����s6ļz�;�,WJ���v�i�ʡ+nH 	�&�	���[�������,J�?*��;��Ӿ���O��7q�'��4�v?�B�����'B��M=��z�lG�� E���CB�Պ�Te16�(�Ik����$�˲t��^sL_M�]���g��tbJ�-�ó/�u��入)�O�7�c�6����jәLF�buCb��0�f)!��z�)GYk���A�.U�ͩ�_�X��%)�_ªlfM�T++�s��qqy��#ڌs�M��Xm�O�"P�֭8�F��pGGc����[�gXW�dh�k��$�M71�w�����oÙ]n�꫎t���ۼԈZ�t��ڮ��KG�b�-6�Ǖc��J�)�v��Gy�����=y�P�=}�����&���m�B�٣	�'WRF�6��-��fg���Jf6�q��%98jx�$��s��kH��C���ʡ��%˶*�D��x����C��isS�vk�ca���_�0�]s0�ȅ���ג3AM�# �U�������{�q��ٳ��}��C�X1��%��|~���rW՛���զka���c�R�9�.�;<iɜ;�����9����6�`3�nt�MuHB�q8H�ė�C�Na{���j�XI�A��۸�ѥ��1�qG���:8s�~r�sۙW��U���u�2��\��<��ӱ�.��V��8��n2e���'�3�����������_�L�'�f�Q�v[I�j#Wf{�I��Ϙ'jV¢~R�?@����	v'I6lɢ�/��6F��)�>QR�"s<5Cꮗ7Ao�8��qZ-\���1ߝLIw�z��S@N�?���Ƚñ�w��|f�R>��b�'�����,]o�ֳfK��f~����w��,S�qC���2Òcăo.�_���Z����1�	�pU���>W�640���xn֢��8�!;���A�ҫmf�\��x��8��޼y	#%�+�@t(;׆�n�r�쪶r��캂5.�:96�uMED��`0 �Z��/�F�ߖ�<n�.r����56T֐�s��(���*O*�kn+���S�`�N��߿�[5t���Y�kJ��ЦLl��9Po�x6��ܚ��w��=5׊��Pժ[����q�yu�_ɺ�F���Bx�"=z3}���Y}�mi���~�xu��YM��p�I]�u��Ƴ�P>(���f���
��T"�>If�y��A�RY층R�A$�MW/G��3�*���ѱ��[D
�s�ǜ��rCM?S���k{Q�3R��
�,�OU٭�S��x�����~��OɍEj6�3�ؚA�j��7_=�Z,��`���$bݦn�u�tX�%-��,L����n��t&����tn��N���/���tX�۷�1��o��Q���(��q�P�Վ�a҆����Z1�a�০����B&*����x������ٱbKZ%NBK��2��|�)�l�X?&�c�]�G�ͺn����1�i}�_�n4��.G��¹I����U���S�l�᮵���[���DJ��n��ޮWM����Y��D�a*�	�il^��_/n�ǳ�x
�x>�(�l����ͦ�|�NFX���U}9-J7��Z�$~����E^��sݩ��!'�����ٔ�}}b(>|4-���	Y���� ��?}���]�A2�̓��^�Ũ��J�f�t�˪mm�O/���k+�"5EX몱�ΦK�Oр5烱��䄨��B�z��lW�є��������eK���g�Lm&���y:.���y��ە���l�꽷N{׭��$�7��A����QHձ�'%�	8,KQ����y���VQn��x�iG"Sv�(0ȝ<�N�n��O��nu��C6�=[������h��Pɏ��J-Y�&Qq|Ʋy6�����]�\[[.֫5|�MUf��n�}G��\l�z�Yq��ϟ	ϋ#+�˅*��s.]�Gb
ζ�aN����p-	��@�*a6�O�}2gFoc��|ʔܤ'�r�tK��6!$�Y�θ۳qb��4ɳ�ب��0J��w%���j2>�)cϲq����?z��ɝ[�G3s��
B�'˳طUk��<!�<�I�j�K𹛪a҂Dڃ�|KPF���އV�@|�ێ��۫���oVI��it���!�A�+��AZZ���Y>x.'b򽖰t�|M�U]�*����F�#���s8:��	o���í��
���H�Q�!��	�f 8�ǟ��[����|d��\�m�)>aT��ǖq��e�4��d�ԛ��E���fU���$�~����o�Z8Ѐ��&AŶ4�tS}��}Y^���yY�R�r�6ҡ�jL�qx�X���������#ۺFE�w5ge�C�Y���՛װ�E���]�V+DUu:�X��o��?T��(iӛ�9*��ɏY1h�lڤJG��Z��;����U�	l�rz��x���[W��w����I��N��e{vÀ>֎�C�g�ۧ��͎v�nAYْ�%7�EiIv*\�3���)�(��.ٸ���x��յ�K��3�2êL��N��z���a+r�i8��`���u�4҈�Vx�,-w�F�E�P�˛���x��]�8w��+�q84(�bkߐ�G�p$�`O�1aP��/��y8�p�,��"���s��`�/��Xfˋ��M�a<y���q�gSh�Tk>7-��3
���3˪����v�<�B��]Y?�i�/�&�t.�O������&�����}󽊅��,KC��2�̡���F�]�дn޼|�p��R���:��5���Y�GS�Q��e��\��$"錛AI�R#�R� < k��ZN�=�T0-�������Ͽٮ8"��a��Y�ggshr�͌��q�iu,�ɱemG�
C/�O�c��F�����2s����ż��Y���������}���(���\~��߆��(�Q:O���x$�xvvΪdf��V��U��F��a�R��#{;]�n:;
�yh'��@��ΎbBمNX�9�j��R�1���#��j��*16�j��cs�ֻ�[�� {����jO��Ývmқ�''���:��֝��y*!F�%',T͆��F��޽svy9@3�G���V�����`'�vۑ@EZ8�}:���&�q3�rզ��\��kx�p8i�kk�����,��m����C� 7���y �զ�b��L0�!����љ�l���o�5�C�JX7˗�~���{qg�?~���:����+�+��y��]�db0[y�����.�[�z÷����j�ѭ�K1��/v�ކ��x�B������"��~�����O*�� f���<0zJ+�6JN�":O���R����f��6���-gZ���Hx�� %E��N*."0ǰ��-��C�(������[�}��� sI$o�T��W"YO�,q@��JA��M�QZ��_"����M  ��IDATŷ(�K��0�TA�j̔��Oa{���gi�ƣ,LP
gީ�0�u��z6����~N��{���!�&�I���m�����0yP�a<۾�H�d����9=*�+!��;��"eC����o߾���믱�,6$�GL���.�n�@
�ԤY,��G�ݘ�Q��)x@��e��(���줞����v:>w0�J��6��Z��ǳ� �t�55	\�=���<}��ݮoݺ�O���mlѸ7�N����<F1�"w�J�����#>��5�q��i��;ܠ~��C���bQ�-�����(m�f����b��=?���CϣVFw��P�Jk�:s�R�v ��C*���Q\_A��Q/��~z4����ȹ q��Y!J�rQ��0
S#�r����&h)��&v9���������c묯k#��bk�*E��ܾ}�b ��y]!���Xݑ��2��3�	��-�<�k#�����Z߼�8���E(�@�L�"x��հGb���;��V�*�m��#܌B+��$-��Ձ�ͦ��)���[o��r��U1ώ���,����4}n�@"$�}.z�Q�x4�p"��b���XR��t7��UB��X"@�
K���%����@9%�ZV�t\�`<B_�Ѭ�e��Ch�ܪ]?|����޺�J����<�IK�#X�q�զ="[EึC��E��Qp��s4{ί��&:�z����(Tg�5�!��㘧�c-!�=���Fڗ�ua0���.y��=	���a<*-1�Z�*Ă��c6�`+sY�H�k$��5s���G�@C���h����ִ�Y��<�D~�,�2A�r�]5E�{�_]ZÈ�&0�G�z.�S���������O���X$X��w��0)07fe��#�4�T��b�����;�d!fq'b�W*<��� �� �����j;�m��+.�
���8�e÷4����yY��t�E������/�7(%-��v�y��&K%[�����\Ƒ��M������v�t��81Ѓڈw3s�<�x�h�{���Ӻ�a`�oGGb\�l:��垺��+[�=��.���k�>߬�͵Gʋ���#i!�]����r�ѣ�q]��1�ێ����S$�M w�"���k�bN�ŋW_}��r�����9�Z� ���I���":iaԃPf7<x ����̮�Tf=�#�J����fa�B���ZR��d*�pC�)�)�N,��@�>����#��(�m�lՂ��rt^Ľ%�G ��ĩ�� �'NZHn��͠�Z2�߹A���Y�Ϲ5�ڠ�`��������.��D�*v��"V�Jg�6�K��U���,����/���R���2�k9c�~���9�x������̒'O��X��Fn{4婄֒)�)�ÅV������[m<��D��d�ʇ��m�[ 9Bvg>��BB����қx�vٴ_8���6��9Y��M���H�:��K��*�>EeG�g�%<v�Y�/F3����`��B�dQS�G �L�={eh)�S���-���$�q��
 ��81b,��*E�J�<L��4�1ď�� =?�����ߩ���y���?��?}��g�m���o���c=6�R�����H��� Ta2Frз�$i@����O��n�g��E�4P�_�4`	���H���OdZ��I��onp ؜[�xj��Y���u)�FcT^o�'�A!X+�[9���tvBU�󟿋����ߧJ�yL�<K�R��1�F�˕�!�2�	�{Im�"����-�"��bq/�$$�oQ�Lw�Y�J�7E�������؄�4������<�.�IZ���mǘ�G}h��}?�Y�4��]��7U�ejĦ+�e��>���@@�#����p�_G�����3�q�0�����ˋ7�|9���]?bY�}�~�)��lJ��Z��N��ԧf�Xt�3��s~p�&B�.;�م�<�d*�\,7/_]��P���E��ŷ?���d���r�*F��q?�Jq�0�X��\[L�k�Q���y��2<�Qq݌��!�t�*�Q+,�v�x��:�Ӈ/�M��Ãk�[R%������h|���Z�|�
���ྑ?�rz��O�O5^ق���yh���C�Y��-w,�0�6��ES7����r��m.��^��Ǖ97PCf"M�./�L,䋔����X�U����.lWW�q�pY���g�dn��ejڲ�:d7:����7T�75����e5X�d[��6�u%��jq��#X6�2Zȓx�
���i�&��5�����{M�.`�*Z)+9�w�E4��w�b!3�̽�C7���bH�����D� �ۏ7J����k���{p;��
Q��x�r�@��>f�f0T�֙mI�l���5�W�����E<PNDi���6ÆoImD@��&�6�Y���>��)QGG'�	eb��a�1�Y,1Z����&u�K��W�o^_e�o��\}��G�y���닥:���ղ�C�,�6��|���Q�@��Nq��@$��VЭ�H�֔p��D� �(
UND�9����!�>���Ӗt�,�)���
��3�� {�������"0�<�6Do?t�H�NN�<�/����� P{�ӡ@%ܧ�o�I�5c�T��!���a��Ղi��F��t��@�����-��]�dḧ}i�!��Y'o6�Z��j��k�ڝauŋg����&� �vW5��Xv�A�I
�i�Į���4�v��X������i��Z'o�6���ۧ��%׾rFi���d��X�:#��c�����ĭ�
ʹP��3Iy�G*�C="	���z"(�o���Z�s�o���y����q>��v��.8❍J�ΗI2�
��+���{[�vS�%�����01:d��Kw�޽�9s�����7��D�)�\Y�*P��穈��.�$[�}3ϟ?��ٕ�h@d(����'�)l~d��L@��2������/�aT��9s��6j��:��ĭ8+���\Y̼�U\5�@q*w�H�6�RiMհ��K4>�&�q��l=m� %�癊p۪ڤ�/�"���t:28��1T�B��6�s�']r������jK�4�U�G��62H妹��M,W(����e���A˱}$�IO��` H�-�lg3��b#�<l�`�������69	�y+*��g2y��q��Tw���Vj`�$���Ix�St��M<�i斫�t6V��x�����j���\��;�4�`}�R&���fD�Q�6W^q�9���o�K���x	�K`�V�O?��[0&��$_��%��h�+y!�9|�ݻw��-�{��Bp��AW��X�&2J����GêB#j�5�q`]^_�[fG'�޸*o������Ѵ6+�`�����5�bEI�L�Ç�}�]�Q4�V���<�l��{f�e���sé��v!T� �g�w%��=�V���-��4�8�0����F��{o?�B;AZ./�U�����e{��2��D��'͹��'c���?�)1���(/���
5u�f����z��4m6�����#pKt	�3�fy�j�:c����!�j� h���s�pl8��s4sw�<����� �m[!�Z͎��RH��:�ƣ�4͊�Kd.�n�}t�p��Zq���,�@��!K '>RH<�25���?��o'��b]uX�$!����.q���=}jT��w<9�9�3US�bzu2�eZ\kJF�tT�#�|}����Le��p�������߿��ꢧS�\mF�����?nݺ��O~�����!N�c�,����/>�����޵8��DG<hd�������[e�ÒC�Y��X���b���bLe���C_�w���W��V��>ಽSպH�?*;*�y�]_����v�f���ËB���V8p���p�����$+g��tȈ�$�)m���AZ��SBj2kZJu���dv�ν���G�_�-�>�����̐"�b��A^FY�gϞ%ǣL_'��إ{�{���'+��S��m�W�Wأ>� [�+LFc�����x��B�^�qzDdL�~e��S���>�,!a1xtѼ��!
9��4�e�Pi �K���@�/��c����)�YY��R��I���y��kT&���q�MR�n��l�Um�QCZn+2�T�ե-LR��[o����֝k6�uǙ�y3��f��{��u������f�c�����3/X��u~Xk����Y6��H�枌c���Ĭ�g����jo��c��	�eq�0n���4t!-?�iwn�C��J�QqC���@�՚��{s���O�74��K:��ɴoz�M���kLH
��`*���bT����_��i2�쨩&1j�j��F�L�nj�J�#�!P\�	Ǣ��-���)��0V�F��sg�t��:`9p�$����B}����[��x@�X0��1����2OE���$�J��ln��Ϟ���O.~M���td�7i.8� ���� Vѷ:��$��݆�F���g|�R���<NCv��F��5͋����@��rG���bl剢Y�ӆ=������M�G|&�U���L0VMt�e#�)�E-���P�Hy5B���ФQ)�W:O�B��]*|����*k�x)9@T;OOp������Y*�ùK�0�c��|!�_L�E%�d"t�;�n�0�eEvD�d��4�1d��D�y���Q0
�격/.P]�\�ʀ>-叶���w/�1qÝicS�T���H*r"x�����l$��!*�n���m����g�P�9u�=D��aU���� ɟ��EcA1b����<L{�8���\�P�j�ϛ@@�x�OU�L��J��<�,`6)*�n)=�M|��~�z͑���_%��%���K�	����#��R�%Sc#C<ɵ�5B�0�wg�rLAZ�N,=������`>�X�8���hk��@T��AD��ޥ��Ѱ�+�>C���*a����S�Wg��6!4�M�I�mR@њ0�4u1����ba����P����:�|a�L%S:f�^�hkzQ�8K�p�Kߞ&������1�4�6�<�Ңk���w��˗����֌�L�6����r|�rɣ�劂u����n<� Ϛ�=�@��uZ�MT<��_����ͦ�2��5��d��d��q&)�OL>==�s��`,,K�a@�AY�;!?�t�*=�y��	B�4��\���~���!l�����O&pk�G���J����:pI�;#� Kݡ�^��!L������<l��fb�E�:p�N��*�aeFc�Ǆ��}����X=�N���W��1���g�&�8�7B�5%6XIK>3;���C\��u�"��,���B:)B���H���Lծ�M���u��6�Z^G�1ۑ�B@��y|�����)3H��#Ģ�4� �U5�O��9�\<maµ�u$�S�>�CO%6�:�F�w��dcl�ChM��EH!���gQ-�Z���&��|aê�ԧ�F�[�{#�y=����|��|����c.<X~h��eYd�����)&��`p�0"&61Y�F�Z���ܮUƟ+\���� O��lJF�{�!��uf�H�8=��S��
�����X��l��I~������ݦ�s�o��op�q?��#Q܊�����#OE��[����H&u��ZnrM�cc&Y�|���֍&����(��!�6N7�qpDc�9��VKzD#����X\�W�Nca�T<'����kbY�+��p��rod8%z׷"ȱ��������9��co�#Yr]	�[}�=�ʵ���H�-5!�D��|$@_�m ���܍�$Ei �I���3+��Ȍ�׷�=�Yx�8�D�����̮���s��G	�4Δ�6W�ŕ�/�ڒ�"�AYF��tS"�u�R;(��Z�}��/D����W��)�y+��I��Ō���3�"�����w��.fb�K.x�E��r�l��S'��	����G
5��������g&�/u���s��I��-ldGtB�\��l�b��>�a:��X�\�.��Y��w���}��+���I/'iBK�I�ٱ�I�-�(���X��|�J)TD>��w�Dr�������I�S�z�t-y�u�*�����>�<jy���7_�txs��#�����;�n��������o����Ӈ�m�)0͆�G�N���	ihtM<�i�G���nc\'d�^�2�j�NO��џ�"t��RFV�z�$�x�����dy,�j�۔��<���°>u��C;t]_���J�������s���M�9����J[������ZsoL�͗s�"�&&��v�	-����=�=2h��S�y٨4�6��/� t��36_ط��ޗ��|��m�^�u��/�+{�#��9�:S&Q ���V>>zG���Xi����~���0��⑄"Y&&7a�a����55�t�h����yIܴȵu3����-��d��Qg��K�j�B`�ǣ��]J䃬@�9� y�]S���&��c�W�F��޻w���Կ~�
����Fu�rʘn�,�b�s�z�ɴ-�x�&��%a������<�d#��Q`��f7�B1��M���誸�1���!6a*F<�u�1:��L��s�n���c�Q�b�}��]���ӣ+J)yz226���7o�<ǈ6e*�^Ќ유O�ٱU��0��5`��f�i�����^Ϛ�<�dxB`��^C	������N��n�w��J��.�D�2{8���:��<�:�w������sLJ��v�PG2�������Q�F�sW��FuĽ���R���(:kU�s�gE�aO&T�1�5�<����U8u�@K�b���z��NX�
#Jͺ#[�����&�`�����Y=��^�yuz�d�nR.$_,1~zՇ��͔���#%���d��e��D��ׄd>��*�V̜V� �p. �����~�C2L�dU�M�R��d~y�������̤���]E$Ѡ堷$E��9v�!ڴ�pl�Jc>�L6�|�yQpޯȟ2�ر�o��7�Vr�����.))z(-���c�*�-սrs�;H�@H�|zq>�Ӆa�Z6_�<0��X]�!�5!�BW�i.%_P�\��)�O׷�(ꊁ�BG��G�j�,q�rtL����o��'����{��g�d����̬�Xl�P�\����(�w�*�/�Y���[xV�, �h��`izb���6�����4�@ۛ��Uk���ŐPt����U+��-0X�B�%���ቺ�tMB�v���Ղ�߼��=�<Z�p>Ǡ7�R��;���L�T9��A.�X�H"f.�s�1d2C1�������WY�.$ٖ��zO�.���ǹ'��@+Z7���z�Ͻ�HC�J �Hd�1�m�R�a�����z�-���=���!
U����
��#��;.���S�Z����a�A �bi��X�\���M�f�:37�\�vJC����UI�����x7ϙ�%��b4i�g�Ax���zQ5��nZ���sq��EX��Ǳ�UgЂ��s��������VVN��gv��:Wߖ���ʶ¶��t���k	�A>�\(l�"�΄��0cVȗ|NO����|1�4�bNյ�Wn޼9;��^�ш�����	Ԡ���&�L�G��5[���*�0�o�4�V�~"��f9�6i	�9�W�^���_�Cv������2�I�#+�j���R�����T�
 �j��uv�_|��o����I�$'�!��##�GJkB�}�-�������n��Ϟ�G�$qv'Y�1eǋB{��o�ն��n�V>���!�luTM��j��Yyp9���H�)3χ ��B���tk�[�;��Sm6��G/"�����ƒ j �z�,N�M��r1���-�7�v���k���n�<y�d4B�y6�g�;��E�
uP��@�q��c�����R���`pzv�%�4X5�!Z*E
<#J�<h�iL��k�X�t��[��LJ{)�UA�ѳ�J�y l��ic#m�P�|���/�Gۣ={�LQ�rX*X�Tk(�*�ħ��َ�������>{`"}���ϖ��!���֡�Lq�V�n1��Av�p�1&I����)�vcJv4gj?�j� �9Z��Zٍ(�P���SR���Kڙ��T%��DB��h�u�?��3k`k�5���]��a7���ӗ/_q��D��������D�<�I��ǯ�����aG���S��"?�N��͗�sv�u������9R�Y:фDKy6$6�wiA��M]�ӕ)��P'[��^�ɟ����l�-lq�zN������\g])��>i������M':|`%r?�� �I����S�C`0�Ry�XTP�Jw��Y(�]����e7n����>���7�T�Ğ���7^޹��7����ç��M�+&�çϞ��n�٩��W��j�%���^s7zp@��y;f���B�WGGS��#Y�5�����ݭm`H�'���j���)������ށ�"��""W��A�O�%3�WY͇i�g�+�U{����ک͟㼶E���~�j%�]�E`�W mO�MUҀ��W ���	Z��N�ůY�����$ٗ��-���>�\S[[�IMޮ��u�?�
&��H�T�������{��+F�]{��������?���.Ɏ�^����������wك�cw}2��8��
~~����)_^���X�db$?>{�@���񞤇&�����^�|�i�")�y����k{`��fUɀi�b�h�56E��l�Z͗뭭rkkǶ�`���.�	���Vv8HN��� ��9WUm�[�Rsz�`�4pԚ#��n:[�7�1�e��S=���GG����PΜ�Z9�>��4�����V���I�~k 9���`8�Ɛ{ v�y$"Y
�J؎���-T��榪��{��4=z�� ����V�zuL�A�1�z��f]�d^bG��L�,��w熷�|�	�NRDeޢdz���~+"E�F��5����a�3Y�ƾ��w8D�����ss�X�Hm�7]��f 횻���þ���7ڜ���PA����n���������ϟ��_�嵛�v�޼Fzl�$���nhA��%y�-�f]˻L}�ѯ��>�V�\�,�K�ڙOo&XC���ϖ�����P�$p��U��I���->�G�߸~��]�/��8Pp�|��]�a����G��.���Ad�z�kv�t�������S[�3B��t2�=�͖���劮~C�1�*sL)
0�����sTR�{�?;[7��}6#IsN�]��o,	�=�\9�	�5�s�D&*V�>����U}b"َ�ʕ��[��a*��.�#�V|6��/ROc��Q�@�ԇ?3���G�R�-M
��u���wGrRr.撔[i���1���U�*ˏ�Ǟ�|��(���H�;�S}�"��'�
+3:�3��0A�Ue�tɓnU�L�~I�~D�KC��T-ʐ��7�L����m�j�.i4�Ci4���@w9�ZR%�1��A�b#~]���~��6���D����&�ָ��F���1V��J�Y3��p�?x?�S�l&(u��a<5|��y	�jS�ZE-ԇqf0��dr)��4�@�X�`��H�o�_XD��^��!�f��ʫ��`�̞��,��d�m%�.@<���6>{�Z$:C�(6V-���Zg&2Tn��5L70�A�b��0�a�T#��
����hb���]#�n�&�B;����n���o|���&����*k���T���d
�|�� s�Tu�v4ɕ�Gԝ��rTDu���6������j2J�Q�Y�y<�˾����{����ns�Z��0&L�-����W]h0Īvix���%TN�g�O�:����C1j#ˉ��>�"�@�v������GR���k��e��DҨ���How���d���'�D)��{>?� (�)%Y��,L`G�x�`�^�o��{Az(�ʁ��W-YG�@��PQT\r��m ��C�`W8�3�bS���� �����U�8C���l+L�ʫ6��J̏���6t�-�R�{k�~TN�By����u��[6aV���&uo��܇~�IA����~������v��� ~>zq����L��e�UL^=�w����[,jǑ��3���y7?�Ν;�n�rDx}���O���p��i��K��tm�â%�-ә~���6��\��e�d@�ˊ|��>����͘0�����L���X�yΗM��P���"��6a��mG^�xa�HVO[ӑ3[(�_t��9sC��\�e�l2���T�^Q��&���5|�ᰌ�N����&��^��Է��ڢ�mgw�6b4EJ��9F�
8�s��qF���9Ue�Ȑ3Um����Ĕ+lb8dٕ�_gx�����itb�"6 ��o�C�BTlլ� נ-P!Pկ,̦t$���L��A�ph]-�ԲQ�R�m�
v$yX^�vU�ɺ�<檹>����O�]
#i�x4�l��пx�����P�'�,���,��T+zY�Fh��ւG�a�pD(4���9I�����>�JIF�`IR�i�����׃8r<#���)�j7|R����i}{!�L�l��:,ZW�q�f�uݠt��~��D�%�C�d9�Z�)�E-�}R�Z��O�q�R����v���]Ά���8�3���S�I�N�o�������:d�&hޢ�ert[n�]�>_h��K&M�H�N0j��ډh};��+��/o;;���$t���8�m�ޒ@��P��@�~���r�c�o���ݻK">>��M;�/�L�������<~���/�wXI���$BK��iˮ_���6��ٹX_e�y�iB��8��e�������ʭ�-K�ӂ��Wv��b���#	�祗I{զ��Z��5E�I哮�U���_�$���W���ђ�c #�Щh���̠D��Z#s��c;���7n܈.D�Y���7����~�����?����ۿ�����w�t��<j��ѥ>&�f���^D4m8(�H%*�\�v��Z�Ȓ�b$g�>`�@���k��I\�&���IRoⷷ������&�<��θ�a���DS�P��ĸ0��)"��{��/ȩ�Ctvv�<8��o���H�ZPΏ�]
$�$CY�Dv{v�1t��vz������$&U�}$�	�'�-fO7����}�ӧ�M0��i��	����@¢TOd�nck���seM���GPV��� dLr�|�\���z&֍O��,�-�0�jނ�	��$&8�x ��'a>j���9���s�h �ݻw�����;v'�!���g��?��'?���+W��ܿ�<�탩����m^�ys��L����u]&o�H��*HbG������˖o�9��D���<�/i�]t��呐���~������B���=��vϔ*;��B�^���|��7����[�)�-�ܶgi ӛ7�0`O-�}��[t��4n��Ա*����y���j���]5Kj��:�$�4�ed�C���ݚ��./Y_�C&`k
xti��V d��gj�M����)Je\;�Jd7�2HQs��K.����Ӕ����v��x�0�[-*3uU�`�ʧ;��f^�@��--�H�X�6��ԫ�6���h�΂�
ɯ�dޙ�ly$8-��Ș�����.�;[��M�+
��3c1fگ�ၸ���o��`0����D�l1��j�P�n��v��#���7`�pU�:
R`=Fؖ#"c�n��9�u_�|yQ���qٚq\)�]I;��V���^	�{l�&�US���5��R�%n�Gu��Qᢅ1:<�h��+���J�b�Z�^횪7w�dd=]��7v�)�^���n/�33l#mz���KI,��Cs�
�\��6��b����k�4�LA�Rq�4�<�6�d�Q�t���p����F��Ц��������p���	70�=p��Qw��\���^`$����e�� ���2�I��L&&:Q:Z2CR�"v�K��su�y�� F3���(��l�cߟ����
*�y�燜���;��.�H�@
���N1��<;CSh��?~ubv��¼4f!ͭ�-E�%��&��do� ���Q����u|zfH�Ѣ��ɹ#fsM�� ���W���w���� +?��o�5��s��`�204<}�l�)Ue���K��-����R�A�A2V��>88I�r�jSV����YH�6]��Gܺ=�-�}�\Z�Q��s�P�>0�:����g/ 3���թ�y��I	WD-��}��`s���4G���K˵8`�7�0��,�Xa����ӓ�1�)�M߭�.o�����o�,-�"��?�Z|��Ie�3_5�U%�b��Ţ�MN�����,48$��8X6n^9�R�櫛��\v���������V��d��O�4a����$v��U��֐�FK��R�6��|VՋ�Ҥ��G$�qr���l\5+�8���>�=�Eﻻ۶�&χ�/�G�{�l�����Ν;�Egϟ?U.[���;�U��O���[v?��/������6PiʈكX��1�G/Ntr�4�IY���C����u,D1�M�4�R���3(�p��|�����u^��i�1K����϶��|�A�!��O}]���ja��ɲI���8��B�:�5�ދ<n	8g��Ux��z��ƪh���0�"u����4�H�=�2S�U��e��)�����5g�\��e����)l�ݻ	�]���T�9��+�I�"_|Q��Ybښ	G�&��TO�.�^�yi��zٵk=�����k��)&���N�se�z���N	���,1�8�Ĥ�^�yz��=dg�]���1+12�la�/��K����M������{ν��}���XR�c���l2���ܳ/M�('�+#
S\`���6��I9�U�`��ab�<%[�5x�z��>4�N�ݸ��y���9�=����1jf�TV�$���u�"==5�kwv�֋uU;����Q��)�oڮn�+�$,V�Xt�U
s�Ԫ����VO<v ��ٜX9��c�D����Ny�8����T�[�P����h9����i��v�4�(/���F��b�@*��;_b���x�K:E4�lMPkY�mj�����B\kf 4��"��b����f�ۑ8#.�����N׌f��g�9Ř��'�3S9�pT�/�B�9��� )�v���,Ľv� `��PE�/��������1r�d/���Y��ȇg\T��p���oU�׿�ۯ��P�eY��n�ݝ��њU�>�e&l{�Ҳ�ɞ}��p=�8��7�T�6�>Gj��j����<������k׻+WSX�����_�8���P۩�^&ׯ_5C���?�����|ut�x�������m�p����я~�sg���W''������wu��žż�v��)�����zq||b����ְ�'��[4�M��S�z�ٯ����9ܼv�ӗ/_>~��n�%� :fXT�C?�Ǎ��DE��c�n�U]�@c�6�er��m�S�o�|ɟ�!���
��P�Ki�A>��ڣ�k�՚�m��:И�����^��_��?~~x�w�>V���I1��������_��W�χ�|���O��pk2E���ڡk<_P��ƈj�$%1�^�I�6д�ԥ}V8y���\��7�d���0�Y���
0+����Խ;w�w�F��E{�d8�ы��$F�t����H;�y�L�Yd�Q{Y�2�Ѳ>*{�����H[I�VAl+��k{h
�D�������&'ϟ?1o���nl�h�>c�~zp�o{u����0R5��98�L�y�:�B/��D�.zS��S��D3+J�+�&��ݻwc\�ZE�	������ba�=4�hk[�pB!���ޙ�� 8�8;WX�(������}_p�^%���I�lu!��4�dc���C�9e�=�l�8==��|txh�=�/�f���,�`@���Pi���iY&�	 ��U{��-!y����S���w��2b�eQ��+3��ܾ�s��ִ��G�1������v�+�ƀ�YG+��X��+>Wo�sYr���<�i�~��񋦋$��|��K �P�Y���!���J�ĳ�М��t39��DYnų�� I⧝�?���|BVn�z�F�z��i�������*��O>���{��I���;;�o3��<��ަ��4cwuu���Y�g�/泋Y�Ҏ�r>��ٹ<u�3��^7�!*�����G��&���	��+�Eɹ���L��/+WdZ��*��dp㡪�.���ڕO#nQs=U�s����m�ǶGz����
P䦙L��ٱ�K�S���D7��k�����=��l�KT�R'e���s�UP7�^ ԝ�)�6��~$a~���)��)v����<F����g�ߘH��j�iZ��MF���;\�h&#X/Tn���N�TIH��t���w���\�V����>f�����22���Ng�r����y��m�B�a���]V����R�����t��HK�ǭ���-FG�^���=B0!��%[� ������o�ɉ�6�f�%���&�*0i�B��?�DT�׊yT�8��Z���b��J��=��Se�ժ6��p<���?i1�b��������(W����s'�J{�)�,��t�Lc(xK���>�&t!)YY��(Ø%)�d�[a��P�i@?���g��$�p���"��Ϟ(�k>�yϞ=��R�!����|:e� �	���d6���N/4�Y�w�Ǜv��8�E��Z���n#j�U=?_ɥӬ����N$���c-��6�z�D���,��,���`H1��v�Ia�B��4K�>m��\�T�C�D���M��q@t�&b$�b-JO=�sʅ�5�²ӰK�!Ҁ.�+r�VZU�ɤ��>�<����0<�c���ۥ�#�	Y֪�~���3H�VM������%`\�a�k;�ƕgfkb&�C��,Tj</��NZKmh��!������%U.hYj ���¶�|��]�ѣG�g'������i���W_|�Eə0{|�a�A!4�y�4�B�:�K-������b�u��k*�#4�m���{��Ӆ$�EnR&ȶ5v��cbuԇ�?���M�Xm�C�5�?��K�&BZLn��x	�d8Є��o����v,�c�����FR�y��N��3ƍ��J��u."S^��
�[�8=�M��|F=����:\��,m�Ы��آ�S�ٛ�~���Ɍx�Scw��5 �/S6��������I߮&T8�Ѳ��F�����õE��kɄ�U�o�քǶ������/��X"�$��<%3K� �/ˁnF�$�1�B��c�Uˎӗ�	�#���*Om�y<5�k�����#	c��٠R�m 5�1��왔�0�3���I` قF
{��H͔e���a�/����'�ӛ�����_���:��R�|��	��FIQzf�,�&�Ϻ����2���z,���0o]Ά\&����1�����rlye}`�b�8gp�bJz�*��� �$`W%�:�E�k���v���m����L�v�zI��:���9�O��,�{�8�MK��Nc^��[��G}�w���e;�־��s�YD(&E*���F�d��������/��$��[ם�ΰ�8�f���~OX�����kea�М�v�O�1�v�i 
�wT����}��wn޼)8����禮�_{޻w�J�#�_޲�3{�ӟ�t1����=(�`O��y�����l�����|�p�rNO��)��׮��	�|-��tƙ��ӧO�ܹ�N=�y[��l�9`��e�X�}k�����ح�x�B��b���i��Kp��-�^���=�6bI��]�Ôj1�E��ʕ+fX��yj�\��8՚����D���,'W����3>~�8a<8$��k��� �� ���-;K��������o������a��]���;w�� �"��(��g� �7�G]H� �.('�=JUpf��*��2m�k���pU�j�������"��\-����y�Rz�E�ܶ��NI���������@�)��V�e��v� ��+ܕ����g�}Fa�5����q*����i�$�}�p]��эk��mN��3�Ԝ:�i�Eh�V�ߨ���/�ؤtX�X��x"�+nܸ�w�w�A4l~� x���0�Z��R��9&V?����Y���J��4Of�ȣ�u���y�;!!�:ąY4:�y�r2��e��ÇE���m,���}�/;R��R����C�T�H���5f=w=ǁrV	�3y>.�O9P4�m��~�0�N���_:�6�G�]L����D�(Q"MZhLJR0��6�6����:"'7\���!�wR�dT5��n������V`@��of}fS���6Ԭ�S��+�}|�Q`��J��H�����$��g�fL,��� c�l�yoS2{ഞ�e��0/~0�ꌠ<���ˁ+RrI��5	�\Vp�`f݆J\��_WM��=m�,I�NI87�/�d�;���!-�ޔ8����r0��S�tz7Z{+�y���LmX>�6�$OЁ_7~�vh2AU��"d��r1[l�Q���b��)���9��Z@'d�M��8U���b�Vur�Ja���(��X�2�I����y6gkTc6�u]W��s���!}^K�
�x���F�ۤ�#�����8d��Q�u�S�.�\���v��bɢZUU�L�ܠ������@�$�9 ��g7���V�
��Zy�BU���
5Ot}I��y�v��y�P�̛*�`K�W�}1l�޳`!���T'������Ud!�'!�*4��ռO{x�5Ҏ�o����F?
0����m��ǌ�|�WЫĜ�R3J Q�Qx�ʞB\�� p%�ԗ���=L[�M��5�v�#JR��fL��n��*/����}矷�L��&�B��ĸT��+�"8u4"�/�����t�M눍��DU����b��rU��T;�'w:��M�L�b"�[,Vd%G��>l�ego�g�X����pP� �����].WU�fl,N20+�b&y��R��i�$�ƾ�<���j6Cj��V!�Ѥ��&�%,���r��l�J}�&�&v����˄Y�&e���L��ɢeYֳ�u|߁�ځu��$f1U'�\�yե�0���͐�΄�����P�x\, ���;{r͘ ���M�C&����-�tYۏ��� h�d(-r4�_p�C6(˵�$�������������ۊ<b��jn�b1#����Ϊ:JzwrV_��Ӵ�4HjQ�455���3(��p���}ҴI���GF�eÁ�r�G��H�J,�͌l32xoXj�2�l�r^�D��J2�<��T|n_� G�ʚS��X��!v�H73q׮]�zU���9�ͭ,r.�jt��3�?8�A��������[�^�q�BY;S�0mt<�l��`*��>�?�N�,�Q��R��)9+S̀��Pr�SAC�0���b/�ټ����l��1��8�]`��������T	����^�f�Ʈ�	H)�4䝜M&#9�@S�W����g4�H�+, ` ��[��wb��D�U�h}��HBk�}F�pl��Y�S&%!�P��lwL�|�ajLUP�8�T;���,�P;�"4���݌��
�gg>-�*�=u� �1���S�ߜA�0?6o<1G�V�0O��������G1i1��Ȃ#����b{u����LLs���ǫ��������0�������?��ӣ�'�J�1 �<��-fw{�=�|�ΙlT�u��(%�{8|bH�f,�� ��v6�H>6P�K<��p����z+����ϰ�.��S�����՗9�F��w�_��:}j0��zS�y�`�\�g��C�!z<ZQCƜ�����QNSr��h��.���ƕ��4A�fc�	��,m�� }�\�C�a����ׇ�q��B��G�(I�<Q����[U�Y]����	�YV늼`E 8�ȍC3R�L��
�M�Bg�.g�J�0�sr�oܸf�>xP�i��i������s�:lO�� �q���@uM�|���vD<<�V��>�K��λ����TP{q1W+VUc0���JU��
M�f}���=>��@*m�^cP,����~��n&F�A����͚A�'�b ����� ��R'4D���. �ߍ�]�������)(R/c�bk{:7�_�8;u���f=.Zs��#�U+3]�l��͝��93fF�2=;?y��ћo�i^b�Ol���LVTY����&I��ǟ�.�ڝ�K����6�ԓo����h�l�ε���[[�ԋ��~����t46AW+@�	S���|_����VD�t�	wm¸�,4���^����(��ryp�������4��)��k�"���l>;7�nNL�����ZZ�;�ٮ���������W�_䃺kcꡡ���w�<{|��׿y����K7��� �y>���%�T�P�쉧�C�e<"�Z	 ��) ����X1e�n�<�&Z1�'�{���_9�ꫯ��������&N?�џ0�G�j�$m?*Y�,�gv�!2nZ����)�����q~v�М���W�}�F����?~mk�N��9r�Ϟ=��O�w�/^���oV��eM�����u||j��yt(s�����LM��GuZj��RTʳFA�<�YF	�R�J�IM����H�γ:��W�l�Sc�Tj��$C:PB�_�z�`�4�Y�W�N���>���/�@�c�l� Ǉ��#�b�$	�z.��$�%CLݫ$#���3��ɫ���
�k;<v�M�Um����*P�ئ43�����ñAa�4�gO���vxM3طl�9p��	�6��ޮ��`Ah�-�[�����1]w�έ�Ϟ�|����q�FwZX�RS�#'CR���	�T��UȧT��u��ۀ4�����.v��(��@u��xCg֪O�ɍK�0	����>\lf�9���X�~K����;G�����lb�jG)�a�=�	y��A�1P�y�F�hh=t _��/�͟v��\Β�Ĩ�]1���@�HEh�9m�x0�%�bK�<cRӪC�M�:*�G�����0� �5(Vk��Q�g\��� ��r��%+�=M�ȆX���d�)�Ьϙ1I��N����
̹:v(�:Ղ�K�Q&D�����.jF)�,����R`�H�0�}hA�_���ܫH�B��T	2�nj۔B���=��,\�J����	z�.e�"z�6��0	�EJ�{9�Wg���w�X�L�"�F��cB�Z".�eB-��ʹN������waB�j���@���ު+������(�,�R��'q�ҫ�+�����T����k�K~������f7�fr�^t������L�ȇ~8,	̬)$�a�ٯ�ѨV�(/3�:�(��uӒ���$dY����P����aG{9�D�Hc�@�C�q�1�f8W��@�P/�jSK� xL/�]]���}�6f~0_�n/	Utnb�K�!D��u�����(Z'�6�u|�t:��!Ҟ�i3���P�ox��4�&��%��aO+G٣�h�2v�<�=�R�������61��5��7T��%���O���1E!o� 0����t��F��z�dƷ	�|���붳�y�����bw¼�h�f�(��À�"���I�i:�:K��u�[j��-�� �7�r�WJL=I��d��>y��Uq���k!}�B��>f���}�X�RV���qW:���2+-'J�@�|�+���G�D&��pYFx�T�X5�����p@��|����}����\�	6����×b3�!%YIbA���ę����w�r(�=��G�\�n���"7q*=��~E��,/.���j������2ql�h�=/с�-�1T���q/0r@����e��Y
5	/��y�31u�����s;����h�=��bE��������(o������v\�/sո�W�rd�*=���]�&̩�G#%�9�����q��iI�$� �+lk�J�/��@)Ci4)h�p����4�P�od��˧ώ�9J4�mmu-�.Ó�������@��])j�6���~�Yxn�B�:�j�k�qA*�=��I!�L�����n��<���� �`¯�5Hud!Ͱ�a�2\�0RAU��W�]����3��+m1��A��L@O��*��4��> Q^�2=vNu�j��6�-�6NOW` �O��^��R ]c�A�+��Z�i��s;���	%�u��Ax�ȃ�\b�|ES�yBC@&&���(�ڮU ^�R��o��Y
������"�W0�i���z�>L@��t�0too�n��K;�G꾗3Б���3zq��w���i���&Ig�G�O�(rYZu=���gZ`�p��0)^6H$ M`��OY�;3�����xk�H��� R�/?�����}�,~��*�5K��;"��� 2�Z���-���J�QÌ�jݤ��Pꄛ�ˌ0���ua@D�4�>xq�/X�2	>�l=��B��%�%,�i6[4��'O��'�ݻg_����޶lo�>p��mj?<<��]+u�7&��m���G�����i{7�a�<>>�&��n�tA^r{�YH�>�{���^{�mz1c�	�>��R圫svr,��~��l1:�Z��i'a�+2A/b𠛨�y$�wsg.��#���j_}�UTb��}��:�?�
ǧ�H�oyQ�
^����:�X�q�~���ׯ������&�F�?۔��>�I׊����eI��׹���&����ۇq�f.��*�ӑ�#y]�e_�m�o�akbo��d����~���-!L[�E����I"<F�(!^/�/��uw^C����h(q�����������,��ٹIΓg�@�;��~��!(Xv�t�w�����v���Q;�>�:g��R�݁�����j�ձ��|�D�bt�@�rVl����!��$�s�!��$���,��J������������lS�$��q}QT�zF�i����!��A�����򑵥t!>������W2�!������'JCo�]j����!I��4��1浛^�c�������W��{�`2�͑����ͳ�^U��{��)�hb�6 �	#2#�<3oβН��7��s�y)Av����KG��4$f��}��R�"	$��Ƥl�T��ѕ�I3t�N�l`�:���YƉ.ޟa��,Һ�v�t�ԩɪ�n���Ĉ�O��󈤖��i�'�`��d&�4�<�U(��п���A2q���g�vW��]\�:���[���c�W�d<^o�abi��v	�|a�jG���.�Xn�W嬥�G-Yv�0ߕ�Y�����j�t���˔}�H ������v�͕I��J�����$�J�Y&0Qu�E���5����--N扢Syq�F�Z:q�3'� �z��-�갞L
Ѕ�]T�[0Qb��2��bۦ5/��`Vŝ�Lc%ʢ�zV_��GR[L7�� �̀ �D�r�\�4i�<�x�,��xp��r%}� �g��v[��=�"�,�v�2kg�mʶocF�+���nR�s�&1�Esp]���n�Vm���^����;�?x� �ӐǤ�z{�bT����dC�i����\�JH�F3�zX��*�a*V̝����:Ĺ�2cʸ���vLFn�j�O{,m���)aL�)��܆���A.���#�FV�
#2IAOG��hc�e����̎g(�%a����b=��p`x��y��_a���yM}1�omḾ9?9�asc甚�C��F1��2�Q�e�ajvf�~,L~h�ŀ1� E�fEډ��Lo3z�?	��ih^S2�j�7\g�U���f�ӣ�b��	�&Lц�@���g�?��u]��ΟO`%�h��
����q��@�@�(�*��K��Z$`3�gZ[��A���f�@8��x�pt(�S }���ӹ�Qv�4�N��0d���'X�˴�ق�ְD'�i`�&�-��ɐ\�Xg����|rz��\�� �n��p�k�L��8z�mMk���ϲ�����u}�:���#t�1��dȵ߈P��>t�yx����j;{L���o糚+��l6����Y$����굫J�[�渵����.j����d��oW6o�ٳg�-��M���ԛAƱ����*�yn~ؔ���`�(�3�b+�R����وc�+�B/�����7��\�A�415j���p"���b FDީ5G9B��K�R ���ȭ�P�u��}sUu���:+Ն��Dh�C��u�����j�P;�|*����C�T#B2)�4QU?Q߱�e���9k5��,�h(m�1��'_!�M�~.6���q��v�h�TKχ��]F#�ah����ae��#DS��4�G/�NNg�����7޸������o~���B<��tlʓ�$��K� �*�J�Q��bX}¶���e��n�j��$�"˔�Wލ�Nۅ*�]7Ӯ�D��o�����k3�[�[v(�[C�#Ow��t�!�מK�k�ٲs[v���J��[��d:=S�zϽ-[���F>S%�bXb܏<F��L����/�G������ �j��}),˼os?���X6P�\.�Ԇ����3�|����u��dmm�[²({3��g�5�O�� �y8���,r�H�!M
���c`:xc�f�]�����G������%��\̔��ʈ�F��lY�#��и��۟��� x�������/���Ç��ܻ���'V�A�wи�|��j���P�ؑ�lk<�A��$M=7g���9��|�Iy(3��zR���Q��g.��LT��3�~b�SΞ�r$M���*���oN_��|u�`���U��ƍ��W�\���{��З_~����+�.���w�1�z��S�,��{�"M"�`�\�/fv���h�Ԍ#�=ȕ��j�x����|jC�o�=�@}:�e>���$O�/N�M��:Vj8ݭ�G��)���F��%�1�_�)��!�tK9���¡�	3a��sh:T(�ʉ��)ROy,4�T�`���g�)wdj�"���k��&�d�Eu����|Qzm��{�^�:��X}��um�������z>�����r ��߻c�`'�]�^�<Z-׮\y8ooo�WO��#�̀7v�b�J����I�+�Kn^"��D�����&�-.|l*7��O>�d�n��ǯ�g�4Y-�&�G/^^��h��r�G#k�M�ЊcI�C�b���"X+�#�9���Z]�e���z���?�ן��ρ�J�:h'�Ӯ[W愬G�A���y���&��!��ղGgX��*ӦA���@��`�#;?G�<L�&�A�d�|}��Jy�J����I��l����"�Dݛ�%�Z?��l0��'�RVd"ݼy�������}��h/�}�'ư��h��~��I�TE��8Ǡ�Ҏ�W���
6{�%�#`~��k����� ��nz8��_
2'!���sڲ������l����%z~b���k;vW7_���V��IƼ�	++>�)˕t���Y���W/y�	��̙�E�!�����	��CX��t>�byk��|�C�,|��Z����?���8����i�.̰�@��BԠ� �{B�X��u��Y,���^�޷�L8�3BMYLw��}��S/s��%ʣ��#b�T��gGu5�qm����٢��ڧP�mU��\(-8�׶y��|��YkA�f�*i�б3�L�[f~�S�3�����r�����WՒ9x�dn�����jv>	Ї.n}��]��d��!#��)�_��<f@��0�������ԘO�i�v��(���(OS��o�F$5[�ߚW��Q1�����m��~�{�M�4�#��N���o��Jk��E��'ܓ����0&/P&!�����u����Q��@��0>�3bNM���;T"VK)�6���0���Đ���_zMs�c"L�Ƙ$ra.3|,���W��h�|�;�2�u�g�Qgz��mx��:�ap�:��W�xJ0�Gި=�D븐	���{W8J#|���y�X���R࡯у�3���;��=��؋,Fr�	J�bZ[s3{���+�Le��M���Rx,C��V_����q��P����@GUa�/�D�-]Z��4>	�*b��w�D����y�&�������_ga�,a=kSu�\Z=�F�
��y��A���P;�+�G���i"ݐ{�N��Q'�^�q�}H$���L&#�k\�Ċ`���p�K��7���[U�� �?�Mǽ��2&���B%�OO�#	g�z��Bu�Lɍ�%-��V����Id��L����V��፨J�I�$�%�tN������|<J��Ts�c��[懯���.�'N��W�g�e�t�ď��I|��v�o���vK;trt�M�:�H��:Q���<���ѻ�{���W2o����?d�W3�gj�/YʐmO��b��a�����\[o��Z����ٻ���l�wF����S�=��vϞ=�0i�H����Q`׵�M�a�M���>?�d������"�&�#�I*8>R�����.���d2����W�pv�~^�j�a��Ww��Y��� j)����]�EY��V?G�k�(�׶�ݫM�f�6@�06:�yL��H%u����H�,6��&�������#\�Z�_\D�k��Y��mɉ�����ì��V���fn@��k�+7����9���P�*�C��D��F��4[4��p�����~��Wi�K���c5 �<}� *���;W�5���7��r_���x�S�=�t`q�=�Z]��4������Ȓ�H�����{���7�����߿�.+�i���m`����e<W�g<<<���K���N�N�>��L��&�hP�,p���dW`�y�A?z>�Y(�ˋ�Ѧ�O��pPDOđ�a�eG�G��H���҆���v�=�,��V1=��i-�}�7��f.[^4H��1��g3��7у���v�ޑ�B�U�@%�]��a$qL̅mJ�D;����t��M���]�ژ��ׯ���E��&��߄�fT�wV�,]���RD.����^Y�=I[ZԢPtIE���h-z��sf�U>��璁Cw�D.}�Iu�����H�� ]�+�/fru4�ß��)|a��+�֧w���Y�9��T�yCڴ���4DK9��޼y�������IT["��\����} $��9v�Dm۠KT�x|�g&��I'�X�8X	�,M��SN7V�����������T0��1��rJ��L����1�q�5�E1D��/�79��
�l���{ �?z��&S�7�����U9�����7�<~d6�a�.���������Km7E=!�mp��ymY�c����B~�ǶiȆ�u�&!���tƢ��i�����~��'&}�{R�7lXQ	��z�eԄ�f]Q�����ɦ�*� ��=+�M�c���~�c�;�`��W��������+�����ɺ�q�;ѩ�I����(��"	Ι̢�$�ڪ����z�>b�_e��DjGP�P)3���W�H��`>��mC1���<Dwل���R�t��;��jL/);����}`���i��@o	��J�.���75#$�r��^�@[^��O?���u ����l� {w���Ē��#P#l�^�0h2.�����"}�����vcr|��$�0>�9�*s�x�^M�CY���|* V���y��U���D�I�J>�]�!�@���K�'�����������U���Ыɠ�en���9����+n���&�< �o*�"�v�^�I��Ms�ś��'�6�����=Ana��D}s9{D|\�+�x�׶7�DJ����V@�ECd}֔&�U��6�v�Dl�Ț@���6�r�Q?࢏�lݦ�b]�ل�� j��Cr%-�,�*D��R��\�9��R�9ڿF�j��V��KV���Љ�=q �rinQ�y�&�Y1�����$�9Ps�*KL)�J�VU��{���"�;7�7����+cAP��2�z	ө��j��ڗt�U��DŴJ�i�k�*�BՁ�;�z���j���_T7������"Pu���G���Tk��&y �2C���u^���m�֧R^�	]��c5�8��8i�s�8c�k�U<QeJ�/���o()�C�B�s3�b����^�:������ʄHa��Z�5�uJ7�$�f��!2 �Si���z�(	z9�j7����=�r��,f"jש��#�&Ϲ �c:�w�7������R<{_��fNF��`ۇ��x'�����+�.���rNV+&Vs�-�@��O1.J��������_�?zj�x������gM��|��{��a3Y��s�&��DB��Cuۀ�D�P��\�Dr���+L8���'#���������EI~�)<�&�u*�	?�V/-H�^WfX<�B�(��8����caVAr�Da����Ԣ�.�(��i�KUK\�!��KV�!�t!'�l�Bo7�(	�����Ml#�?V�j��ejC�)B
����~I�:{�%ө�鴭oLfm��???;3mE$_�Z�,PI௘�Țj}��(xf�^}v6�Y��G$�]߬�K��������� �HM&�����X}냽��M�DoCɈ�����r~��/�"�F����{���#%�����2�W��[�n���=�LmN@�y��G�*M�|�	_ah&��p�R��ͧ�T͎�9��e�s�5�Z	�TN������R�/'���"�ړސ�г��Wz�������z��IV����VQ	KZT�77E\Qv����ϟ?�*��_�}睷�z뭊s9~��b9k�z{gjϾ\�Cm<��3w-L��8i��W��d���͛vo�E[faNtt���{���i�1�J�j�F����=�,�v���i����o49d8�B?���R�:�R��Q�&�5&l��Ijgj����s�d��mIF>���J����������WoL�����ɞ�O�h[�S y���E�eȋ�=������1�g�7�7�����_��_{G�yQ:����.���t�tol�����3��L�Uq��1G�z��eA�Ѱ���"���c�Ģ�T�-Y�ɰ���h�=�	�����|��w��I��S+������������Ҙ�c�I�,(7�j�W�Z�2�uYb�<���]�4����� D`����P7�.FJR���Ǫ�z�P�K�'��|�,4:�mW�Rf �-�Q��n��!h�.����ݿj3u���P�G�#,�i\F�8r�'�� ���~��!Ǵ��k:Z���R��%�Ye/3�r���s��H�y'��7XHr�0fA�+�ԅ�$b${\ ��^�C���Vd0rl�{������k׮ي|��g���lE|��B4˵�9V�X�:�u A��o�mb`D�W�a�1�+"vY��u��d��`���4[[|J�%2�ҫXN���3T�k���_����������������޻�P�=��>|��;��g� �`Ivm�8�흽�|�zi6u��YpZ������jB����o����rt~~&�c�w�����Cb���ry��J���~�=�8|���W��yk��s�����-���F,��×_�������D�L�l���|剪��:3M	*���<C��o�rx�m����,��O/��M0�V�d��~V˕|�PQ��/�<��Ffv��ujo��n��kI���'�<H� =ܼ���{fXW�g��/�lK׮����iU�ZB��'˥�Mz��L�.���3�@�@�H-�8����BA�]ӖT�}����g�''�h�\�go3#9��H��{��稢9đd�'��f�+ji�-VM�$��[ �1���v�]n"WǇGǇG�<�/me�ģO�(��c�W�Ĕ�J%F���ЅI��}��`0�rU5׫`�>L)h؇��]+�%���L��^�|$���T�HB�utoh 8��w��"teJK�, �9��1"����{�������.�5�*�eT{i B60
v�kI�b�uR>|�PCSfWm3��&��. T��'9�H��[���c���F����4����rq���8�׫Œ�б��{������N˜����i�&{T�X*�ږI�&}n�N�-hOrD#"�UWy[�p�<]�Te������[��>!ۉ�t��,Oj�2i��M	~������jY6Da��u��A�\�>7}`Y6mY� ��MO��kξKɿ�j$S�<�e$����)
ZD ���]ͧ�}���}�Zb��Y�$��l��+��k�A�������x2�w�������� ��D;F��u����h#wd�sa�1����Ӊ��l�%�E�F-��6+J ֢����!�'L�L�<��uըo�2	�u>�!,@�N
 ��x����O���6��n#S�	_
;�E�J]U k�
�Ր����|�vS�����}�ը2��$M�]�r!3(�H���b�墇ԇĭR9U��c�h��|r���NC3f�e�W�SM�D�)��rΓ c癉RU��tқp�{����I���9�.$�e��T]Ȃ��r�����b�m��B3N|�~��Fa(V�*f��뻴�yu�HCVw䏚�k�p���%�fNd��K���׎�ӳ���m�-����I���	��Ѱ��	;�M$�rk����h��.�Ĺ0M[4�JXd�˛�!�se�[��E�Mh�`��5�xV�g\I��<�ʪ=�	�艢�O��oj���ؐ��=��ѣ� N�.��������K!5��U��׵u��)޳:r
Fa�*Td� Q���W;�Juh�b�QW�^w��U����DuP�Y ���.Z$7��g3��<2��^��i#��z#/�������>�. p w��[:G��J�˔|3->e�x^W�<Y���/|�-D���Z(�+���uR`F���`J'/�N1�z݌�*�d�q~���U�<��p���ϑ�t���6p�8c7�`a�\1D�H��<K;J���7�oo���j��F��~��GC�_̎����׮^�y��\Y��p�&b�s�مf��ؙ�V�x�Bx^�!F/������j=}�o�V,-�����^2�yb������\yC��x�\çO���2��飦��7�|S���JmU1����Jw%:j���l��sL;�d���o���믿n�lu�޽���B_۴i�)`�/���؏�-KD�$�6k_
S��
�U���B�O�:2�5��9���s���Qtf� �YKc��g�
�������VN�+'����Ji#��"�A����y eη4�+�����q*�@�},���dDK���E�&L����`�����?��,/�~�ӟZ4~v���6�+�ΐ�Q�[ï|R�e��Y��|D*OZ�V�����؅2���n��� ���1���7^��n�j�u�Ƶ+W���1f�,��c�"�����{�?�bt�	j�iae��6.*�2��.E����U�'������V�Y(�> ��.Y�hҸ�}���IXGh|�Q ��,�]{�`�Y���<�Lr��m�Xh(�b騭d�P�[RC�2�j��0�,8}���o4Y���?���[�NE�=!?W��8hE���bF�D�L���^��]x��K�wӂ�|�RSG��1���Tl�W����;�s�Ν�<����Rqdɫ^+��@�Tj3"l*R(��B�6p:kYb]��j~��_���lۑ5�!�����g�n�z������~���k��]&	 ��L�\���E�{�87�9qq�����vY.;����?�䓮uf�b��@�6�fGr��	�̓�j����m�LZf֟>yd_4�K���GZ-�J!+�4�}��}j����!ޤK&�&�Q���!r}��y��i���~�-����|`����c3v���#�YI���\��M�d�����P�0�8ɀ�*W#�����9:|��z��^O����ݯ�ki�$��+��Uj7�wع?�C��m����ճ9���4D�ZA�8v'��8:�QA%�m �d�4�����p]�l*�w����g�7O-q�db�Dz�j�m�*�@�/�i��O�����x<R�Ѱ}���+��Y�O��Y���T�ڬ�F"�)������(��/� �����#���S��!/G��������Cב��,�ݒ�;m�w�����;����Z/�:��b�Q��0������rC=�����<z�h36��(�|֯	�|1!�G������.	�����t��ɓ�=t���aNݗ�}�_��k5��SX�	A޹��0�e7�ou�j�|��n�Nw�֒Г�g�Z��<3��w�Se�enx��WPd'�i�F�W������Ƅ�^�X��g(�#�_]�E��TU���A�6��i���ܑ�7��M�/[l���2l|�㶊]}3��~[�|�&�|���5�/���!h*�{����>&`����.�d:�	�
2!'YGl��.������.��8�C2��g�~EiWz�<Dz�k�d�4pi��2RM��Y��ㆺ���hX�C��ue�T=�����-�m�%C�Қ	f��%?�r��D<"O�yd�r�������g�5��0�Y��l��mm�����Y�&�x9�Č��$<N��a���酄��b.c.�+��--�	�J�6%,86�_�R<�G���Ͻ����X^d���wP�� ��0�;�'�汁����!� ��Gy
�y��oܬe��c�1f.S:e���@�� ��6t�fE�6�����q�m_ �쫥KF�`�/�xYh�P~T�B�M>P�[�5L�}��q���j董���?xI�9}���qPIJt�1��P��T��X�4��6�h#X��/��$c�v�d��T+���:~E+��
�/��KM�R�:º�\�j��9u�WTF��<���W-6U���b��H	)׍l��u�A���##�Z˞��S`�
 4�H_!2w!M���#�2I��	Gb�?�>\��,�H|�,L�ڣ����7��<�")�E�k[צd�fv�^�+��OB�Z2}ʵJ�&Lb)ael��/m�ir82]J���F�п��:R��S3L�e���5@��L3(O{���E��,4��X��(��LBE����0A#��_՞��͇ůd�D����ؑ;N{�]u0���O��R0t]S����7bb�Z�J���JA�7��ȩ�iӋ�2Ӛ��!t����y�
�����&t�d���+�Ar)�ܪ��]�w�ӊ�g��3#�&=Jvy�KupI��m0"i:���X�1��+��D�{{[���.ɗ.�Qe�p�.o�\(*؝H'�%U��	W��bv||���	9��ֱG�^yi��ʢD�j{_�N
���DH��UVTh��Ŋvٔ��v)=���_����/~�����q1��Ţ�X%M�I]4�p䊀�4�ǟ`����	�﬒��C)��2�J�쏴����'|�� ���"����AOD�W#�hd�/��hg��r����\�!B�R�]��B��ޣ,Z��O�?��k��rT�N<0�Vl�_CJ� �AAm� �Q�M�&��b����5R=�~����Y ��[o}����v��d�lY,'���H��4|�+�X/�ѐ�&5��R�<���ʓ<���{�j��7p�N^X����xz��e8�I^p�����7��m�a���P�Z,�ta<��p�g+eK���_�0�M扳>A��è�%�>�kb��e ����^�$丙q�>�� �`�)�K�\����o��U���p�(5|9�r�y��D�}ʾ��[�&�������]�eǵع.]e���vf@���H}��(�/?���@ 	���L�.��z�}"2{�����Y7�='N�; �D>2g�OP.6�0���Z�LĚ�2��W��Ns��$ՒA�����7��AV8�S���rQ- \y<�h��H���B �%��ҞX��q�:�
G�s��a�ըph ���>�L�T��2�³(��.&�i�B�9�1W
)�f�����)��ϟ�v����İV��ǏS����:�2��B���$�vD��b�E�PD[lfEo�:挆E�^�~�/�t�έ�\޺u��?���1��O�+<~��?��b6�����%� T���ju��mC�j�g���%�8�ξ��Vtc�������7iq>��s�§������\_���c����p���S|�{���;���ߊҸ�����������5�j,�s�r~~Nr��YF�_[���K�iP�F����)cU,3�*��S#5���`W*|7�޸>�4�_�����Nx!��^�Ku�%mw��p2�� ��O��}�ֽ;w�=H[L�^�Q��;���o߼z}������[���ʓ0�%�<�x���s���Ii6 ��Oz�Q����N��`I.�l�n!���%�~����g�w�:��U���O��;�?��{.�����gϞ��;�Fr���÷�I,��P�4�\�Àg�W_�~�ר�����(���_����Hm�Z�X̨c%�f��^�,	��ڵk�r�Jy9�ԂӾ@�8)87|Ikb#�<K�F�Ŗ�@FK�������y�]}��g�M��?��<;';m�&R���tcP����r��2�6��]\�j��L�#�n�O�3d"]h&+2�����Y�J/ח_~�^b��7߬�-=~u�/(�VB��p��)%��-�b���P�2G��7�)y��)4LU��Ah�c���M�F�Yv�e�:'^AHb7q��>���$����,3�����ӥ�LI�f��L2�p�����U���BZo�f�f�^�H�C�"�����Y�4ɢ�tV���q@��Ȃ���A`I�h/a�FT�6-P���q=�T'=��Q6%���u������9�FM�d�%�dn�`��P2$2W+OW�����o\�)�� ŧ�Lf|W���/.�f�3i��'��g�>���{��쌍D��lȟ=�Hz���/P9҉fU��u_8��R%�ܻ�g,��6sFr�]�M}�z�Lp�$��K*�K�JK ��D%m6gm���&�_1�u	�Aި�S��T�Z�u�l�$5��Ҟ-����POK�ֽk���1��2����h>����W�5��b͘j!���iy��af��F�G��?к(�uݫ"��G��
:��뉧�a0b��n�������JHK��R1�T�e��N���#�w��8��3�Q��Q����>P��>q\��*��%ʌ��J���Of��d�L��=[�i�[���xǳ~��B�诜_F&.�LȒ����k Kf�d6&�UP
Ua�C�u�2��>��:�~����bz(1�&-M��=�ɀ�������m%Q$xc�D��X��*am�43f%.f��T�8���tgx��҂�jy��K�'¡�/��R�Tm�Udka�|���5����bg@WY^��gNǢđcKu �6)r�e~��N�]u߹��C�������17��+�`�U�V��S�#^���2�cjKJ���^_�Q����;�j�۽M�N����s�]:�@Q�m,Of�� nf2�4֒/�F����t��N�k�YfB�O!�y�ݯ��)��@�	�^2M{�j�>�oу�D���H( S�r��0�`h����w�J]"Ke�o���,���$�(�W}A"̀0�����떕�:���L���
R@�s�[�G��X��T���8˞�Y��G�Q�ZÉ�Xq�y2�����3zA,N��ڈ[���lV��ə�;��Va�R|��M��^��ٓ���q4X�rp0}}|5T�PԿ��|���GR�Gg����ڌ�뵆������w)*x_��tF'��������?��&`��2�f������ؔ�@;��.r�&`�#1�e&��t�m�fa�8^�{����Jݕ�An}����s����n��y�:�\���XIJ"Z�'9$��.�!���j/|g4f�Q{�X��p��6O��3-$I�R�);$�Qn-���7�ո�$%r��A.8."��Dn�D,/_�-�>����ә"J�V���pb[\c�ȕƏU�
'(-"UqǵKj��K]���ya��C����?�Z���5���d< 6����</����<��a!ʦ��\-[�i��v#띹��+��({��1�07�/��/���`�EKF�Kq�44]�jY��&���εo��tE�ۦW�5���#�����2OEc��b�*O� ��X1�ȃCn޹���ŋ��T�SD�ح"����JМ��,��ͬτ�!ҋ]�=��	��&�s+C��E�\:�!	L�r|�(�>�42X������Q�r��䘣�x�Dc�=�¤|j���ޏ�bn�s_�����85�WC���xG�>KB�Bg)�`�\��N<W�fi��&!�/�KXί����O>!����@�7T�{�旒�u�4v�͛7xpB�(`��?����.�@1򘤴���&�T��e��Z��/��/��/R���'~���Ɏ�������qA����V����ן}�o?���Bh`>~����h���<���9j��q��k�p饗�H"<J6Ze�x_2�@�]EQRK���o0��J|���>�CI;�$:Z���eg:eXG_�:!`�6$��R*ay�����[q�&c]��B���/����O����|,QH�0/���)�덻�H�Op̯�c����F�Lcv�����IÂ�Ī�r 
�ŕ+�xzs*�6�C�>���w���I�m<�Kp~�(B�zX|@�Tص�ϟ)��
+3�^��S�`o;�N�tB�Y�"ƴ�C��?>~�j9Ӝ����R�ވ�N"�t�f8�]Z�[/V�q���0N2���)�늟I�@;�]��<6�]$�*62䡌���޽KE�8)2���\wZ#!>�qv~A+���_�
���N۪�.Jd����KЮ,��<�	�J��FC�/>]�#�ِD&h�Dw�X���#�d֧�_�Y.B�"ؔ1z�L�Jꆙ�8�P�����P�@�*f췬�.���ZE����c�]h�*�i��W9S�͐�/���y]���ֱ�}}>J�h����P���p����z�,5�A����#A�������U�Sg-PN�/�:ӥ�m�5_yd����v~Q Mt-�
�OV�Lh\_�-(Fjh� R�|��(����1�HDk����{�������|uñ6�����I���`&z�Q䒴�a�½�R"���?6��W��u_��]�ri���x��CO0K[�(z�Uk���h��ǩlB����Ɠ\�尡���(68)EdN]`�h ��&�X�N�9�@x
F��r�M��D���J�r��C@8�7�j#ND؇����c�J���Ȧ�{��K�V�d'y:[��k}B�L���	'��%ԨIn�V�2�g숊!�p3��)m�����}Q�%61Z'�6d�#n��wh�2a��<�Bd�Ǭ\c���8@�Ax�mJ������#CX8�#��%���Z��
�K�y+K٥ҵF0H�Mw�)	qWV�T��{(�r�f��"O�m���C��!1y��A^0����Ǖ�7!&[�`0�O�>��DQ�Y���`̛lޤ���{i$ЋF�z���՝�wG��d4�KɋiX�]0���*Ie��+q�����1e�1H{4�j��-��r�
:�hW�R/��_.W
TH׋e��/��	�i�/������%>��Ao��KݔU�Z.7�bL�5^dN<��r]�g\�h]4���\���A�$�j��8��!�g�	P�Ph<�tj9�w�%3M^�����O;�}`�LZ�r٣����s� ]إ:���˹�Ǚ4l"_�P�P�4���y)}xR��e�"6)H��H2�a�O�wt�&�٨��q�2�ʟh%��[pf(��Hὑ:���|&47�{�&��7��d�\�vM��s$��[s�Dΰ���
!��$1��tO+-�Cҭ)(d�T�Dj|� T`�qB�F�8�R�~��Z��E%4�z�b� Չ�*1.bD��k�1�A��G��V`x6LB�Z��UszrNFQ�=�0<��T�)���ї+H�HG#�ʺ���ԇ�؋��|�p~O=�f����¸�(b[{��+F1nG�ğz��J V��^sp���Wi՗d�R��]fJ^��J,����@��������<F�K��'֡HW�#�A�eݰJ��e������:��r��%眲�	�Y�BE��k���\�h:˲�lr�
����(YQ��-����X���uxn��>F$�����C\������ko6��q�6���[,f���o�t�M���E�O4��-�9k��޻�"�&:�*��ٓ���G�#�����?���ϡ��(Z6˻�����V�^9:X�W�x�����͛��jDz*�L���ѷ�r�B0���u�O:���%VX5���8�+���v�u�d���֟�w�k�؋���b�޿3_.Je�ÛW��r�i-J�WZlC��E-�����ݶI�~0;_���i���7�j�޶^e���o���В ���SU�]�t�t�H�D��j)�}����0�kI� |��拺y������U�Bȟ=�<o���$��w$阦~���|�:�zm�l_������(aP��`��Zi!�Y/�ș�)�ln�Y��٪2��Յ#!�;9?��m<���̙�L�N��8�~�0Ow
V_ zXa��Θ����b����F�q��*�BT+(��ٝ���E̮OI�L��.����쟡+7���"�a���ȷ�J����En}��-�ٗ�<ّD���6U9,򲯅_)mNĢ��)6�c��W�{��i�]jxY�q���D�0X�4e'6h���9��b�Xs^���ճ�KM�^8?;�}���í�M%�{�����Idh#�\�*���q2ɠW���$����Q��)b��r&G���Ch���[@�%Aஅ�si��V�Օ���@��b�R�&����#2"&��z����b	'i���W�u�{�����E닺"�R��R���@�7^�=O��3��慲by���	㫝��Y�5 e��mC_kG-3�)U@g�s�r��#9�´X�i�3�)�XFM�/��/����͛7����7��������"¦����Ym�v������th��4�E:*���%=��[I�ś�A��������+�w���$i� Y�=��>�����p��33���׫�����}F@��Ѿ<��"0���{�m��h\h&�J'"Ad ��`W�6�޼<�<�V5�z����r���c'��N^_;���Z&bAB>��D�_"����|c:�ZR�����0=��	^��������'?��,ܽ{�o=z��pwBT�D"�yY#pK��2����l9L�m��m���d2(����ȯ�<��	�_-�r֧�U�Q�Ǫ�
��O=BZ�rU��� �C&E��G��w�;=ܡ���Y����ɵ+�7n\^^6�t�{X�J|Nl���|O��B^�rA�Εk?�z���>��^Ԩ��1���"y��C������1����	�NG����K�ݝ�|ͦ[�{��iv����`�3�JOW��-每ߜ�^Ƞ�$�:�Hhx�e�Ѹ��*�N)����?�8�{�EP���ҹ8x:����[E�i&��%@A�Y�/>|3��|z|��<|?�q�'�(��-��,DXf�몭�x,����럙e"͕0���}�f��+5m6��(�rI~D����ty>�$s'���S�X���,MM%P��Z+ZP��׈��*��Ub�5�{��dI�6u�aO������֞u
s��E1�Fñf:l�4|Ӿ¾�����L2Ϩ�T�ؗ��$��1 |q6���;�%P�b�F#D�Jo�Sܨ�����v�O����n�?����˙�����ZNU�J�$��S%�w�l[�Y!�q
��A�Ӷ���b2��W�JLD���ڄ�B~M��i1Oi���u�^(�m�A�A%�#���F�r1��]&5��5�wN�}�v���+S��,�-;����<�+�� '�Y.��C���/Ņh�܊>~1&;�97�ٞ֬K����2�'ڷk�G��1�[#�6�%�����H"�ωS�6FRc4�T�������Q���&'�n���* �{�9���5��78R�U;����z��F+�ZGm�*~��&~ҥ�\��x���3%�I�Qe#��8�3����@���>���d��7l"Gat�}���>S�ZBHo���ݲ�~�	�E���W��u�pق�J�D�Ƶ��ܶ�Њ��٘-\Q+Q�:R^�q�����("����x���ɷ�t��Dl���\�73�_��@�a|f�>\R�~Ǒa�8~�~���Lu��\��ш��|G�E����n#��5�hyV�{��d� ���%%D����c
mq�K�¬tˢ�����:A��r�1�D���n�����5�F�0���y���/��`C!�8�8"a�-�@�)��UY|�͛7�ɚ䝕��B���C��\A;O������p�+�A#19V�ۣS��3"d]�ȴ���~k���+��^�K�����C��>�HV듩2�=N�
�$w�6bV*7��Ib�ҁ'��PͶ`����D%�"��g�+"�I_�tu�3;��Fm��w�Ȧ?�5q:�&4���;����U�83�8(|��j�׽���ɽ���N��S��M���4�����&��/�RphF���01䣛���
�3|Vk�����ʼ+�
₮���v�Iw��5?�th��hO�x�o� I�q�\���B����_$l�U���*��>����7�قKA�<3>�g�GIb�����kG�T���OuH4�ݻwIMH=����C�s�q����%rD�/2�x��+<�N�',��,�Bܗʦ�����,T�n�!;�Q��5�M�Y�<�իWy�yۂ/(W��`�j�(V{e_�]*�.J�����E�$�Ժ�`�9%j2R�ʉB�8��c��"�B�CHj��=���=�=}������?8<��Q)�������jYAr�6�����kG6���1�5��D��qce���do4��͠�g���	!NB������,Qk��znₖk�mqV�����R�m�%�_)�.!�W�%6q��/}�Ѣ ހ O����7����L_�+�q�U�&�����M� 9�Èm#�Ct Ytg���3�a� ��%B{v�%�;.]���n߾������E/! �;=���nݺUiO/����_��Q¹FxS}�!�&�����4"�)��>�i� L�9Q0�x h2&Y蓷z{����7��BO�m1$A{���=y�>�ڲ�p�h}�J���ׯ�x��g��]�H��:����GC-]�U��3��M�ϕ��Z��nY���5Zc-'j�����u�ʳ�.\E-V
�"&���#��i�]�+\���%�Q����ܣ��l�?{o%��F`�z�L��ӊKû���Ӝ�b�3�ԥ㝉�i�M�ߩ��N?ǣ}��gd98==��p���>��eJ�"YN�:z�"�$j�}��܀ɌGؿ�R%��>�?e�����^���6zY�3սk�#�����G����?���5$y�������@4���[u�:�y)%�̑+�s�ߢ)!���4��GNsiNo�a���٩�<3R v$�6��6��	]�b���3��	�h5��u�6�yT�!Xfs#��!�U_���;���i�{�=I�M��hh=����l�

v��s
7 ������Ce^�-`�%�o�A.��$6ďIa\�Ih����ɷx�V��'O�@~`"a��� �y�	�J�)v
���DM~||ʉωvRCz������w�5.ٹ��\vj4P��5A0�S�T�-�C*M�jSmM36�[��?���C?v5E���������5$��n��:򸻳)?�������I0�&e�8)�4���u��Z��)���j��Ƚ>j��ڳ���-�2�G8W
6�P��q�|�����'��9�+O,D̠���	��Ԟ����$7�7�w��XВ�ٌxv�Zq0��⹐�>���:͹����-�"jU%�B��$K��TEH��W�鎰�ɔ�R
��8s	D�j�O����lQftv�\���8է�AC��Q��'g��6u^�K�_3�9����������|��!��މK��:ݳw[o�����J��=��Gz�Pz�a��'n��d:�5qu��gk�a��!��CB:?l�I֨���6�/M��R��:�ě8x��έ��b�gP�Z7k�vkj���-���N@��J59�e��湽�a0�V��X�.��Pf~��z~���U��i�\BZk��(>%��&+�{۝�d3b�G��-*g��WC�d�=�AOf�|f����}P���:99����) q�b���S�a��F�R?4��wB�5��Kjߪ�Ӛ�ښ�+9�(O�9(��$-�k���������!��k.>��\X�&��M뭜��er��
��=g^.Bi�d�K[��2��U�YF�4�# 
��&�p?�Ƃn`�#�ŜY<�4�
�!�Ɩd���DoA����.����z���"���Y\�$���[{�gN�W��W��c��ʲ��IY����-<��=����(u<�1�$Q�3"neSb��ކi�w�{h���Bߔ����HZ0JR���"ޣ�0.����Ѯ���]�����m�E�[��&6�RP�F4x^��EU�M��f��0W��g��A�e> ҕ?�;YO��ɵ������Y����H�@gѿK�f=�^�/���x3s��f(��Ý�Jz�Z�,5bv��۷o'6w�|_��x�����Ut��?��O��?�\'EK��jUD)9�e�8G�AK�q��f��+�?]
	���p�w���1|�W������?1�C�s��<���07�G�"ӶR3@� :ɠ�8E�6d��Ӷ]�'W�93�>�p0�9�d�i��T@�m՗M���>M�^�8������cDA��%���T��,R��y�D�����-V��j0��Y�6Iצ�� �wRD-�k�V;y����7��j7�K�����Q�b�����Yi������Y�)� q��d�z�ٱ^_}�ռ��G��'�}-8��&
SwiR��ޏ�)%%BRT���hC
m���ưA����I�؈_���ggg��Y<x���;w�\9P]�ٖ���6K���r��zs���R'�\��^�z��?9y��X�\�2�÷`�`/x�ON���ś*?�W��믟={F�O�Ko�,�w8ϗ"B��EpCɔE�D�T��FJnu<�V�t�*46W8\�~ݡ�m^�~���k<��]f0��5M�Q|��C&�߾s������7R.H���	 W�����Н���q����c�J��C%�7�KP].W�@���-�C��B�cu�|���k�\.Hא�:���Lg)P܀��V�.�-���_�'3H7���Lu6R�gG��<���myN&�鿵@Ҳ&����>"�'9ib|��3����C �~�M:
��2X��v�H�v;C��#1:��v#F�Q(Do^�v#UjU�9S-˜ͧp���o!b!���~�ŉ�M�bl�]���ꌈZ���eK��N��i�tg^�U�24e�l�Vd]q6k6x�ѣG�/P�X��:�Z�u`ꐵmw�2�H����$��s�,�N�+��|�AӅ4^0��s�V���XZ[���'t�	��_���88G�n@&)!/�=N�{�_��88��l%ፅ�����[�h�-���5U�-d�G|�L�m�\��-�m��܌4񖔾��n����7��*�p<YZ�����~����������Rt-̟-�ɵE�EǦjc����	�#�Y��&WqP�d�{G糓)����A���']��δ�q�	�}<�mOd�󳧯<�i~�V	,���<u#O�:T��_��S�'i[լ�� J·�@��5`z5���@��t���w�:��BK�=|@W#��`����z��TIu�a�@{�o����'](�M_4���"C�,�B��J�	Q��8'��E]�[>���4֨�X&�5YO
����ED��	ܖ�i�"�̋��K�d|���k���`�_���Uu۹)�U���b
d:o!���˗lς��W�c�V�6�5�R�E����
���-JmFm�ss~~�����ݑ�1�wSV�Y�4lԬ�3���U+����v���K���ə���]�������[���(���BSƉ�mS%��;ّ#)��N��Pz���]�$u��
�X���hKЦ
����߱���7J��b�3��;&?�v����Q�4MU8L�I|*�S3�\��ƅ<���ec��g��!~/+�Լ,������d=��'l�N��`HF��v��#����:��ꖕ�)�k�j�Ě�Koˇ�˒XT����"�Q��Jo����$����΅o�Rn�x3��ng̕�Jw6}>�׺��phkY�h���ڸ����,�*T�Y0�
�/��u�d6��1��`�9r��&��yCت�l�_���1�����M�ӚI�����|�KE���tX��Xqp�bCZ7��"& �1F�l�����k��p���l�ħ,�r�k,i�<r��x��i�P̡ڼ$V#�{k@��c��J�4<n#u �&�����V�9�a��R�]�H�M�:+�(x@
�eg��uS��`��"sgq�����%A� ��.�SPk���Uj����`/�^�%�p��>E�������KV���e8�X+eoӮ=4%1�&�
]l�6�TO�����у­�M�UB4�@�w��ݓ'�2��5��L��05�k����n�F	�I*�Ƚ�n`�}nL�_S��t�������p�.�3]�Ds�5ς
H�sg�1^��[ț*��@p�adH���돠I��ѷV)eQ4oX9�ۛ2u�<�ta��7�')P�J�߸V�UmID�s�=#� -!�B�+�p:Bf�+H��ϡy�ܕ���D�ڸ`��j9��&��ggg</^��!���=���_�vw(�!��pή!Z��x_���j��~��>̭x�Y�^e,g6\�E����6��q�Zg���O	�dX�����aYXpj?�ϐ��:��@��l��Y�2��T����.���۷g��~��[likpQ��ؙ�8s�7|���2�=��a�kN��Ԑ/TZ���իW����9֌a�6ni|�4�.WnV��9u��9�.�ŧ>L���G�ٛ���ܘL؍r1�V\���G=�]�j�5t�VqJ�J��ޡ�g�L!�+M<�ZY����ڋU��Ot�Ck��qe}��5���L���@�a2�C��Um#O���a�_�|y|,���/g_|�K����.As||���S�-�5�;�.m�z�z�����7�Pd6�ӧO�<a��7_M�0��ɉ�~�O:~�PD����e�RТ!�kl�:],Z=�V&�!?�o�q��gݽ{�&��/�L�7Q-'��¯���t��'�������7�
!���r��AC�/X�������zYv���C��8�<;��J�&;�h/���f�CT�P}��
��g�<1�<Ԛ�s���$N#��؆ ��1�pp�5�w�%��="t��,�MWh�U�LR6�Q�&�l�V<Rmlv7�30A�����C��*�Tע+ ��!�Ԅ�u�P�6���"��������5y��H?G���j�j������O��(>Ŷ3L���x��Z��,"����F2ߚTFG��T_��IQ����f+A��60�����q�jRcʩJ�V
����>�뭵Y�1�����y�?��¿��U��u� f9���C=}�������"?��O�敽]<�bi˶c
/A�q���T>��6g�R��)Xa�7������"Im�"�����ǔ[�Øo�����Cg���ր,�����6ʶ���R��X,+�r�Wt[�V�,d>��2��W���-5l��	[�����]��!>��6D�G��ry���fo��c �"����E�W�i�ϐOl+�E�E���,"ɫ�z�z��1e�Rk�5�5�f5fj�6a�c��¨��'����V�˜P.W��<T��	�*���:Sd)z[)K`'%?�[�	y�,ͭĂ�g�k�,�#�r��qҗ�8�|:}G��lԵ�!����M3h����k���C�A�\y��fl�r�;p'u�P�Ui��28[w���$���oh����E�!�gt�!��V¿ih�F�����^h=4�)�������G���Q��'u_��^���z���}��Gc]ASS��L���"�n�W��M[��������Y�צ�`�<Wr�z�<F�;�	��g9Lﰬ�K��Bmsup%{ֱ�Q�{�ߊo9�w����K��X3})]q�I�E��(�"�����8/���X�B<K.$�Ix��t�0��T	�$<��d��q|0%:��'V�S�l�h��Dөx��F�c��I���-����;��P7��c҄[Τ�F�Lz��Kr����,mw#��0�(s7�>�ì�Q���Ю�^�&1���2Nc�Gm\���|dVH�8i8Ć�-�KK]J^�kZѭR���Ħ<���nV��x8:����:����l�n�W�	k95k-�2��u� R��������)���6R1�Z�@[}q�Յ�vZ:@5�&O;�lu�+B�K��`���LT��K�_��㈸~4�p�m��j]�8�@�-��9)�H��\0ܕ���=r�E"�B;Ue������67�0��z�{x�]wFy0��t1�׹~d����V�h�����q����|��h�΄�C���u�Z��rk�\�R-9���ѐ_����4�̦dl�9�ֈ�$|]�6v.�G�r0Qo(�s[�2�p�8O�?}٭���+�'}˖�K]�%��L�]/q,��ti/�^��چ>�l��K���@ˇٶ�Ǆ~��iC���y�H2E�]�,�/eP�֋���z�e��H၍cv71ˢ�ā�j������u��Ց� � ��Va�2�P�m���s)���u�H�j�ajeg�˕��v��R�]ϸ�ĔP`_C����x�L�1gDϛ�{��V����C��[��J����,�3,BK������T�PS���>�Wf�ο����/~��|˫W��"�
LO����z���K4Ё1f��iA�;�oa.�v��&���\�O}�3���Ψ����X>��/�81gi۞��Q	7a�Ze��@q=�P�y1\Y)d�V�0�$�a&z>�Q��L��c���w�����ӸG(PĖ7n�9���iƽ����br�|2�ۙJ����@RMʩm{��*���M���r�X��h��3������Zz蘼j�����Ѹ�V������+W��z$����b5J8*D��8�^GR���l��	��Nk��}*��2׎���~.I�6�ZEAT��ŋ;w�8�7��Q����V�DE�����8Ν�G���#����J����FQ56n���{x�j��MhT���޽{����������)���,IR�n�Ĳ�����~��p��Zge2�a�������x��uu�ڟ��GO�<�'qA�ۛ7'왕D��|���y���kPP�I)1SQ�����Ot��ūW���8����5n\�:�Lɓ�*7�.���֊ P��l�Z��6W�ٜU�L�!�������5�>�J7���
�o��'�Df���t����v㋋s�*�^="�>����Ƃܼu������F�C��pt��f�'>��vT �=�e�T��!o!$�Y�`�p;e�m�Q	��u��Z���K���Y��@Q���Nq���O�D�U�r�!*�nݺw�>�D9[j:W��L�7�*�9$��b�)3f+O�t[�@�{���:tZ��'i�V9�S����e]�d���P��_��_(�,� D���Ƒ��T��)��8��?����|�Y�V��X�/�߻�勧ϟ?	t{l,+�0_Ș��Y��K�%X�锵A�^.�d*qG%X�;ʹr%��姟~��'�����ܿ_ ��22b��c���h�TA~�rB��>n1+�Z�Z�t8��dk�k
3�~�he�s89�qåX�h�gvg)�~�:k����f����_-@�W@4Z1���S�e:k��^s���s%��I/�����3��~]-�d�R�.o���I�H�V�AXi���ۻΰ/d�(�\�aB�j���sb:��g��f�U�T�dH��}W��]���
կ����
���C�˲^�W��x��!>�9��
w���n�ǘi,����N���ui(7p��a?����7�^&[�P����gl�{G�x��OOj����aX����}�{�W
F	�.{��^SE栶��9�tG���3��(|���;?��;����H���at�+�PN�V!ʒb��L���&�@����.']�>������7���^�Qine�l��l��R����V�-�l����}�9�R�r1K���F����}O�Դ�$��b6/Wk�_��z�X���pJ�۔_�o�$������e�:� �K�YQ��򚦧gŢ�U���s�~����g��*�f��N)b�Ű�`�\#�m�Q�)��I3d���_Z�5�
s�o��H�e[p�)���ü�rI� �f�x,�׉$������i�-'VI��r\EG�_NK��n�Qݒ+|E���7���8������~�	J~����:�V��������oj�"�
���8�*�ߪ
�rd�k�d��[�5�ś�C���`.ّ&T����3��b������:�͸�8W̾w�U��RЇ�OI�|8� }/��V�2M6%�jYG�Pcz�C���Ϳ��;0����^&�?k5��D��M)��vI��&���þ�K`Y�q� "�}��.k�K�!�f�R��Ny[p�ES=�YJH��"4��'�4���	~-���^�Hj�̂J(NeMW����L;�<t/�-�ڛ�B8.�K���-���Q��Ld6i͹d�+5 �p��O�ܝ8��bI\=��p ��V��h��M��6jUݠ4��� ���u||�Yk�fK;͟f��4�NcX���f�U�|`����.���:�f}!�&|>_Q�TM՚`R��r�
>��ЎJO;x�ޛs't�3k���PJ��l��]D�c<օc�Z�"�i1�i͡Rz9�!3�����q�z�\�㛲�:	D�i��-�i�R����#����~�z��ŉ��T�J,߅鴠��>��+P9�V!����|:2��M�'�,i������73a��8��Ʀ-�6���+���x|z���M:>43зZ�w�>�5�)�u����l%��$�X�;��0Tv�R�g�K�Fݵ wwG���6���,i�+�=��^��^P�O�_�4��(jm��s�#m�O�]��U��ɪ�D��5�� ���������c��ͧg�q�I�I���e���S62�/�	���	8��Fs���u뜽�/?4nMu$bG9�m���x�0N�V;�a��7E��W
���z�����(�~�+?z��,E�a$��ݽk�bS4�$\N�2�}Z��vwE�W�
'$�W��,��ש�)qx�['v�&������U1֦ru%#�r%����m!eFNA�}(���/�fn�܁Iu"�{�wnʁ�;S��I6�(Z��,	�r��p�n@4j:��S��j)�[���PKs�Yg<�y��-���b���������߹s� NhQx!m�������p5���rYp'�$ل�ѿ�6|��aP,@��g�}���(��r0}�}Û��h����}�����o��w����E��*�e���G}��'���KN>�l�v�������,ȫ�7�|lU ��������k,�9�za.��~IoK(�"ҘM���(^=��Bi`x�o�}׎��N�N�A��v�����E����=��i��ÿ�:M�z;���H(F��6�v��s����a�ߕ��ak�db3F����cOw&�'O����8XF���[��+3#�j���O�'(W����8��%Z�&4g��[��g[��s}�Z��m�D�Ϗ�m =>)(γK� ��F��)��:�+hE�S���6��M�c�V<a���̩�����p����S�^�Z|/�����LB�mSc3%��{����f H���3y8sJYtϔn��/�ܛ���K��ZV�w�wϨ������޽{l�
[�@$��o�<3�Q���<��M6E�B�_�|����jx����x�ëY�	9+�a$'C���K���F�\��>��5b�f�6�4s�K���`�N���d���١P�1[���B����pl�_|��/1NI�������Mb�B�*�ٸ�����U����O������FX��m��a�M�}쑧�b"��J�"d��J2s�亂k�kMb��T �1q��m=������A�/��py�>��/���+���g�..��"���0t:�6X:9���n<���� ���UAnh�za~�k+.O#g�{�����6F��iؚ� �6}��������nX��2���JҸ�9П�@g�޼z%�"/����k�9���P��y� J�٫�~۽�D�8�����f���H��o�y���m
S��vѺ��~�����se'����j-^�p���B�cϒ�l�Px�D=�nk�)�0��nX�>��F}Yxlҝ��R*�ɵ�+!��n�A�RC���$�M5�f��1�Gk��n3�]j���\���5}����3D��WC7��V.���j�5Һ9wIu=�)��5z{̃pC�-v�bk�2?�Hk3ŹV��ۻ��)�n郱�ct"[����+������ߟ��~Y�Rj9�u�n7�I��/$Mכ)|�]���ڷ��V��>�N�[���*��ݻ?��qe�_��Wp�x�&�q����l�|�tE��~�,U��d��B�<�b�ܛ�U�'��������'1�3$fy�/�X?xj�aY�j����g���H������ٵ3�������c�X`)C�6�����	k�Xl:g*��jU4Y���'�;＃���~�����dBU����oҐ@��Z�D9������,�+�h3M��M��܁����9�[���T3J���<�V�yq����<�܅���:R�o��{ww���;�)����ʢ=k�MR�N�u�q��\�$�*�@� ��{KXHc���GT�vs�� 2� l�Y�
�G`t-7@��D�HgJ@Ud�NF�]-�j5����+����\f:��%>����^�����W��M*L��?�A��N��t���]�+��h��zm�=����Ս2���?ĽѲ�����\U,	pt�[T/��t��{,�1�:�y|&��ufN5�ڳ9gv:�����d��QD��OoҽM�v������ih���g�Y���[����/l�IbkjGbR�-�N�c�nz� ���%�t��C<�AYũ$��>TL\{rr�*7�x?պ�z�Ȳ�C������gp/<`5����{�=�@�͛�^w||rv���B��^{���Ê�:O���m����p�s�@*�g�����l���)��^Uz���iyS��u[�Խ�!�����!"tB[��y��0�f�Z�i��5:�N��.�
���vN�3X�˽�ƸY�q��D�����SW��A�g��wp��{0�
�n;��'�_���Eb��L�����>	(e�W�;p��Z;鰑Q$�Or�{Y�u��M�ZqO�`g���I����%������bU�f��_#i��G�2��ε.���j�S���E��%�4Χu�;3w��HD�L7"��v�L,9�3��`��ڵk7n����=���b`C�8k�����hXX�	����v�������˟� �ۂ���<��+�0�T�-����md�E/�.�{b8L+ӚP��F#E�HA�ǚ�b�F{#R�=*�0�ԡH�k���GxA'���������C?������g�Ë#��j0@⑧���PH1s���zX/�5�|���,�y�/��Ĝ�R�|�lO�y��IT����zt��������;�������o4����S~������X��+�F�Cq��kW������P�F���։N��U�X�b��|Q���$[��ۅy��rcߎ����n�P���?�Eh^�v�ĺ i� ��Kqޞ?�+�����}�7cza	��eB��a�!Vŉ ���^+(,�#)�����e��Mh�n����N���?�(���#�&���˗3N�a�#��V�����&�g�0{0�{2�+˳<��]W�%j9_  �c�@�Bm?�裏B-wb�o�m����Z�>�C�j)�x���C|˵�7�F�	��������#�s�ʑ�|�۷����4:�:��͛W�����g��Փ'O ���������$p��{[/�/���pU��NmIA��&���߿�������t�"|}x6<.GafFI����|�_f�[�b�#�G3�x:�TM������CW|��j��,�-�.q��.rW����M��n�AY���p�+!e��ry����b����s�����᫙�J�`1I$���~kh��hax{��]���Ӌ�/^C16R�`�$�/�����%	�D{,��}/)�\�!���46އ.U���r�Y�M��5���Rf�1C�$)	��x��Ň�Tj�J�*W�YS���ŵ���_"������������/�����?�u����$$�<w����0����\��(d��g��r��� =<<��G����^�m��mLuy����
��G�'��A�r�M֗���8����>�����z���7�ř�}���ձ"��;�kF�?���4���k���B�q[���{���0H�Hq�?y��� ;�u������9AEN�@��KX�T��)�^+@
�r?A�����t���}���5A�ٲra+�����7��_�ֵ5�ǣ��6B;ݝ�z�I�/��q��e	�`�NR����s����Q��z}�,��eU���T_���;	͚��]����8ד�{�k����N7�ꐅ,�[ٲ�'�h9�k����)Ԍ����C��|.�Cv�����Ϊ��L��9D>׬uxf�=?��t^�d��h�����b,2����K74gAnW/��ł���a��K��I��4�����Q�%��t��gqa�}a���W/<�IX`�c����*�G+[	�wg��Ե�%3�.Qg���M.km6�gZy�����qh����`�仹��?����9�*��Y3�!h�\8�������dD1״c&(�YfD��Hm"a�\��n����6A��u1G�\���%V�VXGz�!\,�Z��0��C�v���Ѝ�����e�r:�s���:�=�� ��r�.���G���!r�Zc6Qɏ@m,H��L1�^<�9�!��.�����R��,��Y�t�am�El��WU���wo�2�H�ѳ/��5V�I��������}Y(7VctN�����.�8>N��:�c��!xX��s�B؈N�L��^��0]gG�N��Yi�ph��3[2ߵ�}�s���Rcs�2�3��"��uVu���־��2wh,9�y��:PW��gQ�=O��M��S�Ji���sX1x��J�}�aBT�;̢
hK��:�E*�C�O�W����"��f�S��XF�8�4��ح��z����jnW���Diyi�'��,�IЩ��Y-�v숝�2�����Tsʩ�ƢB�O����իW�1�&!)���Q���M��)���Æ-h���{��=}�t��t��ك�)0��,Q]� B�b�ݻ��a�7	���O~���3~V/�4��$�:,�V���jA�0�����/^�����G��0e,����m��`��t=*�3z���:r��cY��W���;P�{�$Q�+�dzia�͓8؊c�4��jl<2�Br�3t�f��Rc�Ā���u d�s玎gY-:>�M=+��lS&F�RÑ��@6=��*�}����fL�7�X��V��w�>��:�u�S�vp�w���-������		�3����j�ܻk��Mج'�q��n�x��. xf�R�	-R�sA�4�����x�ۿ~��?Qu�y���
ea�7YTpә�-������'���[@i�0_*���Q:-�O2��l��\y� ʒWјD��!s��8渓�}B��WV#|��w���og�|��� A�z�&7n��ۿ�[|��ʞP
��$w ���lҁ���+��+M�����i�u�t=h޿�O'v�3��`ש��}��}��4|���D�駟j��&~a��^W��+t""�D�fF���D&���2���n�՞?;�Cb�V*�����ci�i����@�j��o/7p"~�)ڀ)i�M{7C�>��2���e��0�:p
?��7Z%(7����f��0�Z�w�Zޡr8bGp���ErO�J���:��`�/^1$!���}r�dgD��M"ʶ@����w,����2�H\|�m^|.������ݼy���@2Y�k���#�n�����_�{��|iO���
0s��W_~��_���b�����o߆e��#uf�|�������2�������w��=3�BޢD.�57෈h��R���Q�дтxښ�jl�:�qm����>?�{`��ӫ��bQ|$~Γ'O���b�b������D�e��bt�x3��2�.�0�b�0��z1_G���e� O�Q�;�ަ\���ݹ�
@��	8��o~c�{���G�5�6�#<p�� h��C�5,u ��~���dd:����Ǐ���K2����F=�e�
㻄S�����D<')�����Q�\�M��$]��2�Fw�;��#.�7C�-lĞM�D��/��裏(�C,W��� S� ��ݖ"�:��R��`u�@+I?PN�q�hއA��H�*:��-�2	����pkXOw��w��"��A�!�M��ؽ'�D"
�ɳ�t�p�\s�0�?��N��@�����N�X�VU���_�U�,����;�`I���2�0*�BC��{N����΁x
U���|�z�Q��F1�������� ~'��CW��$��~�?~��P�4I#�˖��_���GM�q���'��*�P']l��C�H��kR]�]H���K!�m��Q��c�70�7@���@=��ԉw����m�F	ï��/]%]2�ծ��K�_�Y$F��`n!k�Vf�dUP2�������Y�sf~�q�>�Ȳ���ɘj�7�a������k����jm|`���?5�Um��ʆ�U:�[� ~����P&V �Ehw��tG|/��)T�y�r�!����nU���E��J ���Z���y�:.ڮ�j=*f���H��]���=|��;����i�_E޺~(�[�@{��@�1��¢��&P�˃@MuI6��<1�`9�NSli��rZY\�	GJN��0���ɵ�rPn#G�i@|�p�%�3^��Z�.����S���0P�g�DZ�a�I�W�3X�l�zu:ڽ�jY����/�W� ��hH��f�O������ֿ��nG�e5?����D�_�c�Z��;_1W>Dl&M�ѫ�� ��D���sS��
T�f�4�㴇��|/ �l���@q~_0��d$csۜwR����a��=	�i����V�לE��+mMd|�Q������C�Z�i�|+CP.�1�}�E��[�JQ��ƭ�t�sH`ىwU6���Km�M�)9n'��d-�\�'v\Aj�AZ��%�L��9��a@��ٳ�w���|g*.
O��2C����o$F���Ts\!S�kk�������O�#�������T��M��x�"�\R ѝu����]EP�r)؆	���<��>nV/2G�]ۚ*���/�Pl,rv3\��(�4����2�'��Vkl)nS�k�ǀF�!=<}�U�[!��'x@��DG@�<����ZJ���g��V��b9C���?�����?�9�!,B�N��9�zM��44�(\�����#@���/_z���7;�0�t�0-~��祦ȅ
 {���7>鲬hG���j6�v�d�_�}�����ݿ#g��w�����(
f��FV�(=�Jp�� �؄���@[t'�,����2�<�
�W���B����^���ѕ[U�U��J6gY����/����9��xM�z�������K�P5AA=��\������V�4D���������څ6���^�듰�;]VMb9��nS����%F���+�`��5pe�H����*�14l5V2���R��s�Xa�j��[y���&hM0�KK����.=��Rr^�bҩB��벩�T�o��W0�C����I�=ugɓbf#��3ŧ�m����6��Ê�L[!o@}��ɢ��g�I��N�F"��N4��ki_Ԋ⦡�ᱲ+\L8<��,�w�������l9���/����۷q{��߹y���p<�Yl�������e�<�hs�}Z�NS ���&,��H���LI{x^���8�[�B�g���Dӂ=.����N'?�B:�f��n��+����!��ӓ�Y`��޽���{��	-���M�}��=���i�z<u��n8YX�5�fN�MNFc%�������2+_u����9�g^��k� z5�m��}�E�����xqO�{��~/ޘL�L�28g�- �9��:ý����$��gK&}�a�>�l��&\�6�2���g����M��Ӣ;,�`�^�y��7d��#���%Jا���$B̲!��;��Y���=��ѱ�Hj`�i�.��#b�y3k#3a���a�.?�VsC�hZS~Xj�Ǩ��E�ሸǽ�:0<�		�F�y���������;ׯ�����A:ٯ�8�r���{ׯ_��zIݼ�~H,��|��G�G�Ù��|�3��tI���1-+��G�6��,�q��aJ���FOx^xV�*x����RJ�f]{�wdy��ȍ{��8��.<4���o�4�*O�C�j�:�\�b�53��b�ɇb�;�����D	XO�Ij�x���-/^��8\���l�Gj>K�f?b~H)�4�z� ?���������s�N�u�]m[y��9�����>��D��������7�\	�,�Z��|��_���"\�7���b٧�y�i��fW��CY��m�M�0��!��T��ī�Q����޽#�������f���з��gϟ~����ƣ��r]�H��\�����Y�����`.a��� �T����[�\U��?P�	��I�9�H&fb��2�4*_Բ��]("�պT��e��a$4C�^�+�<6�\��M���a�7��E�Y��7�O����Y���z�A��.��˽�D�X�P�>��E�������ܸ}�O���r�3rv|���_��o�>�M^��U�lT������U�8k���
��H�D$����ZI�j���C2��=Q���Y�)�R��Cv?�آ$�s�ݽ�ի�Z�0
�i.غ"]�#��ײ�C#�!Ϣ�f�KIn���\㱚�@3� �dg��P$���[L(�A�p�kX�{]�2��^��$}j_��n���M`%���=�H�n}�t�p��&z�)�K�P�u���ϗ'��Mj�à�c�fի���H����޺_�-��-Oh'�$ib#V<�w�����8!�
�A���7�g�=�mqo5F��h�����d���իW�p�&�ȵ�op0p�<x�h�ZCI�5�3&X�7�#�u[���m
[��N��2��]{��"In���S���!g��^��;�@���ĉ�+���"�mh|<�8y��-�L+��nf�lgf�dX	l gs��-���[��ĝ�$R�ސq�2��II�.czN$Q�5I-k�J�Z�𐰿?q�e�i{�v��\p#�pw�����^6�!73it�
��ɧteܟV�U��8���[i�+A��t�O<��
�lod1K��q��p�C�(bc+R-�q�p���JK6mhF��G	3Y���y+P��`F��c�i��N��Lмk>;!	��8�Ru�T r��ۀ�u��P�P�����h�!"��xl+�|k�(����[N��J̰X��'�j�+IQd ��xg�/�l9�������Mm�� ��Z��S)���&c�J���<a2�����j5����&5 ��J�`��v�k��9�h��AuD
E�ye���7H��s�s�26���/otA`/����! xdhQ҃��	�|x��.eV ͌����6u#��rk��%�<<��؍���G��n���]�J/$�lP$�"�� X�Md�*8�K�h�o��o>��3���gt�H�Gz�J�v$qAjګU*j ����YA������-ڛ&�@� ���n�͸@���`)�D&H��,K�vpu�w���ݻ�zB�O�=q�P@Ā,fM�&I�A���41-�1Q/BP	�� ���+|:�>�@��]�t9ĮU�`�*QZ�3��>e��#M���E�P��M?��K�Y?;t$�ׇ���M���AS�NI�~�@�y{"$O7�\��d��'7d���Ěj��h�HR6F'�ٌ&� �S��x�8lM�sρ�<��������N��/�C#�^���38SK����AM:����qj���:�0Ҁ��̈́T���2���OC;_?��T�k��m��v����������>������Kňͯ^���;��ɟ�	!��S���dM�!'� Ϲ8�ǒ���������||kh�+B�Ùi���#���;#�j�����.�$�[�Gt�ꑪ�'�2 t���Z;�J�gT#\Uh���D2CZ��o��F�46��^ž���u���l1��466��LÌ,�˺��d�6QA��޳㌹H
C�X�"�%jz�9"�%�ϒYؕ�Dٓ�*����#����Nx_�����ӧO����VY:*d`�i6�9M]� �7�?������c���6��2��Z$F��[�ŉ+_l(��RFv�����������;�oF�(��&�$l�mHx�B�K�V���8�13D<���Ç�|��M�'&�D���M�H�F�rmćD�����EX�ꍉ21�f��=���+ʯ�'�c�l;�pe�q{��v�:^es����_�xo��o'&�vd�緔aY��#�����&Zy2���6Fl���\yW��4�
7B��hU��-2�t��ԙ��>�SV[�
U4o��j�趸)�V�Bܭ��*�x�'��7��М�o�&==�]�W*�|��}�����%Q{?��O�ON�_��w�c�������㡮b̒� P. K����	FZ�Sag���B�a\"��H�2����c�V�_�9�%�⮻�#]�b��66�;�����;O�f����_��W2g�wp7n�	)�{�G�F��~A|�.3�|���c�ɍ$��x�*T����㋼XlP6�C��Hln���P�@}p���2�!�c��iC�?����c}�x!�2*���[5L���J�#���&��:��-���N�}�ŕ�zk|E�0�۳g��!�*�_�c���VHPk̞��6X�
�(�ѷ�c�{�1���O�U��0�)	��7%c�����ГW�^KsXM)�tF%��h-M���7j��`<{�4iH��$���S^��]@��Z��T[��ݲhC��H���(:������p��D�*P�k�Ȍ涵VkU���������77����v��[sqm܈��q*��7�PO>��px�R�~bnؿ��J�-��{k���V�o�?Չ�& 5�D�àR����y���5Y�ƿ�>��yy9�!�����F�Yk�+�����\�� q�Sx[����G��/	���eD��P���r6�70�&���BM��p���z�G��0a�ѓ�M�ZV;�i�l����|�6�j\�� ���aS��pW��(4<��bN����)�ްI�g\v��E��lX]q�qeA�h|�3������i?T"gh(�a1(;��H!�PG��#m]�@�Ah�%|鉐_}@���E���'xQq�*��y=H��.�m#�,3��\Vi�B�6E�цTY��O��Y5�ۮ��hP�[��0[$��'g���kb�\�C��� iwX�uői��%���A�
M�>������?����q�㫿�+�r聍G��1��L��8�M2
R��Z`z<�<nzf�n�Ѓ�J_�W+ڏ��];��c���(�&�*1��0���~��8!��^��-Q��+ �,�
�!�QIM�g�6� �Kf�(���Fi�Gh��Id��[�׍�:�|�|��e%I�捍H�?�޴ٶ+������nߨo�*�"
�E�;��?}�/���"0�(!�J*�������4�_�G昙g	���r���k�5g�lG��9��Բ���[`��Lň����! P��q
<�&p�����C5�c�v���1h��o���7	�Y3�.�����|�Z�T-�a������2��׿&�^1)��Xq�,K�A�F�QU2�3�Wbs��:��")GhJN`�P}�B�Hh�F!=q+�b?����X��WbpT)�%�y��pL�&izJk�M#E`NȰ�H�.���t ���V��j��ɳ�r���!+��lqr�%i��w��PI���z]�4��t�XV�>����Yequ���A��z8~r~�}���m�}��L�=�V!2{���HV
��-�,BS��8�k'����)3��$�k�����;� J�Qs�$�ցA�M`}���EC�R1gp��u�X�)ní7�~��_������X̘�BH��h~4p��T)ڬ�d��Xl��p��~��:+����9f�U��h��芴F����A0�jWu땿����	�ݕM���>0�GLReI�������������;���(�z�������<̈́�!��^C)X��i��R_7"���d�0]2:c�1���qu"Ǵܼ���ڤ��x�܍���pO8U*�\�4ϟ={����'O7W���V�؋��U���_��0V�x����P���)��O�-�,B�Q�dS:iU.��K��������x3g�~/�/m�8�q����@�\���=t/�'����Ӡ0��JN���i�_nL�	[���8]_$CW	]n"�����)�B ?h*vPpϧ��8
��A=:��$)�n9��ݖ^J:j�W�ߊ�	2CIk
�9��O���K;��TFE+{�G}T����E* �OEC�%u�}���T�X��R3V�ڣ;��1a��^r�DV5X�X��3%��c��0͆؂0 �鱮y��g���ŋW�M<z���O?��/./���v��_�j�(ݪB��=ǌ391�\�>I��P�	Ҫ�Y`#+n�cݴdN'���`��t���|erDB4:c�)B,ȓ'�H,�?�56����H�	��:e���&���x��.�?��q3����jKMȘ���b$���&W�F�`x������6,c.�}��_*�gF�̤-ϯ����E��Ɲ���������M�̎�:�C�/2Զ�b:�1$A8.qx5R#,_������?� ��'O�����������NON�1@�rr���4Hu���d���=d�{�<r����*ICօC��^x���H �DVYa�Th�6�L��V�@ū���r��n�����M�n;y/�S�>D��/C�I��$h���gF%2/{�ݼ������n#��_����~�գ���/�ow>_u�C�����$�4 z]��ިG���t��2�u��@��dVW%������c�6�/֐p"�4M.:�(g	B�!��c�v:����Z��ryzv�<<�LR������qōB��ѱ �qN��?����o�gp���o>���A>��_�Ƶ�P+�tjl�b��}����!�Xy&1��qp�41q=��UO�)�"5?�U�7_}���z���!��ZA�:�yhd��r�W�b�'��#�qU�1�@@z`w"�U�&��'09��{�F-�y��F4��j��6�u�����K׹��J�F|1��L,G.�Ġ4���d�6�ƅGm�-�j6:��~&U��^: !W���� fr�����s6=j�������&�+3���G������\���x�����4���~ѵM��[��*I���cZ0zoq<S26��Ce�׬IT·=~���x�K����4��1�RQ[Þ`,�����W��Hä9�;Z&�I����L�_�͟�L"3m�$7{�&�5�h���֝�h6�v!L�1�e�q���o�	A~��kq��6sDϗ?Hn�W�!(5��� o�vS�}���:M*������4L����	@�pz�329:Z�F����5"[n.#v�\�	�<z]Qs�	޹캆�3~��kS����*qS����Wv����	C2
�#6z�[��'r��ïh�:#�'{=O_��J�?z��\�H4����4'͛�I�v��[wg˰S�`��������~X�Q���t���7�h�Q~��6�Ǌ���>�Rt�pٻw�rS��%>U���� �9�:*ZRx�0;��0��x��poZ��#�W��8�a6K��(6!>r�@������%�c*��4
���VG��n����w�I��<Z0<rkc�"ԕ��(�-r�zށ�9��e�#(QX�.�m���+Gm��c�<K/�
�#�= j��Nx�/^`�؜��$Y2��o���Gjrv�&Zy�(E��a�A�L�a�A>5�R�,=����#F���x��?�X#��rz8��iI9���LaZ-Q(4�'�@�=V�"���i����ϟ�5��'7Z:�U�0�M��N8
� N<���8%�8_��R�o��kyC��ԟT<�r}k6�$i$�����q)� <f��O��/��_���^�|�;X���ע��C7E-q8c�ZQc8k1(�����;\@���V��i��V�q���5�x��'m���jM=��e���:F/4I�bY�:��j �է���|.�R�m`��X��l��{b���V�砞 9@U���J��el_P��^�������D�B\w���3Ȍ�PwF;�'5��i�Ƞ�В�ɢB�.�o�l�����0��aDZͰ�[�J�h�4�����4�4��O��`f:!��I�|�m|�6�>ڤ�KV���ل��%����N��{�������W�.9+��:���섵��vmdR�>�����D��s����>��<\���T��_qc��D1�IV1GO��Oie�V�$��%�ѕNqc��9�=U�Kc*`J1�%Ā�c��ȸݞ��	#8�L���;������+{�D�P��{u}��LS�_��
^%ʙ����cm8����LP2��\�����l���8��AMa�B�ྮHpF?�wN�D������أ�d�'Mm�"�d���7�˝��QW�������x�7���C۳��ʠ����/!{�������}��[����~O��k�f�������,Q���ܚ�N�J��[�fm�p�!`��F�
��N;7|T_��K%�ꎍ�t�!�nV���NՠŤ)a�֧V�?�i����׽a�XT�Hs]#�Y)a����E w���ɂ�@����)���F�QB�7z�����\�A��s�G�{Y��G�++��1�^�Bz��ݒ�!h��6�N�
k�O�S<���wh�I����Ѝ�|�7�x��w�%��#�%�̀�l���{��C��?���%]N}0�˳�[��<�<Jc=�D�k�u��_-��v�g�g����S}�-���d�}Y�T��
�M���xjb�ܼi�@m��p^�z�O��Oy��m�r�#���:�(�c#�����~��Yu d�Sw ۏ=�n�N�]���P�m�,��K�$�Rׄ70��hU�u��pM�,N�8?�L~��o��������,78�37\c��0J/$�5dr����s5�F\�bM��U��Q
އȠ�7�H��gF��������,��7���x�!⦇Q�2/���7~U�L f}�w�%s\�Z��$�U�V�3�Uß�cenj,\(���OT��$�������M��ܜ�1�Na9�i��	.�rD�������)*����%�=��8����P0!�V�k/3(�;و��}\U(� Mc�Ugb:�)9����8�V;������k"lp�]ǹ�qf�0_�����>:��HUC���Y����IR����g�m>�p!gĠ�7p�Yޤsoh��Q�i��2��u��Ua�"�bHbcL=�y��Q�L)]2CsY ]����E�����ւf�Ot$Of4�/P�Q�L�baC�
�fUO
�TΒ0��<?�s�;-��pZH�����9C��+�Mq�X�ẏ΀��!h4"�{-]�&[k{��Na}�yу�ͳ=�>.��J�GG�5�z�#��TOK�1t� �8����2�<W���u��ѿ�}���K8;U؜���#��Ez�o&�BM1�/���yl�k�|(�BDRN��^�S	�[�kȵ�w�йXs�o��W�,��
*�)oLE�E��ʆ}3*\�'˳3X���������R��u��-��-E�1��}/R���+W���Y�6��>3�Ɔ��u��Ia�7�m��ީ�8c�����Oz��-c�Lu��K�1��""�$A�ɀ�v>P���8�&�u�b&�C��U~�7n�����ʾ�-'�5m0�P��s�<��a$�����'�p�=���i*I.J:K���&di�e�|v2On�X	6�2�+;�s��ķʦ�f����؎V�_��d
wsR(��BYe��g*��	J�l�c��y���1wD���W��3� 1��Y`ʘ�K��I���6)�� 0g����d�����L���b]�bL�ߕ*(%g�����������	U@��|����aj�� q(���"�A�e�b�ɠHW� I��<�+y��`?x��jM�O:�R9���:!�i�Ĺ#'Uc���s��[o��k"���R�X�c�k%�BV�Gs��z�'���-n����]��#�eJ���%��t0��8	�e���n>|���G����(͊}%�<y���d���Q�\]m�Di����S�ٺ>���0�E��ϐd2o/MLK�^�z��}�OC�?hT��3���w���-��A�'�Q"�yS��	�Y��i**4�ژ�M�R/l�#[���n;�����"��j�ސĖ�Ĕ�����< �ww� Q�di!Onm@�����O>����8�������ފ��M(�^p���+���_�|������I߉b��!�%9)]�D���5��$�M9���<�Y�sR�1s��8u��6�^�wO���"'Wb��|TE�.�&��o��zCZ�!����o���.�W�i&[��]�����t��+9�u�ݼy[�5����gV�e��TZBw��;'�)�>�ΡJ�ϯ<�3����^�\��}��oV���ϟ�|!X���x	�P.�]SE���X"?;����e�m��|�[,�%i�L(��$��k{l��JO0�`�9��g���Vo~�{��yL5a���Ѥҩ+�����}f��<��3R:�.y��7���*Og3'�x@�)}lO�9�ŃIj6�� ���&��s���Ӆ�Ǧ6�U�\V���_Axɖu)��6��[�1�������_A�޹{K[�+��N���G,�2�3�<2�-�T_\�i~'?�?����?���#mMH.������n�v'��J�G3���q��G�$�����7,���)�ϳ��_}���]��mS�e�8������ى�r�xFF
�c�.f�Y$cu!X����DiJ����O��B�����6����rW�l�NS�ئR������k��,¼���U�� 4q]�$���*��ݺs�Qz��i���Y$;a��iܨ`5�����փ\w�b�V媪5T�'��i�?�|G=-�>���ݻ��|�������,cG�l�)g�zs2`�;�sC�;�DD����Ţ�h�K���2cz����"h˭����DH��O�U;�,�[�cg?|u�
b�ʽ�.;��K�&��'��r|=|���即�����9?�Oqe�*��xi��哑�[��(�����w���񯷤��_\\�,�6�S�wZL���)J�] D3�=1@=uG���;qwO�C�<<��v���=y��ѣG��6o���#w�F�CAD&ڿ�.���p��K�(�=� 7�Jb�,���r���>:2�  ��IDAT=�����~���������7�����sr��V��l��;&���G�C��)r��G۫�t���j�*՜y$g������@�S�O�F�hF�"h ���{��ޱ�s�J���%S����U'�B��z9�� ��Y. �z��Ɖ�`̻�Tm�ȍ�<�&�F��8ٚE��P���z���A��ۄ_ȇ;C\��Po�r�clzI��5�͆F��$�#aDi�b|�̠j����v����Aug�������`l_���g�\���8ɄΥ~�q#�X�P7"It���P�e�\�.}�<dMlZa���c��J��b)�_Z}��y�Uoe�Tf8L�Osk�(�dƲK��S`0A����S0�����#����O��Ӹȇ~�{x��)���hί���]`ZM���t�2��'�M.�)I�@��f��OI���b�wӣ�[��#���:�UL�q1�;|�A����)�����0\Or���O�og��J#}t� �����]/�\��F����YHB�et��~u4j��F&߉��c�KG�@M��L��ւ���]��5�Y1;FF9E�-�
!HJ�LN�0ީM����v�f�_a{+ͱ�^����өVnqM����Ʀ��b���^�k"�T6C<���#���Mv��n<c>���箁3��>�Ryr~~�7r�,�`���jn�
m�s|�!�e<S��� �&q֌j�l�s$M�i��;���Yl��	¢[��^�Ф�
���o<���@rG?a7uw�<����|��3&
���M�li�&��pXDj,{L���\s�����%�6�bl�Ȧ�н A��b慊`��^C�lk	��r{rrĵe��ڏ���FT�;ؠX������C����CN�LA��K�	���<�^�w�9.�Z�q�Y� ?��e�Y9��$�������ү<�Gp�n�B�h��U^�|�=LSϿ|qɭ���²CrQ�y3Ÿ��[K�|۠ݩCl����Rp.���de����@�C:j;�5�]b̏Hx�s<+)إ{:�DfB�z��.�cqO��̐��ơR�O.:�Q&+Bt����IB��tU�>��a�an�5)'���/�U���%�KjS���������[�����X�yd1��L�]i.�Vݯѥ�x�Si`�4&�8�����&���U@�E��`��j�U��`��J/�*|<�N�g������������XO��*jr|���f�;����wf�Wӏz��Rϖ}岒x�'-�p�EW�XL� ���� T����9C��q5H�L��l�RY�ꭚ��@T#��q�A�,ƈ���N���:����x��[N'>��-N44ǧ'4�B �G�Yz��}�ׁ��X|�be�f����"/�Í��7'Q��*q,�N�_
��ʭ;����F{��^����	5�g(�?�O�cPh�Q�݀��޽pa~cn�V"iY����Z�2F䃏 7�J� >��$n X��2�J?J�Ql�w<Wcl�]�Vr�
�m�;J��px~�Rd��;O�����#0��^xjZ�1�%��ݺuK�O$}	��`\�_@V����B��P�9v�z���K���.�Y�b^�����������s���bϠ�g9��|�IQ&$�HuT�6F�TA�%DC/���\}�ͷ�=j�?)menSwE��~��x���V��;��&�Gnkς���,%��l��?̜g=�����v$7\�� ���m�ƚ7��qjCc/�7��ĳ�Y�%o��C�j�F��8���;1R�t�㑬�a����J�p��[�{�?��?����y�����ќ��^\���NF�u��=�iL�9kn"�a��3��Ϡ�Px�O?���%
!&�<�N�Iܕ|o�	�ϳ�5��\o��F9�rVe���P�P�8aO�� �]��fs�%���f+�8�|F�e���/�K�&)�(��G4LG`o�?�GA�ЍH�]�Ï�$����o�
�g���Wunv[��t�<Cg���d#�<E4��L�e�!R�A]O��2?��״~���˿���~���(���/Ne�$���y��6T�3L��
�Vǔ���M��s3��NMM�������^l�V�5+w�Sa�/"��$Rf��4{���ӳ���Ͽ��7��4���Rϛ�yzquq�4B���RC&�|���j�)l�k���籪���P�2�R�^�	ec=b(?�F�kn�E�TI�]�Z�.llXp:�oЍ�l
�ɿ���Z�>-�`L.���F�?��ɏi��[,��aRbzݧkƙވ��fW�T^������K]�����5��Ӛ��e�/F`IB	i�}��big�ũM�vm=���J$�@�ȏx~����s?9��t#�|LF�TG���`b)��3�H��G�qrʐ/X���M�qK�w���k�Yg(͞e���`~�_�`�0�j�fg�x��Ll�odbWl����ߌ ��}(qe�BK�u���?J��)3 �}�U}�����b�g���BjA�;+Ld�_���N��DS�9�w����cǎ�����ݤ����̰9\QؤI�f��,��`�K�v\�H��9��&���G&��\\�o��J�wY
L���R�����˞S�c��b�)zZL�rH4��t�����d�b ��6�6"s!eͳ�\�B�*Ҡ�6�]:r;Rё�?��	�<�z��NKs�+��Y݁�x֞�eb��Ad7Op}p5��j�~q���rB&�� �Ǔ7���	.�����c.U֕�5 �gggx��ߦ�+��� �	+����/����[W�դ�ļ.��]p�ln8]ҍ��A��b>�i�t�kel	�b�_A��~���Tic����P����q��ۙ���f�Vh�j-uH��=R9S\Y
��!��ɓ'���V#������J�nP�%�>4E.'��3!$"����׉��]`������JF�<==�T���{��!�C؞X�ǉ`��v��ތ���w�>�n[��jc��C��v�b-�'"O>�w*��1X ��0�*�M�E^��ͳUWKo�.<yx�y������Cߴ�M]1%�c�x�t��r	����M�o����hq����4Z��u=�۝������{����/����~��f�Em��༤9Nټ)�C#���I>Y1$�"�*��s���t>;9;]ǩ�����T�*,�'��R9�5aN� j+��-�}��&r����{,�p#xj����g�����$�^����OO��}�����!��I�0�o�\�N�Ya�^to'�Pϫ%Q�ص'aA�i��!W$�'me��2z�����ֽ�c�^�G��y� ��2]��۪���LB�̩N�t��[�����1��+����ʣ�N�������[7d
u�S:61����X�î>l���<1Rl�VT,x����l�9�fe�E/ھ�ޝ��L$zk�{�>�k��a�U��iO��x�������g_�z���8bx�Ǐ�/�"�cc����4��������ಳH��Vqv!�@��"h�c��`��|��ʭ�Ń�ޠ��5g>��JŽ���V��QQn�h5Fu�̽��"uTG�P�$����%���H�c�es�!$��"��+�v�3N���],���z���)�C�w(��i"6�١��9�b�k�O����c4Ɍ H�=+g��Z�k��>z�h���_q�
Ց�ԍ�;�n�J���$�F���Xzk�g�V� ��X����/����"�R�2���|�	�d�!����(O&��y!J"�
�����yĳx*ٳ?^����_�����N��RZ�4?�I���=w�f}�p��ړ��X\�Y��M^��_<O�$K!H�2��CRWCu��e�l�N� u������i�Ӊ�Q>X��tjy9a���?V%ٴ%��L�Jҳ*�F4�؀�`=F10L4L��~����#�!���D,¡���-tJk�E~7�3#���(]��o�7<99��fW��IIt�W�2���<���� ���2�E�H���1��F��+V r����a9��C5��Y��Փ��'eZU�n5�N�n/�)d��i�}��<��T�#��z�ѐY�7n!T��їRh,�G,�	ұ����؋���!T�����1AQ�4H
�g��v�8��D,�j_ׯ..��~#��_Igt��ֹ
b9�N앇���\�NK%(���;��ZU�;��rMAdU3)$�o�v蓦��]#��捦k�"��Xm�|���_���C#zR�Q�&Y��lz#�I�M�Q�'y�Eqq�n��#�'�,�xБ��6����j
��J�Y;��5�|W���-l��^�g�W��(m��Z�Ժ���j[st��q&on䃇oS�SE�Yoi,�UC��$�v�z�n���k�;Ꟃt_���d�Q�eX&�=0ͬ�M[�C�@|Gf<��3BW��wQ�"I�^���\ͫ��g���FǨ���:���g	���Wˬ!7X��z�S���k�`���"�h>��6)�V���*Lm���]
ĸ�`D��~5�M���H�r�z����&�d 0(z�q��2�lMy=�81J#��F�e¢Fv7��J�`�
�	y���t�>t��]���Y10����x\#@qj4��R���3��oWU�?��M��#s����\�8,5�/�*8mk���^+��7���q{A˶x[�4%�)�����j%-��M]�ܦz���Y�M "~pW�3�\�%V��Nn1��� ��
ꑍN�g�E���$8m?g�zv���tn�;����e��?����ŋ���}��)����:^ "���3���������=Z.-��)��#,�G��7�|��f|�
Lg[A�5�?DS^"K4����$��ND�.��w����/	�������/��r�������)%�7�S�C3j3e���<x�G��/(E��+/~p�>�G���#\�q�`EU�1����Ը<$��tVr���u14e��Jx��#��Mt	{N�.%UY����������u�[�i���%9��!���T4:Ld3�X���"�W����$�3SNSH�'��j~&�6K�q$B�-��@o���зZ_:�=?� �7��qC���/_�a�zƺuB��&UJ�kD���@W�2����ۻ�K�1�v�´|�fl�6�0�$3K���C��::�+��4s��P�|��zsE�'^�{��!ݸ��p��qF����֊�W>)��+�]�� ��<��'O�?�%OBJ��-G��kf��Ŏ36\M]AE�c�[�ZU�38=�j��k�R����d3JZ��o�"�}���$�{^2�B%�ۈ�zP����w����c6!)��7WC<�F�$��u��MyȑYL�\��O�;Q��T�&:�j�L�[�6Į*�p��bq�1�A�r�	�1�F�H�Urg �HFi����8��[���H�)��R�5�L�\��b)���3��}��/e���oScK:Xg��uhQ���o��5�aQ
.>	%78���U-�G,Q>{�>��o�����H�X\���N�;;;0Q��:1����
�b��gy��>$�6W&��M���P(���TJ2\��R#�5cZG`�Z�ɋT�\��껐�L뾲�2y)��œ�1	U���J�ǋ�^���Yj��S�3�*^h-�'t�j��O�V��	�x���|�W��|�Ab�ؤ������Ԑ����'���W`�~�����_��0�x�����fNE�t��^xxi�����S>'6��Z�'��&㌹7�06��{���b[.M'S`txz�s��K��6^��F�A���Y��z�;ݹ�d���)�5�0��d=,lg�;�1P���]�I���Lǡ�z=�/;��|�m�L�Vz&�����r
�.!����S�U�Y��Ł�Ȳ��}��5�R8©������\@��\�4����!�K�xܺ�x_�gAW)�"Ž����!�2V�LZ�>�+�@]�	H���q�I��ʫ�Z�R+$�2,-H��[�����P�VԤw��]��@�d�F�OG����	�h�,�Ji=���=�l�Efì��\{:c�,B�Q!cR]����Y	�v-f�)�)��ț�D�8Ϫ�	��R.W��<��LA�̙���w��MAj>��S�!ӜQw�`��r*g.]P2!Ƚ�Y��l�#�4�Y��D�9���gH�T�;X�;3(	�����ذr?Ȭ�m���u�Qb�r�����A�H����i_Ydd�#�On��y$d�3�M�e`���%�����6���`H=���HW�
]�,����Kv�H�9�R�HK��/o޾AYe�O�@ƗԵ�Jl�q��C��t6,��RS�!!|���w�O��T8�8ݨ����u�z5���`���p��YE�U��4���kڗ$��]�|~/KDʳ,
�� ކP��n(�y$��a��h�f�}'�Cڕ����o�ݾ~�UȊ�R�WO;F��tCs���0d�'Q�ӄ���+�U�f��n�@�!I ��������8�,�F](���+��'�1+ÿ�����p�g>,M��������}�;Øx�����e����K�dĹf5A�j�&�q)G�1����6j��hn��G���"��V(}T�㪰:��i�\�a�M���&���7�o�
�(�;칀m�Y_5��P0|~�|^��!\�:_,��`')�B؂zfc&���年+�K�(-W��&Hl:<xY���5��k.�g�T\
	��>�<cuh�
��Y���P���aȒ�<�B�TyV�w����:Q
��;＇0�=X��SQ~��O"�||�P/]��G��sQ5izyuurv����˵����D�n�I7�8x�̲K҂�+j�s����f����5-�g�<��d��ʥ+a`�d��8�]�����/�]V*�(ը�S����*�ne�% 1=;���N�(�C�N���/O�z/J��v��*�Lz���v�S�0ʼu�vk�Gs�����ӌ�;�rBw<HÅru*��[��/^>��ݦW�\�`c��.�L��$���'w��f"x��t��R�	��0�7o��������v� 9�QO�?Xx,��N)��� 7��Y�^��ʰ���p�$��q�'��1���a��NZLgG���R�G�����
�r���E����fB� F�He�(9#����,�æ+��g?����Dl��}�&��Ƨ��I�ޓ��c?]�*˧8����O�-����/t�'����[k���
��p|tTN#���B )�<�8v/N�ٍq�E[���2/�Ά�Z�찰� ��,��5n ��F�.���j�&E*�bGsH� ����=��:�j}Yd�)	"��D���?���Lh%�
�t6��j����:
�a6+k)�&�\𒢬���i�+���l�L��8��M&�"��h�Z����6��Np������;usX�/��Y�2���-�W�I�WW{���&�g'D=dC���f����Օ�CX8�9hj�6��&�n�5�|I[C<�v���`�����z~D�r���ݻ�t+��{��v���4,ǈ���w�>n.�C�8*�}��T��8;æ|�N��;＃Oў�'ӷ��7�n&Z�
�$�r��r6Z�CZf%<�LSw�/���j�<� �����<;�{��r>�~�:�������̷n�JtԱ�:-o���i2�ϒ�g턀A��%V�ɩL�;[_mptpϸ���n����P2�x���,j(�^�A�p���9�yzr�&�����F��W��v�۫�"�fY���I<h�w�ZB�:Y_�ˤX_�~�\�J���B�E)�-8��p�m$�i>/gG��#1�C�+��b1E�,�Ɲ$�'X�����VM��諸/�y{�1�K8fY^ɤ{1����:����9GRY�+/�VX��j�.T�AԤ�i�����uu9S2u�j�r^@���|��XA�}���8�!e�[K�;?��$췻�W�/.�����/}EI���K�B�BP���]BE�>99��|Β$��x������?�7_}�h��A9/�3����d��t����s(�5-Md���a��#(�8�}�ݾb����SCF�3�9�`-{Gs�P�JZy%UO7�0D^AoĚl���&�^���T'$:���l:�g�ͦb��r��U+�!v�t�h
X��	\�B�z11E���⏵�ዣ�i�u�a���QmВ�Bas�� ���pvv3F���l���m^�y#خ��b��w��/�D�Vk�;Rr�D�F�TF몣��\����o߼qK��4I���n���?x>�ӟ������/����D���9�V���}�l���w�ߕM#ۄ塴L�k�n5K�ɦ�:�$YZ�M��� �ſ�aO�������뫁$�=��I�����p2��y�f�:>=�JT�Pi�bO��A+p�����ie�0��F�p���ڧ�=�R�>���R�C(l_�X�*j�r�TH�!ThYO���}+~�|�EV1�[�
�P���v�ryLp
�x'��z�̋�fV2O��^0�G�Š��zd����/X�#�-�L�2瞦��]����e��a�͉%�"Q�A��VRe�~��3%Lj���udR*��	�X>Q�o�r����}����ݻ^7����P*���`�g+���I���蚱�#x��B!C��Ӊg��90;���2.K�c�'%����髍�@��	9O��V*5���6�����\�r�e�'�&�(�Y�+�=��'D$>������Tnl�p��#)D��n���:)'��F���;��=Nv�,p �$O9�k��уo&�i��+Ѵ��� �u 4t*TDJQYR�����i��7��y�T}5[H���j���
xLp�a���fS�}���pe��� �>��<]�����[/oݾs���g�����(5�b�a���uv(t�C%��T�v{%���}�byC�p 5���l+�3��j�9v?0���O�I��l2Ǔ������s,A� �o"U[���	
 _��K<�j��O�w!C�Օ��d��z��/fy�?�9@��0j��$&��z��VK_Ő�n*o�Dǡ�ws�!ĳ��/�����f��ڼx�j��>&P��:�h!�s���-gg���P�QV̨z�f�*�/iuM���>�@$���wu�� _|2�.�D���	@���n����;��b���a>��R�K3�uŗ�c꺰���(�ա%����`5�[� MB�-�W��v����� IϬ�r��¡�)��A'�>�	��\�"h�,M 
��OI���<���3��n�G�c6ˤ\*D��L��@$�-�@���uq�ײ�M^�?� �Y��с4���!�#P���;*O[Ed���y��=�I<�N������h0:^����P���<K�OG:�1�F��6]�W#��c���$tb����ֈZǱ!�炕X��u�|�A�F�.K��7"a�i��f�x;\�#G����L'#�:�Z�mFD*y�g�T7qg�;,�:��C@ӕyJ2�L�]O�I��جi�7'D��]����|o���(��].�~���5�O�V]�op`Z����h������r��"�@�.T�q�C�٤]N��ecN����	�����1:��8��ӓI�b�)ǐw�Lɚ7ĢPt��^ba�Ў%V�)��hg��esV���I$��%|5�7{��NF�����1\	֘��h&�8����A��}��m��2��(�����k�x�_��~��~�h�Ab�6�đ� 

]�@SjE�^Ĉѭ�:������k�$�5�4J9��H9O���K5�Z�mGCW �p4?��#\�4��^���5&�a��zQGE
68�Z;�yِ"��Yc*A�k(�m0i:"��[��tq��;v�7��\#�&~���E���9(@�y�hIfDu/�k�����'.W�U�*Ezͪ���չ�����Q��ё��g�4^E�Vc��g��7�|3��n��yo��)c���I�
�=����v�PUwg�I���N�pPy����hU;Õ���$�M�8S�6�z�Vՠ�&���pL�JK&�凚�+7�x�t�p��8[ 	��`�P�'$�c�孷�J���FU���j8�<�$D/�o�)|�����X��Ex]��6����{��%��n@n���;�W�L�ע��ΨN]-�RXH��g/�Yı���ŦG�U7�~Ób+���cǧ���HH�y*R'�w����s<Bk���ޤ���c2)��4qCb�$��X�i�%�*�r�.�8�8l�Q���DO]�'K�|�ڒf�5O��c=�e�:���̒P��n�`=)��c-cȮ&R&����z���n�z��ɤ��!w{������֧O���w�N�M�Ma�Sh�~uT�����@��r[Z��!�~�d(z1"Ft(gKԪ����Vvy)�����1h�NjEӅ�ykTȩ���@���AW��%�y���m0 �>a2��jf㹻�D)�N<{qYNG0��wwD��Дn��iy������._c:�5f=������-��陱��+nk�Y���~�+���W�=�i�)_��ݶ�Y&R�?�,�9/9��`厏��������,���d1?���$��Aԋ+&�N�{Њ�W(z��Xǃg^����3��n�6�O8Fu�Id�-����n+}��fŋSG�F�^���T�#�:ma�H/W	�7��^X���(r��S�"1��3HBg bw>�p�����t�<ڐ&p���$�-�KH��1���x6R��;��I��'����W�п�&����FGC��:f7K�pv<�~�s��h��w���-d���EZ,WQ6��ɳ?�*�>5�_q���Q��.�ɡ�@j�jb�w��d�'�\�v651�����Ɣ��e���/툞�mb0֔0����oO�0f%Rg�I����X�7�M��`�M��
#V曩W]���y�����7u��ݶĸ�z4��ֹ�jLD�9���g�!���O���n����n��Wxgh��K�c2Ŭ1xa �~慛8�<�3���?(�T�\���� ���ZE��b������	��XB�;�"�K��S:B!ǄJ��1�m�s1"(�£l���]�뙨�>f\@Q�����X�^�F��
N8^� ��n�o��h3�w$���Yȭ��1i8���7g���;33�V�����><-�׭WB3�+o~�՚��)"7Z	Vh\_kZ�G�d����=�|k��A��r�ڝ�H��&Cu���
b�ݿh�y���~�$�:�Td�+�����\͟ʣ�O�Kכ��
�����c��{!�O�F�.��rM��� ��ā�D���ȓ˘3��ɞR�T�&�L'��Z�8�V[t�mk�bt�ēD�q��gu�v3#<B��Yb�dZ�vD���l_��5a"c0��Ά����Y>�L��-�|�a�~�DZѤ��l�O%�L�0�jĘ�v�
\ن��J��%1�����ça4P�y1$���GiG|1әn+<32��<�x�'7bJ�_ҡ��q`�Є�;�)J.��:7q�w"8�J�t)�����1$��
J�m� Ӥ>4�a�8��wߡ�`<#^T��0���<�wZX���Ґ�7�sbС�د��紸J�v���3��Q"9�L5��ϧ �
=6������lz�`��A���j�
ͅQ�%V�ӟ�_�ƂL��M��u�RH^\k� 4eSI��,��/�rƽt<�L�ɋ��Wx�bڔ��ͥ��f�ܨ�EY�)N�n���Q]���+H̖~��'X�E���2���ȩju>T�%'���
����A۪n�z��&�@���B�S%��m�J��`D��l�a{�d˅�?!��m6n,S����s��KQnǈ�N�)���z���]�hǃh�g4\]!����Od|�ʯ�5�y�y1)�6m���e�'�t&���;AQ6�%�y*����f4���h�Rm�c��m��	��a�Z�yqﾪYOެ��#�؝D�J����e�RzX��ޗ�п`q�JV��wW<� Lt�to������yz�i&��L��Y'Ӡa�.�輣 �P�+�Z�Rf�I��KI���Y�{�?Ƞ4��)��?2�U�Ё6�`S�������+Kcb��]34�1^��é���j��T��7o���hY�'OS��̘T!���d:�n^6�����RS�u�j���L�F��W�����c����Iڷ�~Wͦ�����ꦿ:�Z���S�F�����Nj�\�}�]��\^^@�dS��	�8Ĺ��8��\��/�&-���d:щ�8����џG�,��5,d($� +V�:�x�%�}�dFf���ǋ��_G�g'R	��m^��*�	9Ckϑ����<c&����նR�Yh�m���/��g?|��g��n߬+q?da�'Kݯ���[۠��el���'id#ѳ#ݬrgS,���9S�\b�[�w�$ul=./���ǲñ���1vaUz��E�a�Ԅ�d1j�K��~���~D,QϬ�x\�_�h����q�ߝ�������#��l1ύ-��}�,J���H�����8�	�A��Xa���!b��J���g���Jn]=A��gy��t6���#ܯ���-ސ��©~#[q5�\�:W��I/���L�>:9����K~��89|�Jf��i���k��>Nۍۨ�{�5�V�����X���$W>�;hY�W�������=Ƈ���d���u�&&3#��CJ�G��$���w�y����ׯY⅁Bh#L3I�0m��5l�.���b9�pWew�ޯ�����׏?�F�͇�����?���Vn�9�\��f#F��:���,c���p.�Yo�!:���Vt���ʷX�~��W�!+��w�}��<���Ғ����k ��D���o�z6U�Ox�at�;��2�wD�aE�'��=�Z�U6�D�@1J�A�J��<P��ܰ���Bڡa�����߫�5�Dƃq.1��DN���ƆQp�IS����lbC�Y�r0��w��I���������T7�е�i�O�҃���o�ѠU>���8��"}Q\a9�Ɛ��م�wE�� W-'���C^��1CAL�A;��������x��*���"<4f�6�:��]���D�����O�xJ�ߘ��G>3�F/r8�*�k� ��n����G8>5=�0��FQi�6O�s�,-S��6��Z�21���]ۺ��MC,T����7�H�T�^�ӡ�������W��<y���c�����dы�d�\|� l:iWI���d��n�,#
����e���5~g�y"��/�g���l�*���Ν;R!خ�?^J'�ZS�oZ��1Ѓ.�$I��-)K))�it�9e�T��Kdد��P�AsD�(=��Y�s��dt[�E���ooc��ռ 7�ڧ��k�驻�^��N����E)k��:����-s��	���|)H��Ҏ���s��IG�f���+���TěE��ʶ���g���t�+�]��71�ůhm�@bs~�!5���I"�'�Y4��06��$��\��*4���U�S׉?�!߳lioȃ<v�M+��a�=��?�K�ۼ�A��q���]�(����4��U�`�,|W���D�Y�eU� Vyբ���5ޡ!!�tD��nߏ���θK=�
#ğ�7�IwP1���o/��"���3zɏ��ԛ{ռTc�����MW&�N9��l�1��#�:�MF���R'�p��j³�+�݊�P��^N�<zf�(tA��g��'��y��Pc�%~P�������-4l��\w��*I1�F�� ~��P��tC?�8�Ӝ Y<���(7������{�G \a<�7�����"&K������;��w�g�egH�"�J�z|��Nȍ��8���k�J�IN���F�5��|� \�)>5xo�X2�+4�Ԃ�o͡!��ߛ�1��F��$��z�]�[�rV*L�����L?O�]� ����r%�U��c��8s�s��a�1�:pg�x:�j�w��X\�7��+����6x���v�BPM�&�Ҩa:m�p�Lm,�ʭ>P�=)F�嚚���S����&D��b�Lw�᭳Y�<��SN�L�AǼO�=UI��/���,&5�"�ȂDOj�V�r�V�e��*��1+u\,M�{]��=�)Цf.�OgV�=hvJ-��~�Mw�ȍ+�+<t:��i�빑��t��Q�Ȟ�;[��.�K%ʃ��������&��f��s��Uj9j*��t�"��|��U�@��p�8����hQО�� ��a���'�=`���'L�ryU�F�>�^L�#RKI����e�;������o2�o�Pr�:��da���-QlJ����gE�a���#�*S\��'��"'��͓�0��W�^�3#�Y�S��A���e�\�mܦڡB �~-�[��u� ^.�H�*��W���_���_�m��=�]}�p�Q7�`׊gu�\�Z��
J�uo��W�8����^B����C��;#�Z7o�ӻ��,-�z��R2F�n��p����~8l'x��p����L���I+�� ����i���T�'��F9���aZ�)�Y��P�{д��x��T���u�X��W%�}��l��8c�A^$z�ġ:������yk �;��OU���u͙'�I��m�y��E���-��s4zF$'R�w��Ų>T��߇%!ِ�35��������x�����#��tR�Z��0i�m�{w��&Ϋ���S+@&F��oN}�䪡kA�Nʺ{��O�&׭6r�����"~�T�$!ZM�d�B�JO�!����D4�v��Q�&�������ӧ�kycB��n�My��bԺ�Ĝ;���`���i�4$Vc�g�Zݓ �ͅs��gy�ݟ���M�"�
/t�&D�;�����qM�*}�T
����?�pO	�:�0H<x� O���0���M��H��d���YTqI��x�|_��=��T'���pq�/�y�w�����~�������?~����?�Dg|):��,5��l�T�{eA	тf�;k��Ԓ�E!�ic�,���R?w2^�FZS�A�����ꫯ�"46�/������}
xS�c�)�;�~��5�SsC3IQ��oǠ��TKk�!���)c�QZ����#M�m���/��h8��cձ��/���:�5U�ObC<\p���������b����ӟ�¤{��f%��%�Jcc��6�/&������W�`�b"�p�E��BJ!$t!p������E������j% KHV+^�z����(�ﭕA��D�;�D�+��4Đ��ÇIےi��|ՐzN�͝]%�ž"�T����U�h�ȸ@���!g��@�vt������Z���y�Φ�2~�8.X1����];�k��[�MaJ$!'�=z�����6��7��k6��{�� �r���fAJ�DY�\�q���zC����1U��!g-D��"�]���^����	ig��p��De�N}`�\.Ho��AK4�.�Bt�n�c�н}?>�eILa��p���D����|T����P�!�r�����6I���}��d\U���Wg�|�I�)Y�e-�dF�m�2�q˅��e������vu`!�푄X��� �Y��yȒ��R5Q�3j՞�l`G�;(�yq�'p�q3� J�`�\�S��1H,��[����z!)I�Q�zpK�`���>�v2Tx~z>/Mw4&�,<��@j�� �%
B�֣����G���[����|IF�|gw����M����͋x��"�ft���������ɬ,&a�6��$vl������#���j��S�����_�@�~i"��"\���y����D�߇�����RB��+��4z-�y'��D��`X.���\kS�l6��0Q��A�:ڬv����4YIm��ĪEψ�̩����Y_�D ��χ��<���^G%R�)���x1K&��iQH���n�����ہ�I�P�/���L[+�љ��Ī�1t��>�Dl�t�J��V�7�){��eJࡣ�Ju;S�#������*E�E��F)B �=�£�'�ݷ߮���}��o���C}P8��F1/����7�@H~����I���I\X=��'M���~��p/�с��P���!�	���6��3��4&p]89��r���!�e^p���%�%�C�&�Z��Ħ	f���S�:�@n�q�"�ܴǵmwݘj��JR�H�1w��/��v�~0�Z��� ��� �����q֏1�6�~��_��Ӭ���q!�N�i���*"�C��<�P5��IԪ�8���� �y��̕���3"���p�
�L:�Q����J�.M�a�o�bk^=��v�.6�q�����%��v�m�C힄��S��	VA���T�~8�ȷ[d��
#`<D"�(�ԖAk��JY�0��s�+~b.� �,m뮪+��8.p�6Mu�;5Q�A^�fn�4=���z�X�����S��qW���?]/V���ٯ���$�^�?^e����N�RP��{�'�(�Xu��u���g����!��N��&ke��RKH|u���4���Y�y	�c��L�<:�!���hr<� >쮮`nv
��~�:]�L3�� �}�ֽ�ws=�|��H�v����E�Ϟ��l��щKDҘ	l"]#�XE��QL�Љ���봢�W�fi^�?fn�ƍ���{w���A�tƧ��@Tzgf���ի��j�ͫ{���$��7�y��m�0Im�OM4�G1Ñ�4 -g�,�$��`�g����F�6��~���g���(޽{���[x��od��'��h��n'&Kf%<r.%]�q^�f�����e9�X��C����	==E�́���^䝵>����̶S��	�#�Ofi1�sm
Vf[Ag��?�/����j�<:��Zgy��}�w���V~�ZXk^Lʙ�7/P�
�u�j �t(4ҕ�Nc+��LH��vw�=z#z�C���o��"!&�P귵k�)$3[�H�:� ���=SRaJ�`�bq����$X2�n�4�l����\��+\ay�)���w$m@�u�;T���|�R�A�(���d���	���|>���o�>}���}6���Kt�c�)��0//���C�x%�����d«7 �G�p���D�+��p!�o���P^�d���~��?�<����T�y�!�/�[�9��S�Ⱀ���D�ٳg�}��DC��9+Lq��B�F�'.H��^B�{�����_����������?�O����M{xF:NlJ��v_^G���M���x��aSC-y��J�aci|v�q[���dd����}�X����
��?�#�jf��!�� T�m�YW��ҙ�0%YG���
�r{a��fGK�~&c�� x�0�2�^w�gT��1���WL�EJĉ�a��u7�X���4S+Q�	�Ȭ3��>���p5Xᡏx���i�Ƕ~��2�d��>Xi��^�~ynb� ~x��D������o�ǐ�0>DD������K�D.�5�M�$ĉFpԅ�bT-��b��J	!Q�M���lV��D9��Z���/�Xj_sצB=)^�@��d�	����v'm�:�<h�7(�+�x�~\I�9����z�O��Y�B�P�L�4�)��|2�����AK"�[�}�l>��K��L|�dz�6�"��@G��?y�t���Z��і�ss%O���`Y�0Q�yM�F�1ީv4y��f�%S'�"*�)�x��a���V�;U^�2��#=�;-���<��UJM���(j>1f�U!�CdV�R"�Y���B�VZKQ��w��&��O�ym#�*��{:Q!M��1�ȥT>hl�5#^`�Ӟ�B�"�R��H>�y=G;mc��D�E���.|C�=}w���d�(���-�4�(���z�r�O`#O~o��0tcU�9f�*���(��X�}��L�����j�1}�A���a��oj��Z͙�b��\;�C�y+~C����~���ȳ��h��8��g�k۲�O��|A����]*�+o̓�Tp��𣨙�8��W�W;Q�!�mb�ʇM���S�uS��^*��83�/��'E����DR��
�Ц�pЧȹ���Ψm���Ѥ�i��������CcNXoX��i��ks�UۓݪRG�����bO�ԑ�>f(�:"]�W��T��v"	�`7K.~X�]�$�M��yJ���*�ҦI#c�` �qڝLzl]�)�^̕T�q�������.�Ъ���#�A�C-��ۙ�#���A�d4�[ϑ�|:h�Jrӱ��*���mA�̴s��5h")��g'��'�X�f���gA�ڲj�����gp88�(���v�	����(�)�;.8��KI�[��(
&>
�i ������n��6�67l<n��R|a���f�1�PB(�OF��q=��!���>dm�F�SF�)����H�ȁ�x3?E-���E���f5�hTӫ�Ĳ������}R�Q̈�w��4��������=	�ߩN���:��6�N^��Ex��x��0�۔Zm�:�!n��B&Y�H00Y<:ڜ��(]ëW�]K�U��t$��������2�ad]����q�x�PD�byz�̩Mh/�u���/�s�1v|U�=�rfx����b��hC��������"�Ȟ�A�rM<�1���o�;aD8Q����g?��(�ZT֐�#�93Jϔi�a#ĈZ�Ce��5n��l"(�D��a�TK��F���(��&T�XA��y�W�e�QӦ�;q�j��߽��q_ŝ���`�-� �8�g�9�D�gq�}����C� q�4��x����78͕b+t]�$����-� �X']�Za�/ίH��|��YJu���B����ЧP���s�#�J4���\���kN���B���b	K��`�L�`��0ZF����2�+�"�^śW�Ȝ@��!�`�7Ӊ�w���4�2�̝7=��:��y%��:�,Q�浺����.�fYIY��\��:,)��S�� Jl%��D��4��\��w��Qm$��B	d�l3�it��+�_��Ǐ�F��3�'ḧ�y�E1�]�K����Abi��H0��aMa��Z��\_��o���ABa��"�e}z����o���R�;�[�I�ꬃ�=�����"/�DB�(|&%���}�]��zk����s�q��x)"����޸)�G�w����$Ex��G���x����WWk<+�r9�܆$����j���.��P���c�[;�۬`�3������f	wk���~����g��6
��6�)��Hh�:�G�Tj�;�*�+�ת���L5��R���d R��F���G��\��"P?�Nt�=IJ͟4ҳ�D�z�46��h4"��l�+�1{jMl� <�c~��,�#��1�ىu����V�����½,7�Na[}����uӬJ:���b�*��R?�\O 'x����ǜr+��D=@W�=|7���b��<.�ta�D��	��e�[֏�^�5m+�E�3/�n�6f39i'�,���7��
6
�A�"�zO���&\��/_���'���ϟ
�f����Q����K�Qzd���vI�V>����e�<@A����O���:ҰD���T���:��l�k�W0�un��s������jɫ�ej��a�rD�%~|�	&p���->��BQ��k[�~��������Q�y��ߣ��̱�Vw"-�A�q��`{=Ѽ�Lx��Ɉ�7f<��Q�Үi3�9�L��������ej��E����Wv�Ɵ�����65Q�Ay��ؐa�}#���l�Ǘ2�]#X�u,A�k�]��4�A�.��f��Cg���H=���%��sj��6�����㨦�b)\J�w��+4t�d�b��"1�G���K��;�i������ʭ;�̓+�Խ��2ĩ��`	�~�PwU�����X���E�S��[k�	�C(�v�@ ��w�H��ԝ�-���#�u�U�����/d�x�E*��ϋ�+�sn�S���O�&D��D)r��Fw������\�,`���AF�Շ��aZ�[Ɇk;��6�j/tN�ˣ}%L�Q1)���h9,�S*�Gm:��}[v�i�<�B7�7�\�m{��K�A�3|�릛��H,ܥE��V�ƒ���ҧA��<�v��# ���~vv�0��"�\ �.�'���y�d��|c��G9F�I�)����{Zs���8SfS�`j����6:.y=-�j�i��7z'��O�5fK�("(�~�I�r�������������w��rIۏgO��g�s��,���PIJ�Nh!������z�^ɲ�\l�����XU�V7{d��(5/mP��d=���'�4��Ő��,[6pX� �!��b7�]U]Ù����ߊ�]}���>8�'s���_�.záؖ�jeT���4��T�Y6��i쥖���Xs=�jEUN�1,�C�Y��{*�l�[>�Lr���l�dl�����L���>	I�9�%�m�-FkF���c��"Ŕ�������i[���I_��U�d�C�켮o�61�!���h�p�9Zp�P݀z��K	p>�����rD�[W�m�I���p�7��'*;G��}�Ԍ�� �L���nv�3�Zڽ
g6���\�h�pu�k�Y�e,�Q�b�M�̊up���!5�O�� `�j8��L,ɓ/��|�g�^h~"�nJ����y�n��@ā�@�/��F���`���!�n����L�~{��/��8��E��3�>[��#ݔ�v�^:��@6So�I5kpp��b��g���p` �|���U�ż,F}����M!���?�4�M��6@��J���栱��zGw������� �(/L�y�tnsA���r2��`��q��5�فcX_�5�l�lԶ�6�rz�O,�>%�:���S$�R��-���1.���D�cL>���k^�\N
����'��]]�߬�O�Dj��
��fP)����7�Õ�7`>i3�-�p���rE���f☵=?ٽ=96KΙ�������3��V��L/�^#e�>�N ��}�\�e�&`�uro��d�1�OI��l>�&)F�GC>���tS7h�C{`V�D��p�$�����8 ��x̦�>���k��0혊>������������I��Ms��+�"+�i��h�d%$�u���\IrX���I�m�|uA��F
P��<˶$��E {��>!/�'��\O@k�N�'��G⼻��u�0�\�E!���?:�t�i2yg��,sx����I�AhK����ʅ�$����ݣa�W5�t�p�:��~Xu���8`�ҌO4�--���՗��d��U�',@�@!"�
9o��o��� ͘R�"�O&W�
s�㨏��@����]˷@���qy����O>�����SX�+.�	\v�;ɭ���c U����>�$R�䐜T�8;�Q�I�8��ƅ�������&�k߿g�:�p�FB�e
~�݀_h>��>��/^�}C�����ݳg�֫-)Y��iI'����l1�n��:�@ԝfU�D�F����F�Q2�tiF�NXDYk��п|���,2��_�w�O��d��$fڹ��Ѷ����-עפK��!�~C��`�F�]t�*�� �V�\���hc�8����N�<S8F'�܊A���&~�J���S��RJ hZ�"&݈���)�y�ɘ�ۀ�1ga&���R��d�\�؊��b�[ʡJm�up[E��%���ZloXG�qT��N�ʚ*�	s7m}��-��������t>��Ұ�3U$�a��	?/��^ ]�bvu���rui�!$-���4�/�����۴CK��'��6�j�V���[���Z��$�hb��`�F���K�v����QI�����+��X�n��(H�|�٧$�������5x=���F|p�Jیl�fɝKYFj//����7d��A`��4�X�B�.L�H��NMر�� w�v���-:�z$�.� �!�#�UbV5]��|���&Ӳ�̦f�%�I����c�h!;�N#�&������F�2�N�C��rR��pH0�s�9ɉtE蓈K����	�{���k�,�v\O?Gw�ܗb�2�^���kIO�K�,)��G3�A��|'���>0_1�l@�o�@�MF������k��y�v;�5���.�R���^n�[��?�G���l�L��0kAat�6x��,�|���Ac����UY�
���1(����8-1��h]��u��_B��5W�qXmz'���B�۰c���7_Ԣ�q�@Ei*���ў�+�H���]�mQ��ԉ�̋F�\%�a@\2�\��H�m@i���*��ޮ��>��t��ۥ�v�^��C�$�R�w�\	��ec�hƖVx\�@'Q��1�.�� �'ͬD�όB�\�`�,F(�i�=G��e*���G�mE���mQ�x"�k>��(US���6m8��&�2�y@�nS�rZ#͠t'c�$��O�r����;�'KՔ��+�%q�@�t�1��P#�=f��(�hA�����"Sڇ����իǏӇ߾}K^���S\+h�
	~��\�����^��f�!"`.=*2l&�P�����Z��Ҕ�e�z�F`�@�TE�2R&07�"�<���0�ś`{�no�i@�';�)Z�(����]=��4�)�G9)s6��L�3٣֊-+YpP@+n�HS��!7 �S���)�r�K���t��λ����j��� %��&��Ĺ����Wxc�Mm���s�&u�B�L����j�A9`}��RO�Í�m��#Ö �G�a�mfY�)���Z�##C��	غӒ!'��!��m�#��$��BUN*��h4[�Gki:$-zz�g���8��D�&�H�g��P�~"-M�����q�� ��^��5݈F�(0�8E�����
��\�9�c�y��������yrc" ���ɓ'�B��)#�KJj%�0݂��ރ�n�z�G�U��LA}uu�����/|���<��Q���nes�Eh�V��
W`��8�D�1(A��yP+�l]�\!�4j�I�IJ@�/o��w8�x57����1"��Ґ{bp���'tA:)�h�>���2m�i=�D �����/�������Ӕ�����~�3Z�ׯ_����W_O'�&�����Q�hL�aZ�&���&�S:$���f3�v�Q>��@���˳�w���aR�5�"$�WVF�u��R�$��5န>C�Bt�pnwɐ"5�lqZa�;mBK��C�������Ð2�" �Z����:�	
���<xaOf��؄*���w��m�M���X���&�e��֏g��Ǝ�� |�t��K�����? �s�7����i������\U�[9���6j�2-��>O�H�^9��1�Q+���#,f� ��X#D͂�+Fwh�[wm�O>���O?=><x����LB{��X�Y�CqB `$���8�����HR�K5�o"���JN�W1~�|푏ϥw�O~�G�oA��������_��wG~�^J�ie��n���T
�F@�a�غ��Y�^"0�����(E; W��4zdI��je+#��ez�V�c���
�d��������h.`��_lb�<W�%��}F�W0B��_L[W�Ġk��b��9�����X+#�Li���X���U���E��3{�|�y@��2���3-1'�.rυC L���i?V�钨جWց��f�5ݔZJ<a�a|		`B헩��[�ɞ.�k0�Y։�XM���C�F��D� �K�0l$�Cb'@����xh&m�aW0u���ؚ-�C�M+IT�k9"(��茚��i��<�KB˒�;<�J�(�Q��N4�}��q||������N�'����(`��.��j.V�|R�0l<�qY������!���䄑��	��Z6��[A+�����BuA��&�,LaNj�Ze���wP�a@�<!^+��akY5O3�����j *�lu�@c�  g��<:k��S<$�l���&r�TDޅ�tT�[��}���������&�t6��M��E�@޽�)g��@J������yj��ā8'Z��&�/p�!t�qm�%�M�:R�:V��jQSid�0��6B�cZ�0�db*�$T��/v�b+v:zΛV(��rj���v��l��v�L[}����r�7֏x��ˊ�\b��h��arA�����d��ş����֨��,ߍ��SHO�Z�?��u�i�#�Q|r}�� �qe�}��N�P؏���X�m��8{L�^�굀��=-�`#�R <���6�*f�Z�d;V����@(8w�7���\{�!�3�(��e*l����^���Q�}.5tѕ$a���l'Ҳ`��b
���N�␈�Ri����dZN�1�đ�½`���"IA������ϳ���M������������!"h�u�~�%i_�?�-^+�}�b��yd��'R+��_&@��b���HB�$��Z;�7���vSGiGE�R�z0Lq��Ia���a�xF����[�P�놋�gd��S�5)���
O�0&>��1��,����2����;ff�n:M� �eix�r{�j�:�O�LC���c�4��Gb�� �������@�����-�io��;�n��*�V��@��n�?�@�s4�K'(us�R��iC$37���2�5}{2��ڥ1�����κfzڛNL9E�E�AK<��Ý�'�J��}N'�����:���M�E_߲(���w�gQ;�Lf@	ţ{G��p��mSJz�	d�g�0����B���V�ת�d9���W��ښφ�h����ܠI�b��ޡ��O��D�M����c�a��Uґ�A�۠^U5��D+l�B��I���z��xxx����%�9�$�(�鱝�Ow�ˠ�ox���ޣ��8�5�I�{���������	�"6�f<�_H�a<B����1�T�MT��(;m�7�,�fq�OIdA9b�ӛ�&�!r4gH���'�m���D���L��n����޼�ӛ/~��kEd�����lZ��Z�1w&NԮρ�d;j"�t2��@�+x+N�]����AE������jUo�rFb��?=>�d�}����i���!��g>�u�T��������1|" �L���K-{�����ܶ)���'jA�8<8�Y��gEJ�ᇟ|�'������?>:>��BN��v]���ͺ��Aã�COG{����t�KW�����oOi�*1���c�Wh��#���A���b<vZl`fٻD�)}<Ɇ��t��f{�����6�8��l�?��i>�w6�� =��`������'��Mkz9��d6ǁ���j������(�:e#��[d$*q
4�t���U��0�yG�2	�Q�OA��a?;p��+���*Ntɕ^^\��҃��a�m7�Ç܅\2}����/#�Ub!D�����׷�}H��좔�0�x��߼9}8�G_i>2Y�����5��QW������V�ҒX~²kR���Y ze=˴ak|�T�{�n�uEF��L{
�u���x���?���?�䓪H�m(>�v�&*(�\���S��6V�D�f�A�����+6͍�3�^Km߶´��Z6�ڹ]&�G�2yOt#:�>2���cB��,K���?_<}������Vj��?�Vi�&�o�&<�vx͌ªD��6�S^$%���<�,qh��$٤�iUN��L'��c�a�ɕ�f��J^���Yꑝ|=u�|�2��^ l���L-�<�
*���3-���êG�h;S�q�g�9S�A�w:%�DFْ�2V����i��T�J^��¯�>���;y��-�Rj���n������Ðt��P��=ᐚ
�J
�i�Jm��؉�@���U�Q�Q�Sw�O����˻Փ�i���	2:$j�<y��&"��,!�SH���r�~��>�L�p@z�_J�D:t5�Hl���@�0�RL��%���/�ю�pqyF#;����ނ���+�N�C  �h���8Stt�6��O�,@!* ][�`Ǚ��+�ȁId�Aj&�ݻW��?0��l'�T?|��%|N�ʄ��@N�̃�1�y���G"���\pq!�����9)��/_~��+4����|L
���a���p�����2��䱧oq�ܔ�l�ks�6�S�QF��$L�k�uܸHz<�Rr�Ȅi4c�⁩#�Hu�8�泘��bA2UH} �ecy8��������;�t�AK�+X���,�#{ O��7�Y/��S��̒�+ːr&�-�˫K�5�<��D%\�<���7�O��ȀAK�c,�è�ZH��jtn���"�T�RJ�Sc��!.ӗ���o�צ�N��r�#����d��q�6�y��Ӱ�ci딽K�m��Qssf,7�iKx)�����-��hf���1��+ {�4Z��lw$��Ĩ��{���3M�M�[e���R���F>1��6h���Kj���`'��z�D��
�~�2IZ�i�=�I+��?~� $��a�!_7�N��5�/�Q�˻�I�R���W_}兹��7�;?7������k�ض
�:i~�2�d��~�c�O��S ���*K��<���fR���7�0C�M̹�$�E�E�e�ŀ-��YF�#۶DX��H6�e�̌�B���ID h��AI{e�4�Y����a�W�I�/�):�)',��S��Ʌ�G��6�M�v�G�Gi:�}f��� >x�����׫�X6�)�I櫜�7ef�	�۵tj^V?,���t�� ��I:�	YJ�	jl�.���=d�"�!��� ����aq)S
��Ja֐�4���3T�#��i=���{��f��G�G������q�:D��W��r,@�j���3���wh����Ƒڿ�)�rB��_�nmYk��J�8�nԓG����%�J��>������-�57��Z�b%8z�Z�$��
�ö�j��G�[J�ѲS��8-c1����tƜI�I�̏R�;sܥ������ 0�ܶ(]/�TLC`b�$$��	B��k��F�,t�mTȀY3;��v��p�l��e@�G-��]EF_���R��#��%V��V0jL�&ߔ�$�,~�����@��aDaޏ^�$�S�Wo�x��A2�p!u�6P������2�;"������b�y�7�LT=$K�m�(6�T���2-,�Zd��B5.�,���^Qz���AN�8�*b��ю�AD�pb.[z�RԖi��E.��r�
�����E�����<�FVJ��2��>w~��~nW[�����Y.�EQ�Hi*\�=K#�>�}�����)�����R8���p4?A�9��/;�M$�1Ou:����3��ҹ�|`��V����k�ԂyH�n���2��,�9Wf4�q�|��0�-��)S3�*��ÛI)��g�&.Wd��Hx�^d�ޠ�N���C�A
����s��]����1�?+�D��C:Rt���sZ��{\�3�\b�<�8\H!�.fUJzE	 �/��^��D0���M'�w���g��	ΛOkׇ�赃6"z�b�z��]�-O���Dӧ�9d<.~����'?y����;G�c����t����g '���#KV}LUAp�͏�� =$m��o�N�z�7:::��K�lT�o	(_V��)���f��.�����N����A[W���
��.Y�\1t�^	�¨Wf*hS�)S�oVa�+`�p$Ne�$�fND�z���v��K���.��$1���y�'��p�B[K�1��ݎM��s�^�qD��xu#j���������#r �~o���66�
MBԏ�gDID�{��y&�̠�ɝ�q8u��֐bCF�����p3)@��L�Z��f �B#͑�%é�>J�6�x�V2Q�]�f�.@�hc���ģ80�~�p*)%ڮ��	��`�$}�u��ީ�#�J�b�M�)r�-����`�!/^h�F�K'����O?��˫s��I:1ϸ;������Cj��l$LTL�j�����II^0PN��1$,��a�<�_��K�.j4M�;$��xĠ݋�����L�>�tp&{�����kS��l�DR�X���O(nI���=�h���_Yif;В����f5eJ�=(��k+�=H  ;�z���"�'3�ܙV��A��IM=Jd�C��O�>]L$0��.���'�`i�	�R\�i-�J��%�Q�d��=�7��W��}������hD����_L��3�$�N��̰V�h�����VH�̨�$�Q�ڑ��I��O߽#���h?�~(X��n5�W�	�n�n2���:�&i��c!"'U�l2q�4���kF�`;)j��bU��h�ݱ��6� �aW��ZF`���@n�|�Ny�i-��P��ܼ1M=D�������i��>�«H�IxQ��^�rYb��󐘉��&��ݶM|ե4^jMb�d|���?�+<���/�\���+xNi^�%�����M��qL�;6 x��E���r}vqU.s:���Í/}����ȉ��S-����%&��J���@��zӷ|���0
�����i��ܹ�l7C�VâVa�%�(����%!;mZ,Ix�$X�cJ�8����E�[ӑi������N`�Pe)���d+p���'���m��A�r;q�*�@(���N�~��V7�7i�Q/���WH]fI������Z�N�y�j�PL�	<���^}ݰ�~���lk�W|v�D~tp@~'�`�= )'`
�(V�`
��t��ނ�C7Z�z�i&[���2*@ �w��̘�hEU�FQ\�ܳ4��5���7��͘25�$���`'`�%=A� �[�e�Sh�D���Ir���B����Z��Bx���Dʢ`L��4ᩱ9�wp{̻�t�$�ሿb����ԁ��ACl����Q�DM�k�)���yz���!B�Y!l�A r���l����s(+x�g;��tg�5��6�f�a�1�i��I�%B��f�i�7�1�Q
'pk��b�l(��w��T�t5��O$��ѾZm#��),��,.���b&����
�3�d���g�0�@���2�)Uqc���msyyzx�&8[iNo�7bj�8�A��@����bJ>�K�����:�P E�u��R�o+Y,o��WQ)#a�F�d�)�E�%��ޚ6���i]���W��ƾ�I����n�٢x�p+����ږI��{X�d���c�uo��v�����o*y8��W������K��۽9����v��-ݴ	 �a��U������s�G�=I@Op����7qPn&�u�K9t�����|�Q�Y�9g�_j4b���wp*Z�\�c�C�����g���R�ݥ�V����Kie{$�?��s����`���8]̣4V������r%�d�ZL�tմ�rW�����v� M�*M�i1a>DR0!��l
�+�i�<�JIF"�;v��n���FQ�����1Ғ�ڔ#&�]3��
R��l��\����$��/EeD2�fK�̍�x{��&���N��]��d4G�G�a���������B?d�p��ء��;�)��H"y�B��l��D$s��
qR>��E����`�d˥�E �3�v,�*�T�fMK�N�^�:c?�f�"У��w�%?88�N�M-H@,E.��Q���nm�/���YA� e�t12;�.VEj�nG՚iS�F�gQ�6��������n�'T�e2�M��Q7X�N��9#�����_���Ň~H�>;D5%t�_�^�z��.N�FY��I� �)�	v/l3�xc�yH_�$�L/��R�6 mw%R��H�lVk2�H�1��H8wM{ws�N������d�=~����ߧ%&�ɍY�x��џ��ҍ��o���w���ブ�
�tJ6hc3M�C�ÏàQ��DD3_9}��{���cR���n�ʿ��Γ^�X�yM�㯅�!�������G�?����M�z*�B*����m�y�Y���6O��-;&D(K�N��dA�Ap����t��P��)�Q�,5{>�{èQ�DZ��G�!cl���T��ۜ�;qD��5l.�0�L <R��F5�����7X����r����*���۫��=� ���ThU���_�4�4oh�K��-oo��=z���ӽ�=:\�0�'f(Π�|���|���J�O�����$�hl"�<h�&Ҭ1�ZiI�Xv;T����|1a{�|M�٥��z��hؼ�7	��)~3�욑��c�)�R/kf�X.o�cl �b�u���)ZF텨mG�꣤���ɍy�k������W��MI�g�`r祤���m�}5MUq�f����e#�����Èn�5�$v0�%�r9��-r?"�Y�01��0���:��a��p�C<�C�۫ѕh�|@[A��2��΁�T(�g_[�	�.#�_$���D�/��������̗ea�}q�<P�.D&�m隗�+ؖ{��Mwt���F;^7�5�0P��6*&J�e��G�w�)���rS�q%g�5n�����%���6����,�pAbZ΂P.K�ޖ��j]H�Z`<N��.e���~F�aԂ:j�rTR�lTn���N{�Q�`��g-�޸�րDEW��+�r��ʵg�/ܘR[L���"!�h.M�j�V�	����:k���
�k���6�H�`K�-�]$�5d����>\��F�����E�f�u�oo��`#���|�1��Ή�,��G���X�j%�Ji�yx���tk ܊2��
�|��BR�t)����H�D���  ĨKG�P�J����JJ�Q'AX����A���"4B�����'��Ҁe�������1@�@�B��&2�LNb��=�h�G��^2�x(dHtXJ
1�^�"� �%����N��S�s����Xs�����>yqqa������{��ދo��}�Rb`�<!��4����6����a��;d�KC��<1�i���"�ߌjc��3O	g����{�J�5VZ�u�*'��g����X[�	M�#�iB�3ଙ��)��)�b�U@��On�[<��{P0W(.�*�x���Bs�0k��A��*W��5�+����j�'�Z��+y^���t
C��,�t[��H&829pOYj(�}9h��	� F< m�A����1�T��_�FG�.���̕+#U�e�fp��]/V�e$ZL�@�ґz�7���+�-�)� O�@8��@V�W�Y�į���d {7*#d;�����U�\o�����G�$
!v���,��a�'��6��$��:��x�	�M�i9���Y�D���@�˳K�!�ڨP������ 6�3ޓ҅Is{�zL2O@�ϸJ�L�q�}��H�*���A�i�j���f�0�����t,$� ������:�-4����$Cv"�%1�w���Χ�=���!��g����TP�1��<��б�l� �P�!�d��̩ZގSU�5��܎됼w�(r�>��É�0��)
k��!�+�8����[��1X�gv�z��-�K�<��A� ���f�&�X/Ph��ap>0{c���<}^�9�Rd���Au v��`<���!Zݰc�*��׾L��R{m'� �Qz�O݄C��L3k���0(��������94ZE�k똨In��Y���yTS���k��r
�C�����׫5�ܻ��5����ΞQ����)!fs�1
r�B4D,���`�H0�h�A�¶4d>��m���|�8��PW�9�{��%"�{u.P�L2�P����?����Gt����\]�;���_3{Ɯ߄�����<xpzz��^��5��[�\
fI4�L#C�ѣG�;�I@ޠı�<b˺�͛7t��|�}����c''���#�ͷo޾}K��g9;??::**6�H:�EJ��?������ѷ�Հ=���'�+�l>����֣6Pc]��Y#Ak91��fbK#s�5�@�IYA���2C��"`��� ��r�Xi�@�H�?A9%m�1B����}*L�Oy��A����5�Rq�n��~#��#S�`������33��C�e�uF���(V�F��CG����*�h{�N�È Z�ʵX>hGM��Hx��km7�����WY_��<�/�������>���UB'x����d"��q�<�@���I(��մo�	�.�/2f���5���nye��^�Bΰi�^�p
���ٟ�ٟ����N�::�O����i�V}R�����ȃ�g�--\�S��p�����O$��S�d�`'��i�a��1`�؎��D֐~'3���L��\2lHۇ��T��\� i`sWM���=)x��
�u����y/LBx����b&އMBe�$ܮ��	8�8G�����R�2/#X㯤�� 2{F%'�	�[\Ua��_z�-[mD�cV��,B��	|vli_~�8[:�MGz���k���L�A�7�*�Ԥ��������d���r7y��K%	<ɽ3-�%�8�8�fc`A� �T{�)�*քx�Ȕ%�pF�09�7�����ϣ���^�z�fd#N�8r�MV�j�֦WLߠ�uqD0�F�-�I;�g�8K�t���+,�N�%g���zEh�Q�'j�s�`A
�5;r�ܜ���&���!!������J7��s�^m!�D[j�$"����$�D�r$�z�6�Pɸ��v,�i|�6�$ǆ�X�+w5Ԙ
�C���ً���n�ԙĶ���_p�{��7� �z�@��U��D�V6��FS]�c�Y%d"��1JKAR<���� �N����DϐI5+�	X���^�n$I�k#���L!���F)����Ǐ-i�j�k�)��:m��H}�����G�m�B<M���u�����	~/��;�|���)r&�<�	�k��1�GǙ�z�2���s+���gGǇ8ڴ�?B�s* U&X��b�{1~�c'���#���D�K#Y轥��i��S����k�E٣�L��"�,(�k�n�M����g�����rC1����JVn�FZ��ͺƟ��mC;�C~4�z+���R���|�G�0;���ūgHG�C3���=O$�����K�z޻;N���0�ίo���[Q�1��~�Cf�,��<I�zy���av$�{*���^��xd$H�'��,%��@&I ��*�zuv�01��ix[A`�Z#O� �+L��3�\%�I���;�!�4�HK�ؽ{��1�4�g!hZSa�9�'C��4�g�l��h�R�7��j�Kh��ض��� ܘF���;�i�jm���o�lf��oݢ�Fj�l���x���{,'ч��s��#b������Z M
͋��j�u�0��	����j�J�LZ��*Oy������SIw����(��M���W�=�uH ���J&>�ԫ�s�o��I' �ퟤhô�u(�[��"�"8�t,Y��\�v��&�UT��O���>X�j�N	$�l9^]�mظ�"|��̕�C&Z8v��o���Ǣ�8��e��AX Rر��j�V9�ٝ�V~X���#D�=k|z.�A�(��E��K-,6�sn�l��[�0�1�G.�.���v�>�A��p,2R.���d�4��8�d�͆g��L��$��:ZF�0�N/fid
�ڲ �e-�$\ x�v�����F!uÜf�u��۽ee�6����(!���!��l��t",�G��o���h&%yP�}Z�j�2;p�2�CӃ��y(hKB��T��c�#_�y���k۴�Hz��t۬�򁁙��#`q7j�.���!����6KD��dyS�!z����2�桥��06)�R�䌍m����·+��������G�����	Y�(�u�I����$s>��?��?�������1RC�W(S ��b�P&��O��������}TA�uUÆ	����y�8���ռ{��1}l���Lf�0MuC�����_�Xº���~�_���Z��J����g4fp��3���������#�� ���Fx���9�j�X��|���Р�n�G"�^[�q��<x��>@�'��$��ٹ�w�7�j4�j'{;xf�z�5��qsL�����������g�q��R7w��P���mz�w6+.F��g���Dݦ���3,ۙfWX� ��kN�՘WeԎh{�f�/v;��Qڐ^�v�	Z��n��q�ve!'[dnl0��:u�%�`��A�Q_��7���q�����:U}GC*�h��R�������?��7��b���	��D��[/p�*�[%م��K�'��A_�b�x�/6
<�������=B���j�@;�������W�W��ܫ��L��,I�(5��Z0�;�Q��J=�F�B�уcu��pߓZt	�qx�g��Ak��.jBoHT��5� �[�k��@6)�!������bhqI��L
��	�����kKL�b�KY~j�:(�ae��ߍ���%)8zS���d�$�'6a�������� 	<��Y��o�`Q�q,V�]��y*�VO
��� ҹ�qۮ�uܴ���MS�zE��; ����v9t�)��Tvh%	�]�,J���> *'�#�S3���;�l��0.�K��cױoF����e��E��,���(qmF�s����QU1`F����m��P��A�H������;(�Q�N�l�!*��1C'��_�,�2W�L����X2�l���~�k�|�Q��+�¬���q�pm�R1�	w|��/�"CbC�
��IɤSB�v����Fv�[$AE���\�6t�4��F�r|7M1�ϰF��p�rw����@�qFפ=Or��Ç�O8<׬WF;�5���9����~�!+��kw�0���q7ض�|�h(0��Rw�;�����N�P�o�J��Ůb�+��y��L�G�. � ߻Sؿ4�]��eJ�-ǖ�E��h�3u!d�@�h�$+ǵ��׮�j+܅�ž�L�a�s��d ��;b���و���n	N�7hˁC
ѵ�y`EV�5��ѭ��J|CF�=re[Ae"a����@�}ł�:��NA=��`�VIC x�2��D^��a�w�/B����go�}�ki��e�h���~�1�I�-	@Q@�ô�&-;���S�ڮnОH���5	 ����}��D�!����y�(t���1�aP��'��U*��JdD�aǧr���-���E8�;0�W�m�D��&�-$g!�=#��A� #����xΔ SZh��X&��V��z@ ݬjL;�&@
ᄚ�mZ#�P����%}���Jd��8#u�VD��jԃ���Ll8v����:蘙s�P���e̽Q���J�I�z�pt ]A�A��4ʽ�w���i+3Eh��[:����lg��IUIM/�*�Z�v��
�A�����,����n8=�v�뼄8ڵ���Z��� ���%����ylx+t��J.�=��U
�p�6
�b�J,r^Ӎ �B��K|p��aq��fk(	f�Wף�b6����v���9�b��&���t���Ӭj7�'�� ��S�X���x�ͼFx���+�m�5{�:N�&��Yp7tH;v�4�7�UB�하�N=2�|����.z���v�+�9��Yu�ҩ��,8��7I��$*G��DܶrF���fR�CN�l��G'K���W�*��!�d6̑�6ֹ U5ʂm��i�̭��F���U��F�A���I�DоA)ͦ5�b�T""���!|z-��	7+�2Rb��*<�eV^��i� ���5������}��t����5�"��Š���4� �a���\6xt�[����`P���Gd&�9(���B3�:�Մ\�>�������`�扈 -:m��oߢ�0p��i<�E���??��C���6���ٞy���o޼At��4>����3�1�!��do��0�QŌUn���o��x����5��+?�������Ǐӛ�]�����������֮��]P^�C^�j%S֬��a?C;[���i���k{F�I�i@7���j���B��;�C�,T����(3k<�ޜP�{��W��f�?�)�ٳg/_����|h!�.���N΀<�#luԪC�4��t�ZBn&=fS�u�)��5�3_ɫ�nr�i�$�Zk����.Ø@<��@>q
��G}�͝4�cgʢ��ɮ~TboF�׾v&�l�2��R����qyq-��o���g��_4"N~��*&eβ(8�t�Hr>��L+�X�H,>V���ky��SKG�(57�c~�*Ha��͋��@�@:��-I7&�}rRM�F�{x"�}k�ヶ|ὧԷ2c��uJ�,��Nj R$�.0�������.V������a�X֍Tᮋr�xXPTu�/<�1~��D��!ɝO�����V�G�Q�5+36�y�_�H>7Ƕ���֛�^C�:��ySgXP.?�a��*촧�����^)hKm�c:��7L��⺖�'�ʤ�{!:˵
�����t#&�K�"#��+GU�A�|u�����C1X��iⰑG����D�l�#��Z��7�= ���v��DX���Z��l��6�î$
�zstCL��h��|ݠ$�A�,&��$�Ro�Ғ��V�#=No�Q��E$��ď2�YD�0��JW�$${>��%�6�@Ԗ���p�f�b��c('���Q���Ҳ�%:�i�礿Jx�s=}��@jۑ|݂��t>��A��l�3f�4��TK�ć��+��"t��rY.A+N�K�z.��Fݲ�>�`��Y��W �dE���8 _ L��$X���=i�JH�#܀I�X츉�EaF���f���z���;g0��;�ca�E5M}�r�O�#6L%���\��Z+�i�n��,�mKPN'���A��ټ�+Y����컦k��y/�f+C &gD� ��"�nH��ҜBۧ���3X,��W��q���5;!T/�FfQ��F�(l#�=x����!��Ǆ�Z�TkT��Y?P���}0i��v�q:Z2�Lɗo~�GFV6,F����e��"˘Y:����~��w¯��赳N:��K���L�����5lP$?�JEIt(*k�.�{4f���m���O�%ͱ���[dN���<yBc��^
��G�^lTl0�mzP@�'ŐI�'/w��&=#�I��c�����+B���B`��G�H�5i�i �9B$w�i� ����{�rܙ+�`�a�Y@�x�Y�|z���3��`�<�L�c�p��;K��!q�G���$���|;�D���+B�*�g�A��t�\�n���1c�)�Y��m�
#�#6�F5ː�f�o��p�^+�E�`G��9��؄�3p�-D�^H��7�P�8��$QZ~�'�Ԋ���������8@�\g�?�8�Q�@� �'��$� ]��Lt��4�c㼑��|�~Xr�XF>��2Z�BzX�J�$	H��A��8��s�0��I����8$dH^F"��̧�QWɻ��.�0�:�(qLQ�!NڧUE�8�5�2�Ҋ�X���Qs�gZ1�9�"�/(}l�br��n������R���J��P�V+�W,9�J��yҬH�4>h5�R�[�ҔL�.]�}c?�V�p��N��hժ���WB  7��|,�'��6Q�.[l�3��Cv�͖I��!a�c�Js2�1@@�;z�9� 7�	`��M�������}ɔL6a�9�X�m���m�XJ��]�6K�@_�I�P�u[�h����-��>\����)e[�S�H��R�E��Vۘ�f��8�dx�䌦0Q�!G�\&���/|;�}�K/p�B]���f��et�L	�&
T6xW�Z��c����^�d�0�I�"��,�]KR�+������cN�EϐU��Y������f��qYVa{�vn;ҒONH��5�t��ɸ�$�
A*��e:�n{DO�ڍ��V�8hP+�B);mjU�j��z���G���?���H��LF��Z;	P�) #���,�_d�̙�>��C��)�) �M]����0���Ơ���{t���kPh(G[�Fzss��W�F������^�  �~uu���#��2
���='�l3\^�����������������I9w1W�Q��/���3�d�ÎH�SX�('�H�#; c�%�RʰG�w���W_����t���>�؍�jٽ��h��)Z�|r��հ��0�ƣ��>;;�<��Ҳ҄�0�G�(b���˴�4LP��X4?�wݮlsD|�w@'[�Z��io��ڔZ��k��)�
!f������g\p9E�Y������`A��͔R	�`����i�N�EĈK��wR�U���4M%����&p��Cp��� [���OT�-�h�z��k�&v=�*��-޾�S���h�5~ZqP|X��
��4��K��`E����o�X�=��:I ��z�qI��N�z�x�L��x�J�+�}ޒF" u>�!�eM�h_�~�y�)���<��Eb�ܝP���`��q�ⴰ"lW@ng��M�Ȉ�ג��i)�?i�~��.ŝ1�Fɑ2�z���$Y"����hr���ʡ��t�2A��]�>ا� Y�Arx��)*��]��
��id�La���M� �R�}��~נL�j�P!�'\S��,�	�SJ(��6[��j:~Ƣ�_�~��~^�]	eO/�*e�}�[J�xgd���\*iy�Cf��(�_�DG/\�B�l��H���p@NN�Y2zb�zB[@\b�!�P���%��\�=c;$3�f�)_��t�8�gq�lӓ>6��K%H��p�Ҟ�&kX?p���)��E�p*��e����Bu�����°�H�j�9ye���cgp0�sHY�T��5ol�9	��}��(�� c!ķL�ƣ������E�p|W����^�?�t0�I�8
�k-��dS�܄�c��v����s�l
���G�n�J���t��ߑE����gi��ЩqT��A�CTo�nn����\c���3x���@�-��kSp�����g���P���J�A$S��"�K\
%ƖU@���<�مw�t1 ��w���*�=�tkЄR�\(�nDo~��7ϟ?��}cq�B��<h�^X~�r~pp���������裏`��z��^����A���ŋ�1p`�\2���߀v,+�Fͧ3Ҳ�>"Yt�W�_�w�&��э���N�����;ib�N�1��H��.���u�)#S���i��1��_c���\&d�! �ꠕ�<��,�<'į^�z����t$躚�|� �#2��^-W �bG����>@���P�.����D�����,ػ��l�l����ђ8o�XLA6�Ӻ\n���OD_��EX�rJ���I�w��O�����φV�/2�蜮�f"s�C��e��q#y�uYlB�C�"6$����8�����g�Pp� 7�a��d�]̙K�{'���+K�3���o�ۨ/X3ae��	�Tc��f�6��r��i���J�0��c��!��$����TqxF�v�̣��*m� ]�vm��]�`���~�g���>��_�d$�薎"H�-�ä�J�2&4ʴ{R�u�W������Ո����a98���H7�HP��i�.��w(�AR���m7 ��2���noo6��N�<���*k������O+kL�P�3Ux��36Ȗ�S/�����єС�KAO ߉n�uc�b����>!G8���p'�>n�!� ���1�[0�A��$]IʥJ��M�*g*�Z\Y�ȩD�  `s����KW;���lϱ�c6�34M�����ߓ�t#O&W�b�"�R�D-�b&@�.��� 5>I0!2�������FH��7LmF� d������>�,g2֩��"hd�d|�f !b�~D5����8j�3�`��%���W\@&��L�;p��1���z��0�a���4�{�V0а�����K�o_��jY[�vD m�� 0�A\�3I1�75R"����7��d�7Ҁ��Е(%�H}�q+/D�K!;Fm]��������͛77d���JT��7�-�Y�*�];�%�j�
ar����s�aQ,,�E��Bc#K����fH��s�Dz��5ᩭ֌�����5H�_z.���T�Ɏ�t3Gѱ��c�OR���u%��?(�Z��� �G����y#����}�����H��<鸌1J���韏?�������/~�1�� ���G
;6J�?�v�803z�\��2��H"�S(Q�5M���-c����:�+��y�j�\��Z�ã�	U���t�#���kz��ǿ�����OJ�MSA�b6�y��	ȍ*̂&�s-�@�>C��	=jY�9��	��X��c�I���1�97mp�0j�
	�k�-�?��^[���aTbwZ�	�s���������*ߺ�����@�᯸2�p���~ ��%[#��E����������;U�kA �G_�>?�����H,���td,��z|uv���_��bN�ĤTL��s[#�����9t���	66ʕh2P�!�������&�T9]���@�u�J1�Zh�ז2��`��v�)��[?j����j�%Ҙ���h��B؟�$
����A)��r�h�J�0+�խV��7N$@Q1�A9�����Nl&��e�'ɀ�lf�8�a�E�ش��([�h�Ǣu�*�,��x��#�h���v��sn���F�8腱.F����+�}��fWpvZ}
�k�;c&�2|�����[-�d���n'�#4�r��{s�������5����p*ok)������lC9e#I��?4����|\k���TV#�
���s`��}�6�U�n��j�|�y�
i�Mن�}�[y�xY�q�~����=&e{����,�g�p�$���P�ό�ٞo"����6o� .�jP`�'Q���3�P���������9P���CL�О�zYV�J�dt#TP���*�}�p
�#�h���E�l��0I�g�\U��ҳ�/�"���!J�('�����gg�"W{�v�<�=M��0����˳�	Cw�!�}[��EIn�lӡ�W[��4���)V\�=d�M�"�Ӝ��*�i�nq��}F;g�۾�;ضk_ǉ��<�����P�Q��:=eZ��Ւ�%n�B�Uj-7B���ژE,xgi�]��ȴ�C�W��oѓJo�W7׷?��ӷo����t����� �U�!4�� MO����L�j�]\_,��(;;;�s�\��`Tj�NS��v#�d�=;���{��A"�
�D�J�\{���t"=�f&l����q�/�u"��ʙPP�Z��) �~*7��Y�н�����H"c?�v��|�??��h7.6���
>߬�}�u����2&C�3X���rq~.�^I���M��z��o�嗿�[o� ��g&.�:Q�� 7�R����B2��_������9�t���v�h �_C���U�Ӵ��W_��G�rz�
Z+�ws�u�%��'�w{�DA��D�BZ�`��hk5�)jx�X��k�[�fY���oO�	0d�X��ˌ�k�g��<��t�����
ã-��ih������7�m'�R�	��Zh�h���%����]�nbլ�#�G�9���M�$HE��C�D���h,xe����闡���`S �4H����t�M�"s7Ҽ,��!�H�F8h߉<�,`=��L�q�@�?�*}���h�{-��{�5듴P��a����L��@�s(�93�$J��,"����}�M�&#�H��E����F�v���d�$�q�AE���ٹ����;|��vQ'ǧ�([�Ӊ�Y�:�sKȲ����k�J�.gF���TY��;����\!A�r��H
�xϔ����Ĥ��",�)�Ku-��2<Z#�niŁ�AVw��g�S0 b�xӂ�m�5%�)B$Y��n�W�<~p|� ��3
�g7{���$�k�ᆲ�y��2t�~:-W����{�d����E߬�`m2;��՜N�<LRJE�?��B|�e��F.�A��+���k%�y�r�ƣ#Ġ��z�.S2&�Y�W�	' Y�<�[��=�8;}ɼlm�}n��:�~�,�֑H#	ww{vvN�N�ߐ��;!�'
�Я��rNDk{h��	 |Le}�*�I����=}1�u�ʱ�mF�2�uno����{�{���`c��{����͸�`�ԜER��g�w�w$�H��*d~��斞������YY��:p=Y�1,�$��\-HH�`{>?9WVe1)䭆YmR���&�EP{٨^��J�n����Z? 5]�W�m� �t�}�jZ�+'D��2��+It�l�OA
A��N4ui���h2M��.�+�����K�K.��䌡�q�b��)H؜��#hծ�^*T̳r2��h�O�,�Г!Zf.��p��r����b�Pp�$n�9�vÝ�!��M�LY��۲��IE��g�I��*&Y�в�l��6�SZA�L[����d�]'ʼD��st@r�E�nf�X��6�g7��G65+�5�5�c��Ǧ��$@�����o?���G'&ӂ�����[2��x�l�m��/�5w5��ʡk�//���wdsf#
&��*;<<����������K���f	g�=���{�}�ZtI�:t�#U�����{���8�{w�)�%;(4&=�G�6k>��#���GO�^����/~���3��W��������hF)��U�������ѣ����ދ߾�6�Ƀ�Oh.�,Yb�[m6-w��ǸBm�@��
�I0�䲐�12G�ʙ>psw�p�-'e�3�Ye��],���G''��ǟ~r��!�����^!B��"���VB��v��,�t�P�}9ao�H3��0dO�+�hx֪��_�|I�0������7�i�1�&1X�\Y��bٻ`�A�A @��f�)�0X4Rk��fSy��B!6�AF�Ϡ�hJm��k����88�C�[��8<,8\F��^��"�J�"��e4g+�'�&�tt��,%�)���r���J_Ī'7��a�P������=��� ���d*��� �r������>����~��{t�B�̋���������o��w׷k2�����O����}˽t�..�?{~vz��-\,2��o��5�٨6QR )�*���>�0�n}�������?��^gˇl77t��*�9�����ˤ�4�W=a,�p'uQ���Ͱ��d�sD�����1_^�Xd$/HFrG�OF��l���}�yh���s&+K�T@+�@[����[A���y��C\-����eK�� u�pRb��!�yptDE>]��f�F����2�(�B���Q[i�"+�,�q�b��ެ�q��9�9P�����d�fmy& ��R�[�-�@Y͆�%ぬ�պ+J�p�I&�g�W6@�%}y"��
qKR�)�ړ�V�֋fIy��zK�3�كEF
��\
N��t�Z�����%-]3�߅����#���-ؔ\Kڐ�%W�n����s� �K�}���"K�u�ˣ*��h��ap���R��$������� ���Y�8�);14����B	�ԹI��'QtA*����&j�&|��5�_����|bC4WG��p��lj�J3�Џ�
�*hw�!1�1#-��M�E����l��QA��/��!0|�!t^1������bO�Q�O�^�{�ڜ�i&S:B���X�ՠ��^1���r�/��R
�6sԘ��D�ȹ6��e��+,
�e�䔘��H�z}}]
�o~g�B��<�#m^��R5&�j�(LVT����r�R�Qf/^}P�`+jQ~<uh�s{uK��?�c�h# :o�e�~&1�q8o2�;J�j�a��Nu��{G�{=m[��DVN� #�V�_�FOC������z2)� I��\��q�Y@���(#̊A��������a� �	��!��~���-�_��w&ϲs�Im/�۪��t��x7��i!!r�-����R~�`o�D���xS��E�s�aG䎑A�t9���pp@�B�7򒸜�����ny�^��r�Y�i'�}xT�9h}	��5m�AK2������tq�X�@ɜR��3�P��M��0��u��Պ�	��ȲBppR	�U?)yw8��q��9��(�쯻�����}�Ə9�+�-�DT-K82��(����I�YF�{����:@�q�r�$i!���X��� <X&�q��1*u�n �/�}F�J@�!�aCt�ߓ����NP�lY,��0&�h�x�nD_9~w0��a�=B}��wo".����
��9%X@y2[�ҍ�������}.=�f;���/��`@f| ��{��b�:�tw�Eڏ���[���?����ױ��6`��%f�We�&�}c\��AS5$���4��"���k��.xVh�.qIV!����~zv!Ua�wK<`�x>�]Af��z���Kh rZ�x�%�N���W6�ܮ �s�':a�+h�^*�_���x�?Nb|o��˘��,�@��8�f��^j&�O��\�vpx���{�d�^/^� ����!�	��
���at���d?�&CLY�u����8zGylĐ��Љ	:4�df#�t�񶿀ULN���i^P`DI�kWR:(�ȍ��A���7T��/�͡Ss.��bj!��^av�RԪ�N�H�x��̔ߢ�66�ܵNi��|��l��5�����RF���妍�l7f𓤑oIjg�&U�� �{�iW%p2B�N5�!o�m9�$ �N{�&�E>?h�d�mf(�8�qB�kIf,S ����~򓣣��O�ƈ�-nno����2,a�ӽ����	�=�j3
�=zrL�`�&�� �4it��0���\���Ǐe�w�����Qq�{ l)]����!��E<>�v�r���#&yI���~��=_}���Z�͈��\��G��x�C&_�=�	�֔�E�C1o�B%��K���mo@Ho��w�8�k��%�����p���W��E�!�_P�=�!������7i����	��Ͷ�U�fC/1��S dPl�:��t�l�(�(U�8V�ħ/(�U���Q*MJ�\x}|��*8چ6@�wɵZ/#�(�v#�t�~�+���&��ԑ�[m���8�4'�ц�ԥ-�Kʫ�ʕ�ۂo<d����4��R8GT��X'�K{������˗Mϻ��ޣg$��&�;t�#~�3�ht�)n�+�fH=6�P��I��\�Bc��+w�r>JM�4�{���*������?� ���z�Q��Yj�-��� �����
���'�ʁ!���!"�i����9�@3K�Q��Hѿ��w��!��b����Ս�#Tubsv~Ĝ����7�܀|@��i��.B�ӎ��?S � B�]�W=泩�������[q1?�2=\��w�x�L	C�<�C29Lq�9�;�!�A��Lyys˜Qe��{�IE �Y�5�me�A�i�o_���M�R�l�c��eU�Qv�u[q��8�)�ϰ?G�2��80j�Y3ʡk�<Ў��c|�+���� � ��z����a'��Qrx���[��1o�*Ey� �i��^=9]R�1���d��o��L�Y�u�Ȯ@��s��`�)f��JZ��1 ���fSh��y�R���%0���_4=]J��nz��$���np��(5��]a���N-��2ߵ��˘�g`.�.�m�"���w^+F�Ƽ�6>�c���
i�Z6��=��MQ*�+m\	5t�t6V $�rZ��f<"G��2�L!t\ҕv9�OF�z�@�YYzf��,L���4,�כ:��[�����u����HT�2ZH�����6�l��K����htA�+�=&#�pd-ޭ$Y��_]���[���W��g�)\�ۆ�[v>����;�͖�D4%�ӄ���L�7+Q!�nY zVS#�v=PZh����seG|�L�l�M�)Y�����V����QUEg�{��4���t��տ9e]��{{��h��l� k���v��~�88Y2��f��G��("#̛��
�Sp���\�}k��C[Į���{up�GڞO3��jM ?�m����Q�*Z�^�5��Y/������X��eEL��">�e��v�pD%�'!�p).5$��J�Z�(sR%B	���ZNXn���(��\'j$:�t�I��s��� ����B�F����� wy!ӵ;�)=~��=���%���D�3��
|�3o�g��e����T%��;^�^TU����`@΋�F�`h�f )oynavx����}�e������K���O}r`68Aީ����л ���Z��α5嫪�%���Id�Tg�r��>��__�!y<�Ų!mD f�$� ��d��ޒ�ZD�Xt��>{�9���+���2�A��b��R!H��z$<۵����G]�y{L�[��+ݦ��O�R�P�&f2hL�BB8U'�>G
�I �|:)��)�8��)�ɜ�̦�샶�=d���p�K�9ʤA��HT�(
[��3I�{�s�6#bp,�m�!W�ɫ*z7�Δ{tw�Q�A��7o�t�_J?֞Uh��x�d*	j ep/Z�Ǐ����~��_��?��Ӓ1�w�1%ru䷠�nC��F�̦�����d�2QK����������hb�) I�XB�E���	���/�/co�$Wr\F�5�ګ�4���V��zf4#�^F3����z��dF�1�n&Qd�It�ԂZr�[ĸ�	��6�/�	
�7��������d����p�׳F��i{�!Y�2Z1�`m�ک�������$l�`um�F���?<���Gף���vy���EXH�-������b�,���Jx�0j|aQ���}�����9�Zl�F-2���&Z�[#yU�T�X!�t�����#5�K��l�86��>U3����)�AE��ULڗ���3m B�?��#��ȳc �6}��#�^��i���7��:w"E�>0�`�=QtgO���#�D	Vک�Q"�6]�����t��+�6M��H=O���� {�@5�T{�s�Q��:�jI�	���^]\<===]�t{�	���匬
ɇ�f:������]������,���<>������=��Nx�����=�++�/S�����ӧ���,�q��͎��)�H�M��N�-�L���k'U�H�`�B�&9?��|T-��o�oKΏ)2>}P���~wp1�F�{��:)�w���/��Un�i'q��PC¦˔D��`%R��@`��#l��l#g���T�0*��i񾍰YW�*(�a�6A�5�T�������,���Rd\���*D�\���^��:}�ʕ�Rii}��7E]}��W���H�s�ޛ\&"�Od�~���l~����z}}�����g؛�G'��x��ūo�������w�}'@go��>�����qL"��:�����N�Q��I������/�r>̻$UDAbQ6۝�n,�^��|��P�&��@�7ޣ=�1J���K�$�'�I���|���t�o�lv/m����ܕB��{hQ�*)�a�㹢$歆Ҕ��Q����lYs~p�|(�]��:}�|�GJk؟bdZ�ɓR��dP����B�>�!{�$8����a'��nP֭�%:�UR��C�-�,�I~�����+�%\�
�I}�}�vۖ�z~6�9ʣ8���$�W;6=d�h��ل�;lo�r(?��K3*��`BD:��ɹ�����E�Sޤն����6I`P�۵�L�x�:<jh�i��.Ͻ�o�ق�0w�)p��F�~q�nF?�s�I�ɍ��ę7cP�nf.�t��//�u3����:uw�u�{#���pD��=.ԷX"O��S���0ڠ��!1zR�a-sM��2�I6��nyѶ���a�:9�$듙EF/T��);bm��ϒ>���ok�L�
�QE�2���`�x�A���xb0-��n쾋�p7VT�A�/z@-�n�@a��u�noWhsYUZH��ǅl�����~K�e�a�<�<�M�v̇�����@Obd�Mz���C�n�BԪ�YLq2࡟�	��p�m�P%�e,~>���!���O6ѡ&HBq��*s�GCc�r�oɍG���;����=�}�&�����4'-�!���J*k�$��W�N��T�~��
���/�28 ��Ƈ��]c����ТԖ*yApz��EHqدV�V�	W�V��&�F�w��?2g~mh?)}:����Q1��������K{d
���y�Eʢw�B$�U1�,�,�p%�E��7�cd�0���y��X�،0�f��R���ro|+ia���ُ�c�LD�z���_�%P:�`�9ug�(��h�6���!=p����BT��yd�@M���I:�`�)ϵ�l~S������8~.�s���z���, ��y5���3�[h����s(G<�^�ñ�"ϬO��ܔ �hD]��L�r��]sR;�뙻+��M�y�8 X-T �Ȍ9��u��W[���L�����
4ޙNr��"e3�TQ7���k�\u;�g�A�]'Q��Q�q~~�o��o!�����Px@��Z���tO���f����d��;e �S�3e�Xih��u*�J�B��dpl0A,	��J%ۡ*ez�NxG�y��M����g�g��+��CDǫ:�e�v�$�Z|Wjs3�r��e=�^��R+��9<(���K���+}���������T���ނ	�����9���0+�J~'�u<���-��Up�p~Q�j�Ө�f�*��gJ��"��|̳sj�90Z�e^�9��
�ym$b��'�v�a�!��pЛSW��u�T�5���'�����Gz�N�)�r)f�������B���:pz{�š��g���vKX�y���6u�,r�ف�4��\�s�<es��$c �ń43�\���}a<�q�L�Y�A�nxsA2H�[-������?�C�@"��z��w����k��ZDf�"�����Y�U4�S��U�vÝ�!C�G�.s�(�/9o�"dk���>�y͍Ś������EϞ={�
�d��i�"% Q�z�}���<}cx�ʑAf�n~���PЀ�	����l2����O`�4�)�� ?꣍ecX Fl��nE(Ǻ�5�C0���Z��H��>X��X|^������Kp�ӒއZf
Ѕ� ��UP3�����8Jz%�A	�����n�:����:�`��v����*:�3.>��Z���TE�Q��=���u�Һ�����������Ǧ�L%���*����@���U�K����zH�Q��uu���U�x�I���$h'�O�<���x�ɋ�/_�����?����5��6������Q�����������i\]�X�ݩ���2-˃Y`ʂ���Ŗ�5J����Pi7]__������@T���lPDUe�6�R [#�se�&�� ��X��2�5��6���v@��w؀P�H�gP\k�)�fzA*$^v��������&�и�M>m?�S �m%���#�0��F�Z{OPY9���DU#s���kI9O�3&�����������=-�v���S�z���E�N�ET;g�%{��9z�Xl�s���%�>�IX�a��~G��i���9z˒d�n�VX�`/ M6ˤ~ǌ��U�Y��gt�CVN$�(�_X&�Μ��-��b��C9�8l`v��*lʇ��,H3�a#,#Xd�iY�ܼL:ba��IMy��T���
�9���"OW Wj��>ڊ���k�+��[�j�����f��F�~'�y�ug:UV������.�^�r�chf(5�)�B� R$����E;tZ�54 ����]Z��y�НNj2���+7���f~�v�Yp��&�TE	;bY 3g��go�)����H�O!فU�ݧ��&����85�r%ń�������l�"�,����Ї��vj7��5_g���>B�W�(*��d%�5Aŧ��?G�L��7�I/�fא��/Y�?�45���F�hH$]��U���(�NFf��ڢ�����MR#������:(�����ۦk2�M�&�T����|�T*��`D���L��F�7��FV"��q�$q��p����+�=�e������,�6F�CzOOn�J��㢰 ��<���V�]�<�K������%��1a�����Ƨ@aZ��"��`� �������(�(O,7��J�݇Br�W��s0�"�5SN�*��p>e_��D��B߃�27�xb:����S��Ǵ�Ԯ��^� �1JbM����q[ �T�)�N[�e}r�;�lƣylP{����Mu�*�Z�nR�YJ�Z�}�Dn����(��`p��؈$��+&�F#m1�s���@Ƌ��	���5�әA�΢tK9���3��G$����MNOAa��،ơČ"��V�SZ�`�p�=�Bu{������Ȕ��f���r�0��C�ƆN`ϔ�w�e�1�[�EOk`g	��{QN݅4����\2଒�R�������1�`D>0�"�����t��,�Y���M��p���eqR�D�p�"��Y��N!:�ɖ8���Rt(S�0�	�,R����k>۞��d3!�á�v�ZH����#�!�|��*-��Z�9�UO�",..rf��"^߲���kXgKԥ�<hJhq-�l�B���ŋ��|B���Ͽ|�촓�i������#�=l�^�޾���g���,�������������g�
�ÑL��F��B�**�Bh��b��Ue���ؙkp��e
��r4{:\ڎ�[a�����?E�O��7�7�w��n�ш_Q;��A�F�:8v�����AՁ+NR�$�Z�L+���(�������[�!����@+��C,Es
��5�nL�"����J��T%�B��,tMpCh�(�C��F�2uzU�ɒ u�[��#��p.0��^���-��2�c�b����]��B�Pv}�+�$���Fm!4���
�#J;�EK�kumJ(��+(���я����|�>�b@��`{횊�F8�I�In=�w\k1e��s��ǖ�Z��%IȂ}��qb�E�Ħӹ����*��Xu�F�.�^���y���HI�
D�5�a\-�e}&\Q��X���d���ˮI��S�ԕ�{��y���/��A
��_߿O^^^J	m"���M�5w���X�߯hȏ�N���0�/�/o�70�� X�m4B�	e��;5/���������<)꓂h���	m�-��\�rw}���o�+����ٽ_����˯��_>{´���cZ�h�L�_������w�� �{���xx���h��|�2)��m�e�^.�J����V���)�do6]��`P� b�����2��?-�Ԣ4���(�k�����]�@�c��J�#���rqT6������~�La�R�Ӌ�����sm���ZWk�	?[��F j�� �6�4�1X�!�Ը}W�=ک~�q����z�v��G&7W./��D$8�ƠSBm1�IЖ�� Bu�.[��J����2��s(E�r�z�����iZ�P��ӧ��+T�U��<���7k֪�Ĵ$��L�J{�b$��o�M!�C�MG��m�ê�C�;��~Է�n/..��!���� %��K:)�� ���S;� @5-�A)J2�����
�V:�$,�q�
��ajXX�XC��K+\0�4G��iD%����q�6�=$ qgK%jG٨/s�x�A�6�ƺ�^�����h�E�������у� �)��\������WϠ3��7�D�2�!u���p6�J�s�Nс$UGUY!�S2�>f����L^,���D`��rh9�#�L]i4�kLdT����ԇ���O'e-] �eeY8}<�O���i@3��C�A�;Py[�
ç4 A�` �cX4b@(������m�ɤ6K������H��?=���F�B��)���� w�/�*%�O�p�����e*�LFad1�"�4��K����䐒6Y��B
��wp��!N"���Ş@����hh梉���lbW�ǆ�����8]����3�kɄSGM�s�X��ڍ2�F�������A��8�A,R#��jǌB��:l٥\�J�����+_Tp���:�����i/�8<��0��e��"����@-~�u8�`��$����y�8r3Q�����4J�� �=�'�X����G�ޥ1�k�'�!F�2�Y���om�M��W���Lx_�4��H�E�[.��]��%ʒG��k3��������Hf+�����ߠm�Z:��2{<;bzS���GX������+�ROޣѪ��W��0�����j�tD�]�󉠑>'�x1�{Jv�a�}��0Et��U��4�{@�񚌩O���Xu#= �!����.%/RY�p�i�9��i���7"���)D�u_e�W�����zc�?����B�=k�����	;���Y{t��5���Mqa1�����ف�� �Hm4�LYT�w�i��Sn�PT^|�G}���gسRG����|+LJ'��$^�,f���#]���)�$
;�D�l�f_�^�Ȇ�)&��c=��Z^���t�+�����$PR�{���v���I��t���)�S#z"w�6������閶o���T��q�5��]�Ǆ��5��ƀ�?iS���m�膏���A�d}��\UH�W�ԩ�N=�3yo�W�����N?@�aH��Kzϐ����f^�4W��W77��5�@�7,9�L��s��i�pm�
�v����s��z�7o;i��٠����J"�wP�+���?@�]��𜟟��|ۧ�ʏ�3�I|o�W��UI\�TY��=d� 2��޽����'�
�hl�www1/je�t=��A�v���Y���,y��N!�T�
�S��\�Lj��z�n�Z��IԫD�()jKhT'*H�2�`|`���<��پ0�{F=(� �[�GrK��4���2��Ƴ��x�>�!�	{s��LjCn&j9.�1̴��>��M
up���URЮ/�G�^`W��K���I7���kФ�%�
'l
pPE�Όlm`.��&�_��LQ�Ls9�'��+�D�hJ�a`�'��%Cd���;Hs���-96��c��y��ț�Zޯ_��2F�	�f��\ڍ9-�������-]
�}�P�gM��wq	�׀8S��$w����i5�<y򤒶����v5O�U��`���F�S.��]��/��(}�Oi����]O'�B�/�ᤙ�5 9
�MÝ2�e����
����S뵍x��T�\�u�\��
r-ϲ]��$9$���a9��A�,�ǜ�_�C��`��_o7�<f�q��́	��.���P����t������}v�2��1�F�����M�my�1e�ٴ2M�<*��+=��%��r��  ��K�y�'�L�� �r����Ryf�Ȱ8��^���?���a�C�p�����]�%��'��"�A���;��Z��o�i�k��8�^�i�+]���hD�`(� K�J�!�/m/c���U5"jM@��}ۅ���i�����9Zr��V@6�g���l�Y�#n�G��,����.*a�+���Q+&�l�b�{��ݍ�����N���sԸ��^0S�<m�W��|�Jn���	g��}�,Qv	�*�>����q�ʾ��۷�^��L-�0�+�܏цekE_K�ݝ�A��$k�z>^�V���o1?fk0a98'�$���:˫]�Q|W
�~xr|�^���2�#�ؒ壹W��7�x���X��WE9)�2��"��Ċ�N�J�1"�=%/�ZH���ٔ���;�],&��,���̔c'�L�$kU�j���i�U9?_��IG�l>��eu�7hk��]�=�m����r���m,c���9S� [m��z8\�W$�q�j/m���kQ���LΨ�U$)YX���5և�"�rY���,b���`T(��K�\+�С���33��jF�ѡ`���!��Z�ݾ�Xfp�'y���$�� �{��2i=��ʽ!���8����6[��X�\�=��ȑ�Q��o4U�B�eX�
m;���8W�V@��/��¹MmI@�+����@���q�ㅼ4ϳ�0V��`+�r/���e��p!�׈t���0���v(3�����l>{���]AB���Et ��E��A��:q�ـzŤ0�M�&sn(v�����~\j���F2�����l��[��N��z��,p�"4�벒��+Y{LN��*�n���N�l�r�[A�LKjK�XI!�f1:=� �}v�>{t|@O7�zQ����	�g�Lq�'�y�v%Nz��:�/���������Q������A��@S_s���	ҭ�l:�j;�3��,'��}t�Gw`q�2K�Ï
��#PBA�PQ�ѓ�D
UK�1W}2����}[����lK�XF�\��|���1�EH���m��ʂA���iuyy�^��O�)=˭n��VV��;�C�v�A�y�yaл�i�&1G�ZR��SL&�n�nv�^��]R;��`x�e��!Ɩ|PG#CAC�q9�`�AX�Hk��E#]�)�ku�f�'�0�2(�ws�]����1��(�D��x�c4�ي1M�eQ���;Y������ �.�"���� ��Vd4����b�������Cإ�%X#�L���S~���g`���� '�d�/i�B�$�B�e�ehOE[��U��C��ׄQ�X�73��C���L��B���f�ޭc!id?r�@J�uT����.Z�DAl3�����_j��Q3'��+󌉡U]��4���S�V�ل��_�R�f�=�O)n���F�����m�vߤ�[>
�/�.��6�w8U���(�[�5<C�8]�2?��kw.
I�ee1�B�u�FATS�-��U)%��&�/v�$������)�X,O����m ��e)<3�"�_���(���!̽P��k�UD &�Ȃ�z1
hv{�c��v@�mdr�8主{ ���˗��,ӎ{@A#��kkOĠǧ��i6l��;�xC�,��55�$n ��敮�A6�K���_)�-Ao���A*�������lp2r��F&|{��PY9!+�J=W����p�2Zұ�r�z��F�Q�@�Dd�(m=���B�hH��F.�h&�4�Ez��큏f�B��D�gg��4�|Tud�Z&b�V�MS���)�2��!����Js�w��u����R+i���9��Lj�F+��OG'I��e�`����ڮU�y���1�c���1��ggg�0���As�a5�~��ׯ_�E�NNG�dI�Ӌc��*+�V�eadM�3釷o�5M��d�P���s�\�AO�g��ÁbQZ$�T3�1szrvtz��/-]���<-$k[NX"`�oif��|y|����w,���v��.0��,S/Z4S�G{_!޲
�e4�%&��|Ԡې����Jj�wRa6GLb GcC�� �6�y|�f�����Nb�"=�=�	l��y"S%���|�L���-�u�^p;��fn��`U?w^;.◹
\F-TGz��� �h^$V�%�WH��v]O�������FqV�/�	3l@�[['�L$?̊��U9���Dhs�I�v3J<;M�_lHa�qfaЀ��d�<ר�ͥ�������7�|sz~��_B�#�gbV:)2�Q9�v>&�m�'�ˣ���
<w��Me�V�ٷݖN֦��џ��2�x��[]�xy4���uz�����	����U�[I;.HE�1Ƨ
��h��D�d�d���K�
�F��\� RV/�"�U�y8ͣ�k�3�n�����"����@!�"�D�7�.��Y(S�N���űeC%�&�f;��muA70���l�)7_�Ǆ�c�_K�
㾺h�=���x��E�q�^#�D��9
�c���{r�0z�GM�ph_�_�97@.a�a���r`Z�>���Kŷ���綧S�X�G����������������Dj���� �oM��Cϝ2߉$C��b�Յ}���{�i�;H��4��S!���ř�bO�>++��ؔ/�c{uD�o��3��"g��m��ۨ���`���#�# ��>����0^An�p &���p�� �z@�i�Lô�Ä��^�O �_�zm�-/� ���E�O�<#1�^a#f��ne�P)��"�Ȧ8յ�9�M'I���KQsR=*4�~Ǫ�rQE�B�$��[ȷ�DD1�.)��9��z���=l�ZA�ne;�H� �7�����F���L�����cܓ�G�Yc�VHt'�W��w�eSD�L��a�M�T����R�RMn�IQ�`XT.�Ч3R�97�����.�P��P��VI<Bhi��b{�"\;��o�m;��2Xf) L��jX5##Ϙ�Q�C�9'�N.n��*
�=`�f2���@!�3���Ͱ�ד����\�r�=S��٦fE�� A�2-�Й����&��$tT��Mᓎ�dp��n�����l��lw='W��u�h�{T��*[˦���6q^B�sxm���T@p������|"jE����{O��I'!8ð �F�:,������0ty^���Е�<�
N�9/�GB��EK����l����Ba(�H
�з�mǈv	u�Ԫ�m=��d�e{6�,�SZ�,eH^��G��_J'�Z�-T��Q6��+�ɼ�vZ��^;�8���~��7Z�  �Cc.H�0h��|�ށqߏ�.�<}���n2�7-1�!���0�����/�My �L�`RV:����RL�6̩��]C���6���c��r����`[�1e�ڠ�hߌ����~4%�E��KH�P��M��蔪D�H��N�r �bQ�d��r�oF%��te�ć�d����ǆ�uƭb@�-��]{'�H��rU����,��G�Hn��)�wP��A<ӼH������I�-;���ɛ�'r��#�d��,��pe�JF���}�����P� � t�2�x�ޫ@�������{�#MjZ�BTpx1�֎�Z_����S�%�8�I���ݻ�B?�q�d ��2�#�X	���JL�(u���LK�m��Q��E���8��5���9�z����*Re�\|nT�g�X>*�BPj����٨�1w�	o�K�Ϩ�\�+�Ո~��J�أ`�G��8�뽊nc�ya{�A����ʓ�T�K��X]N�M��/U��0QT����I�$-	�ˇ=���h6zg@
)۽S���1�\���⟰��Av�}�� ��i�D�|�>}zxxHN8~�M�4���(b��F�������W�^�c8r3�tZ�o޼9??����_~�%�����r����f�9�ia�4�������vP�,�4��"���>Fh�ŷ�4��j�4���M��O�Ӌ���.����{�) F��"�����]�oAd�E�]nQ�`@ ��iM%=#7��������T�͎3;ӝ�������T� �!>md�O�-4���O�	`2~��bF�7re�a���h�J�G-�jU����μ\ħ����fX�¬:�˪Q�q�a+����|x�=<n������a��Q��^;��Y:��g��*3׳����={�B�x�����ރ�u�2�e�� ��[jO��3�v���
��xV���Ib�<3��&=�V�_�� h�EH����j�,���fV����u1�܉��˪N���O4����,��{��P��b��-ժ�b�m�>
f�Nf#D>j����2n��1�XH�D^3�E\�� f��3F`�זL���ʶQ��A��M�-~�x��uk�ٚ�3=�R�#�|z
�Wـ"�� ���|ž�W�.�[�X���j�|ԕ�T�p�A��mga)��/?�A.jV�Ʉ}<�/q)��^0d+�F�eT�
(ǅ�I�w��˅n�1Zi�:$m��:-Cڮ�YQ1l1-��bZ�-�}�LH�Y�z�7�W^������M*�Q<yE͒te\��U2t��������e	��.�ꉓ*[��>|��g����ۅӊZ�g3>���|R�IGa^&h��V�q�d׊�(0X\�������
Ժb)/糢80�?�"��'�g�c'����.�y�,�Fe6�b�m%�wdm'���L�b�۝����Rљ����tL�wr�dr
Q�
����n#j9��*���H�-ҧ��e�D�e�}hf�D�Ҹ�L�bA	 /���Ʊ S[�5��`�`��B���| Sl�dI���,�H�ӝ�o�^�@�h�`#�3�cè���o}�G;��6���AސQ$K���_\�;|[��K!d��K���;l�q��5,ȁxόȎA�Bh�;Fd��k�3��Z���ܔ��t����7�zө��9�U�6�	O���A�"�F���6E2Y���	.BO9���|����I~1��v�G+�O�]���7̀��0r��@�c9�\��a����-204]5����&����{����Y����.w�#f ���%�@�f=���h$�_x�I:)�&�=?2��+i�Ƃ��S��Z���-�Ppw�O(`>8X���M��Ӝ��*�t�~`VZ.����wC暖|=�R��Qb��ܗ1��z �t��^��JԣZ�� �p_��	k���b��1r�V�9�J��hF�i�b_�������K�X�z�/O��)G�?^���Vd�O��o޼�ɲ��ɟ<��f��Q#�ٴ])���	B�-H\�� 4�^�g#H��	w���r~b�Nh�ԥ@T7��*'�������b���o���<?�����p͐s�i��������Ƭ.����CrͶa���T���={xt8�~�[*Y��"�C���3(�B��Fo��P�LI1p5� 7�t���!v���Rd�5��>4��O���f��A������v�����1�L=|����)���sE5tD��������\��I�"25� MS����fG��Й����ˤ�<��م�HJ���d�x�g�B5�+3����AJ?.�����@�VMMUf'���*V42U�0��[!�q}}u-
&)�������<��M�q�#� }�\���p�I�Ďx�r+���nê�C�">�p��,颦�*�I�ZK� K"�� 3=�SW�����<;;�cW�)߉0h;;��m�ݴ��.Υb�`	s���ju�<�����=�7gN���j8�f�[i��S��U���͇���!�Wቓ���W�^���ݻw�]�f��U׷�ͼ0N�Jl��E�����>$RԆL^B*��ŰX����Wb�E&c�>ES��p�&0�H�4YZ�An�塸����P�a\�+U�"����PN�k�/$#�0����ND|���Hv��R4h�B�L�i!1�V�X2ʳc��"z���XJ�e�X�: 맏,@�a��N������4V}\�b'�1C����F'y�89��B[s0�fT&�k�J�"�2� 6�po^�
!�1��t�S0�}YR��j�����[�*嫱pv/�"I�$���{���Y��B����22������v��l��!(�^p5�PQ{�\j.��"�����bq���ň<5���4tD6m�cN�T��e�]Y(<|���������7�|��QP��#o߾�����������������7��ʏ��C 'PE��'+��0��Z&.��&�����zUof����!����G7�A��]C��9�ӟ͚F������B E�ZYW؆t���cڪt��g'ϟ?/kVQX��UX=б��� bl�
큋�
�-�G�1f�֘�c�����Y�	�9(3#ͦ���*o@��f�dM@�\�DpW4�kn���_��Ky��$��@Nɹ*U����>Q��`�2�V�_�J�5y�m��,��xo27��P"��D��S�&
��TX?���#P����=x(�f;cd0�>�� ���o�T�Q���\`L\��rz�o]�1��VjӪ`�U���1>@-���(F�-�c���C�������v9�)���K4pTFZM�>�� �J7C�vyy������K�Me=���АG[c�*bq.��N*0���+�������+�h����_��A�EV�7�^�� 12�S��h����_���=|�9
��~)�����̕ʹp
���pr����hI���&�e#4g��3L�)| $#���a��qN����r�ʄ�3�h�p)�0A�J��Fy2�1�=����೑�7i�k$����d�#�R;|��y?��h�dlO	K��Ç���\��.ck����7�=Ψ�%o���[ڵR�\����a���bZ?Bb�wz΂����U�iUFz�V�_��j6�UH��f�E~h��0$t�'/S� ��H�R��7���S�?����v�2�hjk�9�
����mA�$m�� �Q6j�sG���<�UI����R�^��L���N۱��)���*��յ�d��}bdP$����˥BټO0��-�ρ J�E4�
���'�����j����^գ��O)6�Lg9h���d@�ݝD�P�DV�6����%)��{�F��1|�u���K�\|�����"K-T�y��	.rM`���*�R$x]f獽��D��e_mO��ѫ�iV_6u�H`���NV���)w��RU�V��� ^N��z�y�V�Ơ�ǥ���_j؝A����r�nz2���L�����Pw�I�囱3T'�G�m�c�	Y^{�:I���e ��ل9�N+��g���y����%C=�'4��oMU<!�j���K� �2�t�77�E�̖��S����5��}��:Ra�u�5AުZ��Y����2�:�ٔ��^\�������yoӳ��Ź����
8�yr3��X	�ʜ��$C8���,�����o~�4Tr�r9͓�لn+FUm�r�D����U\2��;^f0���'''d�~��_-�,SM�,�	Y���gG4,��-0�_��
Ixa!m]�2Y��F"�B�k���Z�W8���l����N��(0&2��1]�Ι�����%<��%�U�~�J^>e�"�44�\s�p�^�Ri�Н�UN�%�+��'�h�>�35N��E*ۑ(�Y���)�桏7ғ��uP��?��>����	8�Z/�H?�a���#0Y.�z�F]V���E�={��������]R�>K]��T��umœ��=2E�dͳQ_<�3L�r<S�Vˎs�e�_O��2Q��� ��̹�ń&(���%h>�qHF?c~�����p�tE{��Z��4t���w�ry��*A��I�a�T	nRW0r牤O?��߱��m.//��POp)/d���v�2�=2���4K��F`�DH����e)�9�K,<�w:��CY�E���ؒ���ɒZ�~��v�~Q��X�g�1m2h��y���M��-Y(�T�kJ<Ӭ~2��!\Ln�Yop�AT�3M}!��n���ꫯ�ж�F�����Ç�8v߭«�qP��BP�0�{�:-'�
��X���~>��m�xIx�RU킪��#r�Xf���ї)Y��ГK����$b ��7/QQ����љr��!|||$��'���LV
�{-ن�
j���ާ��Q�	c��T2¨�⠂k�B�}<ͽTt�y1mCZ��hi�4��̸
���i�CN����5�^�b���w-�7�4�'�,u��
p��٣���}ߕN�dMe�Td�+u�Z��?*[>��L�v�6Ĵ���pG��0e8ȼg@b��Ɗ>���S�/Q�p�x�!蠭��R!}��㊢q��Q��c)7��$��`�0���-1.9�~���:�d�7��-}��hyvvF1����f�p"�i�Ҽ���y-6��=�dLll-�2��b�D��P]a�Y6���d9U@�$���-��,������vR��D�8��'��z}�`5��y�h�ZGS��2C0'��r�pBc�pP2�!�VYee�X���V�~�j2��a�b�7��ɩK�Ѹ,(�#�M����l���5�<����y-8���E�G��yҷ�,ӌ��/^���'�O���ۦ�$��ș�&�*���q
.GH���K���۷���O�^Ĩ�Ǹ�w��׹�QI��fu��Ln[)�.�U��y��딖8(O��G�k��/$�At��]Ƅ۠��iw��H�٭!�͚S2��!ĳ�A�]u��1����ikϩ������;N!����{i���F\?�{_T8������N�p&� ;�����{F�m�.���מ@��C2��.��I3��y�tZO���s��͠��68���cI�T�GS��U��8��O���M�I��vCc3��
����0F�������c+����i�yB.����������t�ӣ�_=���������n:���|^���{Y��*�H�γ�/���tR5�U�ϟ�f�KnǤHV�w�p�P:�'�"���N�˳i��f2e|���Xc�U�$
���ؓa���P߅�V�(��r$�f�v�F�닀�X��p3�l�zM"KI�Բ����r���u>���}QB1�5�$�Yk��̞�q�ݨ��͸����nq��EZ��C�P�۾�͖>��Rp�w�j���;]r�:�>9��"9�K/���L3��u:ްU�N��4x-[�1�O��r���O�f��(�Y2:�}ν%�#����Y�:�lp(�!ӎS/�T���/��4����u�G�rL�{�����|����m(37��l�A���1,�p�!:�Y��|r$��r��v�><<�䓧r��/Η�D��\�5ȗe%1nW'zu= �
�n6��j���`�(���W�?���RFl:%�/E;��:t#)7#�lMn�d7Q�dl1�w�d7��I^0��ٲhw�v�n��V�_��:&�o6���3����([S�/
�.0�)Φs����(ܮi����V=��]��P�@d>�n��]������\�㯒�q��].���L�ʹ�h�
��)������#/a���oNOO�c<����P���Q�Ac���|�Y�!�5�RFƘ(��,�#��n�;#w����5��-,y��~!�l�i)r�8�]�!.r^��	�Rwg���?9G�����b描��D�ՖkWyuE���h����7L��\���]�����m�Z��,���m�C/t��>�-6vX+:�e ��h%e��B����ݚ�̗t���p�4�fl�.��c��gϞ��@���	9\����9h��N�;�(�������p9�0��೓%��`!XO��pX$��1D�`L�Q��2�l�t��i�]K����jSe��h)+��ͦq�����UT��_�*�RX�ڔtF�b�]%�3=%�2z�����p0��"��\�+��ɓ�����;t���z>�Ԡ*@K�IĤ�@L@���C�-΄ݣ}G��g�٧rD�.Ȇ��ãCT�q�o#�8Z�����Ԇm-w�3��u�[ɻҶ~rzl�(��S�qZM0��0���J�]�x�@/G^�GM��+�.u�>=FH֌V��*+���t���|>�ч����vM�L�,��YD�������]]�$4z�������:�	Y����L��h{fmG�-�(m�2� c�|Z`����A��5ԕ���б�ِuE��nh�|�y��Օi��L�K�" �Jk���,W̆}�YA�TI&�-�t2�Ɯ��
ɵe�0t ˒�ө6?C�uj*�V}�HU��6�S�U�x�-�E8�����5�]��R�b��1��Nn�}�����@'�������_�~}uuEÅpZ$�3nHs�]�.�q�V`%\�K�"AR2_jp)K>9�x"�&j�g�*b��  ��IDAT�)���������(p1o���Js�e�Du1:��\�a��<M:���X7�\�M�-zk��7���� ���잚���Ǽ�	$��ŝ:�#��L��ԚC���O��5��X�߄H(��r�K�iTr{�h�TyRE�Ʌjq`"rKh�$��E	���ڲ�f�����,��n�5S��e��[j�;�X�3\D��R����SCCx?v����}?&�������zީt�xaTɪ̖3��� {�R!QKA���?�|yI�����bZ���w~`���"߶����d2c�Ndv]��m���h6�"��|y��^I�("�Ӄ�zʊ�d���W:��^��7����?j�ھ9(�8��2>�7R��6�7?�ܑOU�|:7���^���TY꿑�	�P��cR����F�%0���is���a
l�d���z7�Ғ^���pT���O�0�&�
�s��k�ځ�5a3��?D����¶��Rb��h�_�J�������0n�T :jw|2a6���BQf��(��@�A;�M�sJ���DGЭd��A�dچ��>ř6��Gj�N�TxՃ�}m���}\�z�9��>Mf��n{pz�}��n�5�݇�n�hlV�̒�b`]0N2[�3@��#T霡x�����-����ӆ-�%�"%o�,���q=r{�����v���,%�Q����tΒ'O���+�4��۾c9i�­�m��}@ZI���+��̰hKz�DZ��C�6\\��R�Z�i�vռ��i�c��x �7.��4�SXʒRQ{a�q߿�;�����)��<�.���5��ǥ�b����}E��T�!2E)]�������H��O�ĸfRo�z����CA���53��6߄��n�ȶv`W�,�{d�3	�t�����S�Z.��#����T�aц�biڷ;�d���瘆��K���)vt�� �FaX�|34� c�xP���l����Oi��>�3��j�ey!N����C�d���F>�B#���>�l#δ�}�7�#|�V{-A��9���'���jx��X&u���b�Н6����5'�+� ���w�ICwu8;��|�=n�Q�!7˱�Q�={��FQEp3V��#9�r_H��&6�C���NP��U����cP*��q��i-��	.'9�l �塘�Q=���}����یy�<e�KS���v�8%KR���
������t�!hF
�-�Fy��o��ͦ�m��w�G�jS��m�`��|co����!���LGC$Z���t����\���<к}x���)f
������a��ܤ���p%��ġ�h�3�>e%�D"�P[R�Q٢{�=�n�`�
�JaL:�!Y`��x^�NY׷��(@�ܥ(�����E�7؃A��Xi���G@b������_qNXb�(jY��Sy]]_K�dѡ9ȼ�O�؟0d4.��R6�f�t�+���6;�Y�7�P�����??8�b��>һ�իW�����oAgp3x�v!<'Dc�c�W�f/J�r�K�v�b�) :S�e8�1�g�?��ٟ�ާ�2����f�����f˒�N�	��t�O�<��o��ԱY M	l\
)1�N�%�����$>��E�R����R���Ɠ���d��̥ Ď[s+�k�����������J��N>�J�.��w���p�p	�	�v�[R���J�9��n��[�H�[!��.13/�(���,����C���
��u�&�OZP���� ?z��>�_�~�:%��{�\�ؓHQ1qX�|��NN����w�E?���n�O��O��x�ڞV/����Y��)IGg4采�?|ؔ8�I��K���UA�p�Qc��E�s�f���H�y(�/���k�����L���`��Z�w^u��f	���=}���1�U��4�u摼`1�"��Go���ﯮ�b���ڛ8����e�b��B��D��[$/��Z*2J��
QeӉh��b =9K��}��Y`B����bn>W!�\�n��rQ�\C�]�1D�F@�]�8wZ��|���C�
��J!��E �ޥƠ��.mϾ�F�d�ɼa� �e��6�2��R���ܾ7�	��b<���e�N8$9�����EK@n�q�%8фx�B��H�����"EBv�ȳ4��N~�6���T*����5�J��;�k1G��L��l+����'�(�&7h+�l�A����h��1�����ҷQ{�cn!�|:�|#�_�lʜu#�٠�mj��q'c�6S1q�U�i�'g@�w����U<O�K�GLSo�F�'�0<��QIW/1^��]��3�T�9�/��* 8�G���.�7����� �P�Aٻ�K]������$H���OAi�cml�� Aͻw�~�����|c�#�]4R
:�LS�D�������%��^���t�9ȝߞ=�3w�����:VY.�H	�����gn��P*�>]�ɢ>}�#4*�y1\~슏!�q���� Evت)A���Q[U`�̔��������f�r�JՃr�����lSO^�������e��`���q�LC܉�P��X����Ω}�2#]����P�m�X��/T\��j�q{�x� tZ22�٠�\y?*���n��k���1�~��Y��(jf�x�(�$I;׌m� �$�W��"kh����]�������<�����Ǯ�P����bn!!������"��P�=Q'E��)��� 8V������:jR`�Y����v�Z�h�*m��2<h[�����%L)Ɠ%�D����}k����N;�JU!�H��<S��,*L�KB0�錖�!{D�x��u��*�e��5^���;T�F�b�8-�e�(�6���)i�?���QP�t�����Ѿ=6/~T�o�����1&>�V�F
[�Q��Ɍ3��D|Q@�1�֫ά��gb��������R�ⳢYs������v�������Y�?0?�3�TR��oO�>M^�0FL23OHpe��wgy;������#���Q߮�KB�in��*rV�~�O���ܱ)�4êz��O��EP��8ޝ��Ow�slcS��4	�k���c?��G)�B�{�*�	_�p:�rͱ�9���v۷E{=�9���5���vAq��ྌ�,�YvleD��T*�k�9��� �{9�
��Ж�$ �y�8F8���u�e���i:6�0���>H� �o�R_X]�{{WB7jV�9�H��c*n-e&��1����c4a5���w�5�P��]W/- � JC���E�'Z<f�猥N����k~�}��\�*�y��/�?�����y����O��f{3�L/θV����>���~�_�(��nӔ\�K�@s�ۺܻ�±V]ۅ~�^�L��~�NU��U=A(�����ޠ@�A����aINC]�L>�9��r7t;&��YTk�n3��кӣ������bR3�k�c7�ԓ� '�}�rF�pzrx||L�����u}7��R��ͬ8��ܤΊ|8>�u!_�?�q�ݜ�O��~�$�g���r0�x�1�(�I=f.�)��V�H�V��|���-��t��ɓgO.�Qk7�v��]"����Q�]M
w|̲)777����K����t�2�*n�5����UQ,g��m���q���Y"������U�v��]B��֏{M�)x��	9��^��5բ�*}������?���hs/���s/r��咥:������5��jRKfh��d1�J�0[.~vvzHN��bIa�n�9>�m8�?����oߑ���;���ց��=ϵ�b������g��GD��iPU��Nh-��.L>Xr�(��N�M'����/~A�����+�����ZǪP������|ֻ[ZEð͋���<��D~��!d�zZ��Gg�B���Dr����[�3x�Y6��,�*�F
@��㸝��J�N���U�����,??9��VWD���O�O���g���V7<_ƈ��t88�#�����/_>�Ѫ5���o\��.�����㼘������v���T�q�C4-]�z��i.
������S@�\.�O8�G��L͋O���9�/���|Y��f�<�ȫ��74�5m��Y_Fr�ͯ���fw���?���rxKޜӐ�H}�r�~FC�ûK����̿�}h��hb��0�ɳ��勯����o����4>�vC[�E볶kh;���+F����aǝ:#.���خ�w�rn��։g��#� �
�/ݤ��{�i+�Atrqm����@�����z�p���p$N`2�R�r��rJ�ȥ�k�UwuuE�y�X�L�g����:��-�|��`�~R/��g�I���/��t.������I{��ʽ�cfq\�<�N�|�~_"4�B��5�(�}A��\*�<;;�P y_J�K2R�dZ�l�"1��[��<n��;Hg�I�O�u������I-]�}n�t��@�@8�A8��Qt%��Sj��1"`�e��1p�|K��B6q��v ��4J4ÅaD� l|;d-H�C�|��6�倜��+^S�V=�ׅTq-��z��3�i�n��2��$M\&��dF�"-��([���*���UoB�	 X�Xr�þw�S�|A��,-ر$tP�"dC��1*�$d��fy�pRp������]�ƀTr/z^Li�ӱ��\X��3]�~	D��΁��i˰��\��=<Y��ʹ�b�YRm���'%�&I|�v���/..��[=8��g�e"�ǲ�d>�싫�K��oo~dj��.ȼ����q0_��zd`�t)��t�M��o��`���W(���2�z�v��@Q� <���^�����D�/x�߱tq��R鴥jb�M�tl���p�+yuQQ��b-{�|!:� C��m[�EB+V]���9�t����J���bX)��aQ2|$�h&v�j�����c��8�����Pn�e�7��$�Tn��M��"�y�c*P5Sc4:�͔��#�a������3C-�ž���C��������9��f�dy״��h���M�LX������|O+��&��'��M�����LܞF���u�*ҙ�m��ʇ-Er�wNU@��p��>�Mw-�C*���]LX����E�h��c�e&��S+S&:,�%���i�����E���[ܫ�'������0Ӡ�x (�|m��D���nM�r��k��§�l����4W�Ԧ�8�d*�Fb�8\\ӥt/K�<��PF�D�cQƼ�1��E2��	ޑn�}@��vV
$/�)VW�DI�Y���A|�����e��DYc�Qq鄋 ��$�V����￿������Z�;^[O�=�M��ҏ��=p�Ā��*�q�ҵ�μF)܋���j۰j�6۳�e�̓L� ��rD�0�� �
:D�sT��r�ň�?6F撚:�˨i@?�
U�ǎv��f�2�*(T1����1�Ύ�@�w�Xڀo�t�N|X�&y3vD����	�k�9+� �g�O|�^:^���'�����|,m��������ldE����	N\ٮ��]lz�G&p0�d0�ȶ�#V�A�?��b��-&�q�g�����Խ� 8��j�C��`���_��_�)/�vC�@Uh���">t�
ȼ��I�=�j����k�&��3v�G<�w��Σ�����[�遙p�!�&�O���2/g�*�s)���fv���N&��>{��%yo����[8O�3'ɟ�j:=y��i����O>���ٿ�g�MQrz��A0��Y<==mz����p��� �U�H����u�l��7�f��#|�3%cN10}���Ŋ��-9�M��	��O��`yNq���C �����@��4~����Q2oSn���3�2gn��&h�&���t����5pȼ��CU�~��z��u��;z��}d}����rf2j�K>�]�M��a~qK���L�5c4�8Ο��~������^\�h��x�HB?��O�%� �HM��UH�4���ɓ'�uha������ի����o��wҙEW�;���%�����M�	?�4�5�+����kp(��1�N���9㚾,����CU��m��d�G�FP%]R��%� ��4kϟ?��Y�d����h��_����"ht)z�۷oe3n1�4|o���P��q�������K����Z�J<n"��M�{Qt/d�4���{����a���I���&4��Q��"�?QY���0r&����Ω|���G����a�K�!K��k�vV/tHhogJJ�'������=�Ϡa_�g��Oo��#�u����#Q�J�q�BR����+r��yK9-w��'9������O-D�P!hEӧb6	�nt��b�m''�h�M�HCqyy	-�x��I�8��Q��C�)Zړ�l}��$�R\�� ��4,��p����c��c�����p��H�r�0}�S)��P�\}Д�0�����#�>��ܦ��u��'���`'�=*�^+ʞh���i���ԩ �O^�j�x��
ہ�b
��Z�`�y>�OR���V��7:-��C�=._B���v�e��>�̹t�8�8�'�AEa�dGv�-\�f�-ULm~;m��T�)h5��m٨21�XN�$F�=G%��7�U=��9�#�"Y+l�%�u�j�&}��)�i1#�1^�.��$�M��|ʣ��ÀA6�`;9��wdI��Ç��S��j���+���Gp�3��<�"���"�����+���8=��j`������d��x�N<F�[�+��P��+K�+�+�J�4JV�Da 5U���SӭҶ�Y�kv�N���љ58���>??��?�s:���������on߾�SL�&ӟ�V������D6��.o�	�+�V3<�aL����z�%�nJVږڙ��L�VH��z8�Gp�W�Q9�n���l�۾�Ǎ�V���D�]	+�T1:˒�S�1��F��N���J�˕�mF�v.~�;�A3�/�~�q���s�%�iݘS0.jA����m�,۳�@����RnS<J��-�-5�{А�q��3�̓ѳX�)��c�F�y�#m8���_C�cI[��K�j|/���O����Ih#<+�����Еf��4ژ�}�J��
�S���He}�S ���kig��`QT��Zc�m�ᯋ�!�>2M�fk�1XN��n��>��,'�Y
ډ���uI�,�����2�0��aB�<��G�n$�lN�	 �<3�0S��rl�gg�22�f�������M.CA�;�V���(:�h�f����΃0Y�5�`�[G�y��ǖ�����j�c��k�t�6�8���/UH1�O���	�"�K��ݹ�J�K�ư΋>4tߛ��wo�#;��=$H��, ���l��:@u0z/����1�"K����:v���7�pwǘ`9]�B|�w�^=b�f��4�]߼E�:�b4� ���w����0�g�� �:��(�FǧEe21C�]��_�˦���kYD�*��|$����s���C��d�hz���mr��j3#ߘ5�7���m��`��?��̘B�>w��|�ݐ��KR�9&x�#	����KI�Mm��n��i��h~���*�����|�<��\$����8�n��%�ݹԔ�H�&�1�\;u��&�o�Y5�II$�au���BA�5O%+v�O,�5��sC����;E�-���(�#�	ƫ�+�-g�a������0���o��yza�<ľa�]��[�.�&d��z�@	h�m3d�?�Ofu1�-��a3��n2��Kh1��ǇL������^s�_tBG�H��4qFz���f2V`L+���U�j4e��M�s>�g�
_o/�i��N&�D�����~�駿�����_�EJ�������^�)��䶑?����gϞ�E;�U�ͪj�!tj�䙄*�_}�����m��m�o����i9���.�:��g�vC7�	Jބq4z���<y�-8��d*rW��~��_}��$]��j�ۭ�o�章'���rqt\K��[���̹hy�\�77�C���,Y�#�x.���6�!�8�ݪuNkK���e�V�;8�X"�W�(T�\�/�ٙ�w���@��O>yN�?���e�H�I͈���k߮��,�5���c�6k�I�Nhi��_�5�mt��	m�Ë�S�Q㳕����M��lV���p{=��[hD�}�ڇ}O�b5��7w�
y�����~h�ڝ{O��)N��r��<�58??],f���a1�P����ɔYje��Z��Ő�$���k��f�I�y�x��	}Uvx�8�L?:^r����OaJ7��������F!몮�Ƞ%�6���	���V�o���I��Y��_�j���`Zծ�V�鬮Wk����W�>a_�Lq�p6�|8�ӛ�4w��uf��"i>��n��o�g�
��gw���o���	5�ͷ��Z,H: ��{�~��¹�/X(�	~�D��g|�<y��nn����)w�y�����|~qvT	��m�	��j�n��� �m$��hQ����=��h�'(���٤Ƚh��>l�vZ��I8��̓�q�T��|�Z7����p�d�qɾuY@���!���@w�LaM�I����~�B3�Mh�0[g>������ї.ֻ��f��3)`�5�-�	+C�0��'�?]o�+Yr�	���b�k�\�2k_XU�$�� L�_f�Y������8Pc$@���D4(J*nU,֒{�ͻ�~�1����$�s�,fƍ8q�����}&�Zھ��zA��/�7!��0�E�։/}Ű�8�.;}��LZm������Jʮ�AY���PkߢXɤ����G���%y2릒��.���<zq,]�d��#�����%�⺠3.`#:A[�'A&���V�!�=o���G�	�eǾ��!�zqq�jo;�]S-la�Ҝc�,���Qh$�f񌅦���!�jY��UBz���PO�y�D
E1�ok�<9�N�ȕ�1h��Ӧ$����-f��t���Z��u��.\ԏ�^���Nq&����6Uw�����b�GT��iw�ѣP3��@ۍ$�ʘ��JpS�H���}�����%���GN�� Ǡ8�����NGm�2??p.A+�Vt������{��_�)� /aY��<�_��ヲb�I�,��i�e�;iMHΡ�H��J���殄9g�/i���k]n*.C �
~pf�N�U��o��SR��B+�s�>8<����?x�`�����_����߽{�/��/��/���o�B�����$���	9�7	){S����[��@������7�_�-��P�^D�(	 �� +�6��6� ��+��
��
vn��RR�ւGu�����@Tx�+Hǣ�we�x�so��LGCs�]nb�7o�c_�:M7�i����.��=Z�8Q&�/s�I��N�V��* lu��ԙl`�,�N:1,ܖ�)� HZSz"�{g9D�M�62��*"����"+���Z�v�4��@��!�� 31�c2=�<�I�cs�8[Iou�-����Ƶ��1344t�!H���.H瑂� �&�/�������_0��OMr,Q�(a����6l�k�}*��b����E������5k�c���{ܵ^�F��}	$o��8RH�^��z�s�xP{�0��XcI=���Y���W�GbFl�/�;JK�9-2?]9g����g|\׎��T_�^u���o��N��� ��:Kj���&���)op���u-��I�k���A=�@')����ެ!{�D�V�H��]��lwkv��h²���$jy%px�9n��B����S�d�2ܜ����<�O_���g+nd
}'x�% /Hu�	�.X ��b��XE׻Xk��71�n0�f� �$�v�<����#�G���쒵��-�����E�)	��*%�$]
o�q��?#G��*�j��H�>Ye#&���4�}�yp���z�;�礎g�J?�hN�yK�Az�`�^�qw���)�:��A������m���w�\�|T���n�,�}�SYE"����ZuKRUx4l�a�V�5Lx'9Pz'�0� ��{y}� ���(�bd�H;烡lAr|||��f�����o ��k�:_��!��s8��Ƕ�dpg�@�8���4�bn�"��kF�^�>�f�"?99Y�����g2�����?�>���W��WB �;C��D~��6���o���e�5��+
&|Yl^q�s�CZ(�KeD���r-ʅ�ȝF@(N)��z�#��+@* �8Jt��P�Й���������GN!mĳgϰ�^�] ʑ�&Z"�i_h5�G����D�/�g.Dߟ�����(tnpuuutt��ٙ���J�2q"Pw�`�9�l�>���"�d�L���#u�	���;����t���nֱ�LBȍ������{�w�%79H E�0��,��]1��@��Ž���J%M�!$)�J}�^��c1��KR������{�׹�{�o�S�d��;�s��9�$�O�XT�61'�O��D�B��I璯�\rfY���Ǥ��e:Y<`�S�:��?�S�0�΋y���e*
�#����3��k0k����=ZU�8�ADB2D[Yr[�l2B�n�8G,��$Ҽ��hi�*%��S�M��C1��O�î��ޤ�F�5N��?�� ���8�ѭVX�h��E@�I��
��*Ec�P�z)D3��j@4�w��ݾ}�<-��H91W���5�k�,<�b~L��m�A,g���B\<�EP��4��f	�`�m��)���(IT�I�H-�5ә"�[,����u�rP�!'��Z��!/��Z����'��8l¸�h2,>N^;-��n��Y ��4�I�M�EQ�t6����Ґ�>�"�A�p�:}��C렐���#X1�)�t3�P"v��L���ఊ�F(�yĩ9\��Ҥ���}L�8YP.�ZieT`١����KNys�=�[�U|�/���,,9
�4t�ߐC\
'�C�؇�ά����)_J��"(�t�i� �v:�P)3{�m�̥2�Q�
���P�:h�	�b�H8�tҝM�B�r��G�g�Z�mq�Nc/,I��i����e[�	�:�a|u>��-��W����)N�:3E;Z��~�P��H�S#Vh��CK5�ӋN�w�!�V0���y�L��������4���E37w�7�u���Μ��ꂤ�B��n�Yl�D�-R�̚.���{t����E�GMS��zc�~�P��P��k��!ن�%M�������������.2�8_0�`%���ӡ���?�ud�`�O���9Gٽ���B>SY^7E��c�f"8Tp�8�2�b>2��٤�|��c�,N�6�$�Z��4��5�I�M��{� �>-�����;m̂�L!��`�L/%=>t��T{�L}���C}�Xk4�}o�y�D|��~}Q�6�-fm�f�(�f��8�u�6�����WG�O����Uic��Z��i�����jn�m
�+fwB6:�!�����2��C��[�8GD�֖g��7WW������z�5���Y�XQ(���!�{`Rqύr_B)�H�� �٩��RV���s��)�3(+����q��"��N�|�����@a���%�;N��������ϓ������ү��y�@��PI�ZZt�F�����EAHp�o3(b���h<�r�z0XU��ɓ'E��*��l,?���b��V�2,!#�i���Ֆ|/�a[T�6�sV�����H���F��0#�)�S+�|���}�gG�^L1ml��>&�"���v(�݋@l7�`da�
��Yۛ}ēgT��{R%ք���x.�Ч�ʜ�#��U?�ʟ۵po_���q�O'Ѳm^d������Y7���r�,���4�m]e�*We�(_���r3��0p�v��0AZ,�Ԅn.���Qq�Mb?�If��TZ/7��u[u�/�m5H�����������������q�B�U��+�-+S���a&��u��+�e�&���G^ϲ��[<�Ku"�!��~Eo`f�Λ��":H#4��淦�Np�X
����:nЎ:č�Ě��O^j�FB�.b��E�䙂(,t��b�Nٺ�fe7C��Zծ7�N�x̂fܫʘj�*5��c/���7��v��v�]�N��oqb�L��$����K����p8XEN�oL�����ܥ�nK��n�a��s�SU�9M�Q�8pr�]���^��W˦*��+I��H�K��L'��a�=�p�!�-#Hx`|T�R�*�@HlI���V�yK���[�	���)��D�"��;<(�C�y桐���P��m����z��t����/�8?}$j�U�p2^.��^'x��h�ptpt��;�r��,:>����͵�3��\�pbć��t���5�4w�M�F~��['t��Wg�qqg���S0\o+i+ۑeyz�O7�ɗ�j�VJ�7�u��1�o���Q\����yU.�f�Vz�i�ڮ_�]^\r>b4���:�K_&h�J��m��Jר`ⶌ[��%&������pDQ�ɝ=R$���W7kig���1�$�"�dr/�M�{͈,tH(K�q�2�X��]3.2����$[ZV��0�}{o<�����;����7�_�h����G�ݳG)�?8�{y~1�܇��înR��:�,R�nX1�ٔ��y�IB����^�&���bYw��fI�O!.`�t9>�<x�ĢM١l3.��$�ą��f�_� EZ�Mp��?7�-u�-���jy��6s[I�GG3z������f=�/�n��h�8��z�鏦��;�S,vhK�����23�� H��]�6a�E_����Dh�,������o.�X1�TP�q@�Xn�Ǣ��Y���P%�6,��-G�|��lJ��]ߜ-W+ٚ�h��I��Z-:D�g�������Y`xi�f{pS��j?9�IFBj4��з�`XT��U8e�7�.n��f9�L`�3 /�΂p9U햢x�E�mז2�<Q�� �1�(�ᑼ��%�>�v��OC�9$h]8>>�۟)�h{xppx8��Z,n�ί�uHIH�r�U�ަ5�ή�M�����?�Q�A�U��9�2�}�7��_^_^LF�9㖁x.͓����;		y��_�Zܦ\� c��z�^��5���̍:����Ui�<y���n5�`��[����B��oʣ�C�32*����z���'\���s�w}=�����Wr�V�Fo�G{�b(1�
!�n5���..�B�'R��p���t�?^/��j�8�`����q���KF����ﾾ�����	<(��8���.�D���F����I����7[�A6��@QBJ�h��h:�ؒ��tzt���7���o��o�R��$�$�0�4�w�x��褩�Œ\̤*�
��\S��z��s�)�i�d��·����r�ś�TD�f۲�v����v��jh�z�6�ඬs�۶M\!��I�=z�����v^�����3�\)�����s���z�	;�-VK�(I��&��Ѿ�r"����L�*URM��/��֟�5ex"��Z�2~I�,�p/g�4��G�yZl:��;,�"�ٽ�x�޶������
>W�CF���j�r9�����Gc�9k�7^�$�HnMȅ��)����D��`��^J�[\��z[oA�C�;)��w��_��	�>O�ƀЎ����f.YBO�u6��_�J�q,T�~MRKKq"�GgE�l ύ�H ����<�V�+�Z��ƻ�6$Xg��6� $8�NIp�3I�d��V_�I�EhC�0���k%fVq�1И�,�o������`�i\�&$-���d�v7=ªnWۦ([�Q9"h�0��{�|�؇T���_6+��v�7�����'�Y�	���^0�l�̈�,X͊�NP-�ȹ,b#4�\{�l*It�pu����f�eOvq����d��;G�(]��L���\܋ӳ���)��5�֨�I����A�3S�'�5��9�y[�hE����y�����?88��rtg�^��l֋���p��B[�Z�C]���~0 ����fy��u�\K63-婍Hjo���kңY�%J}�Ҷ-���r����p�v{���W���t�h��={�*�W��ý�B�t@�aB^y���֣��zu�&���yͻ誶�cG׫��={£a2O���a梕�d,K�ʋӗR[*H5Y�bvi��͒,Az�t��Di�Z'�pRU�C� �V2���r����  tC�9D�݄:n�jE�4`&�jP���s��l֢�9u�������^0ĵ�H/�.�褬Q2؝ �7:���ܣ�����U����t�Z���x(Z�;k܇�� 7��W�1�%�5-=�D�K(旸ו���?�`	%�$!�0Hw�!����{�1E�����_�0u���bMh��jӖ	����۷��)�����s���G?;���. UQ��۬7��b~���8�q�.x�s�":�aՊ���t�Z��1���+�;R����JȆ�in�$W��0H��˭D�뛕P�*E�[��媃�8)��Ȓ�p�my�sAVnSm�g*Ա�-�'��K�������rIO�Zn��_̗Y>\��
	���� �k��ߊ�X.7��W-��,���:��\5,י;�s�.7i�n���W$�/^�������bغ�	'}	��IzEP3��e�Hn��ey����7�>�Ig��8"O`G��$����B�K���,�U:�Mڤ��8I@v�q[��$�#M�k��\KYt�L�7��o�h�A�[0�IRq�t�(m
�M���9nr?�%�'��pl���HM���lr�������|;��Z]��$(��9m����P:p�}2$m0�/�)�/�K!�T����
Є9RҤ\s�{]�a0��&�ȇ!O�LU�$?BA�+��1�+h��@��Hx�ʼ:q�K%|+M��*r�eWR��RV��qht��ϵ�� �z�1��i�Z\�R����үx�պ$��H��t�"W��)���hk���-����"��� T��^��cﱻ�Z5�E�z�r������Y�wW������zí\� �S
˾�WeJF����9�,��.ڰ�z�Aje<q��d�\��jR��Cĝ��)�W7�R ����8T��#F	~�STb�նվ}���ՉG���A�M�v$�z�рawT)���v#�� ��ݟNF��2=��R��\���cڔ���s̚Lz��bxmG�� 2r@ �����E0��8�k,�h�rxxL�ˠ�ѣg���ۚ|����c�jZ��3��A)��x�!]���4�w0B<�x�.��dK���Mr~��ь�)��h:���&^\\�.wT��+�W�z����=z��ONN��y���%�-���>���֋R�ױqd��irb5�뷕<,*�YO�t7��d@����Cw{u�(�F�}�W(Q���� ��{�|fɹ<�w�SK���l����^|K�'�'��O^��h(9q1#����w��HNPk���y�'��H��Y86.���ٙ�e�!�b�z-����mxa粬���F��������
-Zs-jn��Eg�W�tf�e�=��a#n7$2ـ'�I'���L(QS ��2���T���5�ӱ?����R��u�n�[��L$s�TM1���舧��C�����K�x"F�JS2��c�HY!� @�*�gĄn�t��,�Û���g�� כ)&}A|�%�]76n�At��/ٱ뫫���k����>�s��ݻo��= �M	�M������� �_���Q�O#T�xd)�E��L6�F<�b�+��?�+Q�:�#j?h�u+������2h3���
��=Ѻ��rB���o�����d 1	�� �5t͎�~?H�ƣ)  h5���sc>w��v:�� �A�4��t�H��[�)E��T�[� �VAX�V�A������w����>����r��'t�<y��A6D�ƙi�L����byan�9�-s�YҔ��S��9$&c[��=H��y��߿O����	��Vu���ӯ�����yIۺY���<~Ä����L,�jG�Hz�x<�Ec�P�� 0Ǘb�Y#&��30�k��� V�wtW/�Ł!��( ��9�D64Y�UQZ�j�4Os���j������d+��e��^�r+�+.�E��	X#���ό�qƽ�Y<
����S٘�)n�7��Z_��8��<ؚ��C��!�u�;�.�Ͻ�LE�%*ݑp�z���-Q�6��p�(�$�o^'*����p�7]l:��^�U^_3t�Nf��̻���%�;I�t��+GX��m�E��E8�WwΠ��37ڔ+`����v����;s5���K�O�RE
�Df�G?��Ç�(��"��>��ƿ��o^�z�U}��;�Qɹj��4�a���  	�%��$�A�N��'8GX�L�s����b�`S\�r�&]Ao��<��"���7�|��W7���UE����F��� �~��f.6kN���i���35N��a F�vʪ��1��T���52D�vF�ī�X6�]Msg!���-<�i�WC� v!WRڭN,a^�2�(�w�N�"��Ut|\��Q<n07�C4�Ek����q@�:;ՂkQ�hZ|{��:{�8�]Kx����"A�>Q�=u4j�Spz����A^-V��^���$�hL$�N�yd����V�sA��Q9��X�Q�_�tXNc���%M2�X?��֫���}�]
X�$Zbb�ӱ˖�D���+.�mJ�˫/YP9E��\�a�%�b��7�����&࿌z���EY�����~V���t����c�+�d�X<Z�M2�99��t��A�A�A����?�cn�.���W�����o����n<Y* V�����[+@�i��慚n2�W��|��d:����.�X��b��#�c2�,ǆ��t,�t̷�^��w��Ș3��oṉ�W�/|�m]��TI.#��:��(�Q��J�6�*����4�&c֓�sk9/��u �d�B��}o��	��V���0Ў�累e�y1$�;�Rx�����U��M^P�ϥ��D6�$���_��&$���VI;E'�D�d�)u��iC[S������D�@�	�[e3Q�3���T���Z�'Ѭ�\��ELk�?S�f�K2h5���$e�+#D[%E�i��)]��_!gv�D<���&y/`�A]��7�_M�l;E�v�vΔ	�*����L����F�FG터��A�z��ɴ�����B�N�@L�a�@K/��x��.�^SD�І��+P�N�/_�ĕ�������V�bE�Qs��\ �Z�ІY�y-��2X*Y��|+8��hkaE�_�Q�>�!w̸�XDҖd��q2�Λd���=��`L� ��)�7[P'�)�y�GVUH�G�vXzj�z�@�,Gdߠ���&m�%F?1��#�����L3�Sh������	� ��vL`���"$n��s���prr<�)��k�>}|~���{6p���1��~�I��?z�V�f�]�T��Y�l�q�#��3�!���AX�6�	՘�VQͭ����hj�����M
���������U���Lro�
���� Y�B��j:�MƂPY�V\�!Q;:>����g����?����Ǵ8��ͯ�G��������Z�rJ�U^��t�X��	��\i�y~]ۑ*��"ch	2���K��Ŏ>Py���S�b% Wџu�Y�Ů�!j��1JA�V�aF���3#x2��+�����%'�&�u�!��j��l$�)Z��hwK�z�^^__����09��k������i��h{˩EB�I@�)�A��T�)�N���C�/a)#�d���۷�Qk��O�Jj`�^snSp4b7ʶ��-��JG!��q3���3�1F��>�����"��;�bX�
�swҝ��ƻd�i�PWd�7��y`˛o�I��z(��Ч���[:S(������ܽ�������f����,I�3 ~@��x�\lifhN�8{(3C�Q�&��ЌǤ���v4�U9MH162�c�,�ǟ}����]�П����^o��o�_�7���| �����fq ;F>�B��D��h��넇�j<f|�v:�+z䛥�dM|l��9�<1x+iPzi��f�E���}o0�'�:y�����������ِm���/H����yM�	\46�eb�mGc��l�]��F���*�-��3,g�O�z���Ӣ�WCt�r]>~���,-�_	sk�x1K+�ᖰ�0�WXo�#�1[N�[*a@3��ʞק�d�P�7�י����:H]�L�g쓂�z&"!��i
7YV[��Og�h�����t@�kc��1�c�l,�d��-ɔݮ�N����O�z�:-x��\ӐV$�t����#}���f�w�ݻ8�^�Om�8$m���^op����mv6ݮk�!x��X+�]��3j��2y9�.�AⅫ1��cSW�w&�Rmr&-���y��Mu�'���m�f�,g�I<K�7�B`e�kb�)�ӑ;�|[�:PSh�I�bC����+�{�߾�&�13���|�	��?���L���~�;tc`�ԃ���_|����d�G�us=/����˛�3�fa6�+��b�3ſ%��T:�	y+t���H	#��R����$Q��Ɇ9O�n3�8��/n�JyR��>H./ϯ�N�C���<|DN_������[]�_!��T����������������GnD�K���1�N��:L��i*<�*�4lwg���e�D�\�vv޽�"I��Z�M��7�M�/5�3��M"� {GIFpa&�9O��t��Bi����x�#�$[ZC��[������ �̭� ���F����*�l��\6
����V�t�Kk�@�鰗�t��L�	����.��+E��[4�����FTt�@����lm2��°��l�ӷ��-� ��� �_r��O�<��-�E'�ή��lbBʞ�Dv�Z�A�B0E�I#ąx����1P,��VG��`8��?<�}��?���d���w���������#O���Ab˂��S 8������#h�G|*a��R~�ǿ���ˋ�C�3�!�����|K��p2���3�0�k&��XϷ��V����Ѕ�X[/\��m�evev�ޛ�]�����?�������������?���`�R[�wy}�t&������
��SDƃ�i�ʚ�1e7H�h!�T���^��`8d����L����f_�b�,��ߪY�~V���|ok��V��*/�N����xM�Y���~L+�hrv�C�j���9e�����ffg=7Ҧ���w��[��lW ����3�+,f��l,`�������駟~���M���r8���x��Hش^�6@Z0��K�c�C��A��S�Y�c����V��s��㦚��8]*�$췚v�����~��.g��� -Z��{>/��e�p�3����T�ˎ��>��7��nI�qB�m�N�z 7�"��N�/-C���h�"��a[o�Դΰ�Ѵ$�@�(E�}����85�h��q�z��`���F*`p�P����p��(f§i8r�V�5�#�jd�E�&�a���4}�4��m%&ԵP�@5�]����,mi�Y����2K�t)���h^���#� �B�\!ȝb�`���&�n������)H�`�Q��ޥ΂@|)���C�����-#}5�z"�5EC�a@����¥��8����v���2�ym�Pa~������z����y�m�S�?}�������2�[�1/^�&:L����zoo���T�����K���A|�'U
L��H�$o��߽f' Đ�+��ߺv�`��7CO�?�<<8����'{{���hO����W�����q�r�i�����9�ɂ�Y�>�p&���8�0���	����� #7�zS����&5�s��x��-���M���<;:�D=|����I;�Y�� c[�Y�	�AeW�
r��R%1{�*�����"m,<3=���ٹf+���F}®�S���Z9@���z�:>L��߿����䱡Ϟ=������7TF�y���|eܡiN�Y���Ǐ�ԁv�N�y�}/�\~�i��S�$i��9�]�q s������p~}x�*)�$Qd�0w�%���d̄�M��7�K�N������똹���]��$ڗЛK��4�LY! �r��u�,{�b+A@ù�ME���q�VU������?~��_�
�����!��;�^������� �I
�=H�1l�P|�� G������1���NYl4O���v�F~~d�3�ε�	7�z>����O1�(�󮗧HB�W��:FЂ���J�t�]v�t-2#�&\p:B�bI�����+�����ӧO˚U�6N.�'ri.y�Nf��1���Q��Z��`Y� 	`�9ߥL�@��)F��,i c	O�J���6��7��7ؓ���Z�A�Ln��C�35�w�""1�T�A�b���\s����nh���ѵ�$v��'6aD�V�S����.�!�c�i�	2���Q���faj�Q����#{����$:�ί�ՙN6�����Ag2@�9M�u��ju�1��r]�S&��R��v2��<U�9>z�pb�7Udb��a-�cژ��K[7�@qy�k'�&�GO�M�g�lc� �FaN
�l� �1p�f�L�oe5�&ǧ�>Ŷ�!&;��'��d9��p�>��>~�����˗�^�"灢��z���%�V��I�R��H�Iybg��tFj��qI�<�/_���جv�Y*r��Sq�Mx���`�a�R�����,~ǝ�7�me�sP�r�p�;6�Y�����շ�~Kox��Q�-A�u�����?�P/AZ:sJ�8���Y�5l��	k#�BO �2�	tS��!��*:�g�=8���{���x��V�[J�_�&�u ��l�V����H�7.�Ђ�.��=�G�G����Ǒ��'-PN.�h����T?��U���H�?���mh<�L8�@>��>���wN�z�3�6h��r9��"��1�$���p1e����޼�(=f�(l%ӔI�Lzz2�v�w��Z�-��w5[�[�o�xu}��ux^P�L���̿��;Y�"�@�TE7xt����t�85Y�����O������F��A'#�{i�[�J�/U��Q�=���ߢU�ɓ't�y����~�Gd��R g���D��7����<��1�y��/hsa�7�J��Ā.B���pL�|t��������w8E�y�f,m�5�����t�b�f:����nݢ;��<��о�,�ņ��G��z���=Z���l�f��;r:��V�R�z����,�]�QC��"��2龓�i�I �(z
�Ⴭ�z�,�5��Aj�7D��X�r�d��岃Px��#!N��԰��n#�8x���v�����gS(�(R��������$O�����U�tx�{�t}�0_�p �-E�1	k��
���t�S����I�������E��o�����������ۋ��>��7S������)c��v�$�\U�܁dp���ǁ�Ka��4�`��p1�dvx2Ę_��0 ��R��Hכ��{CQ��s��sV������u����B���`S�� !����>@�� ��Z���Nр5T�y��B6
�T�F��9��;��%i�~�:��9m���*(�F���,�(&B#����RX��bo�Mm��T�Ig(pb��u�,On�N���I'���?���f=��ڬ#�	n��)���t2'�S�ڤ���Ec��ӰC0c������mմ�YGr�V$A��(2O7�ZUҨ%�ͣ�Cլ$kY1�:I�S�ے�y	N��d�^����i��=�s@�P��\:ߌ��l�C!F��x6%�?��{��%����������?�����dZ5���>oqǬ�l���(����MG�P��,�9ќW*�y�d.sK3�dˮ�dxk($�'V�ia�|p$:��^�D�U��C^��h!��>K��g!i����W����{wȯ>��1�l2����b�Ogc0;�;����G�s����Z�M�+1,|YL��N�lT���C�ib�K�kF��w�!l��M慎��&�E�Wi��@�m��0_�_�[I[Ov��A�X'%]��fC��N��$��Rt}p|�t89ا��U�R�8~�_����I�SD�KSnۚd�%o��龻�r�g���J[�y�l�����}����0��9��G::>�ɐ]�Ҭ� c�ʼ-L%VJ�(�}�������H������Q&>y����닲�|�IR3�LG�A�3!*�;��q�@�(J���۪{�Qb�J`�T 0���;![-���d�;��$����g���<o�:	䳻n,"����9��(���?ag�/̕��2z�rC�=/r˨���е-%�]�XHm-���L��ĖL7�ډ������	!-%�N�PF����'9�Y����-V��~�!E���_��s���l��1�`.]߶v�%�� ��}�*bvD����Z�ף�2kPx�\�KZB�y]��Tb'�D�OGFX�����e�7���fӏ>���˗s�2YC��8� UU0{:8Y��� �I0��^tIf�U��P��	��'$�֥|��0#�@u��0��R/2då�.&#җ+6��	�;�����"C'�_k;j��m!`�1�`7�V�툝k��	��dW���V�d*C'� &$���nRa���hE�����A��B��O���o����Y��)%rXcnQ��8^�{���I�(KCn����cߑY����rU�k)�P�p��^Ap��k�ah6��ZF��	��&�f�T�N!؀�`玱b
� ��{��/2]8�����:Y'	P����]�'>��P2=+�B��c��7[���V8��47/T��<EPo'U�;��;j�9q��H?��Re&{!�C���g;b��J�m���3���]Ƕb��}�������>�`&��X�"����]^^}!����3R�VJP����b�Ԗ��]?}��֭ە���9���9��^�.�����+�}R9�O�Tx�ղ\��җ��W䷽|E����!�8�x]��ַw�ǻC�s2ٟ�&��`�����&z��&O��_�=}�l4?���MQ�����~i-L�t^jO�/�l�I?�+�1h���&Rn/�a�� “�:��Q�D1��(/t����$�����&֚%Odd��{a,X3�rD�0H9nA�7߼r�vv�ƃ!�ԋ��>|�wȤ_��:�<�����=�V�(\3'''�Az��]^^�#	%��81����X��"�SqJv�����H
`k.����"#w��zN��A���c[@�7�Td��s.�Q��y�|�$#L	���R�)�$�lc||l�c�#@�M!��L��G�ް���/Z��鰯�bi�_�7ϊ�/N;��F�ܥ�S�l �M�$I��KfGܬS7�&������voq@����\^_��7�Y���{�*8O�W�#��Τ&
>} ������W�uW~�q��{����<���>�>crs���8�����?��֗���Zk�|��t�h��z4�kr�g)�ڏ�<m:w��1]m�����$~O�� 1 �Rw�c�I
ֶ\V����\����R��i���ӭ����rM�LQr�v��I!?H,�:܊�Fӌ��nL��:~�#�w��I�~���
�h� yH�D��l���&Ƿ(<�q�r��^��b�T�j�+��*��
	Y��o��
�]q3$3$�;xU�'G�냜,Nu~ƴ$�1��J<���1!������;�4����;����4D���,n�:M*u)Z�wy4��X�Tr�����|)��8�7��?���62�۽^��Z����6������!KBY�����4}�wqYҬ5�N�^�>��^��غ7:���r�00�Vz�YH�����R�=H��n�eZ����5�K�p��!l�^�.���t���l���%ht6�/����C���)�t���h�9�d+�H���o(�J;�鴻F�b+h�5�����~�Z�J`�
.z�N('PL���g�b���t��Ȫ]V:�4k&��x�M�g�c	�������g�	��[wn���d�q:�2rw���M"��2�DHA*��Q�F��LZ_��{����X(V������:V5�D�>8�@r�Y��E��u�V������(ߛ9�������&�$����f��WeG97c�禊�h�`�ޡŵ��l�<�L&hLW��cv�RT���x-U���1Wh�|��$e���a�6����,n�<<:<:�q���u	�lJ��sI{���<?3� !�7�M�6g��yВ�kZ�X�WX�@-S����\�e�]=`���6=��/,��'���cLy��ɝ;�ϒ�8�έ���>���i���emI���L��8�
B�
�Y�\V-�D�ο�i;%C1��>⒖:��������4��ц漏@��<��2O�H���ztc�Sy(f{w�2���o�Fc�C�p'��$A�%|�Fk�t�2���cc����!���c������d9w��f����=G��'�#���xŚ�Nڦ�"IF���G}��ٳ���
 G��ؐ�7,�t�Ć5f��8;���Fu�Q�P%�T�"�Ȥ�QGФ���������]���-<�3����ŉ��y&^d��:�q(�O�>�rj��_'Ҽ������K�:C���CA�ɓ�>����sT@���p��0�l�2o�Ie �h�)KqLm��ڏ�tZOj���gOs���K�FH=�8�*��lk�p7R��<H
��1��{/�ݴ��xi���d<[��W������"�D��0"�̣R�6$���f��3�i\�,�6���4���FR*�&d���շ�(�08��]�-�D��hA���5��D��4
�ѳS������<{y����
|��ƛ�iq�Y�Y�@��U���%�g(�h��'|�����%:�B81�/[��6=�Y7�Oh��T'���O��j�Ъ��"*T)�a��)[Ź4��3��x��Ӊ��A
�ųT#��L^9��ڭ���f������m�B�'
�Z���+�*g��-���L&`�=v�N���^��(�n����b��W7��B%ҷ������F5R�uh������<��iy=zDz[P�LA�Ko��_G�R����7�L��I��v�g�EU�=%���$�v>�9�;��7�8f��3ʹ�@1K/Ri@�B�=�IZ}4�ΌR	���mt��g�~�{dJ�5OR��8�#��8ݦ�!~ �p��?fz\�^�P&��V���V�����2/���ԑ��B���%�ܰF���1�;Ti�X�b�uq�BfѢ}�H�f8H��I�lC�p�9y����̺�8x���V�����o�����W �nh��%s�Ѳܽ{W�Wl?~���<������o�Gh1 �h�i��oK�S���>RT	��0��[wND�r�6`�`�&5LKqzzJ�_��i��y�����������₻�]��"r���
�t%�IN-H_�a� �s��Q�P��Dj���]j�k��
��ŋ���r|0��u�R�#H��!��QB2f��D����P��ϟ?_
!�r��mځ�#Z4��D��?úN���Xp�_کNQ��RZ糳S>�G�w��
&�.u|t�R��e�:�Gw<o�
�IM��M8"�����tF���vv�ȥ�.� c��kB+i�,/8vRe����,ׁA0���m@zD�5�s���C����P���2r:M�V���0��"7Ed��+i��	K��}��x����xM=Y�l9���O?�!�x.�㍺��Oe ��sȐd9bU����	��m�*`��%mv�1�& a_Ok�'���U ���ٟ���?�n�!q�F����,��oBn��ʢ@�C#'<Vk��i>ҽ��3���}�W��߱�f�mYḄ�+��כj-?��g�c�-�$`�zN���)��Ep5_��\��[�1@�S��p��.�����.�\9���;�Ml},�ɨm��{܉n��p��'_7F*��Ak��&(Qo�u��k�Ёb�6�PPn&�q `۴�q- N�*�LF a��
Dyi�3�I��.��>pI;]z��1�0�=H�	 �SM��5��1�Z!t�˨�[������I�-�o⤋�	;�1�ϫ�٘��x8�ӌKE��&o���L&ӣ�}�ql,�&��:>��A�Ã{�O^<}�Y.���LVN��蚚gI�M�SOy% ��6A�B½)gFH}�^O���U��M\7���2:�<Rq� ���P5�c޴�,	��k�<�u�h8�u�|��������1\��b��b8&�IJ��Z�4������26�P~3�&���������F�D�j0T��%��Ν;t��{�5�Z�a7�4��s���J�e֢�9����@��<4�ݶ���A��:O�7��=9�=ۛ�2�=2O8e��xo���o�M���7��iN��4�"s�b�[�E%'WBߦ@��NF���N;X�,	�q/MSd���g��[-��O=�-�����\�	� E8ȵ%9��-�p6Fie�'''���h��-�סbϼpM�&O�"k���	ʃю\���Qw�JxlƧ�nc��v+�ر��ԩ�'4�e7��:Ǹ9fv�	�#>��Ί�	2Eg8�p��ť� �M2���x~fG���f���k�f���R�3,��\'�-+�Jy]� �9u��Ka�q�i����mc%j������2���932�����hb�Z.*��G���d�(�$��B��+�v��"�4Q��$&�T�ys(����NA60��� =����1j�t�����L���z�,?WW5	�#ټ�OG�O����4%�C�}1p�
Jǟ�߫������EUKI:���U�-���cj��J�[��j-��A&�L�88�#�C��G�*�~ۮ����*�_�^eS��G���j���|B��5Ǳ{��˦�m�;ҾL8ß�:�[�F��v�V6��cw���p�7ե��B�]�`�e6b3�P4�wٖ�9!)vג��3���<+4�h4̂DVek�ľkd�=��N�~���S)xP�4�D�Ӻ�Z��<�S�?h�Q����PȐ�(X{d�U�F����!���E���j�(���]�6&�pۜ��]�� �O����M� ��Ր��T1A����U��W
�!�Qr�ݼF�h�o� �~��|�N��]�d�����)�4�G�h�I��Qq��{� ]�\����$�k���g��Ǿ*�S���|��>"����I��:�ML���RA�	�*c[����՞m����D�I���a�i ��vZP蠟>���B#K�W8��ȾA��P�L� �E�4*�ꗿ~���������۷ļ���"�T_�ϟ��4�-r<xS��)k˪��L-p�H0+��)Ii�_�=�9�����	Ű{��<}���d֑к�D�Y�c@>f�-�WW����WfCF������2�)y��x�턗�O?���!��m[^�_\_\^�pX �x#|䝗?;����1�M2���@Q�A�ȱUd R�ƅ��T(���G��v��tFxۏ(�,� 6Q�a��h�ls��u��qJ�ȧC������4�6lO���{�;o�~����~H�4�����V��޺zzJW;><��F��P~adx��CKG�����`IvJ��E���z��1����w��B��Oq�靋9�EDMuz�����䄜pp(�M�v~�R�����L�ǉX��e�Jrg����U�>�;ep�6C�y�a�녙 m������/.�D 7��3k"�7�������~{�X�!d)H+^�������y��Pk�N[���4)Y��+e��rŷ�99�F���^���3F�K��K@��|:��%,�iVh�~��g�}F���_>|�P���K��h:[�7�7+@Mi׋��|2����=�m���9~ř��[�ٮ�CTr*��{9v�tC~�Gio(�cfy��9��!�,��W���\�d��i���%7iт��\^̗�|��ҭPB+���3/�m�Y���K��-:֓%�9��\����01?��9E���VwJOdVRuR+.z#x/����m�T
�Nͩh�ao"��r�	��G���D.�U��<8���p��\sh�\1iNo
.tM�\,RtAy�i��zS}r���n�&*eׁ����:�3��Ё'��5�b���p���$�#��fA��NzJ�ݴjP,}?��4-ؾΒ��`&�yX�DI���M�ɫ���^�w]r��x���z*ʮ��i��L��Z�A�,k^��{�L�+r��f7֪�zx���O\�t��E�k�h�����r�����[(�Dy��̚��j]�h��-K��3�.�
7R�%eG�`���}"���/6��P��C	�ꇍ ��,P��I-��2#��E]ࡐd��&-`Y;�^�pϨ�f�l%�|d\mR��j6�2���e}݄G�34_"	c��HɎ�^�@-ն�D;�q���}�g��&��(�:�۾`��>}J��kS�_�2��ye���Պ�Gs]�Hbn~0*ӹ���@.=����?H^�����;i[k��@�!�!��rN[l""F0D��D�Kp��'P��`����9f�|�>� =zp��E�m
!��Ĭ�-k���~��t�0F��H lѺ����v�BpR>`>5�3K�[��7:3��>�D˛�*l%�~�s��$�/�<��"���B!d;"="_E�҉���\�+�*��ai�g�#SE�g�$ƌn��2K���a#��K0��V� ���8J���[�?���i,��p��}+��jaF)�r�_���Zg�%�~���sQFcߣ��lfK-Il)���<���H
.��	������l�Ƀ�b�z�>�e�C�6*�Y�
\J3 3�D�#NX-\sJ�8�<�Cٹw����y��U�0@j-�X�"���pպD��p.ŧ;$���p�����f/�h��cW�ٍ�gF�H��B��$j��cX��J�$�!'��7���	�"]R����U�Bm����K�u_Wc���$����7�:��<^�������r";���%ʱ|�X������X5a��Gy�s�)졨f��ϻ�P��rN�Cפ ���A�U,'-��쳒�·�m1���sp�M����B�@Wὢ��s#�D+�F�o��}�,��3��~(8\a`���F�0�Q��{����n��-�%
��ߡ�`��S���Ω���|b��������'���S�-��oU-�kw;��uo��iPݤ�2������C�{�=nl=k0!�("Sp�t=�3ф!h7p@N��JD,#&HtK$�B��a��[rP��ǋN��!�6�@\S��i��6[$�*�c�豱.�V9�po�H�"Cջk�]�:.�v�Zi�+���~�/w�T��F#ê >����w��zk���)@���� Z��j�&,�1SE��w����$�L!��R�t{޻��d"� �t�6$�9KA��T��́Ʉ�x��S�H:��u����%*�MF�k��>�����H#!O���p�`�!���R}u��Z���\�8��8�̑�i�ϡ�˺�~�i�,��������ҡШ��F�B�*9���{������}��_����"���sS&�l}D�� 3�"��4�q�Z	 �*�p�T�(�T!��}-p�2�*�w*���ʶz|�f:��F�Ře���)���v�f���Ŝ�&[^�����O������[�x���;�#C�ᐼk�� �}8��dB+3�����?�=�⻸S���t� }��˗/�r�G |�C�Q��_�Y�ˌ���FM"\+����c���z?���_��N��q?�|����3��q�-�Wk���,d��s�g�A��ji���cJ5�lVɀwq%?$���>D(��?�<�!�gn.S'C��+��3Cn1�_J���_�!KW���޳�{�����nͿ���!%���r�4�L�u>��?��?���鳿����|��tB�%&�@�p��ov~-��ܺu����zN�F�̦a���N�PȤ���Dt�����)�I�E�1a),��:R��>QK5���àI��s�y �N7<����/���h�]-W�Ĕ�YvqqA�`�%f�,�aq�>����O4�m�Q�D-������|,p�l����"e�n!$�U�[6���i{������]5�V�C�G���x#���,��ɐ�]�\�;�S�Yc��띦��Gu���g+�Iڹ|[��ў�hl��2���+�uh9'��ȆP�NY��)Pz�~6JL�X}.L�A#;B���w:��|����ڼ���(A��Nu�Z���evL�C9I���b]��ĩ��|�L�i�C�^�(�ā�ע?̮����ă�Uv��S�Tk�$��?��vҢ�.�?5�xJ������߳�3ԁQ$7�Huis�s%une��,r��tB��vC�6���i���f#4J�ͳ�J��1s@�/��lpO��E�ȇ��di6f�/ �A��^Я�{�>�by��5bm��y6��z��Y[��h�Z�D�7s@q$6���"S��6K�c�y�O������㠋�#x^iI3/�i�B�I��z�A�Rx�\�s��ј�n���4�z;:<\̙�ʋ���N`&eʔSrms[�ˊƣ-�u��=���I$�9�#ט�#c��!�Hw��m�2��l���U\<�M�{���y�qU�\%��[e-��MDN��,XΗ�&�ù��t�y���C�����޽;Ϟ=��Ln���jz�-$t��k���$��ü�R��-���lB�X\��2��0%D������.�0��ו	x��'Ӷ*;�@#��ܻw�ܩ�_r�R8���
F_�5��b���[_H���PV�N���LP�j�pMv}rn@����I����)m_� ���vӎ�����ӫ+>]E�2�l������9��>ZEh+�����͸���Vӝ9ˋ��I��1ꎤ���Ą�S��rG�$(RoM˼�]Sg���u+i�-7��ÔSo<s '%�w.C���8���9E��Y.`�.��W�-��l���%D#M@t-R�0i�D�x�Y�L�1B��Lu��&j�%�J���6��ZF1�<�0�e`l�����<D�֙��=�2�gޑ�������q���p�j��1�q�G�8�bӮ���X�7��X���rF�z����؉�,2nOCSX�D >b�n��`@0KP7���$��}:�ՖVj6���zQn����5-yp�r~��v0����7����z�$qݛ��޹�艐г"�ނ�v� ��Hە)�j�Y+|�U�%�G'�=$�P�?3T�a5��`n��D�\�t3Cwݹ(��B��5!)̧��+6�?��k��f�^���F1p��'�K�=*��zK�[��/r�q � �Q��[C5:S�e��d�.��ۺ��zf�ޮ
<���v�]�IG��|���ɐ���Ls�Zoi-�l�,f�/ЮVk��RA����ވ�.r/v$/$ǽE�����V������		c�H._Y�Իn>���^����V�@L��}�8�2v"Ku��#� �9��j�4�ʘ
���%��!��~��$^�.��z�a	�B,���zp�8H�NZ�V���S��4�i�Uo�p��J���K;�k�zS�pTb�c M�w�;�U�CY�]��P�2	�#	/~gPhq&������:��H�!�Bj�����BV>�3�R4�fZ�^'�UYK|(1�@�ƨ��bh���t,]��j%@�1��
�y
�&�8�� &�t�n'���b��|��P���\^~��׼��	,ON�i1��~��<���Ɂ�3�2����\P_�N�7�!t�)��������t���W�^���;�:�j_�|���јv���p�X�?��c�����t�A�&�I��`0�nL��z8�w���T:̷�{���d!�~������������j~p|@/�|���{��9���3Y+f��xq�sa	7 ^�cXвC?�I�
?�U.�xq���8mr�K��nV2��BK�,���)g
�2t�ܮ�1���t���ů�j���cAv�<��z����::B���(�j�z�{n�t̃�XA���b$���0� ,����03�S�9-�������T��X��vMN)��F�Ύ���B�|Z���g蚨���՛��W!�|������z�~rZ׈[��J�c���'1�D^��� F�ƽ��$*��H���C�u�}��' W�vD9ybO=��X�I�09W�ia22�B����I��������j��2��b���>���3����������֛o�I�fc��_�}�98�G:ꌸd�hBZ�?��?�����W������j��\I�e�0f��~��߉*K��(�횚a`�*$��{D��&/��Bf��2ޡe"z��\�jC�-��'a���N�"���8m�SP�e�d[[q�������˾���v�\���]͗�m��:L�aƀ�t�ǜ۽�o5mg��VqlF�m�-Nu^�G艬쳥N�bV�{�3�Ǟ�6*��7mَ�ג���zCKl;�s��D�Lv��+YG����O�?�#�!C�cմ����/��%����\��"���'��I��`m��ёφ;:U<�sU]�k�\vVrbhI+P3D��5M�:�L���|#[�N���U�+���5^;[e�<�/1��z�Ɲ&�p5s�E�������o��ذ��C��Ŵ�}Z�d�U�y�������U�Zf�_�:�]]g���G?�����4�N�+��ùP�#��oW�6�Z�mb����)уJ��=�
Q::-�C�" w*��A� 7Q荝d�1�	�����:e��aWZ-Dt�A��H
�.��]+�Z *S��o#�}����H/�[���@�A�ڌ�$;�
�3���!mJ!�����+I��eԇ�g<��T$:�)�;P�XZ胳8�~km/^A��
��,dӲ�x?v��t˔�	�2�����Q�>����|��a�U}���3~.aH�H�IV���Hm��b{�$�!��:Y�_�������(R� 1�WR�aP�N�/ϸ�r�G�9>�����}�d��o�|��+f�����/�+cIm�U��^dF��(f��_�`�=vs=��1cT�b�pa#�AiG���ysα\�V�\^R?�5He��A��]�� ���fn}A��H=`S��s�0
���N"� ��un�vǾ!qE���1�_a�v!�����+]H���kRF��̂W�u�����_�A����u�Ff�ZZ��W��4�
��]���I� ����F0��E g�샑�;�a��07�|��x����#�	�Cb��-?M��J�E��L����G��d��|%��Ζ�o20��z��v>�U�8��S]���i��Ty�辴��4`6��p>.=)�%�l-�ڤ�KC�YDԸ�l9#$�qؑ�p�SS,-�7�*���Q�����V���&����7�ŶZy����%��?`�S��qquM>�͒!�f�Ȅ�:�L�]��jԀ6���<�2�xEv��1�D����#���'�]G�t���d
G��[�n}�Ջ���

�n1G�ݪ.�~�
�i� ��'�)��g,�zaG����Jd�(�묄떱P�O�s�Ӟ�Z�D��ȏ���k�۾X��["��z�����2����h-YԮ���!�E.L�`����]f�]z������ f0�tER�)���G�J�C��1�9N5���c��O�*5��I�6�󲭹�9�����|���z����_�)��>kީSlrP��r�~�S[^0��ڌ���B�NNuJ_Ż)���[�Ã6Rd�~��Uh>|���4���$�6ف�tD/T1���k9�+��8��zAc�߿��K00l���k��������K����hHڣ���2vH�P�%;ͱ�~��G�ꈻ���Lv�9==��q�
�����)B�?��?�j~p� ����ӂ���L��t�6�;w�<~������}�6��?���Ç?������|���32Xt�������7k��8�#Ζkm]��`c�H��Hj�ëkcz�yl�A�N6��$J���D])R� v��F/յ�~ָ���{�&�I�ڊU�'ω������n�;���k��-yS��[�n=~��[/]��e��V��+�虃��x#6�^�j�^FagA;6�"�ڝ��~߳m��EHxf�fy.��F���	�FG���Q"�#J#�8���O����� m�
L�s�����	h]���� V�l������-;A�`/u�~��li&�����4���_���w[,����/�'m�Up`EG���\qH�,>]����c׃��	�f׸� �߾}���^"!��	�6�vHħ:H�7їÑǁ=9=~��ww���
t�xg�H������5��6(����D.M Q�u�N��m�v��oJ��s�=��|Gg�n���_��/~���b�[��[�)��~@6�ƍ%���eZB!&��jB&�<
-�l��f�'��g/�q��Y<.��)\G9_kM�2��j�|����l;�Q���VB6��<�h�������D��~?��2��(a���]/q�[)&�������� e]��H춽fT����p�!���vMmQ����������^��ȸ���]��8[�͑�H�RE���m؋&�,x������V/R�3<3�~,�T(�+��Vy�!^���]y�T��_��Uy:I'xŵv��%�B<�d�̑��E�S[�Q���_{�9�Q�A�5��,M�*��?���n�K����Xt�/��d�-9A@zA�H��w����k1U��<���y�[�-?"����Z$�t����D��I�Y+����ڞ�4?ċ�r[d���� 3g�֭�k�V#���j���r2)+ZI'�80�a�U�1Z����z"�S em�I�f`��1P:��@�t�4k�6��"��#��S��r��+�6
�Rxv��[AۇƇAS߱�?��4\�C����TĈ��"�ti�s��f͜��l�;���`���4�LAށn��"�<􈺟I�4����{W(� ���@�Q��(�Y�'�1�d���v������V�sC�yN�OF�0ͳ�*7��!;�m����k�<�(��Lɴ��/6e�T,g�ҬZo����r�ip�t[�e:��6����(���
����T��4КI6�ꄶ��.t�y^K�H�2���?0�?ڰ���n���K�	}���L�\S/..hc���t<���tCi�	�l�ᨾ�I���`o9g�F
�$R�g>���\��'�/�֞�g�!�*��q��\F#
����ČT�&Y"�pS���XaF�1�}ːk��O�V����<Mֲ�k��f5\�����jE���y��9C��dT�pA��T ;�n�b7�oO\������&�h@����9���g�l�!�� �� ��Z�+�	��@*���om2����_�t��츗��
�r�ʠ��i�&�,:�w�y�j�8���o��enA-y؈��">~�Z�?N���E �VŘ��iȅ��s�Tv��-�T�!�����p�s�F�h��+H9�%�F"H`����M���g����X�B,���m�t�Y!H�F�(���l��Y*�U���*��bV�;�	�rL�Cz���*i/�&(���m�U�q�9����I�Y����KN�Ζ1][Wk,/���j�" �j�l!P"�G^������xX���t�pK��v��)�`��jf\�8����L3�+���,K���fM�Kz�6��.�7}>���б�`^:P�ӝ��r-,���l�sF���|�z�I��\v��U6[ɶNs>��'j�O;��Q��E�	B�Z���h<>�?�����.���9/,�Etc���_��OvZH	e�����ʂ�$N��-lj3a�ᩰ����W�ad.~��}'���<ԝ�̩���-?�* �Ӣ�@ f:!�\�+2Y����xy��b��K��ǟ'^3Ezރ�J���{����-���j�n_� M�q�}��ì?������6Cmi�N���v�u�!ev��3QD5��\'9г�%���8\< �#oN-����nيxoY�UףR��΀��H,z��EM#���x��É�f��o�N֊jY�Mܹ�#ܷ�~���Uo����ɢ�k'Ύ�e���$�t2� ݖ��[!uԓ���6�$)2G���b�����ư���"I�_x����ӳ����LU1fH�|Oh�o���=,Ň���*}������L&�NE�y�v@f���)=y���7�)�8�,e����==:AE�\S��;w���kd�h5H�<���ׯ_��7�qrr��o~����ۿ�[���(��׿	�<��!�q��6�+׮&��N�j�+�
�}�#a�����|--�I�����cb��ù�":���>�FZd��{�\Խ�U�7�2h����8)|�Do�Ė��	Ed����1{Mt�:���j���Jt)97^2�t����Z:w������`��m]�>�ͱ�M�M��ZE����K��^�D��MW���񔴋C����z�	R�5���bp6��uR���˅��V�t"c�R[m��ӧ�W<�*������A�=o]�Y���%�'g��/�B�q��}��k��oߦK�L���	�� 3N[�����sϑQڬ�'g��7�����W�..��P��q+��MW��CJ$�	��[xj[H�Ԙ8����_�җ�E�ɻo�����uInsY5HV��d0�0�gW7���Fb�&=8W!��i�<H˰{���W^�"E����z=/WˊQ���a�<�9��~R��F_M~���=yI��L�b.�
����7=�`��F���mp&�n>x����/	���$��/���8U�v�(%��~���%4��������r$8r�8�8�G�8Q<YҫI�e����.��!�F�H�<��_�{�ꪽ8�e�ӛ7o/d����g�}���G��Z��hT���`��M�%>�}��"��P6�6f�v��bO�l �$I�i��!��(kI�FWx[R���Mɟ�����D�Ӱ��=&;�Mқb~[���M��Cڲ��|���{u\�n�s��Wc���B��zF���&QU��"�+]���鴁�*y}��:;�L�2���x{y����C�}fV�{I���zͱ&��"(Q�`_�9l�E(PL����
F�����\A�^s����T�C���{���I����T���xQ�|7-�w���Q��3�seq,v�8�)B��::-��m���2иF�V���?픥(�(�>�����D�F�7O&�.������CI�ʌV!�pHՋ封{/Fpt�n C�����)��S��������:�1����'��\F�Jq�o��#���_y#+<�9A�#�)����Zi�Xr��4�*��m6Vv���Vl�Jǳ���y��n��n*��({��|`��|x&�Ib�'����C��i1�����v�ʮ}���l�E�a�)���O�[_�	��ENM�#��+�	���5ɧˊ�4�	�3����O��gHZY�B�f�]���z�8KQrY���Pn�\��aA��і[�/[Y� P��CS�#i�/��lp�`p��HpCqM�b�75zv�{I�i�X�4p�
reX#��t��5�ۑ��6=���h����asV �)V���E�
~V�\�Ч�Ul l�QԜ;PH��Yd[�c�R�I.ޚ$�Aܪ���F|��[�]������&�OO ����Z���ܜ���ɫfE��9	�:P��v���d�1œ�l�-'��]�B��l9�e����d���?�DG�+xLa|o010VYI��E�dU��V�Y:�b�^%��F2�>J���߀o�$��߬5D[�M�8���07""�`R%ti�|s"]��(�w�g.W�v�պ�#����P���!��,���L�� ��GK� ���ݕK��;Q8b���p��X�����9@��$�
$�?}��c�_6}�Q�{`���t��������y�ڷ ���"�Z�Ta#X�]�>[,-����
��!h\-i���x�]F�E�6
��������.&�/�+l��I�8��4U1(�z��!%�[���+D�S�OAOs�)͵�7l�o�_~ي��2���3�b��Di��kM�Y�m�@�kS�W|�!�p�ч�FΟ�:g���=�dЬ���bJ�ѩ����~K�l��Է�6���T霢��^t�9�ڕ,M��Wx؀mP�
v�i-'�{�Լ���[���Ů��GM�#�"�� Qp>�0M�hY6�֚�ɶ@�����KN8i�>����U� � %��!A�^�~��1�צY̑q��D��̃z��1,]��E��ʲj�cOj̉d�S�K���w����E�6<F���bc��cq�R���
�b���-iI�/�����{>t
"�X^���Ǐ)���&=L�s�1kiōf���i�=9����XzS��1L�#eve y�*if�#e�	�n����$���bx[�V���NAeG|��#�%�CO�ˈ����
$�|�-c]<eI̦�+yCX��P/H"�4�0ӂe�U�7@�	��Y�@ Lfꪱ ��!���&�����3bv>JH�j_�VuD72Op�<��W���:�:ɲ�1��0O�M�z���^���cDפ��Ju����h`��H�.�X	:��E�� �@r����}Ƚ����2=���c���S��Z.�g�d����[o���W'@�=��@��Pf�i�g�]9�v0>f�Q�l���I����}�_�m��k�qgL�7Iv���D�he�L��w�,�(>�����͍ŷ�
�E3�rQ��S"�+��[$%�%�K�-��� ���<;�x�J�'3e%�Y|��dq��a��~�7N �����8}��f:�4�gx�L�����UH~�ަ9��	���#��=���9I�~������g�����9k-�H�HR���8	�Q2eRn���L�iR9z���:�yA�g4`�Y�ͺ,��@\1����x#�`-ʶ�X(�q�诘�s���s��W�y:���b8�zUM̩�����3ۉ0��H@g�g�Z�'��9;�p�.x�L�"|�؀�W�"��[d��}I(8�1��S��B�B��e�ު�D*L�
�x�DEF?EǤ~��%a��cTcNS�TLYG�����:�%w2���?u�}�?Y�D���p2ɮ\�*�"���~h��h��o�W��k�O��6kss�I�R�@D��E�2�v�<�N���N$�𳕉2�si�^��5t�B��G?����zM�"1gz!Ӷ$Fͫ0g��y�"��u	.�_�_��Z��.jr�$�at.�4
�J�����fuy~�["�K�7�	BC�0�+���#T>W�1���7L
�y���<;/W�VjD�1� @���,b8x��.��Ό�	�T_A��d4�����yr��� ��Ǔ��/�4.rW��3|W��K��ӣ'����Yׅ"#ݲ��������TNM*i��3��d���L�"�-fl�y�b���\iAư���aPb(�?i��#>e�S�]����E�S�}ەSf���G��^��I��/f�i'Ő��M?�T&�l��r��=�<��b���ֱ��ed��l�3�a)�� �&?�Kp���Ñj24�R$���R̩���;����+ž��h�T6�x)t-6ٸf��;ҧW��
d��imX8��s'I�|�	@�Z�-J�9'��5�X<�&�<��E,ʵ�g�cM$
jt� д��r�)
�-T���):[�n����x�ڡ���CR�Y�$N�l�lk�c�ͺ�eq`{io���H�\j�	D���_�k�O�����]ƕ$"��ݖ�7(`AObO�ؕ�T8�v'E,şH?��#�d��!r�V�.999�{cqh��ӳ\&N�c~�F��1��hE`�a��b��,��4Gx����9�ۘ���,�yzd���[��yL�z���^Ԃ�K���[�^r��@*��i)v&��h�XTp~V����.w��!�F��ȷ�G����b&N���[c��%�c}N�����Kh�N:�c�� �c7F$���=U����4UU4p�$�I����F����6/�㓇ׯݤu"�MRқ�bN�.~%>	A��IL�:����H�8��Nik���E���I��ɧN�)U��]R�*זd��l�V\ɘ�8mAG�H[/�Z$E�����+޽|1g���ɥ$���64�����گ3L��F����`^�X�~plR��MW��#����Bg��P��!V�Ǒ���ara߁�3�$�9��->GmR G��#��_����;�4
)RU�4r2XFLVwi"8��:�z��]��C�s�`eK
#�$M�Z}��%.�?n���@k�a�,5`�q���`1��.�7�7/h�P�n0O#Ӿ�~��j=�+�R�/ =�[[و��ђX!�'�;p�0�2t҅,��?`u;ɺ&�՛L?p��]�^^y��{�=Yy��z]F���/��!�c28��cP�;굒\fZ�$)j;�V>p�[�0�V2Uq��j�����n�e)��bu����\o��H:rH��Zk���s�n"�Dm^���V禵'��wp��^Ru�

}��'��v��.��e@���A�����LVN�H`e�����dz��_~�����>@��R�5w)��yzz����@t۳ł+X��{�LE��IQ����֑��� �4���>����D�����1���@ԟ���|����n�.B��ްZ/L���8r}4mEG��s�9�L
]�43y#��
�����;V�''�ǽ;�!+���x�p�.�W��L?tZ���o,����m���dN'���;;; �Bt�7 C?#��޽���#!?͕�x�"�ō�W���7�}�}�N�KB��\��W�2=�	�B_!�[��K��+�=<��8P�YE$K��|�F�Lqxۦ���C��Ŝ���Ȟ��#�� y�d'N����S��Ҟ�쒳���QTź���F�>m�[o�u /Zؓӧ�Ex��)-�?�B�9rv�d�G����e���a���K{�%ܷ���z�k�^A����:�Q���.���;?;����LQ[ �7�oR'2٨}�֤Ӓ'N{/i���W���ɕ+{�߾I>҅4;�7Uӆ�rM~ m(ս�G�&���n�S��"U�V�jo7�(�7�	?����G�6����$��8��:��t�y�T�c����Α������le�]�K'(6h���0�E&�R�
(d���9)U�2���ORT,^x�a�K��~�j���Ƥ0�<0s�3Dzu$���G�M���3\ MӢ+a�d��^��A���om��&��s�./��L��v��d��S	=���1A_��y�^����^��L���=�����?#�z��Z�wm����wN{H
��ݭ��O�W '�^���������^7�3�M�:ù$
�Ȉ(���N�o�	���a��S?�oG��l���%*����7/3��UG��p�r�G�K��X��lA�@A���N(�s���N�4(���\^��p�NY�:�� ��^b��I8����I�oQ϶�2TB�%}��U����.�n��%��,�9���P��-��u���l�6[�Bx����<~����t�):E�0�&;;�`{�X�zB��"��Z�
a*$��=&��0@	�&�,c:g�<�g�LKl?�:E"D�E*d��u^�)���lje��IQ�p
�@�T����199^ˡ�2�mי�&�G�Uxn�<[��>@�������a���C�/�����ו��rd)�2�$x��0��G����p(6���ѩ@e����yj%�
z�x��l�șW�+;�XLZs���ʘ���	,u>ҝ��BXm�{F�a/NF����^��f)h�-M��>�ڷ��G{��E��r�ۍj:
Y3zm
*����O'{  ���u�����޽�ӭ�7L�?q�\���jt���[�r�$�x�|�hX�*�
�_ܓ./��k4������]AJ�,65�Ym$���2��Oy� EI�̴әH��n��k����B�-���R1�f�
O�0��n�m�B<��������_�t��8M'�~I�֭[}���}#!hk�:�
�֡�l�n[A[��6v�m�h1�
�Cl�*PJ����ʁ����V�4Zms	 ��%�dPn߾M�F-A����D
<���l�H�/�ll��b��>�ה�X��f%v֧�V�28ØrS[���ִ �tF��Y?\�ΰ�a>���cҲ_;�h�^y�?����8E�v�A�Ŗ����F� �U.��������Jl�!�';cV�kb��i�c��s��]��,Hd:��Lzر�d����1�g��}����[�_�	�Dr?[8'��av/� �Y�X���O E2]�� ��vx��#���I.��幎>�
1þ��tZ˄��|��;�#P�g�E�-�M{��(D�|���!��X0f`�=(Y�ԥ�M햆h+��i�(��? �P����5O/�
��p(d8Z·L��4��Wbn]4a4U�N	�P��xb�c���;�
�u��d��%g��ӌڦ\A�sNa0�sz��=�BQ	��/��0��u�;h��G��cB$�d`9�um�-��(9s;;c"�-��ec�S;��}��
0���O?C�Jf�Lj�פ��t�E��:�RP
ʰ���eJ|+�@�� �\��a_�_����G�E�~2K�i�c���uD�q��l��Z' ���c�{}��ec� #�G�GW�^E�9�`5�ժ\#&5���{}�k���������{coo��o5K 6w�&�����c4�����!{�����N�V�FZH54*)|r �8-3���7/,ؤX�� ��h_ �#�Q��ȔDf�;�����P8Y�F��t���1L �2lS衎;��T�H�I�)Fyt������=�s��LhTn4=�sL)g ���nR��QP�}��ܸq��&�>��,B�]/\5i f���#���SUQ]��#[tjk�,KA�������Đ&���Y[Wq�0�:�g/��򫯾��Q�Sڣz���KO�֟7KgzG��@�W��$`��ݹG����<u�@��	R52�'�:v��u�������(���� �u�P� �O��ë}��A������L�Y>��P�M!Q�D�Obw��%�겶����Y�rq@�kFl�jЊM�,~t�t�#�>�юm��8˥qd�t~��D��_%[LdGq��$Ż����cr�y�rlv�fZ�In��F�#��,�Z�K\d\�6n�3{��gu�D�Hg*S��⸘�ݑ�˓.���L��(�r�l,L� ��9�۱��_��=��-�&.&'mk[��f�קN4�y�\t��u�W-t�""�P˸]2	vV���{�9� i@��!tvW�q��'��'�)?Ѓ��t0H��GT��ÈB���Tt�z������8�R=��ı����_�#��k���*����B9��R�" "�Zx��r2v[��H��yI��Q��,�v�26O˔)d�;�ꒇuR��P��L���T�kd�.�!mA6����)'v&c��=x$�&lz�zy8�N�	���:��F���ˠ8P,8k�PB6�@���5f.7�5��+����a:̒��V>�Z�P�M�3a��=1���st4ގ���bx��]eI���di����;�K���g�g��)W�7�m��v�VkA?ʘ��Ѿ,\�12%.$��;1��5Ww"J*�&��!}���$��GV&�V&��0�����$O>#<bt��������b�u��}Ǐ�~e����?����1"���HW@��)���%���y�jh���g)x���L��;����
���sKqC��L �������|.�s����
�K�^��c�0�9i�r͞�f�~���nkf��F���e@|A�O��)���
��6d`;���^�/g��7	�eUL>2�}���H|˧���P 1�y_���Ud\�(CsQ�4&b��b�,��5L��ӭ
fa2�XiO4�x����&
��=��ɗ��ŵg� �HC�z�mky���K�G��>{��w�MR`Ύ+����X���GPL�\�`Jb\xf�d��T�1�ǧ�T��m�X]o�Q���_[�TѬ��>60v�?5�y���%7C�ME���r7���� �餫�:8�y����)ޚ��]���q��I	!ha��B���@`?��L1ߦ�},[��MGw-�o�u�s+�xp���'O-�t���'�$S<M-�lX�:�b=��eꛦdn���a���B�YDj�3�0V���]�Z���j��#+Y:����IpJt�3+�N��d�RV��'O&�����]T��65�՘s�N "�8��	�{�vR�K`1������A)�劔C�
�e����q�:�U8z��"+gu�S��&���jCvm0��$º-gn��8$�=������i�kE���OVW������ώ��"T�����d��pť��ۂ�L v"Ʀ��L�,���:��!��N�-N�Nd�`k�	e3��N`Khz��%�D�7�O�q.D�X�Y��!4d�ʰLV��?��@K�!�R�Y����JYWR/��Sˉ!l(
���O�Ia����mYT�g��g �XC�34m�=�62}�)S�x�K��a[�ȣGOH.>�!���l<�YK�pw:D" �]�D���)�'
�H��'��Jjϱ��!�og���%�Ұ��|�FB�4��ݎiR��Z�=<'��a�7����I���I(���x,�/�<&O��O?�;M�y	����`� 3���э9rX�~��~�@�Z����
�ޑf�~�K�u��4L�X���Y����V�i[���O)�(�S�Ӳ	�]���=i��K!�CN?�}
�d]��-]�r>FL���ܹs�����񷾵����{�������C-��@���\y�L�Bka)�@7t]���{��V�*�8JV>6�ӂ����9.i�E�d��w��O>���3��8x�6G�c�Sk����r7u[�r�C-@������.7��`I��i�|�ʍ�~H���˙�B�#})�1Qp�K35�	��J��F'�����&�QBN	t<�8��*- fa�Q�u�N%���e�*�hg�N=���)���'��u��N*���R�<�9�Վ�Ļp�/0�I7��l0�t=���5nr��
&���ʗ_����o�9EfVX�#���'N�SRc�:�oȄ��t#�
�)�&���=��==��s��ӟS`E�źE�
z2Zd�-���M$@��8�WJi@%T�p��ⴊ�3��,'':&+1�@z������>b�L�y�޼\��6h�	��t[� �2Ct�n�fp<�H�Zœ�/�r4��{ȯ��t�\�@(*���n�wa�pІ�]$E;����b�X)�����k��/��ð���r�m˽Cϳ��R�Lu_�S#:���B� Ȗ�?P�!}�o�R"��{i8,V]Ej��,��[X�h�'D��#lc,We����~�*ڼ��T�A �,�r,�T�?�
�S'Z�ʙ��'����W��3�ojהT_��{�LT��b�%���r@*��*'i�$;�gds*p�o��&@���Yq8��ѴVJ�}�n�Ub�h�����H-������T&�t���C�Wԑ̩
2�6(��-/����6���x#kF����� sAT�8��j6	R�? Z����8���0VPa�����룣#�Z��>�,GxV�xKd���7B����W`���K�8X�Z�T޸qs�����r��5%L��4�E-�����8�	>���>2�*�p�'Z�_�K��1@Y�2z�C�{�U�x���n���Ά,I&�6�N�-V[:��T�򤃿�C$f ���X�+a%��q(u"߷Y3	6z	�{�b��X^�����܃p����~��RZ���:�{۟�O%�皈+�:s��F!z|A��Xj�s�5?N���X��q6�Ge�T\�>�����=��	���@jԂ=�xv)�hs W1��|P���G,Zkވ��s�����aJ��@��=`�xZ�n�uk~�S�4�i4�4�|ٮV��0�.�Y�)�$S�R�I��>"Z�4T�N��n2E��������un�d��A�,�����q]E�d�W�_�dL] �R�C�R�p�i��-P�,cR]���"V��WA�^~�6B�- ��U�f/�ھ|c��E������za�[��pd�i�N����Hi ��7��K*������
7f�����g74�7���zq�K��?%��B��	�0���ۘ�L;o��d,�S0��&j�fě���t�K�tjbԀQ��P-�����V$�O��٥4�DJ��朶U�04vT������Etw��oP��������9���ӄ��s'��$r��U�Ďd���s�ƹX���0h$��H������ph=bЖp�eN0;� $�F'���[��t$(T�-%�%�΅���O��q�^�ͼ��� ��7m�}�ZV�C8nWPg�tiLe�0����n���8a��cͥ��oQ9АPz<~Jd g���{E���4�aa�|�xRx��ٶ+"Y���N����x�ĳҨ��u�/�15�E�^Ђ��y����R��[�o�>;��ie�r@��J$���B�L�>�y��A9̹55b޲9�|t�	�d��{,c3�-6�����\�tf���g�<w�G.���r�9�ð&:�	�fc-��%Zψ9�Z��n0����t
��cg�OI,�������lw��B�`�Ӂ��	`�p��%����3⻠�Zm�&�@>!�����í[7)��|��W5��lnLdC�ԽȚ��2(��2&��5�}�:���%�-C]+#'l��e��<���Ŧ� �D[�z|���{�y��ÇXx�^Q�^1���Sc��tw-�L�"_Թ�`1�a�$RhL)��{/Bily���^�Z��ó(K��kP,f�\�b�V�2G(�{�:褗%����=����������n�~����M�>r��m��r�q�>�"�~�Uz�����߿Oo���_��h��B�Ћ��82+���@o�jtC�1��@bƥ�܃��`�s�Wˍ���0��IB��Y��:D4+�0 �UU�I]K5��OS%�Gl��}��4u'`F��L���QG�az=x�YǕ���!4$�y�D84q*9	�b��	��N�[t���S	@��,a���[$��trc`H���5��'���?��c�0;�p�c�<y��C&�e��8vvF�(��7nзLw�����?5��$������L�m�M��r���p�(R~��/<��s��;R�*d��AAĹ�ՙ��s_;�p���F �l)"]����۷w�K�	�9TWo�͜IV-��m�\���#�B�ܸ|�%�r��8�f7�6Q٧� V�4M<�� 4�7hU�R�ٺ�tf���^��^IH��`"pwZƫt\*���ri����r�0�E����y�<�\!N�N�m9=���f��^,gFK����x�b�hK�oݹ�b�O�Am�{���\�e���a���NP�y9,�[a6[H�)�n<�������fu�����e kvi�ğ�$� �-�|�(��n���z/9��ph�6�	"'�G�L1��㣛��ҽ�e������8��:����Ǳ.��o�J3��~F�\���g�6�
щ���XEXX9{�;�&��
@����g:P��t�aψ�cx�x����R�އ0�^ �j����b>_n�޽뒼j�bUr���O��qS_��
�Xse���JH?s�3��%�C�(M��|�2����.�4�¥��lB�DB�*�D�^�a&zrz?9.uD��Kσϖ^gA_X$5���bd:3��KeVi�T:țqR�E����D�����l8Z��o�)�I���C��$=;^4����pP�mH�ݹsG�˳˳�bU�b2�G��ѓ�.4d&-q�%����>��b]ٖu�*7��<��5�����M�8X	�L��fq9#/��W������Q���4S��9�xh�~i�#'�,ӦH��A�i"�x'�~
mHI�V����v�w�<�;�}�W_��/~�������q�r��|<���M�]X�0�y�%�΢*ױ�IZ���2䓤��8��������4ժb.�E���K�E@P��y1(�լf�:r�GK�Z�;�U�b���8����S�Ӄ�{)��h�֫��ߖݡ����dP��w�p��W^yrr��G��Ə>��T��k���j8Ѣ��L�fPWm�sIc=[��N���i��D&N���U�MW5�aȳy�h�r2`��ْV�w����fI݄<��t�q7i\�O'iI���t���!7iI�QN&�[׮eiR����x W�����^z��#���GG�fD;Nbpr�d�\LE�".��Z'p���K��mm1	F�y!mN�H�P�z�I]�֫z2�;,F��T"E�I�Gve�;1|�2v�$��e�M���3�7�%��P������(%��^������^��d�s~qq��dU���H���u��e�b#s��tcŦ��u)S�y1y�t�I��y.a1Ȧ�	�����@��\��%aj~&��!�Kn�<:�D6�:�f�	�Ua^�" 8� �d"�j��f]{FE%-�"٤�IU^����|��-����7n��wz.������D>L^���V�d#R|H��w��j��7'і�5�Rِ���&� ���[��Bd��Ee<�ߺ�M^�/Q��N�4������^^��w�o6�Kf��O_�w���p��o��o�"�//���`���Q*`C!wWm����5a>��$L%'%sQװhLgNn2�3�i�2�C��z�jS��c�D����d�3,�0ǻd�B�^��� ��2�gg2a��F|�a��I�5�^:,��͕�q�~�˯�������b~���N�<��m�ʊ��|*$�sc^��	�
5y$�H�<�L��fi�R6��:�#Y���.�u�TK�͔\F`�>��p�\�#ީ,	o��d8r9Kr��Ο�����X��XB|�.W�ѽ��;��E��=��� G(W
��T;����S��s��l�<�`saP���c���^7�D���42b$5Ն�MG��ֲ�&�A]kG&���2л���N��\xęL��6�բ	1�@�b^�vM�'/��0�J��A�T�R�c٦5,F��_���yRsz��G�=2��h]/q
XZx.y����a�a��³'=�ơ�@tb�cķ9�R�r
��#R9��<G��!5�(���~��\`��v�ڡ�k���N?	(ɑ7���O�V���RԄ�!�ۑ0�&�X�b�d���� 	�)`R�R�jT�:a
jqB�r�0C$}�<+�����q����Ea���G9�Rg���g;���R� �%�n)o
������Y=�N�/j=�V��u_�9+��rG�Ңd�X��Ȼ	Ő$��yS.k
7���q��<��s�\׮ҿ�W�^uY'y�	R!p�4a�� ��� �_�Ō��pzbC��VtZ^�(�X�hC�U2w�cW�#�ق�:����O,�k#cb0ҁ�t7�O�I#��t<�����S2�/H���͛��#���rrn%�T���Τ�G��CM?���|���"� �#��TqC�G���Z�ղ<ݦ�Z�v��!!���x������a�֧iɰ�vI�0K��J|0�3�7v���˯�읞���B�O?���{����t�{>�A�{���w�!��^�q���ŢZ��wYڬ��>��+�{�����1�G�sh��mXP׀����5���%�V�E�S6(�h��$i��Q|H������ �G�V~S��:1���M���.;_s�M��d�9��U=��D�W�G���a<�ϒ>'M���U��Y]0s��d�g�I��(I����d�H�ԅ�]..^\\\�r�����'{{��p!�Ą���C%�(բL�A�t%�qG���*�E�.�?1FΤ�kIIB��CM��Jv1�ۉ�L��$�v������� _����<	�/[2�U$xck��j,A/�HTw1�f+R}�0��5:8ˎ)������_���]�62�`��R`�Th����Ha&V��d:8>>y?I�d��i:�q#�Ü4��`I���y�k�l�E�l�h7�Y�"��ӱ��z�@�e5���]^��[7�"�ry��ymw��\��0�����t�ۮ�v�+�nݪW2�χͪm����lV����{�R;�A���ߠ�,W۝�(4�Q�U1�&�݀�]/-�fT���:n�����̩�:a��&EV�����x��T�3��:%�W������G�թ圚��n6]쐚S�������������-�Y�u3S2/M�0Y	:���቙���6���eּ@��?����%Y1������5A,\L���Q���F3���I۬Z����hdpj��i��$=Z(X8a0l�b쁠	J5b蕘�k#y$�TyX`�`�e��-�!�թrZZ�ǚp$	�}�s�%����Q%���q @��Ht&]k�,4(SX���ՖUz�b�@}�V�Ldu`D�ph`Qs�g�{#���r<��bz�����yT� 7���B�_Q���H���0�
�����:o��.}!��.��!�E� �a�0�y����O?������)�4UuȃAH�B/�V��R���(�B��n;0Y@���UKF���ab��K��n"=�AF��w_z	(�_��-�$\U�D�r�q.��t�K�����H!q���&�HUD��5��O���@G) �$r�� ��`�i���,���̬l��tB�������c��P�T���G+Ħ�S��V��$�bZ4}.�1p�׮]����:�g�]l� ��zԺ�<�fd�"���?{þˠv`���z�C �<99��O��_��:�#x���i�&�z�,��r��g@=��=��6��-�v��x�,]$�B��]^.I�ɔ��y1jt�p�7$_/���� �XF�<�2��2� �U�?��?��/���e(�����~����@R@*�?0O[�H�����۟ʌf�Zڠ� 2"�8j$JN7��L8/,�؅�όa-�D+A�pocS.�2��� �15���_��K/���;�����=Y�a;j�s��!��Vi.� Z")�ITz�Y���f�0�9'�� I҉F�Sk�n�#�T�~q�دU�c�Dd�崈���	�d����oW�?�;�--[.��P���FA�Ie+&�¹�/V��	%v���OV�� ӕ��$����ic7�����-���@��'_��Wh����*6	r��OCihN�l�J�)-zC'�,ȳ@c��O]�on�P=PK�AZ8XlD�-:�1�%x�֦=��+����-s��O�>}��]ڈ�7���_��?��򓟜��Wlv�w�ň{Q�1�Dp�b.������l�<�d�!� 1��6P80mKa��x�R^m�Zt�Q~�b��U
؅<|x����u�(�V�>mC�#�aB��X��e��"?�jӒY�aT���d�S�IK(��$�#�.��w��
p
k�uL� �j�qPx#.��0܇�Ȁ����k����2|�.�}��.��ڈ�wR�-�R��IO�.��=�,k�)�6�9�JX���*���<4S4���`�,�e.����y��{s��PXE�}�v���W㍔��]�J�����A�Kb^��@�[�!�[��>��iE��i9	:$��q`YΠ��:;e9���A�����{��p w\�<�b��H�nܸ���'O��ڜ�()�E�q�&���������)���JhU3Nr��������@�3�7��:.�S���q�-��@�#��{g����
bS	�	�S׌C9?���G���W�hm��`Q��̰�!ˈ��3�Ӌ�����G)4Aq��P �NRb�P���G�~@f�L�e�[�]�R(WX�vZ+ї)(Bh�\�E��2�s��ˈi*/����9�'`�8[M[���=��[�<Ϫ`?n�$d�89�SD���ߢ��~�k2� e������N3���K2�:�N�����%����)�m�1bF
mF�.��$�<�z3�K�I�p�k�e׀�<��''��Ɇ�h��&��JA��x�h�t !u&K0�n�z�7rIL�.���c+=R�d7���BQp@бԦߜ��ǌ��R�6��\M�6:��Z�D��M�k�-�B)l/� ��Î� ��-	t���\�w~��Sm��5{��S��Ç��NN�����C���ޝ�X��Ac�+�92�&3^y9����j��5�u?zZ[�p�q~��g�1�>��S$������],�бz��X5I��x8"��=B�	b.YL�!������8-��tZ�\���Ynά��3�1��8�1Y�h����D�T-+��^fC�-�06���� ��>��ƲG��F�~�+W�צ����������<C�ε�ӧ���\���߁�Ƕ-���4���ĖܩG�w��7��|擲�)7�"��|���
ԧC-�>�=a+L^��pE2n�0@V�3�-F'�Ux�d�`f%�S��p!*i���x�m�T�����8m��r���|;9���>i�i���\��bi�ߍ]��+��6���XK�;�ɻ�N ��M݉w�ʓJ�F�ί�]RV��[$F�p-e��y�8���B2���&�rpt�����k@2��ᐢ�\�jr�;~�d��$-Q��w'�yDA[�A^_.��g�4�B���U�����.7OO�q1v�v�l:�8���D���t$��!���Ȏ)�H�����m�\��d�F��#P�>I����eݍF<y�m:A60%W�%�K6�Tە+W���m���%�hn}����ȩ�l���_ȺS|utt4�q`0E�8�@G�[�P���X״��юV�x<����g~�ѵ۷\�\�q���^%��,:�jpY�.׋M�Ѐ���V�Z�3k��~�)��u-�$�u���S��F��S��VdG����Ӌs
��_w
sN�����
a$y$���'�� rL�yB��gg�踿�更,~�!y9�E��d})��.`�hd:g�f5�]�.�׫EUoR���ۡtxp�#�nǋ׶M��!���/VH`/c}�pН">���.,\�ݛd�BJ�Z�������Y�&�}������ǣ+7���k_���_������7��ͻ�|L������圌2;�2���&�B?_^�,Ȧe�!�3J���g�y�
1���5l��Xf@<��=i�a,�F$k��Y�j'���^�`�z<�>]θ��@{6���������لy��s���_�����u�u$�F<{B�/j���ZrKX	��p8��ʋ�?�=��W�ЌN[}�%��ō�ā��)>�9'�K�Z�3 �5}�ɴq�68��&=�����?�ݣw������?=��k�g�Ʀ�J�Y-F�2���p]��1����h��'-K�im�m2`p�E/�H;���%pp�W�����0mCE�����"ج�r��r�n�z�/��/H��?��J����\��zOʌ��圙��yi�� jJr��%�0��q�q�F6C�
sX���*1tl�k�����P훳�4����\"H|���}�K_�?����}�o�ͳ�'�lY�i��*h�u*c7��<�����3�� �X˄��I��� f�$AZv�[��_AUZ��iȮ�]���5����5��,7�G'{W�vw���;�����������Э�:ج�|��:Ǧ��T����\�W�����N�hz�e�L���ܹM��<D�X�
�HW�%�y,[�|װ��N�h��ݻw'��QjNt�|��	�� ͖�?{tv��X�F�%�Vׂ�ʤ?���B�:Q�Ӥ�Ė���(��~�����0H�hU��$P,��J�:�T?�Ht�����Z�ŒX!%��1f|j�m�&LN7���(w���8�#TJv
$�$��o�>�B�N��w�H�*TkܻM�{L�������*'#=�܃ǁjuJ)ޏ(���I�N'j#N�����\�M-YiQD�DN�P6��Si6�6En��f��N[q�q���P##	�� �z��+��@J�CW�'��h�}cq�IA������+/��#�-�������6s!�V������`���B����1,E�����o�z�4{=�^�)d��Z�&�_���P2�&�� Ϙ����uuS�x�c)H; �	$�.Hns���I�`:n0��gd �u�4��>
O�C�0��4 Y��$����Ç< ���7��5�^�0�z�K-�L4�y��H���L
�O�<q
�@&�1$R
9L���
���?O����)���A`/@5�-hB\�\	�o�C �W��6R�`r����F�^z�%���ȸx*:�����$�yछ��H:�����'|Ƞ���ڽ������'7)ދ�����>RM�c���3�:ku[N!�;4�e��+��
K�Y���\'��.26l�K1��dD�x�a8A�@���C������������>��ɰ�������Q��e<�ٖ�	���_0/њ�[��+�����i��/v���X���:���'n��7�q��+�QE�G!M��VV(�>V��Evm�ƗbF���>����)�H��x2�N�c"�|�.�M���̭��B�)�L�<�1)��\V_�y@� <�X��0�������~9��ŷZ���LS��-��e݅fqr������=e�Ŧ���]���z]��ʧO�i)��R�H�r���|2�!�)�&+@q���c�'��c��N�f�`���+I���`y4�P|�
�c<�1�fr����,��P[n`�㈪�7�PR~�h4�Et#�s,�ȩY�M���Lz ���[�H��9�9p�	��]����o��V�b(r���T�H�H���r<$ER2�f˖k�ȝ�JMR$����,#S)��8'PL�L���o��!YV�wZ�Kt<���o)�hv�	n�$@�Y3U��m��f��V�0L"�E��:�o%G@��1�����H�� �5�H�_��O�Y.Q��_�*��q3�A9�c��@�
��YY���`(:.H9�d��/x#���t��ن�%�.�bPpn���n��������S\� 2��MѦ��B�٨uZ�2Љdѿ,/�goݺ��U����B�������<`,�a���G}D�	��VR2/�UP[�T�)EK(��8�!S
?l�kY)@[�A�x�l6�r%)�?��w^}�՟��'?���E���$��`z�K)�I��l'_�U��r�&�yo�t*��:��$5U�3+�nA��U�W �:88A��cx�'��@��f@z��	�T��d��ao��k_���o����?��?�<E^5؝���������T�y�<���WA��X]tjW�a��NXWoV�Ti�寑׆KpMk#e��]ŧL$g9�s�Z�i�_=D���r�dD�m��`4P��m�2�D�,��Oo-���� ���#^�P�@�z3��4IT�M�,,-�D���q�����5� �r��a2�݉%���v���)�(����o���Z�T� EY�%��*�aJ�gg��R)>po\�;?�P|w*ǁO"
������A�!N#A(�E{˷�We�=q�3��z��A���
�ݻb
��կ��^���;O?f��Ʒ���Z�t���5}d���[�L]c�z.�4�0�SMt��`?�oD(sW{�����}�,|S:Y����P$�����ɟ������7��4= W��0�UŃ��L������93�,K�b���u.T�������$BQH����ȧ��(���#�j��_9����^��W����H����	0R��})�5:!B`�*t8t> f0ߝ2�$�����"�2Q��tQQ�إ�a����$�I�yZ��O�3~���)�>�wH���p0��?��_�������s�^�{�n���%=l�@*r���2�-o:�qx�U��9��bU���kn��{��+:ig�����޼y��_s��c�f���=K¾��،5X��Tp�deb�S6X.]�2h���\�P5D�t:�����0w*�K˳H*9��E����OM�,���&�4
�X�
�G�)�~�N�&����Zm��-��bJ���5c�K�2~6�[g2?Ғe��VE�ʺ�p���V������/\�Z�SB� ��R�4���[�)���>JD}p�$��t�j$
��sn�N�/�)�����Ax��m�@��c�{ՠ�GN������S�Ra�%O)�	�y�ӱZ�X�#�+Cxl �k��%P����YB�ʂ(
p������:�$QJ�T)}�P�ҁY\��K�$�t	Ԍ<�7���$|]R���@��֓��E���*�> ���E�{�h)��`6�����F�����D�"��Ō j��7�p��X�<g�ڵk����9�CZR�>����&�m�-�5��������W"in�C�Y7�zPX0S~�ZI꽚!yg��\�IrɘnV��8IC�7n������2~<�����<�gcW.����}�1)O>H?�/xY.sr� <�|�]l6�1�=Б�r4Y�&�y�TH��VX�CR���Ԇ��AG����n�I�������#��{�hO�^�*y��_�������>��o~���O���~HO��l/��ؤ".NfÁ�[�(9��p��l�0���7�=s�����(���o�����V���
��k:��G���㦙������mm!�	O��ȥ���3��`�z�bv��y˦3��w@�0�s\�n���6�: ǉ����Y&0�<�@{!c�E�	��,��(Ol,��E2��N�n�D�3�0�{����N[^pr ��2�<z�(�y�A�Q�//�Ы^�]�xǷz�9�|ȍP�Ʉ�̎'k���D�~ˢ��֫�$'�EC���F����)���a;w4�75�`q���䋷��I��%^<!�%'���[1����j.$�R�Bϖ�qȻW�3�sF�= 	L��[�/vi�^գ�}ݛo~�w>q�iR����׻.��>���G�����\XL�5�Q����,L�Ӫiۛ�4�4��B��`����Uc�WV݂{�l���W'�qZѥox*����{&�:��KÆBk>쥐�D�sޅ�Pȝ�VK�G���Z{���'O/��K�&�qJcl#a���Y[^�����Ƹ�F���C�fKh�-��y�N��Xtz��p��"!
)�,I���N5=Qu�l-"]�WpɕB��Y(��^���{{�4;�U˕2�r;�k�P�E�[��\p��Yo
9ʚOc���T�Z��P���H(�ȋ�W?>���/}�K(��&D�f��*-Xgtǘ�K�@{����ю$�k�m�������Zɷ�����W�=(��9W�VV�|zr�������o�~�5W��w��/��p�i�Șv/c(XI�c ����|���	�U�9��⡚qy\�`���b ��4ɖ�U��(X�ff�lBS�81����
ycMx���)i�a+����&A�;�$4���� ���'}L7��/~�'�p��{��g�
�4�'-��zsr�4�y)�V�y��z�ݝ.���
OL��AW[I�k�2�
��kD�X��������@�YP!Y�<��Q�@��K�1���P�n�t�i����l�x���_�⤛�����W_y��O�s�x�%�(P���[�J��|��D��@nE��-�Y�M>aS�+��U����#���u��O`2>��آ �PoJh�1g��y��Ls����j���O~������\�N���ǩ��w�uu:%����#>�|�:u���I��Dt8� ���NQ*���ͤ�XݦҰÔ�2!6I��kH�d�2ԗ��d;��4Iv5${�Ů�N2c�ȓ'�v
:c����lV''O�]�Nq��W_u���G����7ww&���/�<yB��t�»�A�w.�0���U�L&�aO��a$�SR���b�AԾ�Y})���|L�iG.Sn���k-�mf���]V8�����f��w��^xa����ѕ����<���1yf��O�D�>�`�O�H���/���d,J �,�HR�vu�F0�b;j� ���C� �IGǕ�e�?R��rL��� 3�8��ru(�%(%��g?۽rx��'�v���o�����׿�Y��ˮ���bXdE�YCV;�L
eqd�Bc��Y��I�&):,:�k���[�*�)^�cI�$Jr$v���j�%��>>d��dr�8Lr7�^��7�p:��}v�S� �(��dl����<n���<r*^�`�<'��:��BCLga���^Mb���)������B����sF��7���s�I,!l�9��5�Q/M7}t�����٢*�>����Ȏp�K:ߵr�
%t�^�F��xބ���Ȍ��
�����:�Ld5��tҭc~��ڃ��́��yL ��{�������ɐ��g�G#r~ɗ�\�hۤ����MФ����l`Ľ���eҤ�FboMk�ѯ,_�*�XH��-�\��*
����=&�.kl�T��ȨV�M�,':�Up� v�`�z���h�3��R�)E�]JW#mtr�z�ld�]fd-�t:��;M�F0x���ՔK���Ɣ"W�Ce�i��;��߶dI��̬($4��H�ߘPYei��ҿ�r 1m���Aȁ�$�aj�&�!��(�#�"��B��{��N˱� d�,��l4�����e���]=���U�M����=~�y�#��4��g��t��0�!��Ab��	�!���O
c�.f<��f�Fƪ�V�v��u�̽ٗ���bg���p���>{�����	��[���J1r�('���]�7��΂��F6*h*R�j���^4�pxn��$��$̈́��$�+�<��LAOm{?iA�߿������ �r�9�!)+z���z(@ۘm\*������Ïٗ�zq~9���]M^e�T��"~
/�"4r�N�(8,�-��)���d���x��N?C:���2�I��{�(	w{v~*^���ʌ����ׯ�������{�}��g������B
O�x�~B3�a߭�]��l���ߤ�Dg+�N�� ��kc�St�9�yͳ3�%h���G�ݯ��	k�
�(d�P��Fq<^�U�:�h�\Gn��u]�S�y{?��֓���%�i!��-AF	�do���陥P��NaiAr��K3�a�6�p��Y���������{����5l��K��bz�7�ˌK�Ս��5c����@Հ�Ln1$�|<ݙ���PL����߼�� �7��G��&���r�/./�Χ�HD.��r��ݫv��������r��d6��;��}�(�����<��U��b��&X�S"�r�,&�����]K��0g.��-��)C�]Pʙ#G�{³:s!�7��F��Ik�L-�f@^���P&9�^�.7���$��fv�4(�E�0�����j�:3�32E2~���m'��V�
���pg�e�ȑ�	�6敦>��PCFX�(��F���n�٢�y3�2��9~�&H�ke��(rE*T<�'_o�,Ir��EFu���`@���(��4QF3� �X��d�Jɕ-ɕ�%�@��03=�=���:�
�_�W6(�6x�^Uef������(�`�S�^�0�C^���JYes�mL���~9=?M?5�R��=EL+��g�0R�F�0��=�zYɒh��d�3��x���8���FV�5G���f�i���/�9/���j�ks�߻B�>���=3�����<�������.,F�ŶӾ q���g�%3�T��N����}'����O	�oU�ې2�bQrj�����f0v��.���r{{Gy��0Xv�F�
=O
�F�6��@s��5��H����]���vyy�X�d����׿��o�b�Ō-���Sqޯ0��Щ+�^ya��d�4{���F��J5r�!$yxV��;�:��
á��J���h��ɲ�0\��o;|L�	��^|,��|��o~+�s����~�*���V�p���`f3m�q�:�AT�y-�3�Bn��c�w5$�5^Q	!�0<b���ӹ)��`��[oQV����:]�Z�a~��_+c7�E+�>|�����t-�{lK(�B"G�\n6��TS2x@�`K	��]��b�t�o�R�X2=�@�ڄ��l��$��rX�s�1�Il����|î����?}���ߏquy��J�����?������;������L�UC8�K�{Y��3_��Y�� �/��= 9r�?���tH|�k$��e�Z.�p����Tઅ6�Q��x�C��b�d�d5���rS������pm�C�*pd���2JK��T���PX&2�*�1��d���}���|�����߰I^,�R�1���D����W��i|�?���>|���-�.Od�W��xss��_��ȋ-]2�����!�]1�<�ssЋN̙q��_�׀���s2�������N�3��B!z���KY�Ơ�L@}�G�:t �Roo���?��O�h���f��?��O�Z���6����/��Ar�d��ҸWLx�8�㕵=�c!:o��{�n�ʒ�[a�����[4�2��k�.p��S��nM��Dt�B�	��w��aI5k���������?�l�s�������,%�\�cm�.��C1�2���"8�ɴy)�9l�����J�b���6	D�+�|{�s�¸�`��:H D�@�FFɢP}cw��4�?t�X�)l�&u/} �<ŉ�p����7nk�$����	��=C��@Uf� l]t��3V�u`��5c�K0���3^�"D�>�z�5@]�2k<�(x}�ǉQ&������)��C��t'�瑧�6�4O�*F>>���;1�X�O\1�%�,��7��猹=*#���e��8�+���F�W)���t#���+�=e=i.&/�8�ʮHؘ�3G}:ᬈ�n5x�	�ՉROkǄ�ґ�I�%:~�ˠ��Ü�>Gc�.L�Z��@�������oYA$�`IVeP��Ny�y�8_U<^�V�Wx�H`�}���ֈ��.FDnI\��?����W����g@��܉��4�[ONA�3gG[?�K�0�������aq���ox����~���O:�+gR����)^r?�|�	Q~T ����'�$�(�{3�;��E ["�0-�����V�P�x�1&��@%M!W���`3��w�������{��{���)�c�'�%�i/OO��2N�+��ádr�DK?y��>�:��Q)Q�:����U?�~K��Z�!�a=;�A\e���+�o�4=��2�u��ƋR���q�aAD�\Cm��}��?�яB��)#嗏?~����F��ތ�ki�/OKy*�*7�7�7D��m�ǐ��_�R�V�a�[3�0ڄ_.�5rPN��6+<Z_���,(��k��=� ������7�R����Q����_��E�P��14ăER�w�0�b͂xrs�I8��L��g��@�l��T�!X7��|�&��o�w�tn/����F�Sڕ�����A�6;9SF���-7�=r��rE�9��V��p�B�63��ZX*_��j�Ε�T"wBk�!��ؼ�\z���w����v�4q�d�)�|�q�s`���?�c���!y�����1X.��dy��6�ת�wCV��l/+F5[/XPDs,d�%���{U�'�g����� �l�����TB�C�L9�CO��t�������a�G���C+��)egT"2Y�� �r@����Vc�xbr��&(��A�W�l��6�L|2����cn�� L�-�q�w�1���Y�nv/(����N�8�2���wm�۷7�Ѭ�SB�GZGu|�V�41Q�cs}}'߼D�o貈��p�n>!V{��\T�ZP���Ẫ�vTW��0������k�7�:Շ�i�;�M���q_�䨉��ȷwħ,��^#.�V�-�3����s�p����l���e�o���5yA�7sK����{�?�3�E<`�N�Y�\(����L����O����GQw�PD��_maH��^�C���N%�����c�Y�ZQA	|�Z��l3��r�d�X�L�Z�9�,�|�T�s��̲���Ч���������?�#�r��<z�D���W��J�N��k���W������$���k/�9G/5�f&�yt�E�y�2��v(v���p̹fէ�L����[�_Iwy�����<�s��2�C?�d�k���?Y�������R��o}���S1u�U��oneR������b,��Gx�9t��X7�|�lv��9�c/�Cմ��m-i������`;M�d�K��X��~��5�vzLʤ�SY<h�����?���7��~�C���^g��z�g����w��)�}>���(Rf�yǍ�5?)1m��&=+&I�8m̵M`���C訉��켍�w��u��b�a���![�A%y�ޜ�N0bD�v?��?��_�/���o�����f�Ž����w���������@{�]�,|yvt
�I����1@Z������Xń��>�G�xO�Ҫd�i+�6���E4����9�I�^����+>�����ǿ��o������_\�����Qg6�7�W�_�����¬�����DDy�b	5�F��8��Z�$Xq/�S�E=*l�1�(�#� ��%���p����gO���x��Q�%�����4�;l����?��������9;�8F�k_{���֯_ݲT�����S$NK &K��\h�v�D����poZU[pj	d��$-j��s���x��W�CP؈ؿ4v3q�~����
���wd�
���޿/I�I�z�ô�򮄳��
�Te^���Kt4d�Zy͢�f�hcU���)C��U莾)�w�M��J���w�G���~�vO����aP&]�N���>d;�7����r�q�������ϟ�Of�]��O��[]�ᔵS��s�JG;$�5E����o�U�&�"'N1r5XL�.*���/@����vq��ě뻯���s��k���>��ë�3�+�N��h��`J��]e�1_�1O�b�Y��rw(�H`SQQ�U=2^�4w��M��`N�&��#�pG���@���G9���]� �3�N���ɐ���)��,����i��/�|�^��C%�fuf
�:�rql���Vxu�j�2���d�G�Ѡ".x��F�Ue� ��6�%|r]�$���p����ĥ'��[�dc�hh��P��Ka9;���Z���#uT�t�8N0�|��f�X"�៥O ���tA�#�(]V��}` �L.9��T9�/�8 1�9V��۵����M�����f�������L%�֕��ykK�
��kd��\n��;��Wҙ�剂j�;�1È{��x-9�a��K���sY{��j�'A> k�<),��l���̾��v���ݐ�Z��@��ZW��W��%nLjrQ)lhOa5z� q�ő�����=�C����M�1�m�p���ḿ>~���)L70�H?���Ż0����{g6g\S�����!�RYz��Fu19�/��/Ø;[��c`�,xa
;�Q���~}�و�g/��uu��B=9ўb�L��g�Iw]��;?V�&m�{�[  ��IDATw�x0�c����W�XB�FE��(2XGT����G��kĝ+�{b����&���-��|���b�
�Db�\F*�<� �O>������?��?���裏>�䓙yA��R�4(-<��J��d�KQ��ܿ���ߗ�Q~��_��H��.�����V�ȍ��8̅���������$(�6�l�Ya�!�$S��Z�K?B	lVj6$*1���z�4PM�%zѽ���Qd\u���Κy7j�ݰ��T>���l�ӥ^�L���FD����괙/;uKh�s�,+r�0�o<�UMv��8���*�����`&d�VH����h9��������7MU�H��7��N��k9��M�Yߜ�����;���U�R�WM�ܦ�$�譹�<תsNO��{��k|ڵ�o[�J���!�S�`����A�,�.,-�F���~!�io�����1<�{`V�:m?[-]�\�"�r�/t�K��S�������迿;�R�B�k�ټĘ��MU�C���%������͡I-s�-pU?��C���1�����y��q��)fy�������
t:��Y���E�9���Πd�V�dZ�7���O�t^�4w�.���^d1O���:N
��@.'�����`�,��m���a�H����g��h<�Ϊ����y(}�8���XQ�ܴF/��Qې2,K���|o��=��%��[�QEX����~�K��;�讆/wi�\@�Cf�����I��A�B� PY0ĉc���zK����9?H�Zwh����%���@�%mIRd�*
�"��`!��Ng�	��)$�4�K�@��L���̫��Y��2b�Z��˝�;ߑ�Ҭ�|����r���M�����2��U�7�ebm%��������\��m܉iv�kM�bl3<��e�\�F�X�4�|��W�-r}������ӧ��ˆIl�ՋW���Ź��j�{�y����O��=��ڬ��K]���n�#��m6;=��˅[�BH{,z3���mWW:���{"���$ ��� ��Q�q���k_{�ӟ���/����Z�\޻������e��ke�l�u ZV~���l���N4d���z���%=*q#��4�t���6aS����>�d�����&�VF�9Vη����?���}��$���>|�~���y��>��U%�zB���Do �_�H��.u/0���h�H�`�K�,Ui�og��m��Q�{�~�`� �}�5�>��"~�����/�����G"{��jrs�' =r�ql��]?f�[�
�b��	}#�Ƹi`��)�э|FC�h�=�y,�>X�O�'��ʀEhd��c�lf��j%��ۿ�[Y�i8t��Eh��F=Y�A���1f�Y=�K���8?*Zs�.K�;�l�bF��\�rE��Y�U��g�,2�R�,u� XC"��V%@���s�Ӿ����ŽjZ���Sr�Z�إ;9T�$Ti�b�uEc��/��:6H7��ƃ�Cz�oC"�f��ħ��m� =
��)��ET�#�!�M��[O�����En��} ҈�mi�-.���(��L��0%u��ppm��}�[A����ў�R��A��q��=�Up�J��O>��`>�,�<d"�q�Qi6���p]��/����_@�!��ǖ��� QCN�p���5��rEV}cEX������r�N��?�iՆ�s�[w�ӗ���C�=M�M]y�8	���>��k.x9���!�:�Ĳ�8�Vv&�1#�;P�Ī�n��aS F��0���q�1YǮC�x��~���0�7b>���=��z���y�Ј���3��RB���3XW���U{4�f���m1���:��!7��z�g��	��SI�4!$�q=]���������C;U/�z�BuA}^A�h�W�:�&3δ��-����҄�<��ad��_Q���f^��=w4�tŮ�d�}���|"�?jWѺt�G�CM�'Ux��T���G���0��d]����y|���h�8�I@�Y)K���:7���%�j�ߋ��~�%�:�B=�^(���g�zm�`L %d�ѭ58+��3<�杋a��8���J_l�Rٳ|,�O�x�7��!����h�1�5�Ke�R�u�Xm++�<���T�ꓦ�s�1cmq�<)���m��;:o�F���ƣU�����1��7�x���<V�Cas�<�\W��NntYOz�T\9���9	%���O�K��������>�W�4z�ΡG�K��L�1�/������2`��>W�A��j�W!���.x
*47�l�s�Q�V��	Z��Q��$��ܱ�T����`JXÏ��7�6Ng{P��<�������Q��x�V���2�IŮ�<�� ������=LO����_ÄR�hԩ�M?�?T�kQ#3�S��k�ԯ1J��ok�k53p��Fg���x(?���tU1d�Ǆ���%K����>��@} � �%0��H�$C~��ɘ��́�P�u�"��>��Tqӏ�Cʕ{A��պ�L���Kϊ��8�h��*����!E?�:y���|�z�B}�5^'˕�s9JL�V��2��Љ�:��-��?�ӟ�����/�)[o�{CnJ��[���x9Z<�d�t���zׅX����~A@��(Q_b����jQS�����ɵ\����ǈ g��k�I",cd3tc8�@,j�X��R�R��.��y��Z"��nC����8TI~@e��7����)5�`����I��*rG��B�HUP�/���h������q�k���`�9�ALI�m��n��ꍞ�8���GYH���}?V"��р\���j�81z n.�NUG����*@��"]�Ff�Ua$�z�*��b������o� ��%H�B
+w�OQ63��u:���IjZ�1�W@3���[��E����jb�+`��Lq0��U��l��L{=t��'�I	Z�)O������)�(<�����T�ף8��T@y�1�/�l8�U��0���2��ޒ;ޒ@�$"�h�����|��<���A�V%��HfQ�����ӏ?�y��������z���U6��\_�-��bq"_$��k,z:��W	�P)�[���׍Čw[vv�L�E,0�c��c����3mZ��4�\*u�"���kf�Y:�V��N��^��_��������9`�K5��$������i���ݻ���� h���b��E��W���a�o{WW�l������u[k�љ�D�?��~�ZT�<�a�LE�z�.���$#}��햣'*����/:ms8�lML5,�}��1=�-
�E#��ٳO���������O�YA�����6���`���[���= �L�˳t�<PU6�y� ��u����R�-���<�� UـՋ~5;|����Q�G��) *�J�����u��~���>}�����jq�w�Q���s�1�	�B��S�_�ĜDn�zP�L�(��(�9���,�t��X=��|����m@K�XtD�+�D��o�.�1X��ڷ{�դ-n��*���ſ|��ONOϵ��Ô��G_�b&��)�I����(��`��+)"- #H�Ѐ��OsjZ�� �R&	�%*xaȴ���l��!���2�J�S͔�U��(�]ާ��T�)j�f�w����DL��.�!`	��x������'� w)��2�����3LQ���7�=Jv��?���F6��������4�*F� ��F�O�1����*%�,�����Vy�%@bٳ4��ڡʘ�9�6�z��r@~-��y�Y@9�Z	.�Kc�[͵k������ZѬ�t<����Zļ2��Qk�����9asY5c{X-��9Kz���={�5習�:9Ѥ�l/gJ�֛��u�����[�o�0,f`<�RV��h9s�IP�w\��U��Z�I%����n��Y�JM�5��y{�OO�X���v+�)DU�;���"�e����q�0���c��8�5����BoU?��0�s�3+�^oD1O�x�>��5c/��gd��:1�E�d�_?�e������|��,�vZ�NE��6��
��u;�^ѭ�F���2b��Jƍc�K��+��3�oE�P�11>PeE�ӑ��&U��)��Vh*Vlp�?,c,j�
���Dy��Q�`�q��ӓ[X�y4v�����a�%,@�3X-�5ɢ5��3df[J�*'Ú��� � o���$W�'��\��aT�d7���yC����ݝ>H�,-��T��S�pH�|�	sqఝ���xf�r6-�	!l�,�ǝ�!��H(H�d��ûX!𧵮7��h8���x{�aq�v* q		d���Q��~[/zT4[�8;e��x��׷w�S�RƘ.�,�����mf+��F�p$o�F �e�7U��T�o��J
�@ W��.�b{؋����~��:�ɞ8�H�/
9;;]�=�� ȟ>��s�u+P(,���%������m$����Q� �dYO����)��ڧ�Lr��pd�Y������e�枟+�6�������P����ۻ����}�[c2	A�,���g�� �m<C�ÆO-�Νay
}j��&dF�g!�0����[���ҩL���/��-��|�=���>��~��?�q	a>�䓯�zE�(�XXW=�lWS�%��V4b�M���ϟ�d�=z�L�96�윮��l��P51X�&�|�a�R�ڠT�v6�*L ���<S�`~-��5Y�^�f>��w6���K��F��j�7�����>�XRh~�+��(S�)��P�����uw��)I�ϕ��ٌ���}�&���O�U�CH~ Ď�4c�+0�jO��e��PեV8R� �y���l)�ZY�������������;�?������e��~tO�3�'ZU����C�$��d�vN^�Iz��"닎(6I�=��+���C[)��z2D���#���"��J���t�����(��E"%�w#�=�v�[�6�;��Ζ���j��V/����B���oʥ�]�?춋�x��>��,��!c���~y}��<�fUEw�G��� ;8���R�[�d�o�P��y�P��K����wg�bT����5<ɼV�YƼ[�����h��s���n��-�	��<��8y��> v]|�<��U��:*i ��٩^��
:L�'��p�u��H�����
�4it"�kl��׋�)�V�!!��H~�����o��/�i�?�,�&�����瞚䷹0
*���k���{k�1[*�E1��K,O2(;/1E5��0=�k҃H�b�󼰤��F�Xp,���A���U#��RA�����K��fl�Q?��]/~M�r5��у�8١Iy����G�d%h��^�h[0N�T�ۅ��j?S�U�T�'g�J�f�%�`9�n�[c%V��m׭/}/��gϞ}�����w�y���4ƹVLׇG�O\�U��ŅX^�����M�&�!�8%~V┾����4+:t�s!gv�-na}�d*�FI���j�8�Gb�xu1-��N8f{f�N]���1��X�};�I�Z�ӆOJ��0����S��P���?��AxE���s�G�2�>Ԑg� o�]v8^�f���'��l\��Xg�֕��x@�mp�J���̥�,y=�E.��џ�k" �ٓ��ĕ}�QjN=��ħ�"��gV���u���р1a�,������%�����M�����>RQA���Z����D�pRF���wN��/.2$'8X�`�N�A��1+M�ɘ¤E�6�dx�NEQ-qO��0:��oÑ$�@�Polv
�dx@1���d.�d^�A�ed�����,.\�1�P���\��L(k��U�$��t-]����b/v�K�A�5�'|�|���ó��� *�$����*�E��x�֢^N ���Ϸ:"?����;�M���8CE��Z�1:���Q���`:W��/fA&�|{��z������LH��ƌ`Θ�H�"��	W�DL���2�HE���ұ�+�qa=f�qC�����6�d/���"���?]�^�|	�{�m���a<��ۦwU=���S��֘����r���������i�{��? ��r�
���6m��3�j��]�	�SNdis��ك�]�za�&tׅ��;�5�w����-Gbb��*2�!S@�@�ؐ�C��C{�ť�C�8f �I�'�T,�)�T�$��D�b�P�QGo�gw�<r@�����k1�r�"�Nߠ���;�|�g2X����F���j�8%�`�C��Occ���!�% (��d���1�W�����TzLӹEu$C�����0�gV �!q�	��Z��\�N_:Y�!N���Ѝ�'�Y���
Ϯ7(h�3g?᷸tO�@9w���xBj ?/���c2�͒��l=w�{�2q�OA+�נcC������C���>��ѓ��H��Fd9N&�0�D�%���~�� u�<�����|�S&�������a���f�"��Jp���rK���I�@�LY�8�}�d4s��m.
�֝�v+㰊F}�4Y�f����gԐd��ءT�CٯW�^a��6�+�cu]��v�2��Q�>�`25 �tO]�	�7`��!����]h7(�����r{�7#�E����b�#�/^$Xس������S��E�q�ܡ�o�/�B�K��="�m��`�<_L3G��T֦P�wXLr�,<#��kc�tƳ�\�cI�-��aa| �^�&:%����_�urv��������r��f)��Z,�� �����7�L�Yq}�J/L�n�4��y]LHZ�;$O�+I��E�*y$A�n1�H������R��Xև�m�t��b��-ކ�h�I9����.&؃=�<c<�#�ѥW��x�,�	(�1Z�I���t0��t�lG<z5�5U��|��"���n��;��t.JOB>����8�H���:pF�������o؇�X��&��������HH	<�f�� ̎ς�Ѕ�LCj{Eei?�`�K,}.��h�y+&��ne��\Oa����"0����V������䨂�����#��l)��hj��^@�ylH����CΗ��`a��]'�kW�%�*!����2�ME*�j�(a �T��X-�Jp�d�u.�V���0Yɕd��0jU���>}�
�R�=�h}���x[/�QM�1s�J��7�3n�����E�D!ʍ�>{��%V���ζN�����GzC"�F1�@���z5&X�����v�!��i�~�:$��
$�c3[-�g�C�b�l���g��Uz��E���BzY�`�w� �U?r�0� �v�φ4�Mp������Ϟ�udJ��ݼ*+w-ˀߨ�iV%�\�0������q*�\�4��Q����A��[7*�Y�b���<&�r~�=X�П�5�o��#���؈�?�#��Ƒ���g�}���+ݪ��OC:�I[�٨��T�Ń2�4kc��_%^c.��m��k:k��Ł�m�H���R߳���q�C�x5��y����7	V3�Y#_P�4f�-ǻ�[�լ�i5	F���=U�:Ե*�� �PREl7}�:�y�6�C�4�����C��B�����H��O�)["�{醁�-;�ݾZ%�*���
>=f���T1U� �n�i�����`dz](}
z�3J�s��^B'��@�v���d����Ab���O��ZA9Ŭp*w����� [���YU02�if���c�HK���~���#������Sn<�ON�q���x�~F�#�gm9����N����c�*+�����<���bNK_N(.�d��d	���x@S�b���܁o�� ���p)So���A��Q'���N!W�)}��a攼Q;I�A�AÀb#
f�+��I��A����~#�V�P��c4n�~�Ʈ�8:��P��� S(�����ŋ+��y� AC���G�!j�L�J6�F��7<���D����C��=U���Ϙ�T*ZF8*�7�߄l8�p�FQz����F��l%�B��m���͢�C�,y���n�*M+b��7rX�<r��}�� O-2�$Q��6�4�,i�L��fWK���l��e�����k�l����n�����{���ӧ{q������|��X4����;/��cs-������Q�k}.�P��`��ֹ�6����7�qH�K��g���~Ȑ�dU�i����/_={)�D�'�H�Nn�g,]���(BSm܇mt����G�A����g.	6E!u�֨��B�ƭv R j����h0q�r�EUa��+ge��Y4�N�pc��P+2S��G��]�Ɩvd���r��I�Ԯ�:����?:B+�$��W��5p@N���5<G�*�a0^��ϖ�����i";UȞR��L��}N
�m#6.��47�#�v=vjъA��`���1|R�4Kc�u��q �a��R*#]a��9J�!�c<b	�b`�vJ:���"7��1����{�,�xVV:��W�L���@�N��s����v�rHΞ�&��|r&Fq��#�gb���; .�^1t	lA��(��//a��8W~���<Q��~������D�Ȫ���*<>l@�&�����������ӧO�/VW����8��2"d�gQ)G��Ut� ���n.�����<=�)������5�����{�����O?��W��Q�VI��Ӳ;�L?�sꙈ�����`R���¯�B�k�Df�m��D���<DQ�N/�kh@��-2�����	E�2��	�G�/a14v�d�zc�����ۛ!�b����*۴�'h(��5$d�&(-�W��	�zt-ř�Hl�Loh�`�K�[IĦ�PO����΃er��C��f�����q2�OZLp3~`5�<�<J����,�ND�]�<ܖ�!���¡���sM_��Y�z|�;)��^nG��f����G���L�Td�vm2'��A��D��"B�-)�	R�qvT�&V�$�Oe�
��A��j���+��_R�zƃ�P%O7�ŎJ��pR�_�Ds��w�[af����혤��y9c���QZ�$�K�M*el9�6^�~�3p�����6ףN���
Aj�Em ���T*��[RS�I��k�N��ia��yN�����zr���k�"�M�p9��)�2���t�U�1�#��I
�>T����f�%KE'��%�m�_S�L�C�F���&K�`�ߠS�2�]�^��y�����'�Jy�y
�5�46\��WʴMy��r���؆l�.�ܬ{�uKfv�:�����q{!���"�2��2�z���)���!���#�DA�J�AtI]҄>9;I�����`��eV�+��C)��hEZ�p�(����0=x8q#+r��l:`�X�ȹ`cs�Ia�IpLs�{~>S���W��e����f
`4qy���Np��}���9Pcf�Sъ�#e�;�����#����%�3`d�i1VG�!l ���f�X�[��
��a�[6�;|��B�����'��zT����ݪ�ע�ϡ���00]ec.{��)��zP'�ژ���N\��gOv��yL$��X+��d��*X�(Nl(�<���9�$�(UU��b"L��/^��v4��ެ9�q�]�Dd<D�N�	���R5�I�#�$C�frO=e����8���y�#��`AԐ;��Mę��WOثÈZ};+b�\,P@[Dn�*@���#�޾��z���v2��~|����˓����K�~���%�����$vvkduqv�%&����=<=9S�5�ToѢ�X�H�t�0��{df3u��NC����>�%[�v3;h����R�M�x��{���8�`5T$v}8�ݬ<�"�@]���j����v��L#\ۉ=�f��-z����/��Zؠ�r�C;*l�&��uQ����>4�{�jXS!`��
�����gU[Z��w�.Nn�hښ����������`����mJ�W[��4��<�
T�$j醒�;��*z��u��`���[�\ܪ0{F�ȦJ�㱣6�F;7��h�q
0k�� "Z�R�eZ}	�`m�N=A���
~����/��\��A9�Ͽ��o}���~���}/j����Z*dc?�G���)?�a9r��=�n�UdyW����`P�VP��o��d���m���u�jO=f�(8��dSG<���E���SX�B~�l�4Lq¼m��|Nn����{���>���-w�ñ�<�[;L&<�q�;��i�&ez6c������2Y�Y���,,Ǘg�<Bv��JƏ��d�O�q�軲�"X�,�[�o�7�2o{��M>G�����h]o!2��g�?U&�('����]������}���p��_F'�[����Nѝ.O��o?�A����؞��ȋ�]������v�?�L��Γ8����r��-�'��އ	L���Ҷ��&]�!7ê߈��#�_l�A�!�=���n1��GΩ|�g�}&?<y�D�̄� 勓�p��	y�}��N���Q�~(����t������?*}a���;�x�8a�g0)��#�
P����Ȧ�k)�d�o f�7 J���0��on��TWWW������z�f�l���e
]m/Ӂ]��*�25� ��aS�tF�3�y�ry�R1L��E������7Uz����{a!�,W�ASBs���_��ײ�|�X��G��H�N��}{��O��f�i�o��>���_vU'+'�cFc秜Sh��|��a����7�T\c4Ǝl�O7�&.�t�|Y�V�G��暼2n�޺��H��ƒQ�@6�0���<��ۡZ��ٕPG���ԍ��,�'�O��y�:fF�*N
<SC_X���%�\�%d���u�8YY�զW�:k�A:�E&α̠�	��n;ʲ�4NE}��B��͝��Ot/��ݨ�v�?	N��rJ!���y	��7bn��~u
��a�/E�[��NTG��+���n��JL��Ī�����P�s1V���z"6W7�xT2���Ty�gR�X�!Z?�ꦔ��Cb�^fMߍ�!�|�'n$�Wɋ��h2/*���..��ƾYLs�
1޺��BK$.S|���bQT����u�I���C5Go��+�j_2����r
vh�G��sF��u;Ԏ��y�`�!<Z��y�s�pTY
�Ū�_"*���Ϩ;����v��ƪ��_(�,��i)'�Z�ٔ�R�Lne�~FtJ*���PY�<P�$�U
}ǂ���w�U�)���Ե�r��v�U��Q��Q��c1�+����-�V"�L8骶���G�-"�����ݵ�k"w[��D8�n���ܞ��hq:Xt�u�C�'�$T6
Ž�ߩ۝z�l��s^�����ء��Ֆ���(Y7���Z�}(R��TSw{wvr*-N�rt6�B��\�3q��(O�[�ɆDK�Ũ���RYc]+!_5�u
�Rf�Q������֘�J��4e��&�I��
��|VͰ��L�[�r4�C�c����tuOkЭ�y���n�9��������
^H�ք���a;(�k �;�;'T,+��B'�u�~���C���� f�E����NvG�H	�;%ϓ��;j{厑=���n����l�2G<t���h{�=��d��ȓ�<�Y�!4e�IIYRm�/�q�Z�Օ(�R���r�a���]2C��Rs�)�;�h �#�?�3N���W��mY(��,�7��m��`V�*+��@l�V�(H��7����t�uP��9�ݺ�צW;�]�T
�=�p�v�z��[YR	WDڵ��|�O����<�\����J2��c>`��<M&�uF���j�R]�vh�w���=8QǢY����y�&g{��G��z���4� �Q!; ��:T�3>�*���(&j*�c�)������< uu���0I3�����D�MA��Bb�]�Y�1��݅z^�T�8T��ʟ6��}��U�h�J'Ո\�:�zUhv[Sy�*\�Bg`���h�h�?�MiH��r�v�f:����;e��l�d���C���X���w�T�����q�����趵(9šD�H�w�r���-�����vE-r�:y��a:J���~Xzj�,�f&�6� ��ʌ�T�0�]��Z�L�?�1ߊ�_�C6U3*
F�v7����(�>�8o.�[����,z�0��o����E�Q#V	��`A�^�rN���l-[v����oVf�=f3t�f/C� ��iHv��dW3ʵ������W�O?����lu;�w����Q���3���K1%�쫌D�2h�m���;|���:����j��d�E�m恈�FD@V�J!���sf¥�K��dg!��_��q��կ`4@�Jt 1��8ظ���]Q�Lu=<!W� <+Q5jX�@b{��R�CD �K�Ԍ���S�[�h�B�(�ha�Ť���OX�a��~�q�=x�z��uem��=z�ONn�y�mf�G\�)yj@]9#"�r.��&�[�Nj=I5�<�Y�&�ъg�j���q&ŀ�����\�$ǘ*�D�� h9���d��(sf�����B�@Y��;��%n�j2��k�z�23'�"��Y�TTal-T�Oؽ�,Ƃ�'�G���gmx����CbFh��,��iȴ3} �pK
��͚�VU�x/77k���&��F��Ě'�(��!mʍGXll1���f���H�4�.��z�/�<Y�T9��=�PK�l@Y��?�δMyN��˗/	�&"�����+�b��:ilU�g���VAy�o��(���ׯ=��%(?a2�2b.%}o	���ܵ����h���i�`=��{.kr���y%��뗯Jp!rl./�3_�_�|}8�W��՛CWG���K4��K���<I�S��(��4�p���B����B%QUd�*@�.s_B�S�|CI���u�a�t�}�eC�S�������7��O�>e�B^�{��&j���ɓO>��E�YDB�L�z�&YA����β�j���#O�����dB�$�hs�{�6�ʥt�y���^L��㤗ֳ9i�n+��ӓ��a�s@��*���M u���cs�i%�9�v}�#�1� �]\(�*�b��{�EP9rw�
��\�����x�����K���� ��x����Ɨ���k[��CȐ��YU{򳣱F�x�}��*�rՓ�# ���.����N�����r�'�y�PJ<��6��h���D�b'S��Q?ԔϷL�HW,h���r��U[mp�� ���E1)���E���s���+mP�h\�1�F.G�}�����y����
��|}{��pv�[�W��!z�F�@\C�'�xאOP*x[U���ZN��g�<MC�YX���e�aļ
J����	�θ��A&S�T�[It�t����gi����A��¤s���ʨF����F#!�5��WG>"�r �3�����р����h�JC�g
�z�('G��G.����4W�a��9p��e��G͘�5��?�'t	��f���A��4���N�E|@ϣ\v<9����UO}J�hl��d����Fi:ɨ��8� ��k���z2�Zڒ8#$k��F����=��?W�mL��%��]ι�+X)���ŕ7�z�*X��7< �ĸb@W���0:�\��Y0�˷)f'���(��Q9�1����
e}�~t�� �k�+qw�x@M��K�"ڋ	Q8�0z{�,�����v� H�0���\�\��e����|��r]m(�Ҋu�Tx��~fS�Q���*OV�t���t�+���:��P�|�:.�#q4�������[4�+ݩ!�ۨ=��3�X�6���İS�Yh�M�N��h*��C~\����:����,����U�e9L?�s�ĀG9�z��թ�"�d�8j�=˝7�r�P|Uΰ(�Ȣ��PVq&���Y��nS���[��9k`q�.���V�[��` K��(wuP�n�5kjN�:V��t0����j�ܐ�Ⱦs��D&^�q	����r�ք�<eػ�`��o{�8\ _�V�8��$��ͺ���5���!(Q��̋7fxh���ڋ�K�r�0�q�9���g��&�����fF��Ρ�����L.i�X��V�_�U�U�g���0��%x�ܹS!�R�9�H�9$v��A���/����ڏF��\v}~}}-!�r19��;\T��&OTk{�KZ�W8C��l�S ��:GOP������,B���e��D��)��ce�~�S�ڞ��̎�L���$������N~s�k,Q�R��k�B�1m��T��D\z�'����3�L&���e��9������HD	�%����#�CK 5�3�~Bb�R�
#i�
0��c�e��H�II!ۚ`����A��t��ruγ��3�n(&���f�1���ƥE�Be=Ը��F
c��n=�"�H<���殔T��g�vN&f��,�b����@\.�d�:��]��JEf/r�4�j$4,g7}��0�R#��D'��F���dkb��Zh�3�[�v���bY3�v����1��mI�1Q��0��it����Vso�~a�/d" 5�]��A�7��$> �Ft��&7�S�����ƪ'�n��#휁�������_a��`ȗd�4:~i�p@+��o���ܓV�Z�9�K�b��3��g���A7��������WW�h��U�ب�<����$zRc�����
ð�̐��Q�A�cGo�5:ܰ
��Y���+�ͽ��S��������:��x뭷d7����p��-��i���=_~�%������?G�ٳgLM�~ ץ/��\�0IrY����2,�p��"�PE8�q�U���k	�u��-+�8<�F`x|'u>����D+�;onn���/	��š���������O.��3>�����߽x���*�>��q��	��C�U�=r5�:E�+�(�Q�'˸��	��������g��P-���&j:�-;~��=���G�g�/L�C�﷿��SW���.ZI��OLw :�}�/w��~�QM���A��8����\CX�j��r�lRY䒧�1��>We���܇Iְ�y����` _?]Y=���[͆��&-��t�	,~ǋ2)N���:{�j���ѣG'�9�ę�O-]׹�E���YK��`E���Ki2r gZ-#6Z��G�"��S5M�������,�l���7�֝��o��fn}�h>�E=_7�1F��G6�2�1;0�?��g��VK�dΘ1^9Si�U��ެoq"O�En3�k��<P�輾�N*��(>����q��L�m�P�j�_a�Aӓa)�],s��H�����	*��K֮ƀ����?l7��2"�@��}Z�B��UL:4-FB�r����U�%��@��G�.��YQ�
J�c
�����d���jь-���S]�x//Lˡ�q+�e����H_D��y��¢��>[t��7��@�u�dAڈ&P�};q<_-�5pAg�7�k��Q+�o���`���(\y��E���@P��pK���Dk+E>�)]���r3��3�P_�RQA*�}�@��(k�D�Rݠ~ �Nyr�`h�.m7�p���0pG��ST��b4��Ʃ�~՟���`MgٿtX�dp=�ƥɟ��Ҵ�hu]wd;p�sL1�v��m^��'���5���F) s��"��g���]�qҙr��������ﷇ5ȉ1	ND���ß��]�v"�����I"Xc�-�K"�_��A4cT�L�2#Jc��y�y�7��"[�~Ҏ-���^L��Z����	P%Fx3'{�Z����t�Z�ꗧ�W$	ܸoV"N�l���ON��Z�za��50tiBѭ���F����Ch=b����S��Q%���/+��r��uy�:T�Uy�:���[o�VNv�v��zݮ�`�+���lz�X6E췻����{�ü���8����̔�j�L֭ɪ�j�؀8f0��+FR��g���Lmш�Q��q�,�*"h*�>Y�����j!Z9	�S��q(J|TͦS�T9j������O�߮1%�[��Gxg�'-3V���uE��$�S��bVm���V�1��5�����F r� �!�����^��6��1d��l�FQp=Je�`�0H��AG��B���˲���f���ՂM���$�l�*S<%��G4N�i,]X=f3�<8�����OSu��N�Z�Dq�$��ނL]��(R��aF�J�Ra���k�e�gG�J�i���;>�_�s���$�1��}���'+����-����u4�(��K�t(WoR�+H�8�%���y�UR��L�~����e �T��|~~v�Xj��Y��_T���cOw`nkd�r�Xx��;��Փ��Cbֆ�H�#��X��篕�c��T�����
Y5s)�<��l	�v��;�T�[]��r��l��.���bO�O�U�r�u*����ל鮐���W����mn7�dO������ȰG��N��#O1ۮrg0��`ï<{��B��zYi��]t���R��/<���殸��I�J%Z\4y��`�=]�ѥ�)h%�eV���P����O� $�C]�CG���r2T�>yr���ކ1kK���y%�����rT�6xZ*��5b xd��Tb����x��W ��N���d����d�S�f��P]������ �P�6���hё��0��l�o��O=��-������<|M�)�/�ml���<N������NU���`���$���N`�Y9��<��GV��y?��uU����ڈ���eY��~�2AԙQ�����9{x������֓���ˋ��Ԋܥ�Xԃy~!7�Q�-{N ��֣ʧc��wE�Z�!�Z:Up1K��t�2�z�u���r�-��}H���+����1�3	t���'O�?x��tU3�zo���Yk��W�.��U̪@b�?�\+�e��???y������ɹ���������_l6"��qm��D�.V�{��Ǝ?j��˪=|��ѣG4�\�Κ7KL_�GBɑ��{�E�������sVq�X�_�F���d�m0@�\�H����wd�2�S���o-�^�����z��b!��9�h`O��N��n����6х�DV�����L��GO��O�D���>����������_^���mn=��%���q�y����kp�I$��O�K�{Ƭʕq��X�T�+py����������S�A�n�o_�|����
��|��5��EDD	G���p����"`���	���<�XN����4�	��Ti�A�tڎ�̈́)c�i����}�L�����3T��R�Ӌ}��q3*{H=0��J��ggy���h�;$�p]��)@ԧj���׫@F�GF�ژyD���xxO��DٻEf��nGc�#��x}*�0��o暃}=p��mp��`��ڜ[��R)P�F�''5,En4�3����W����.�[��(ݢ�
S�`����Ȅ�&�$@���;6��c2'�\*��P��	Au/;�)��\�|�,��)%�^DKd���<��N</ɘ�õ�ۗ�
`��TҠWy���Li��r1����nv�+1򙓓3V�Eא���1|�觥=�ל�����Ca0�Xf��H���L�h.#���O�J<�2��c�b�-�JK2\7�_��s�5��Y��1Oɘ�r�V��!Y�#�	o�.�'��ee#��&h�2f��~�5%XB�~�빒���m���+�0��}�7�/�Ӗ��!M��~�7A�N(G�@yr5�[�3�pN���G-�|�Ȥ[i�_g�'I�dw��E{����J0l�DaR�q����9�w�o��'mPA�\�ЫW�d7Y�)�]���n��ѭ�6�R9��[Pt���S��Dfy)n����J�`dT�£����u �N��k��+�bO�����x�G�Puj
�ʌ�W1ü��0N�utHz����,k�h��Pb�x2 ��6.gǪH��.h�� >f����i��[���.��P�vY�l�#�c��8Au��Q�D]��"�0t�,qR��E0���kɁ�����
�C�P��Γ� sr�����*�^7�@��|	�)�������k_�ړ����J#�MЄXGꢝ��@t���_�����)f|πt9�i�����Ć}n��}�<v�yا�:I�;`�x5�,L�B1�дĉ��%��/Z�6vOԳ��N��["�R���D�?��v=��SO}�����K�)�G��3^��Jf�u�Ř�@�$�̙����r>ϼ��m�M��QI6���g�S��֒��-~��������ɣ��@_�nA,&�X��5qR^�)�����	D����O�|�tʯ��pg��1\jnJ�����cƖ�bı��S��Y؜g�|�i������A݅8W���#��企Շ�r}�	�4�(�q|�|w���٬q��2��p�$jP�Z��vZ�@���I]����� YIg�]W�Ǐ�ov�y�]����.�N�����������ߐ�PQdլ 'GGɑE-�:Jh?�tjY(�T4�0a��»�O���5�?�'s�Txb�0�8�M�q��%��\�V�h��\Q{�/_�x���;Otb�~+Ҳӄr6���=��v~�PW���jw����Z�Lש0Zn���'W�/P�0^�}^� u3�7(�f6�Ky�8܌<��%	�a�#A��@ϟ���jw��w��E�$�\4��_l�ҹWT`0l�l��r��L����"����]e�b'��%q�t-XxӮ��������Tq�]3��;&��dE������z� %�p�E��}eϰ��; ٫�姫Q�\�#��b�Y�n���*�+����ZR<m4��3��,]�6�v��Q�@("j���m�h<��5WL8�;w3]�qa��º%<���KɓĲ����A��(|v�BI�qO��=��蚉�9>�&i�=G\��*S�`�}Z�jl�������]���An��=fSs�c�-�<V�ݷ��~��4_pg9C�έ��%ֽnOPҍ���?EO�_��n�᮱�@����LX���h,E8U|���6?��S���=��������K@'o����;�<}��W~�����ٳg���܃�F�O���K���k�Z�n�������o�m����~뭷j�� +��?�������������/��/?����>��S�)��_�|��n�:6�ѱ�:��}���Xi�8\��[z��4T���|��w幾����q�)��j����{h�7ك&���6�G�at�����G*���g�	�6s��w�=��;�cod�r��w�_W�SL[g(Z�Y;�sĘ7�)�/��/>����������|��o�����vopo�O��h"���q�'C��in��PL�T<G�)�;���W�+1�"��?I p|��9�r�r
�N���d&Z���O��1U���t�ʈ�x�`l<�� ��z���1�3�c��蒆�2�:�ƨ�z��2w���\򏃵�D��d4!;�ʬT1���8|7ب�d�f�ԟ�L4%�N�{��I d��=_�&9e����`��@N�����\m(3�^�6F��D�@�b"ꜻ�5N��}&�=��_ap��h�
��<h3��E$�U��Q��^�(j����0����ǟ��`�5 22�)���=��ʈP�E.,q����D�xg[�mx�����;f�v�P]���#Ϲ��؎ao�+]si9�]�M��-��[�4���q���(��jcT�~CN�f6��_�����:0w,7*pZ�f$��yC���\�ʋ-z
k��T�8�þ��p2B�b��&��)�c�1�72�*N�(���S(:@�Z��8$E��!Ľ둅����Ȏ�>m��%���(��ε}��q�_�i�W��"X���=Td4DY)��y���� ��*w^X�4YMp�c�T�]趚�
,�6��pa �om��j������Rc�Sb[u�
�ܛ<��X���1jݚS~�L#P�}��V
	��?�G>���!auC��4L�bvl%�d�-l:mV�2�f4��Jx�CהM@�x;�rm���S"j�}Z���#!O��8%@ı�K�4zV{�[�J�t���C_�A� AN�����&ǧ�b/��6��ɷԚ���[�U�Z�9+��9"?�����n1�@4���-���NjLn�;���XVw�7{�NN��E�X]^�Df��[�ɓf0�sQ���y�I8<�R�D���B��^�̮�43�L�}��'Ke>�P%��W�;ѥ����.i�Kހ���lz���*_.a-��qu�u�ڱ.�a��U���o?Yp蛒����9��������46�b^��R<�f�_���Jo)�j�B<�b��]u�\�ETD���˂����I6�Yn�����TYK��nĀ��QA?��������]�99�����&�M�������"V�œ:p�n�c6Bbt��\4�������U�oֻ����Ë�Z�o5���n���B	�gKys�0M{���r�x+�⃋�����z�ųg�a?hN_N�"�g����X�}!Ϲ:[����=x�Q��x9r���V�U�t�\�.�bq/^�݄!�JVM�h��v"��{Kemk�#R�� ����+Y��� �_�Z�߼YHl���l�j�t��f:�5�}�v�����|1f<��J'�'9��n6wr4��?1��e�W/_>ߥ}��P�d3Ȇ\�U�ĶM=k����>9=���.j� �n���U�)�J��v��8�W
��s��kM9���E�N1�u��{P�޻|[�z{�������;9??���]�?���;@M�S ��FM�0��Tv�>	7��mꙆsW׻"n��E��>�3P��=:]��F3�7���bU����V�z� �U��jՎr.x���٭^��%��~q���`n�H�~۝č���I�h����!ry��S	&8��������Д
���dt3`�i��:��﮻]5�ꓫy%�(>|tO��p�z���ԫz�����V,�r\`gdgS�ճ���ͼ���j�%\yO-�?[+�å��m�U ���5����_�:�P���r���B����_�~���j�5+c/��Z�^��fl�z��l~ڈI�t�޾���E֗+5�E'Ơ[����%)_�z-�S|�b?dN.@<�@�C؇~��%c�����v2o�s��DE�''� ��77w�<�l3%H���&	�U{�.�H\>$M�+�è-l���g�(���Y*֡�ǝ�?�cjw�O��Jv�l^�ٝaZ��&���)�#���ܛ�n	�7�C"~h�h�pzzr�8��|~=[~����ry�:ɓ
4>����Ӈ���z�v{$;�!�
���A���ȼ'�3:��)�����ĖvU�CG�&#S@"c{Y�1w��*�ڍ������]�%�)�J�s��d&��'15[��E�g˹�aǲ�'+Qܯ^]�$$$�f�P��k�7���r0������b�a	M�R�H٠>u{#�)Fe$����NWUL�Lӗ�����p�?���Pc�x���P�u�G�W���O_}"�e��mv����#�G���`~�,*�J� �C����\��<�H�g����K�.d!�j�c�`�<��'��86Ԫ5�j�P��i2.�S����[��&�{-�̙�(����r˹�N�k�b�~�ݜ].�LD��u�L��b�����Ӑ@��+��@OP#�������?��[u�Z�w`��*��NU�>�"OF%?��bi���ɀ�9�L���Z�gcū���X���?��y���d׉>?�Xy�^+bh�@�ly"N��ݍ��Љ���;�z\�E�������O�>]-O��F��u��������/�gyϗ_~)����~�;����Ǐ���~����_����Ç�-ҝ��Ou~�r���ޭ���~���|��R�I�^�xނG�/Y��dIr]	z�x2_�̪j4���F�������5��|X��`k�K���n�*�����{�=1�miY��"<\\y-�2���.�OgON���������љ�z����777eY����tt=��5�M��o�㢻E��b���?`>���+3	�\���nZ�q�_�eCɓ$��K� ��{�2���7S���/o�w��DP�L.�)1tmdb����5D�!�/"<���]� օ�F����D�����Їɶj�@�ǨW�����j;;<�&h�&2�6����/��/�n���8�/������ˈ��z1��ӓ������e8)u��ڽN�>2�(��C����J�@�ݩj�s�c�w��Sm-[U���d�'�'2ye��F�/���}�������[���VNz�g����pq���v���_��W�_�����Q����i0���?�h|>�8
H�*��&#28���ʐ9K~�d��K�u2�(n��[3�g�(�ƶ-2�A���Y��=�O6�^v-^����!^j0k�I6#��Q;۲����z��t7���H�8]�%�����X���,ڦe%�L>� ��EH2�,�(k�Ӊ]�m�x�$J̨���1���m��!Wzʨ�[M�i#��߽{�)v�pׯ�v�Њ= �A�@d�$z�U�s%�v�gt�Ā�$j��܈�Ρ�AiiEV�u'[~cq��m1�v6JK5Z�V�Wm�x�(=<�	j8M=8>S�K�Қ���A�_�AЬVO&\�v�*���R�"ժr�H���j��֦��jզP0�P�J�"�!��� ��X����_~�;
h���*bo�Je���XU�ݍ�i܋ج��L��N��r�<��}2�N��XR�j���ׯo�֚{DR.p��^s�<B��h�O<��a�8M2�ک�����B皊&�B�j�(v2�Z1�4��áA�k��Խ#�\�O��t�:�U�ߟ���qO�S���T�~)Ao�1�8�ǡ���F?I��P9v��4�Ŝy�:���w Z�p�:T��1�ڜ��8�c0ؤ3��%���7�����@K*�a�Z�o��hHL�`����-h8m�<���`����8-��.J��j�}���UmUK�*t�b�H��m,���C�����by&}J�v���Y2N���\}1���i�:3x�C=Į������ٙ|v�+�pY�)�
/xp��9O��/>e��	�A�m1�a3�r˛ ���10m9M�J��P9"��S؋���,��
]ij���5#΃�#�w�_㊃0�)
��	̦�Pyq���b=q;d�d��hf���w�oe�9*g��y~��O���%���ܖ�K�Y(�q:��#���_��^ƀ3�6�LƿV3�u
dH��;58���g�&���� [M'mAS��j[��&�$�,9&\���V�����̘,7	�N�I88���G���.����H���y��d��ɻ+v��z�O)�ο�xD�|�_`�H4g�c��ј�J�C�����][sľkT8�G�,��i��̵n���;`(q�4)�4���5-\�#Gj���FU�޽{H"l31��멸�XU�8�.����f��V���7�c�e��������C��o2]2����4D��ݻ^N�/��esg�}-�+
"���R&��P˔�ǂz恵�X�0��An\G)��/���Z �?{~%Û.N46G��^L(�BumA�V#��BV5�[u�xe]_�{y�G�ư�:���1�:6�?�~ɘ?�	��p���<d�E�,��HcV�`�d���jD@���K)����.�Oa��)����{,S���F~/�������3����bv5$�vU(W4u��Ī���X=�t��fp�����?��H��8�3�3?:�y[���#􌂷�
�Q����݉����W�~[�ח��g�qb��>Ϫ'�gm,��jG����9��>��`��y�gV���%�L���j�x�z�R(�0
콺�S��f�Ҩu-���e�����I�ʖ��~��n�ց.��l�J�Cש��7ڞ*�MQ�+*t�<��� �px">�������E7�W&�S�pl���AΧ��zC��E�ƞE5�C-����7�7�x��m����9|�=ݸ�L.�VS�0/��\a�0��^5S�Z|�vS�&��F�c@�
���{��h���]�#+�~C6����Q������W��!��c�����7@-�Gb5�v����C��z�@?�]:.3�FPjO2 ѻ&��#4<�g��I\+������X$�o}�M=���w�����ǣ,v�D��$kQz���l6Q�ʖp<¬ :sb�\^�l�i��ٓ�������ջ�7��������>@(Bk�$�?��@��?��?�c�!����/��/����~�۟���v��,�A��%�6\^��`.��|�իW�
���=54'�����o���\Wl)5�H�S&���@㺸��`G�M�1�L��T��BW��	g�	���'���d��FB��(aF�{�4-P>MONNF�)�_��f��qױ�DV�͛72���k�4QO��^��]���c���0|���h�d��]��=��ËJֽ=�@x�׋/YA�ԹF,	������v�H<��L;����� Վ��"xkd��uAddw��?���d��7��I��'z���s�r؜*t�	�aʹY��KT���1G�MYވף� ��|vS`�c��AB��zvr����ͽ|�����?æ� ����+9)����!�w���B�^���-����v'fCۆ��^�$�����S��?�8�8
%B�'��v�_9:��'�B����k�"�Kn>�����ZE}�ʹ{���|J�^3������n���,B�փ{DVx$ ���6���X��H��t>��C��'F�f�W��o[���9
H����^6[�a�VA��[�;#D�gj< �'��	`�a;� �E�u0�]{^�����;Cp$&��h4j&��[�l��	0F�{��S�)�m1�F��x>O�n]���.�*0�n[�,sx4��4��Fv�nE�-��E��ޤִI��a�,rꖢ6MbP����մ셣,��f`���Z�����<6*��Ua�89Jo`�`lZd#כ$�Wdz�e����p��h�z�,A4��sCW�m�l��a�]��@:�G�JF2q��	I���~ V/ІO=�ӕ;Q�9wʋ�\�H�h[k����Vd���G��[hA���_�?q�����r��se&"Ɖ��_��H���bǀ��Ł҆z=��cK�X�\��@Y�8:�������G�q �T��=%����2�!{�UH(�g����o:T�R��/��*��-�ѢR�&D�hΰ!����-���.�j
\�u���n\���
A�޷�b�G�����'�(K�Hrn@��}�����@߃�S�iy:R�7��0���qUl�l�`nJM�g��`�:�N��+��Hﻻ�9-v�j��w�ny���u���iW��(+n��ҹ+Km�$kj���d�DdmU*nX:����;$�)Rj�M��yr�r���A%{=����p�d��ؖ�ý�˪�)��aW�b�棑c��Lb*t�3EMB'�ì�Q�3
r�s�=b`c�Je��j*���m����`�h�������4A�l�p�	�(�'�����N//��L��Dƺ�j1=4
#V�݋7�ӈ�b.����*đ��r��°�ĦA�h<�ja~��az�&]U9�/������3���E��Z[j���������l�,�����
O�����|n�A��ۿ�h`ݮ����B�ה�%2���1!r���׃��]*�'�_��,R	:N�����J��=]��5re��F���Ο#����l��z��0�,O���q[ד�B����rS�LOж���k�	�0�+7r&�b���������dcT���i"�i���~-���CWk��@��l����E��C����ֆ�""b�S+'B�u�Y^�Dl��%��g�l�)Od�L��	�P����`q$�b��dc��f}���@	�h�({�>�a��t="�R��0N�QԷ��N��U�K"��c���i��U�o)M�5I���F��^7*��{Ō�V���okqGE��Iط�:o�5Y�q�������`~��i��wa6��޼z+�#ƵB��W@:��6��rv�	��q<�����'��Nb���rg�,������Ю���H����l�r¡��i�	��k�F�zX�W�7���lqP��ru�)'�����Ξ<9>��
�z�h.\i�B][��r�l�f��64��]��j�o����~(�+Ϣc6�31��/uм���V�/���k%C�H]ڐ1�J����~a|0ҤD�be���|���e�_�O�S����&��>,��n�Ap����|�}�m�X��*}ԉ�
����
u-����x�d<��ѧJ�����kW�=�����ױ�{N����uV�N�lT��9 �>�D���"K��QJ_�A^��#t��<��	Z���7�q�.��c��A��ʝiz�ZzLt�,�-�$��q#�c��\���������0e��'�S�fZ9d������z��WN��(�����e�q\cf��$%�{��h��U�����$WL5���6�X�>�zT?�CZf��A�s�}�&~���y%�������e-��Ea.�a��ߪ�p+b��n���ю�}w�Z�EIOR�p2!�(�����b��ct��'D�"����H���'�]�P	�k������dQ��"oqtz�܉F�"ʜ^]^��:�^d�1N�49���7�q9�y��<���>�����X,>����?�����������g��-a��=ˢ���ͫWb_\>&wUNW���LVJ����� "��˗��D�, u�?jp�8�*`t��g�VL �	�~�����qe��ژ�:#AL}ٝ�ȅ�]U
��z���zI����5�����w���/j"�h�1k+�P��q.֯_����}��믿����r�2|�G�[��~�">t��B׸�W5�u��A�A;�w������Q���8W0���,=��ُ����ټ����Ty������J����w䱹���Y�QaONNb�ٷ|ɜ��%Ճ+��l���(W�g@1�>��B�� �H%v|��v����h���a�B;D�g�F�P��]vZ++�ݻY�����2�r�Z���;�=��b��(����K���9����^b�Y~#��~���|�9�N��*��Q`G���cH��Tf׺q�]q`w���qǣ�Ym65�X]`G�^r�nFb��ǩr�s�v��ݯ��^_�H������x&�><��4��L�p���lw<�-t,��"��E�È�]L�m��yo:�a�A�k$&�3p�]UOC����[��H��MMf3���*4؀a��z�CCJF��6�=Z�w����(\o�
'4A�����x7���@|��j.2qJ��D�[$��P;pj��/��\0� �+Q���9QM%�3�+���v�/}��Ry��3kI����/~!n����	X�6���S�o�U��mUy���e1p1{�|,�q��^5���Gۢs���Q�zS��O�h 
5u�+o�6��,p$�	�58�?o�<.�ԇ�Ǥ�x�O:�.�ŀQ��h}�����= ��S�Rل��e#����:Cެ�+x�է.��i��e{G o� �;(�½�y�j�=f�R����986����}}p�eN�gj�x	Q�zȚ\�ā�ׯZ�XՈwk�~�Q����kc�yH¸��Ty!b�.r�#gV��F��D�'�iKզ�����Z�������'C�8;��ܚ����3[�L�d��\/Bj#*��)=���Ԝ�����p���lv�N  �m�F�!����N}�H�Z7�&��m���5y���n����_�1�J�(%Km��ǹVkpٖ[b�0���Jc%
�*w*:��y:�E䑵���9+s�[*4I�ۙO �.A��k�E2�����ggg��d&S�s|||qqqp|ⓟ�ֹ�&!�1)c��ԊJ�����͍����y�bi:8��`,��2J�
�L�*���X�w�cEr��.(EEo�]�N[>�v���ծ��S�~��@X�;�3�'f��k<Z�g���,!�nu������zx����R"S�|L�������:�5M����1wgEGeAR��wp��1IE��3�y�s]V����PزӜ̔���4�Psz||yy9Q0QQ[���N��6[�_Y2��qÈ��;�t�WnĲ:`6�0R�K;�(�*3�ή1E���݃|&�:T���@��[����i��xU)�4��XΑ�JNE"uS����n�-Q5�v������h0�ơ�G��r/e* UF3�;T�6if;ey��C6��@�j:�FTYX���x�(B��n.{\����:62���h��Z�Ԁ2��qo޼Vq<�>B]\u{��@q(]`"ֶW��r򳙶΀Ί�Un���;r<�r�z��kZx�5�$���]�q�zԌl2Ы�`{��� ``�OhUʎ�N5fF 7m͔�V��}�
�h�@�HP�=fT�<h(��N;����W]!�V8�T0��_�D�l�����H<����Uc�Ǐ�w��R(1"`�y8;�^4�@�ӽ18��I�5��������>�EaB��&P�C��0���FW�d��)�'О�;�F˻�e奫�8�dխ��ۃ��x%k,�x:ȉ�Et��;(���'�,�!*=���ȭ����G傽s�C��1�;�!<����>�M&=���[/��|���_�����o� ��VTvpUɴ6�F���#��}�/��`d*��e��K����F�0��7�󫵄F�z�5P���}	أL�=����=DBx�?r���C���
t�Y�ã5�1��ϥmy�O�4>��'?�I�V
����'''%����A�������1�Ϥf�<7cg��j��F,�9"K��5��6��ܩD<10��ǉ���P�T(��GDmu�ż������Cm\����l��.����O((��+x7�_|!���(t��5r����Ȣ]��^�|)��w�Lc�o��2�S�	���t�Dp�ɣ�����*�_IK�R���;�2�ڱ@n�r�r8׮�U�w�C�%�Q��b�ި���5álI�a����=z��2Ҧ������^Z��|V�z�p�����G���R��!@��#_3I1�dq��2�;V�?��{�k��;/I&?�r1����gȶas�ׯ^1**�CD&�����%���pNϙ;�xY,��������~zz��w�9urgn��S}�п79x�X� ���`v)=d[c4��6�|�2���as*}��R���	���|!w�Fcy�,����j��|<�yX���D��g��62�
h��1Q�+��(u�;����i�d��ӄ湋]d �'אk���N�i��$�I~���<��������I�>�J�ZkE�+]�c���� ����b�'t�o�\�ip
~K{Y+o��S�J���N����f/�E��/�K������U!3� ���L�Put`�ooo���Q�֣q���ao��ŋ�(�����c�A�7�,��5b�!�;�i����6�W��d��Y,J
�L{zz�՗/:�-�w�a��|,��J���F$����j�1>ղ&M�A�n�[$�{0���E��^G��w�h��*8cMOޥ8JmL�&c�����$�=:�B�����1mY�L��Y�t��q[��-B;0��Y�O�.@+ZK�%������%"F� U���T�&��2�,�&-�A�::"Ù5���7-����v��yw����y�ۢv׆V��y��f���t��L�P1�|���L����mks�S��-�8����~Ul��<$�PfT���`j��SM��?��J���Z���Ƶ!�ܧ�C�*O��#���H�@&-�l��d�j�8 W������h_d%D��=0��"��(<�U7?����fu;����n�I[��K��dDPk^y��~7�nj]�I���F,�������d�� `��
��H!� ~��NE�#�K�ӥ�F�.��z���(Hc�@a^j��]�IA��F�<%��x:�M�5i.�w��4�gA��] ?-ʓ �5��2u���_"#&���/�ѓ�g�Q0��-�4��!��?Ȯ�h;�p�J�/@���8"�&vJQ�f�	z�jV1��Zhd2��,(�CQ� �
�]�稵�K��K"�߹�����'W�	�q
N�V3�ww���z������ ���S�T����_i$7�6���D�NՉ�+�I<�A&0�I,ҬN�v<��V�u�.ʭ:���[Y�T�yZ���ڛ!Ev�U��������ϟ���4�,�Vw��|�ve�n�r�Gǧ���Ѷ���i�����ny�ڬV���Z�h�C2��{��p��;�?�-^(�wf۴��<��3�G6�	[9�b�IW��o���{� ���lܤ��,;�r�޶�5mbF����l��$F��Xb-D�4�����2������VC�h�����2s����|�v��hO��A �99���q�/��! �ȎC�g0�e��C1(+��
2�{)D�/D�rPPg��ߠ���'$��bĄO�g����*p��9���tv(m�jU=�ª�A��a��{x��ѴZ�_�~u�����L���VOO��h���"sGm�m��ץ]�l�C�5S�U����Y1���H}�YѢ�k�s��ŰBѧQ0���:�9���Q(���|!��E�=<�Ďy���|��7w��`7���Nv�zS<{���jٻ��I��A��U}w��k ����l�$�0�l[� �#3�b�N��7�Ї�P�M�j�#V!�0�Q N�X㫫�<O�˔�!��}o5�'Rn4>�dn�V9�v����v'�R�y�q��]KK���o���a(��Pu�(Hʦ�UE���"�����0������7�3���� �#A���i-p�}Ƨ�j��f��&3�r�Y�r��g�`���������@�`���d��x԰4$zW�[;�Ѥ!�X?���򅃣��]�N�n1A������k����u�`��q-*H�nP�z�z1B�P�^�:��}�ц�\3��}q��%��{=:����1�z
:�"��ǆ��J[���v�)�c�*����V���.qE�_��骭�[%��Mc�>
:���К߭#���8>Z�>���Y����q�"�6Ǩ�j_˞(k��r[�E��E�P�!�E�I�s�G�ރ��wh�n�(Γ4SG�A�pͲ8,I��m��xXt�u��f��U	��1Jbo�z'ſ&�B�-�sDa8g�c���AT&���i6���o����m�;� ��U�;T�sovr�ٓ��~���l*�(F�bp�R�l����kV�/��yǯ�q@J����*L2�eJ�1R�I��}`�m��+s����D�U�#4��Q�_���M��5�IlZ4;ϒ��Tu���������FQ`�J���)�x����;�����ٙ�헿���@�����dھ(��TY��u���	!���v���a�	'�Q�ē�@�OHe�k
z=�,�%l�|j4Q�����!~(��B&�k���^�F���!�D�x��i�q20�� ���a2�.��E��k����S�nB�u��h�o��4�Cwip�Z>�/�|x,��9(�H� V�7z�N�#H!qL���Z.���ȃ&?���m��oo�!=4w���><Z,��[T�'�|�СlY&�A���#�3�1�MH���]��S���~�4��/tH)�53g����1C��cK#����=�T3b�s���F���~%���ceM@%���N��AI�d�w7������勗��>\�U����7���ʣ��/�Y^���sS���d��m��2~����-i��ɒ�If�4��o���$ɵ+�Q����D� l]Y�0�_��a"�*�u7D����N������C'���)'D@��cpТi�lN��E^�y�_V����&�#��-��q@���%�&��J���qn�vu�
�w	-�2���BX��+bZQ���1��Qg�3/NO���hq �����}��[e�s���h�h�lu6FW���,��[�6�G'��iT>h®-o�N���a2�|!��
�ѕM��܄�R�y>�裏�f`�Oş�|g�P[�"� čw�c��^{94cy��� �9b��}�H"�ƥ[����/��3�����o8B�ȱ�{�+tmy�	���{Q@xQ�U�oԂ�}�P[ơ#򆣏O1x�1S��=��vb"z��dʬ��T�O�q�Q�vm�����#\�"�;hU� �s�X��Oӏ��W����*�n��Wj�b�3o�{�8Ng��� ���q��}��ʍ���~���\���M��'�榸�:���sM�e[�D+,Ȫ�8�X�=f�Z�5&��;�ݭ�2m5��k��ȡ�ߣTS��PkpM�i.���a� =E��b#�{2SM@\r����Q���B��"����t�t~xӊ�B��X���ZHR)�)?Ui�'�4�ʘ�|���\%d!�ecIp"�Ԗ��ऀw��r��42j����P�C�%J�1�g|Z����T�c��;�A�vz���aN�W�E��b�F�ċA���Oi
�yA!-0MKQ���I�־!�����p~��X����1,�ٞ��9� ��G �SO��DH��>�:O�5H|"����P�����3y�ۛ�\V�&����\YP9Nk
�hx{�&9dK�&�ޔ���s��;�#`$'F�a�e�m�D!1>��X�6��9�g�1���;Ş��zza���^�e��r�!+Thm��%�
B�QfN&��Y�h���c<@z��gI��/X����"�u�+�:Õj�5*���ri"��' Sb�{k�f��x��٦��h�D`r�����Du��7(��z�w D@�Qx,���!(�d���+�ö6�@U9��G��㓎G$�硠��~���X��E�>»r�ue�R�,�Qs<��.V���op@����j=�r��7{R���� �(��+%#��x��+�^�@�,�|{M`x�����pd5��vI�l��,����J@�]�������K�x��N��w���$+Kb#2��?)8*�q�ƣ��n��O���Oy�54i����)"�[�m����i�3�=�:5�F`�K ���g�|����qUO!�n��tZWi���?���8rMi��ݸ�XrRH䩲�h���m�ŵe�="0��[��<�L�!�fw�j��Z����!Oo�ޠq���+�:�9���Uo��A�[��1�w�j;� C���,�'tBoۄ{�8�e��y��;���	>:B�~�B׾�F��g<6{�������s�0��u���+�7�7ռ�g����n��PN�����5��N�!��#�ٸ�qoXR޲�3{zo=�Y� ����vgz��^ ��=��2^��\̃r�����:�Sl�0�n�
1�d��ʣ����uf��5ێ�.//E�����2ڦҦ�3��u��C\��_��r�:a_���?z荇t汯��VmF�:Y���4�7���kI>=11/Pz
�v�u�q��%CK�>������,�/�����|������b&�����	������(o��Z�zx��I5���1<֪��=y��z�f\����p�Px��pD�ʷ(~����S$�?eQ�ʍ]�������[TK�c�]�H*�=:}:[ʖ��	j��>iH~(��0�<:�k��D�7]��KÀ���j� ���k��U���(�u�����3�c��.��/�A ���FL��ֺ��\Y&��)9f.�r���O�傃���ׯeΟ��mP&��(�V�5�R�2o��L>β�*t�C���A������<y���^��i����wv4}�ӂ�1��|D3t`jN��]�d�[�9�|"�F�-�V|���,�G�W���/��Ry�_�~	٥Q�u'��dƶ%$C�O��}Q)�Y���Y��t���{�
��0�4�lv�t�z�A�$s8bS��_�&1�FƱ,����++T��Q'����E��@�m�ࠦ{5��p.�T�n���}�.�i�N��=��5��ZAGL�jD�g�h5��>�-�r|�y�"�i�Ώ*t`F�~6|�}�����2?��"s>��S��eg�O���1�-����%é�DB��(�ydH3e���ٯ�@�&����t�ud�:�5e_^��|����8i���/=�~5��p�-a � �Ӄ�.����v||��.6i���~�^����w�c���EXK�]��&`8�L1O��b�\E�|(P�cq�� ���-3�j½(���ُ��v ����4��v��!N��:�p8�(o��I5l��5��e�J�m�{p\�1w����v�����}k�}�� �y�4��K��PH��A�?%�?��z�����gT����n8�"�a�Tm��E40
|��ie�6Ag�FU�#�'+dR-�]�xP��QݷUm�(:�LCŲ�	6��"a����bM�k�
N�$�U0Up�Ȍ8c�V��Ƌ�-� �d4�g�1��77m9-�$��<2�,�'�|�Y�{�ݭ�$Q'�![SQf��&��yG'����l�m�lwhш�E(�N�|�+�����VӶ4R�-@_4[�G0�sN�mE�
I��r ��a��-#���E5GPW"�hF�C
�P1�(q'wҮ�[ }���S�K����e��H&�������3D��p}/��.��oo�mj����8�[�
��hED+�S�)�t�� b}��d��)l�$˛�+��l2����6��4���l���GrUn��4Q���p�>�H�֎�����Sn�h�.��ĳ~(7(���Dω3�[>�nn��fhj̓Ay�����F|���+��'S5��M1TQ�Q�L��4�lKd�'"��m�f�O.���?���}F��g##櫯���M�x�j)�$���^�\�$�t�G�qݢ��̅\4�E����b��Fr �NY�@-
�L�I��D74C�(:O�f�yK���4ghd��)�$U.�]v����U�3iQ�d&S�iSX{�+O��թy��L�>:�S����H��s�LDj�EI/B�>J�|<����~=(~Y���C�M$�d��V��um"T� J��D�e����`2]tm��+���t�r<�id������Cm�P��4��aTb�e;em��t�CJFg����B@#ܡ��,����0�2�l<}�.��_��_݋;7hD/��F]D�n�ʻ��*K�t"�+�YQ� ˋz��4�9� �af��dc�Em�Zٛ�X"#��Z��^�Վ��F�#�=���5�Ӭ�c�����I��1�Q&j;��d:[����=L��9 ����6�e��:m/��l���j�o^�8�O5*-�sBV�(aC���o�f�.:�D34���t�8<��m�mOe���L�Q��20��$��x9��UL������.k��9��K�1�x�M�>����I�r��>W��m`�O��y
�����}�X�r��KgC>��ݍ����Ӌ�#����ݐ�*�� O���U��zz<ޅ�OfK��]ǽ���:���qmjx��AT��Ej��q%d~����>ɨ�m`q�U��ŋۇM�(k=b�d��c2�]��Rѡ`���;����cj���q4|�^iJ���uM�/lc
^lM�<�E���1�G���="��.�d��^/�0bBK�^q�����Y��C���D5l䚹�5�"o��YW0\���qk�\���8z|):��Cխ������kQB�����ٗb�'vм�Q����G:���#3`������ټ?�L�Ǆ����my�z�y7o�_�õ����~[��H�8��
�<�s
�J��ށ������0n�r_�|�(�Y[���^���&�NI��S�o�X�H�<�^����@��ʺ�je3L��](��pH}t߉��l�e���б��Vnkց���V}�^v��g#��}����<������ׯ����Ã��L2�b�YbبcN�*��݃�~ШBw�m�Ձ�N�w�m�v�edP�Q����iaM1Q�-0��O��D�9j<ON�`�(�iqt��w�%�(�ן��ժ��_����( "J�XEeܮ��~������{O��g�y� ��<�,�U��%��X[*�9�Lċ�]A���ܴ�kf��<��{���f��,ѥ���f=��^�J����N5��� ���['���7U0�9`��0;����GI���5��P�3W��J��g��%����������6p�/ȏ��4V���Q:V���׌cҲk ��5p:�u{xX���(�j��������~��6R��*GG�dAT��ћ�r
4h5��|:�33s�t~�I��� ��R����̾�~��%z�(g�G�ZGy/�a��Lc[,_�����)�ZohV���ey�2����d������Ck��RR�g�|~ȝLn�6 ����C����`@4,W�����]�݈�ϒ�H�g�w��l�]G&i���x���lQn��a�<Z}~����)�b�J� �g��F�
gZ*>h�맟}���eQ��N,}'�m��1���7�Z�<����3�[�&��DVP��J{Cżm��ц�-P�h�Cz��H���ࢇ|\h�����RK]�H>J;?F}Y?���'�h-��Z����V u8A���x<�#9|����7�b��wE�fo�ݣ��������\�g��X��'�(HR�\��Y��������J\�)�A�Hf��mI�qL�S���w~�_���y����M@�}6��(D��{�|I�
5=J�Z�Zm�;�p��D���U��Y��F�ͯZ���g��xA8�
/y���������~r�+�`RG����g�����U���X1�HE"i������PIc��knM/���hr �vM�Ӂߗ��������Us�k�j�yLw��]+��r�黍ڦhv#Z�,�	��"��Dn�i:s&�\@��crC��lF�ތ����X��N�2�x��Jm��6tr�k��گ�_����Y��
z�`�Jf�/S�ZGy-���l������R��0�IMP;�>�����t����"H���'qd���K��&Dl[\�/����е�3���E�� ��j�t�-WA&�1D����,�)ᢚ��}:�i/N̶X-8�-mW=P��,�ʅA�`��t���"�gS�R�="���P!�w��@�@�)�>d�V?��T�1�#����k�R;����@���D�W�\�3��YwN&/%JE������Rr����G��AC��n�4��l>4�e�Э�
w�O�[��rs4Bń��g�֫d�J��/���( M�X}��(�8_g���6�%x��@�a��������k�m�����w%��cWe�\���)_B��0גgbs�?lzj���W��"z�2JZ����5�)*m��Ll�F8��#Ҁ`aM�� ���G�3{��JD3?9��b��~��	�Gxl�����N�#���hvqq����tP1%n�
zlo�ؒjŉ$$������$șb�_�QT}�Bs��~���k٨m�V�(�gL_Q��JY���d���^5��dε��@��o���iX��x�d@gk'�8pE=r�d&Ѻ1���^�<z����ٞ�`hRU�^n�_'��$p���jX������XR|٫���;ɮ�!���q�
�A��~�����Ǉ@���j�_�t�X4-�p�G˩@���;D�HDq�lv>� һ�d�rp��������a���4����
�`'����2Z�i�O���1p����l�ޗ��V��2`H�8�!���V�[�)�뫗o���E<:<�U�y�f�yMT+����A���b�R�xhDC�ҧVu�<�7�r���I�v4θ?5�և�*�r�uå�8Go�(ĳ���/eT
�֫R'&�3\c˶E&5��mk�c��˖SŮ.���$,fq�)����|}OlE|Sb����g)�ך8�ߦ5�Q����� �)�RU���k��2t��<k�����7X���룳Ǐ��>��"��3{�o��>�Vh�@��z�#�Aj%��MKzטŇ!�+�\�bo��I�A�����j��̽�=��8���qe�|#o:z�>t0Lkf�7��0\�rΡ�S���@e�fc���b�}���{&�F�%���Y�D5m��"���')[�Q�ٻ
/��{�5l,�̡��&�=h��`�J���1��M4����"�ڵ� #c;ۈ_]��ɓ��G�]���a�iow�������v+�q�6�[�'�P�p��\r���{�-4q��A�~�������\А�s�-�0Y#I��r]ˉYc<q6CW���)�`��w9����˫����g�Q�-���-5��������J��lN(V�E޶���\)�:��ފ\���o���k�C������NB^���?�US�zW�*��nr��M��-���Q�
8�:�{{ǟpu��Ȥ�#9i�����x�A�T���8���ӧ2�g������2�x��v&��Ho�%Y/&Z�%>�;R�M����6Wk�z�G䃀��Y4b�؇�;�:���ظ	��A��mhM����]���4@ ���X����b+��p�|L+��H�fV���K��t�.ܮl�8�6�t����P�P�4����,�������������ǜ�V�@<R��()���KP���\vuu+b��b�+����Vk��^�E;��S��=,y��ɏ����92-_}�Տ�j�������f��ŵ�!&~��u�k|�C��]�(�f*y���2��T��W��տ������J�~lI�`�i'Zq��˂�Hwo�q�Ja�v�گa��8y(�<���W�܄r�}b�I#����3j�`[b�(C�<��~��{�'�s�o��5�E�c��%�v"��B��/^��d�y������ю�G��d�t4���^䪭[��y{�a��M0$aJWl�f��y#�hj6��o��������V�2��	\���Ɇ�d���P�]�7}��J������f���B$��<�u�[o(�(�c��1Q�:Sƕ�,1�4m�׸JL��c�f�YMX ���y[�L��:'�:�I���?O�m�ԉ猠����Ì�4)JK�0�/�V"����&�֥m��b1"=d23����lx�b����<=C�}�-�`@������
��l��:h��ۗH
36�Ϋ����`@Ϧr�FU&��hk&�nr�$xw�+mw��lM�+�U�y�)�ͮ���Ā� D�h�c��6�:2��\��c�\�ϝ���d��R�d4Ql������{�K��+7l�׃�Q�,�]<�,�9�X�+��n'�{�*ǒ,S�,�mK��#�ư�x˷֕�KV��) J0I���*$p��#V��,]X��h��R��:��?,�"�0Iêl���z�gq4&6I6굻g�\���ǣ�:��R 15�<�N�D^�yU��fW�Y�j|��a���V?M�|���Z��  oq�n�'GQ�RYn�{戇2�8��CL��(�dE�L��Q���t6����!ҕ��p���X�G��!�ͺP�?©�ؕݦ-�6�����ݨ	��[Lf����l��7߼{�,c��I�R-xq��	U�Rڀ����Y=��Nv�l:Eqeqvzr.�p��D�M����(�)I˕a���p��H�zohiڊdw�Zĉ�C�t�\aA}'6���B^�N�D�$L����ׯd%'�����d2N�����j'fY#��X�uU�π��B�0CFvA��~5�EA)��]Y ����ǐ�}�oU�i��g��������tf{;�Ѵ����]��{��2��\�<(��2Ћ��xv0�7p��H�>�*C�t�8��g���Ky�b'N�,K��b�/t��t��ɶ�s���qT�Da:Y� NR�=b� ��T�����9� ���$��d	fo>�̧���.�m� �h:�&nZ�&�Ǩ��j	h��
�+����kq���p����/7Kz/�q��m�Z��T�,�3Mg6e�.�w�v�8�o`;fc�%�=��5��>���{�/O��MD�k�Q�y�VC�j�E��x����)��ѤQٚͶ�C(׺k��, �5���"4�AONN�i�h;슸0�ȀB���H�(Ԁ���j#CV�t��Ѹ�t*�r^�aL_vp�-�����x��sE�4�0^18F�\mp����GYQuh��t���klR=1����ղ�V�����P�squ�%���+��t�|���onnۺҀ)�� ��l2�B��u�t<=Ӯ/�.�/NK��h��Z>���RK�����o����Ɍ��I������]���l��X���;��Cp��;SllDc�&��Q0�-������Ϣ0���@�\�������O',�)�!N��0��w/NN0�'��n�i��?<���L�a�nm�\��ȩ�6�-�eƌ&����s�<O��K�ݮj�7�_���n�D���y�ʋ��u?,3 @��<�t�h����%����"�����<*ey��U1P�8��,r����t���Jϙ�p�/.�F4��n��[q�������M=�t<�+��4��>T�f�@a4��	�MF>����	�%��
m�)���S.[�j�ۻ����`_1C���ا���x,v48�*־,�]��������QDI�5A>B�����.�y?p��cƅ4��Z�1#\~$�S�4�|�SyG���ō�z�V���|�O�Uۥ��p<�F#1�B�`�| .�k�V兗IM&��Pblu�x�d�PlQ��D1�#����[��2p@Woz<׈�^ɠa��D{9��O�I��5v��?�����xrxT`_�/3؈�����?����-o�8�W��n��˯>���7�^j�'`lB�i����p���n����1A��m���bH�~�Z>�=��ٳ����2:���F�H��[t�b�#�b{���I���<>��ީvI*�noE���^�|-�|u��O��O˦�>��G��L��M�H�2����oD��8;;#�K�#]�T��	���������a,��W�G�$��|D~�����z����F�����֎*�GL~#�.Z����ԺjNڟ���$r�b-���a��6����c����_�!�8��Y����Ņ��,�˗/���e��˵�aQTb�˺��WbN� Ҹ�|�[�M����@Ӌ���!i���u��Ǣ��>q"&h�GM��"������C	`���(�DV��kE�ʸ6[���ӟ�Td8���_���O~����w?G+��=:��O����:��,���J��X�t���(��|�?Sg�gзfB����^������gOԣ�I��n<��m/�_]=�T�y}�ZQ�o Z�?=>��㏭x���|"��R�O���7ډ��JX)�B���x���Ƿ�?}��S��\�A�X�������\����'e\��7.�� c��Uk>1�i4��L�}�ŗ_|��\v{�������tu�'''���]-UҳشS�y"���!�����v��eb��|�w :��8T�|v�B�k�B�j�k-mc��bG�F��YB�a}��(8A	�����Fǜ����\�!���$����Q6���'����󋍘)[��߼����_�	�V7E6 L��G��-���?��U�XN �*�0.��ET%��W̟���ğP�:&����i�зW�2U�y�O~�Y�o�b�eʗY�'NyR��\v�|^�D��BǮ�h5�	�8���В���p�"diٸ�H.9��Ԏ��VĊL�U�=	���M����G�ݩ�|�܇�#W�a��)�sX�z�L&#$QGo\�?�O%q[0~9fe/�� �!y���ˉנ�e�1���	(��l6�9�;�p`<!�qy�(�?�c��j`{�کs�.�,y�è)[׉�,�m�� �����l�����< Ԓ�W��������u��%A@���!]+��W@�=ƚ��!��F����V�'7�$����Dj���6|���ӧ��݃���b���'�J��U�Ӕ���e��#���U�[+�V����:u�Qv?�8PmPZk6����U�e��@mJ�|\�v�6V���`�u�ǁ�g�u:4 �@<��ϲ�u�����e�4i�������^��^����
�1�>��O��Ɠ�����F�g4q_��K�ΐ�lEY���ݫu�;M��t�������l��ᡭ
�G���w�މ��=��#� S�01����Z�M�0� +�-�EP-`�7
w
עW.�u�@�8�em��MR�����k�s��>C��C`�(M���r-��)��-�&N]Y -Ѹ��#�!"2_}-�| ��t4V;F���J���4��ީ`�)�C(�&�U�^�ǲ�ģqe5��v�Tѭ���Ib�^�]Dbv�3�xV�=�L�j����#�D��Fd}Z�;in �)��֎RK���8Y����p䕨	�,�rݥ��ʊ���{U���A�t<1�7�D!��3������E_��b��(f
R��ش!R&���(N3Kb�~c��3��GR�\K�c��(0�ӓconnXnL��*�D����5�F>��>n�c���F0��Z��A��=dbJ�<E��oy��F~�z|`��ߡ\(��diC�\�Ty�t<�{.{�h�~Q/Ȧ�$$3���/m��z�4Y�Bg�ִ����)�wɧ���U�N���p�A�̉̆H*�K߽� ����Vr#������'�����5��O��<cռqZۦ�Y�:�e�"�X���G�Z���c6B_��(���f�*�	��P]NU��7;��4)s�^{Wr�9����E�˘X�ȵ�0.����T�a��U��?�f�q��U��*uZP�2��%�6��]#����0�㍜����N���� �
�'���o;f�6�]�Cr��E��c|�BQ�{��r�bx�sM�h�D������ho��;ɷ�3� ��&~x��*��B�\ZG>4�,�#�J�ZSږP2ث��u,����y3O�1&��Żmd4U��Z�.[]s��-#�t{��
��\�M�x[H��0��K��n�hW,qf����q�y汅��{���F`)�t��>�m��C�2z%w���U���U#r�s�h�b�G��S��fs���<�4�w�駟~��M�
K�� :���� 6�B�Eh�cJF+��_��_�~�����W�� fu�.r�c� �\,��+��
�N٣�bK�� �7��P���*���p٦o�ɳ'O��C�ӟ�Tt����bؗ��,�h�3�F[N�,�[�'azd��e�f���2v��TS��J����syY�_��#�-M�ŻcTRZS���r�Wl�oD����k�R�PA%�xv�z���!���n���вf��mys�c��ՎeLv��\����o~���^__Ƕ�;V�A�,lp�L��=�8r���#�zи���u4����B�}��Y�-�L�C�n�Ȣ��>Z�ȏ���4\�^����^U+/ph��/�����o��o...�������zD�g3>�̧ۭ(8JBي2�4�#����AR�7���+��!(��-?�M��Dm<��'�p�Sc�$�$�-��0����ٔaDy���ß}��AM'�o���l��?�����*w�Kȴ�C� �hHs�g�UE���|��g���d�7��|�M��Y�����p��F�Q��Gy�@;<����ERtDf�JM���/d�80F��2$y뫫g�dTX��OYo�l����%'�k@oQ���[����̰���ۿ�e��x�_�<Φ�
]�m����rA������1P6%t`��!ي����o^�BLc���^"�5*bX(�'��Rnp�L�z� �3}��Z���//3FN�<���+^d-�/�5�B�--��q��|+��B�>8�Qo6pfh���Hз%U�^�C������˛{����m�Xk����Z@���]cU�R�G��ϖ�{�*V�W!s�k"���Ki��cV�w����bCи!4�k�o�wo:��W��|�K5�	�^a�&�vYc���4�c�>e��3�E��s�u����E�K��m(n�A@��=e�5-0�x�B����
D���_^=��ـ�5���_<Ol��~��&��I��G��&������,<�m�$�q  �F��؆̔��f�������_[9�R���E*I�۲�KFW���M��UG�����k�:��i?Hj��<�X"�ai�D����5i\�AZm�q�ĉ�[m�Ɋ(IѸW i!Qch���ho�y��������3�b�5��d�.��қx��d��])�Y�@XL�Q�}��b7�w��)�Z�mN��=v�]d(
�w5lh-$�ce���	s�5m�|��%�um!��i:(5���X� 8�]�*�(KU͆���"��0�J��B�%:�$B#�a-�֡���zt4�����$�*O:�4u�[���У����Ӊ�b>G�8��{��I�݉o�PxXaϤ�<a���	�d4�E#5�Gcjn;�F�)�>OL.FQ��@j����̲�sQ��@Ze�m��t4�m�W������3�fS��gDf���H�%��$����{�+LeiR-q*z��	�sRy�]��=�@g����@8(�6�}�7j�3������$o�Y>;LT�L����d��H#[�8#F�#Y�Z��̭v֖M�L�\V�d�zz�4����i���=G�H�{���x� n�
1�c�����]�D��0?<�6��d5njf�Ur���;P�1��X̋�p{u%�I�${9�J�`[T��n:Fүl�W/�&��n��yz��]۪F��G1 B#h�&�h�Gŀ��郱f9�J������c��>C\�\]�-NdZ�@�7I��v�Z��ӓ�%��.�A���u5�v�U�����GUQ���ڽA�e�:~ؾ���M��
olϒ��Z���<8k*>�|��4W+X�"[�x�^މ�9;�i;�m� ���F����0���^�*Jq�o�n��`z2�����}�gIz�Uۮ���{�ֹ��H�
�*S5D��i�2�U��n^o�����4a�Զ����v��1�:�4Fj�O�8�N,�*Le+�[���P��u�u֡J>����5����
��׿V|(7]��h�w ,���S���z�j�Rf��m�~��/���8�&Q:��`ìeo d��NՇ_��F������%\Gt���mW��Rd�8VÐ��!�Ԃ��^�g�2���N�l>�\�!9���&�NZMc�6 5H������j*E�Y�
�b(h�,up�<ƣT��]�k��A��w�w��<`�FL���H��"���{����3�<���l<�'b��y���|�L{
����;�?E�;ʰ$r�a��!=��HՇ7
����>6gIw�|�e����&"������I{��}��Gc�C+��3)QG��o4�	�	����d@�R>��E��zry�������X�F��� b�y�Q���,3�x�Gf@g�z�oێ֚��͎�h�]z��C[�\\z+��^y��Ǻ����a�i# x1��YRcH@t���8��6+`�Ā|�ĕ�-2u�NOO�@-c���7/>��w/_��S'oF�) f�����ed�U8^>}�t~4ciA�@>xrv*s�������	��/����{S�4���B0�c7��ƿ<�d=t���+D�C��}G�|0�Dj�4����������H/�0�A|���z��<d�����	���/�guC����\��E�X����*����|46r�� �1+��w�(+�L�\ �-
%p �Aab<����?�K8�g�!�E����wD����q�hW�P�>b�8T�v���`P�3h�a#5(�.�R�u7w��~��B�^�5�n[|D�����-㐏�=n��Z����#>M�:v��uI,'@�c�>�'��*���>�LVPas��ܨ���YY1ĎIP�a��f<N���_no�owuu%'�/���	Q<s��U�U��ѩ!�s����ʨxF��Qy���s�b�!^��ĵQb��G?���ƴ"�+�6R��f39� �m��r�^�cV�F�U���jSɱQ&�庱����b�G���0<v��4M��C&O��	�^|M��L`�zw}���ڵ�~�d�8�I��`�$Rv6��������q�h�G�ɕ�I�E�[�c^����]���d��{ B.�8��L��rB������/o��5.k�� 77�,�[=k��5r��r���ǩ�34>L�e�|���+�A�����o�[q���y�lR%םSD��Q����+Z3���e��;���=r�cO��(/�Z�k�	�>#�6ذq��L���lmP�q�9k�K��]�\ǯ��n��a��}��`�ӪR�\����B"&�����Եveܐ�Y��|�;�#)c��[���9
5DʍE����g	3��^�f`�EMf٧,ZG���>����)�鼛�;���5��V�<���/gÅLX����/F�e��ӥ|ag~zG�l��`�����bW�I!Z�Xe���[Ƕ���J;�{l����ݸV\�wc��P.IIȧ��=�GX��F]T7��A�(�t���&t}�����'�ͺ-ˎr�9W����9�'���T���Q=\.غ�k�W6`?������~00`� �RI�63+��w�_�tD|3b��34J'��{���_� �* �.x3��E������}�t�{�jyB�?Y�	kQ����(�B�����z%3�Q{��Н*�E���퓫;��O ��޽����g��&Vq���<$^b?�H��ۭ��7�ʟ?.��,lH����	ƭ�طJ��A�Q�a�H����m)���	ȭ�d�SJoK-�P��*qWÎ5}/�����o�{&�xV�2�W oh�D���&N�2M����/{1b᡽������zZ��;����#a�����ra���],s/J������ �����ٸ� c�����bB��o5�VZmZ��G���>!����&���E�)F_	��	}Z�#�����w#�e�WF�L�ywx0h�#���^
�䩦#�$���EzI*gGH42���ȧ+�zv@K9s��h����My2#������"���:����:Z��^��`.�bc�U�ӗS��G�Į��Ԥ��d.������'��<����7�@����`[��o��� U/;Rܷ�����V��Xߦ�-�=X��Sa*�xj[�7�!gLV\olI����8.�2�ct2��P �ܖ�!��v6��x��"]��e6�]u�h�F��y�6bx�p�����jkmk
���ʅ�ٵH�832���b�P���8��n���a���A���KZK�a�U�3ߒ|�Y��c�j�n�����ɵ�Գ m�P�a��;w�xf�W��ǙY߯`�5]���1�B>gCF]�\�^h4(	h�����[��*r��9�N$v�V���Ƿ��:p2TI�%�;��F�Ʀ+�J�cx���:�V���e�2�	���V���ՂDf���`|A2o��-��X�~���F�iڻwn�z���m�L���Z&�@��
��� 3�w�bQGl;�=~��@�V��&�s����0��qS ɚΜo��	/�j|o��E�������H�gu��d='$UH�k"H5�e�J�#[��ޚ%����	�ί��=���^��Xx.�0D����u�ޯAjVK�����
s#�®!H^��61��F���:�%���F�;e3�g	A��Y�����H�d�Vs��D��H���ќ)��Y[B0�o,2a��s'�����ϼ�����]Z|�%��l�"7�^MX�5���l�k�
�$��^�.F��tpn��J$�1޿6�>y���U�no�������>���=(�1��JȋI�ٳ��yb�[��1��$��E����%������7v������O�N..��c�6{	NN;c�#�_<�6cֵQLFO��9���@��w�O�4!۵�������o���������;�ǧ�|�=2����)�����2"4�[B��Y�^!)���p�=v����ѣL@v���D�ܰ�]��� utcܷ�?�wK���)�Nf+/"_\*K"��7�ٱ	K�T� �@�H�m�u���+�0�2"���{��+$�bGG�⅝�,�x�R�Q�ikx���x��a;f��(,F����0<����[�Y����sɎ �KK�q�Mz�����H�h�<�/�d���U�<[�+=��{Ϟ=S�{�j����x��!I�����NI!�̝
S'^����]�y�q��ك�
�k�ea<��Ug��E��5��W�Q26�ح[�\��%��!�8��Lx~�Hp�s	�Bz<��%�����(ڟ�F�7G(�>I�'���%?��q��C��
bǠ����#hiʟ���,�nz�7X�N��r?'��@�h� xwگ ���P��T�]��O��){"�N��`��.�2"��)�n�6Nl�v^�z��7_�D<���[���9���q�vGB�yL p�!ceUH�Y�<�P�0XA� i���Y��4v\%2*6~g^�yV<q�a�h5�)��=��yI_�٠���rQ'����f�i�m�Ax�ɗ�G� ��y�_]FW�LfB� �Fs;:8Y�V�L�@Z&G�;T�ܪ��2�XPL�21�@�`�?.!��T�� B���<���A�:��aH��!�g�V�.֜����]i�v�(��#�E�n�&.�'ga'霤W���gt�O�0-���5\���b+��ր� �|����W7��h@�j�ϒ�\?�/���~6�.P<��9�tc��jɂ�r>_\^�ǐHf�N8��n�P�ߜ�Cv��o�%���{�r<Τ�D�y"`O��]��0��̂��{�8����d-%7�w1� 6����g"���W�! �5�7n�`8�@�����A��?:<�/���$-�9�"��u#��?��_���[�|�]:��d+<`"��.��E���Bҩǫ�<4E�CL�O3/n�ʻ�'�7$ O^^�V��b��W�����PR&<������|�Ƒ��t�DL|�H�K�:�"d�r?KS.��[.&�t��{���'��Ѝ7&WW�H�]�U.�T�_�vc��WA6:��:Id.OΏ��UK�5�d���{(.D����l���0]��q���@7�-?��yĨ���K8[���[�ˋ)����P*T����f�^�P��p�]������2�k����$#%�j8��8�°&�rC��W%�j6�Q����������YU��H�u����e���)O�l��ώ:�|��hP޴r~�^���[���r�O����Kr'
Z?_������r<6_6.!e<��i9'�s�iqY�p����͌[/Y�3eFI*7���\-fb�;�Q^��!]��F��\~I�M��g��� 5�k-�N�6N����%n�uג�Q`7d�y8��e/��<�7���ܹE%������7ߠ�Ȋ�OW;�;��+�v��YMY9�_�h'x���2��̬��.~k4$���U�:�-]{ׇ��˗U���Hq���79�L�	�s �S�4�(������WP����Opr�ȳ�+��[��w~�w>�կ���jţ��4�ٔ�[�������>�&-S�І�d�q���,q����ph	X�"+�t�牏�5�.��I�Q�G�qNq�|1qn"�ɏ��,�șY��tt:��ug�פ�=[�⧦�)Wak��K�j+ڼ.�b�ȇ�]��i��W�0Fr*W''g���ȵ�e&U	7:Z=���}���`���D��B漬�˷n��Ŭ��A*-������w:�l����� ����y7}p�Vy`�p��w#���F�R�}��,W�M��̫�;7��b%�5�2/��7��҉��Y.j�N�t���;,IcdC��hq+Gb�̖Ͳ
��e&A�R<����V��I2�;w�񸛍I�I�Wu�jڑ�����t^ѥ������uS2|���h�J�esK
M0N+Xa��^�Q�E�N{��.h�������h��7H������r����I�L2y0d��,��ԺJF�ӕ����k,Km4�#������q���A���&5�$I4愓���81�3�NF�{T@C/[��u
qbfQͬ���_�uȬa�R�u�7S#=��jzDɩ�
ZR��'Ӿ9��1��a��S
�T5A�u�G�S1�lȄ)UCƒ�.$	A���2�Spvv���@r���B-�3m"���W7���P'MW���:;.�@�l"3���$w.�!��ٯ�Dm�������zP<�d�Y���VoJ��j�������`�wwɬ?|�MRZǇG[���M쓻��|����%�XL����ՅU������ue���U'�%d,�e2KƣF^ǣ�O�G�����d_�>}�qAb���4�k��1�
�huIݡn6�r��ڞ���s�˻ts��.���w����/2)pr|~u5�����^|�	ô;�ņ�����?���蘮0��t'�O�M�Q�EH*R$٣;9���D�sơ^0��
zYRz���>��������U�XK�ܙE���@:��	8΀��J:����Vb���C�J��`<��SN��%	��p�s�x_�������[�0�$�;������I����W�}��`�|�=U^���I۠��!�e�F�Y: 7����WlL��,��j��V(�N>'��u om�<;;��2�.%_� �`�\�{���h:T��e��H�(�#0��x�x��u�SS��e,�U�dʮ�V�N��� �ڀM��,"/c��?UmE;�k��n%hrN�����mntȓ�l�x��o��vY��y)��]���Xx ���Q�#v�ӪM��*yh'�y��D5�,���(R`��E咏3���k�A6���a�n�O��ӫ�Z�/��:���I��P�!�8��0l�W�C��Ɉg1��a��t�0p/�Im��P�ۛg�G�Wg��F:�U -�.tk�[��ڦ�ס������S��jػ��(��5�n���v��Dr[�<X���pTբbMoh;q0V��`�]W��J�?�.��0v��� U4i�&*����l�� �7�2�iVfM� ������J�Ĭӂ4^.��Hy���z�wr׸fH�dG���@�w���o.G�	h
V`����ɀ����ɖ؉9n$�Դ��[�v�I?}��͛d���}���o��C��yؗ�8��	�#�Hg�58��8u�AM��o������&���S��oh&��Y߮Iw��<��iDR�LM*nh�Uz�C�����#ۑ6�o~X�Wp���8j�5F ���^Y��A<W��f,W�zcנ� ���SpA��,���E�u4��;�X�8�:���!?��F���'�)���P.=ԭ{�o�&1 ˯��6����&�SX.9G'�YM��:�8U.��+W��DK��6�$���ͱV<�f��O���T7-ɉDL>��??�"�J�DQ�HZ(��hO_w������$�f�l��o��o���w�tͿ�ۿ}��K[�इڋc�ם&Vp���pR���ub�F�Q��&�qq8?E[���_G1�����I���FC�ky
x�����+��
+h��ەU���59�ۛ�4��M������R$�u�l���n�a@�6sd���	p~u.����mAzzr"�kh��zfߗ�ҨL�������� �%��ggט1G;2z�(,���KR8/�BW���$M��dvt��__2�I��c��kI��	��D9��3��y�[%��.��e*?;�`k��\ӫ	N_l)����=Ai���i�<Q�����b*���GOǣ�����8��֑��g�������c�ZL���ma[;=>Α]����/�v(U)��`��t/�^�����pVF��/<+��(Mo��_n��G-���fHa�6���w��̀a���$��e<�����R1T����al(�������C�s>�?{x2��bM��|�����g3��*�'��Ւ;6��ON�[��x��Ӣ��e�R�,ٿ�H'3tK�L:��r?,��Ʉ�#,�<�>�`g�̙e�_�����������?�o�����B&
������c�4��D��ph�?��ؒ�i��S�H���")��Z�������t�x�(��.d2�._Ws�י��n�����XrKdB��'c�d���n�?�����~qy��ٳH�".(�l�5�F�� ���5���r||L�U�ӌ&U<A��P�\_6�m"Hk4Y�"w㒘��V;T�b�0f�U��Z	-N���nެ������ş���YD���6���L*���@b�������*W�B�%� ���Ν�Lz��qQ3�\<=,ٝ�}p��%Y��bi���ʁ�$��$6<�I{.?$�tâ�bo�A�(�z�4�@���p��Q�= a�1�&ڬ����m��z�E�Z)�M�G���8u����xI#:��V�q�y��pY����B0 n�U3�b�.��F]'�=����&�<�ɂxxzA[u��5zY��"��"�jt(pߕ�� �"�z��u��h�6T��y¶>m�N���K�(���i֠�w�B$@�e�P�Yr�>���)r5�i�#ܬ�U	��
+
��R�Ka����=He5�Fc}������kCb��+\b��Ҏ��^�5��A2Vm����/�`"}y�r'�������ڿ9����߇�+��pc?�(�a�,/m���Y����ۿ�ۤg�	��a��F�ޅ蘃���/���O?����_��{�&�&�Y�Z��l�#��R&���d�����Me>�^M!�Yh)�^M���!ir���$Ōt�}�C�j�Dp֜H]%sNl\ $��	#:r,�U�a���Љ<j�OT_�z�$���gTB�eq�
U0?҃#^3E�� ]�1�
���(	��:6��G�|�ݷR��C ����a8-xم�}�n�+
����W �&�C��hl�xv8ݦ��^[�S@t��r8�����LE p�v�.D���o�Ǔ���Vh����
�<���'O�<�����I�������~����=RD83iYE�]�$��Qx�W��.N"'�Oz!?�fœ�)A��WRW��,�G�I^+��Z���b�h=�,�w����� �3���[�A��xquE��͗�p0p,#^G�c��1���ǮqV9�NO���+���\ q=?=���-��
<�yoְ�l@�h[��a�E>���T��e����f9��8�msUt}�2 ��97a��@�U@k���=0<��`�F�?���:���V�����Z&���&�@���%�	skL:��>$�lz���j�y��:܏S���Ν;@����=R�Pd'�oWr��聶Cg�� S��V-���)���ɳ�ʺY��x��7ݴM�CG.`y|z&rA!=���2��$�ˌAy]�H�H�U���H����/��j��r.I��Qn��WCn]n�Ţ�����&�v��
NDPv���j�:3�<6��w�}��ágO_<�S#
��Z�) n�!��ո̳�v�-'^�AQ��VnM���1�miD�,Et�� �EJ�i�t�3�ض��ie�Ib����R;�;��z���"��%4�ī�q	��㻠� ֭r��(�3��aq�>�7��Ps�O�t�&�HByEY�Dp޴%��e����p�W+�6Ϡ����K7�,�8�*j�2l���K�"�ٳ�wH7" ��h����1�H~&_CB��@���3����r9�1d�6���{�ũ�wu=�`���|\�ԁ̂w&�e��"�`S�VG��n�k'��}�l��Dg�n-WE��{67��t�Z�;{�5uGQnӺY�U<�4��G L7�BS��~q>	]jю��j0]M�d�o���(��@^*}��귱N���0�G��{E^��j�ΰ�}��e)DrNXDI�5u"�{tM>���IVS�p��?8�a�]�F�JhU��%#m���+�M�\�	�W�Y3��u����f`΍}6�WW�|QֳrrzU{v�BD=ȹ�4�]�p�kvt���{h����f첓Ԝ&�M��%�8鈢���f�����t�\^�&�:ϊ���̼��m���OJ۝r����m�Y2%g��U)X����;�~��{�ч?�����ϦW��tuyy��φ�g�Q	Kq��Ę�aC �u`���X ��L�I��`r�{�E.����b�ӝ:�HJ_!m8O�Y�^�0E;1���ZMs�S�!��~������5���a\�c`+?����N�lks���z��Kz3���#V��e��` �i.;g��s�9�$j����YAS9�;�mYSX2���٪bPp�RX�L�2]ȡ��ty�	�<�G�b���[<\�a~��H3W��:uz�E��x���O�G�����|����t�҉��O���D��!Yξo,�t��R���+rP��n�0M�&0m�wֱ��{h��N�MI�+i3���K]����u�; �q������o�NNIxN�O�
�R�a�V�
�a�t?�W�Й�s������ϥ�M�mMYZ$EK�e�C���X��
!=V Z&@n�v�|A�z$����Lы�zׄ ��L��4�.vdns<�w�����|.F#�+�y��W�9���ݺ�)�d,D6�!(�LS$/���
����+���H���y��8@��n��86�;�L��]\ϫ&�8��H�r2��K>i�1��������e�2s`�!���S�O?����x�kg���j�`��L:
�5���(�vX{!ni��1����@�\���>�j����ܾ� q5��x�Y�y�8CD�6n&�|�x��0�FRy8�M� ?�� �^�5Y����D�"oiM�����%���Ŭ�4�x,��*�@Pd�=��Mb6H׽����wZ�&��2-N�
\
$zH���%I��S�=(��K�O�Yg��~���:-���拺uL?a[f�^l�#c��i_�F�tRҌg^%Y�ws_�
�o��d��-ISO�]c>�f�L���fP�l��� �Ud�Y�8P���Ȭ-�Kqi�vH��N9���_�;�$%���|���I�!>�۽�M��/`�<x����ڊ����;;�b�������B��������������Rx�er�o��o~��A��}��qp"Ht���7�_^ܾ�V{�ƍ��G�z?��ϑ�c��6���1�h�88��)C����C/>y����A����>Y@����x﫫��QH���c.��f)STW;�7��9�s�޽�����p洪�')���h�=��D'8��0����Z>�9� �v�+t��<Of���D6p ��ҝӥ,�:�j��u���礤d��ݣ����~��sU<��3���jЛ�强��#���2����"n:99�/��C�����z!:�(z1$��^k��2J�I�op?t �Ha8���/3���;q4��ӈ��<�q)W��2��Y�O&���g����O?M�ܷ�j�O��O�~�
�s:2>R�ݼ�wxĴ3�wň�*9� s�Ir�`�#"���+L�)U"K2��_��(]��J^�T�y�d>4���f�^\]�����9�)�*�����r�/����?����9��_H��i\>m��X�|�@���?��T!�U���Τ���`�pa{w��]�Z"a��k#" � @��	;G��5ePi[S���'$N���k�$~	ƚ!_Ǡ9�U�G#�O<����ao:�pӔH܁@PhE�e~�V,86v��h�N+N�Н�pa��B:����"�3/�^&�]Yv�7Sf-�d�vE�}���qԙ�V<�7+������6�`�$oڥ�T�ʆEt�_�|�s��A��N�Z;;����q��0�ȃ�cUƉI�%Y|df�O��]�Xj�SX���#�e>�*��`^��1��~��j�x�:���U��A��N7`^L�qA*�B�p�X�j%�m�Ӳg��D?�M/�dR���łs<l����5+��������D���+��E���6�0����<��\�Lע�_f3��s��h�XH,M+^ Im�)�@Ts�F�2׬���$�J�eY.�_�@sFF�Cq:�J>��F�1Q�s�4��m8$����76Z��]�Y�o�[���J�Hd�pN�x��H������t^��E�� -���]�x@���Q���5���K�'G�U*���$����)���t���z໠��!͡��>��;����qN�
��Y�Ģ
��f'���lI�i�a�ҙN�b��D��%)b���O��p���(����g���{�gV
�ˬA:T�$�wk��1�3a��l���e�S��w���\,?���ӧ0tP���	�,AS2�Ri�ř��;yb���hZ&�#�Y�9�����w�w?��������NK���S������e9y?H�dbJ�^q/�Z�I���Q���
���l�#*�,�x�IQ�F-+a���fx�E�!�ƑA+��U�gx�$,""�yq�-��.��$�l<�+�ys�}虯<���DFTߴ+���LO#-�	�'��C�j��H�G��U�'#�F�0;<��9b��0�S��$�&7�ɪ�LL��[�������Eg��cwu=�L4!�ȷ�=߿s���j>����_�jY����?|��EM' �%�ʤ���)��|%>4_$��+4�J�����'%-K�=)�	YZ�"w����x�N6N�5�X�J��P�]����P@ى�0m13+�C�x���)F$����Ǐwb;�4̋qLd�p�ঀ,b�?m�r5�㓠�
ycO9�f���>1���$��s����ЊX�:Б�`�H~8Y�$�!#�ʕ�qV�2i(H�'�?��?��"���?��/������׏�԰��<���R��1 G.�;�8�Ä.����M��l�Q�Ҋ#�K�wX�l5(�DЈ��L��z�ʲ6�%��V`�g�"d�����=.���"�G_��]������W�̙%0M�R[�Z�K�	��&� �5'�C�0� Y��-�+=.�'�d�̛Mǿ��M�t���J\�u
��M�f���h��'���֛o�{&3�G�l
��G ��v#=k�1Z)㰥0�6my����]���4IL�ZUt�=z�I�p<�q%������d�wu}�U���.x�9�]LU�q�rzrI�A)�J�x|��$���띭R���pJ�攙��hV�aӲ$�V��;e>jjI
�.L�}E�j��= ��ݢ=�HX�ژ����u �W�7���򔡙`Y6L
<���b��6���9+���ۋ��W�������uh*2�*���8�2�,��(u�	I�=�q5 ��j_�����0_#�t�F�c���9h_�eV���C���Q2SX��p��8�A~��r+�|Ѓ´'�	`:�ܰ x�D�p*�[weY<���?H׈�OK]0�$��%��U-�8��oޏܾ�ss$��B}&�"9HNNj��#C��[o�S��0����Ng�ǟ�����i�p�}R�!9�|�	� 76Gϟ?/%mI����D/�~����D	`$.�H� m�Ѡ��C ���EY��W���x _��y�޽������/�����kܺ�E_D/>y�@r�wr��|��BB	�`w�{�����Cc����jGE�n�ǢF�Gz�="+�h.�ևԔ0�6��T�㼖�N�n�My�/���ex �N��nZ�M�C���KL����_��_�R��$7������Z'2��P�Ͻh�!S�c��D��%��������yi�=��c���B��Ԛ
½~���Tn=A�1�`�,z}�S�8���VL�J��<+lX^Y�j�F}�m}�����[�����}Y�ܺ+!O���� E�G��#S���`  ҅.��S����� ��S�TqD���G�$���L�FP�ĮK������w�B�|rd!����/����.�l>o�cw��M���iP(\�g��&(g�$�t$�k��w��z�ݐ�X�D�)J�ǔ��YK_�%���� Cc� ./��>w�(�Bj��6�v���jE7_����M�!5�MiI��^Ǘ��v�\d��V2��BmN���.k��ce���|�&*��[���}���|j��>��I!���DoG���`<�Qd|����B�;��"����j��ssg����/�4"K�J��8�[d�<PKN9q�@x3
+��wnQ-Y��僬$�9i���;V��N��H��Z#�Y����{&t|�[����W+���J���]z%`K��Qs��1� �L%���d�v�SV�MAaBr!�tZ��Ł{#����8X���e�E  _,u�R���H;^��6��"�H��,��y����1���7VYu�r�	\Kx�}g%	��`�X2mi���+HB�c���ًe	��|�
�\���
F�4�* �f�s���_!W�.^��h�Ʉ������;������uL�vm�����d1%��i�M�/;]/QI��u c�;̂�Pq����$/��1�g�M�G��VbE�Y�
L47ֱڸno�2�Y�T��J�GÂg�lF�����/�����7߸�����}Q��l�����i�Q�Ըs�P�J�;.���/��.�gi>���������f4{1e�aא>�HB�T�=�5s���ݑA�p	��Ӣ�⟬��N#yl?�/�㧟~�����-�RP�,?�g�'<o�<����{���[7�o�������h)��5���z�O���ŬLb[z�h�O�r1�q.[��2X3�\LP��3 (�duqM/�q�YL�8Re1z�#�p`�d�0�?��ζv��Z���§oߢ3�P<���<{������<v�'r�7�p:�ނt��9�hY.f�<.+I`�B�H���+�EDRJ"K�P���=q�9�Qsi����(�G01��d�e25ׅ��C0����{��������N������	���nq<�v���1y��@2�c��x��?�V4�tٝ�mr�ي�dj��"hw�>Jla���Ad-�K�t;g�Q��D����<ߎ!sӑ���z�M��#�x�"����!9<>*�j�;o�p�]�����씵�s�2Ğ����ǀ�#<�%iB�>[ԁ�S��]�ʾ�P(q�s����bN�B�L����6Ȏy���}Ɍ���w)�4A�VLlU)����)R��"u��������~/-|�����{|���_���.4d��9����6�6�I6�x*�L�Pyk�+�w�6U�(��>�M	�8�+}���eS�ů��

�B�*1Ĭ�nssh9D�P��f=�Y��_���_~A�-�C���]��wY�2J�A�3�N�������>O
�L������V�HJ��`T`��~�ފ�c�@�<����4�{���F���#�$:�Y8���l�8n�i�9N��.$ņVeNOH��������R����~'%z߿��NB����dPŋoGg3���ƃ���E �t�?v�8O����䮴W3������$���wcL�p�67�O��8}�T$hq�Z]޾}��
�SR_t�@���}D��@�om�H�hp�؅@�ZƎ'/�{:�(���9�6�\X$TAp�z�qi�3��&On�|�=���ޥ�*���9�X�10:ؙ�>�R>Ô�~ư!�^p"i�N|��8"&#�яa$cĲ�"��@-�:�
�Hz�U�j%�)�d8��'iZ�ԤC�ll��dނ��Ȗ�H�p�i�I��m"�u�@f2��q=m�Q"����s��*����R�%2�l>�j��B�le�T˭En���9�4��Z�L���"�g���j+�%��B����+DXf��I˜Ì�%Rt��U�u00�N�f��y�a���3-��[Օ���bqqZ�\��s� Ȁ��sC���I}��L6'9Od�S,�k&z�ۆ4���=�yv�G�;+�`T��G��ɘV���B~�V��N����*����:a3�X��偂�@��|B��V5*	���(-H�67�c&e�d固]-�?{���1�+�x�s?�e-���B�gϞ=x��OM1���]_W��x� �����p��_�B�����19-d�Vt$*r���L��H�O2��L�]���T(D���[�h}NO��pr>�ݿ��{���j��2�B�s���Մa,��_|�h1�ӷo�p�x������x8H7Ӯ�M9���m��|�M�nݻ����Jp����z�����!g��P%Sn�y��!Y���c�����=R�H�X2t@h>�~ƾ���D�B,X�O&�r��G�H]������~�������l�Ȑg�N�i�&WW��>�����������}��ɟ�ٟ1α�h�����u�AMr��ȴJ�ŪSVЫ����çO�޽{�G��EX�jv�;��9���@C���̀p�@��q��K:�횋l6���f�����+p�L�j�5����%������@���u���b=�NW^,�"�Cѝ�
A�Ջ�G�g�	#C�� x�Q�֜ţ���W_�zy4�̗��\6{��:uE2f�܃���6�R���ɴ. �0��K�,z��3-���Y~iK� i(%�+,V�O���/��N2A<wд��5�r�9��6w7%!8�߿����ղ��׿rM�����_='��HW�w�y���.)�Z�	Z��.�ARҍ;��L'9 ۤ��p@
����O�}����鱭�q�=�Y�o��C���r�>ͥ�M�#��ܦ�(8�!�#EΑ�q�K6R\r��N�Ƭ}݁+|���$��+��JVc^�H�5:r:�uu<���j ��H�!I�} 	4m��WKwm�Pf�1+���B�*o KL%a�$2)R���}�D������ �^�lZ���\ܾ�
��N�$  S�Bl�c�Y��;p[W�P�f1&sF:eSzO��sXY^7�lZʽ�W�%�y�I�'�1'��lJɵ�S�WW��2,tN�䠐��!rt0	� `�!������l,N���=z�R��d��H7	�rO�Q1�����y��ۯ�cR�E�dD��=�Ŭ�B���5��k��=��Z�W��nwzzIJA3�ǋ����v�A�0rU������#4`���_������d����#T���]hKm�^��4�43�4�-�|0��8�{(�tNS��A' ��7�z�1,�1�$(�.&.��[�����+�C6u�p�z(8���A�?��\���Π���$�啿���I��X�;t�Z��)���lk<j�C&щ��1AN���o�y��	� R�t�P�B�&&Y�O�f�{='�:�n�$b�7r����}(�љ��ӌ�Ck����˪�Q��q���CqZc֙L�B�HB�O>��t:|���?��O@�� �������5=���)���PpܕC�q����Zxp��(׊�܃�p�Q n瘪�|C]�I�t4�U��s�֪wdҫ 93��M��3*Wi_!�&��r@1,��(��m��������`�v9a4��!Y��~���PQ��Y~���!w�mJa�(����Х��?����N�  �TIN��h�z�/&a�� ��~�z��i�8�Աz����^���+�4@A ��K������Y�_scڅFt2��C��^<��B�5�{��x�D��������{7n��m� աS���JZ��HoK�.���zS5��e�zi��L{mq��� ���H��/�&c���a�N*�o��X.�����N$�\z�.�7�7e���%� ��і=z���D	g�G.3������I|��h�WTW�
�oy#� �bPd��@ێ�6���\@��L���43���x��F�àT���)�#w����D$�%X�d�V��z��N���k�`�B܍��#�	�I��'C�}H��ܹC_A�6&݄�/(�L�y� d@ʜ�$�<��4�)�D0�n�Ȉq�i�����>��o��v�$B�8�|����N�`]tv�!zP�C����˗/���2e���X��(�p����,Z<c�̿8�nhӳ�8F��N�f��A��vf��tS>��OVT M��.p^g�I3��<L	�q�5T�M�=]��)��d�h?��<���!;�ax�Z���O�U��	qe�K�x��^�$��NG�ܚg��k�3����1^Q?����PAս1�5+���|x則�H���M\1x��8�hCӚ"�m��$��$�_ݛ�[C3 ��;wv�*4��1K.g	S��ܭ��J�V�jp����
kP��u�a�"����b�qF���:bU\��+�b8b�5�^��U��U��$2�<���h��ȫ�\�{��o0H�(���� @��RCӛ�\���-�M3��L��|2��&���������o�B����!�QvPC��\QȀ(���Y�SpcW0�+��э����7���_^�i�����KS�tc@�{-�cz,�"���ɴ"�I��uKhO�82}��0"��hD�h�B��۷o3W��z̎@�.v�ZL`
ܦ+����CFG0�����܍r��5��p
qϦ��f2�p��`��(�"�j�� ��9��?��>������~���x�b6a��~�#z���.<z�Y�O���Sa�[J��(� ���$ ����f
VT���.�<���2`����� �,�η��5(2�YFM$U��KZ�L�8mo�ve2� ��W_}u-c�i븯E��d�i5v�71<�i��S����2}� �3޼y��p�8�S�#(q�����^u�WI3�����S[�K�yiX=lV�-W��ƮN���/�20���鄶t{�6Q�d(��cXVÍ+��H�+~o"6��{XR܆�R�<�z�㐍Xۓ����>n�y�0vpu��p�+��0:��f
WBM��6K�������ƛ%�zI:�޲��iY�0�䘭�ql��T�E+�)s|��As�ʣ��1і(���-:H��@g�����W+`��l�-8r�< H;%��ZC�K�`3ёܖ���]����=Tee�7�����h/�=��.[�ǔ1ŠIv0~AYS����Т��~g5�I�
��]?Ud�|�V������7���ڻF�"g�K�A���b��u�炝:��p�!�b��f��-�,��K�[��Đh0]z��I�8��ZbHr2��C�\�[OK�	9�:kf_j)���B�6�^��i���i��4�݀fu��k"�������?�=/٪�
�}D�rI�!6��" �>8fdH��2�����m�7���L
����y@p��A1!�f���ty8x�N@p0i��-��!���![��vk!�Z�Z���_�?^ի����w��'��ī��%��a$=��l�l,W3�_Ӗ�b$�,��A+���U�؍F�uy���!���A��&�߭���w;+d�p�thX��J�ہ��~��������C������'���Š���9�Q�ż8��Z�77����Z�6n6���rQ��7muN�2�w2ώX讕i[l�gܻ�
�x�NW���.�U��� ���-<P�"�����fo�������,�/~}Jo�w� = L&pM�D������\2h��Ψ0N�.�4(J_oVT˥=��>q20�\2kY�\��L��S�����nݺE�F�C�&�ӕP��R]*��i��`�7�7X��z���l�h4�x�wn�ڧsDn(���D�������z���#~;IAƷq��2����b1ϳA]q� �čh��   ��IDATd�i��cFr�fkU�$�ր|�(� � 3��4��`h�.�����~�g��#t]����b�5l����k:>�YL��X��\V�����օ�a-#�lr
m`�G��4NM)�	d�Hу����L�č�l�%5O'���޺��+(�lg\��J�_��_��׿�5!������ոIK4�Os%��� >� �ܼ��J���_�ѩ�qF��r֞3�1��+X>�:A��!]��C��@��eD0�� LIU(泲�]y���*'_�R,Th�w{��_�GPNuӒ���j�����	@�û�̋�{}����N"9�t�.R��~�i�S �H�Tz�,>�B��K�X��Ӷ&�,;g^)\X�8��;�p4K�H��;�!�����!�n)�)�ڂlcZe�C�=h/�]�"���Z�Ӛ"�U�M�F{��r���g� ���͵;���J1�,�������iβ��2�� �y��S�22<U�kN@��c��^�ՂoDtb�\Б�6F�qN������ї�/N�+=��7�6�@;�\�Ydߓ�*>�YJc���1,	�ـ5�dq�M�*L�:��k�*^�AR�+��[� ��?oE��׹�5�ii>��A�i����J.�_���Op$ҁK��k������0���M/OO��N����^V�wu���E�����W�-I��o���Ȋ/r�iњ|�ʗ�c��d:r��א�6 �t��'�1%X�1�))u�� ���s'Ɉ��U�F�!�EjIX2�� N����A�TSt�qI��]�#5�|�u���4�g�rU�	�k_9�B�V±�\qZ>�r��AX��q�s���!]��%�D��1�x�d2)�$\_M�V��Ȑ�
�NS��F0c�	$U��Rmo�[�鄦J�ݾVABن~vvv�	�;�2�J|ӛ �|(;{������íN^2W����X��c�������;�ȁ&21�kC����_��V�{����,������ɵ��qc���9�I���\����� BV���	W���H�Kg]H���,Sn�PL�X�j�)K��n��ί�bs`L�76���&���&/���Z!j�1���tB��la_�.�OH��׌�C�y����D���I�=##���߽{� �/����Ǵz�\a�a�a��ҁ��Y�������J����)�nG�ƭA���^'�L��˸s{�jʹ�(g|��������[��_?��ѣG������~����h�Y`9�+مVǦ�:ईO���e� �J��=`ΰ쩶�c�� 1��!0Hf��i�>.K&r�E�i=�
T
��$9�A��6���*�碖 h��\�g�Q�aU��M�&'���!��@3kP�3�
�zc]���qY��Cq����w�{��`�u1wL�x+�XҦ ֎�ȧ7�K��g&�gS��A�~H�Buc��E[2��:]W�,;	םU_;�rN��u��&!�Y�W:Z�߯☸�NO�.+����r%�W"���m	,s�E\�4�{;�X��^�&0��f�R�F�nt�|l�,I�����8�c�Ɉ�Tj����$�冝��-�I�d���A"��
/�%�5�8h^�S���戩�<��'E~J���L(P��!��^��0z��7b.� w���r~���)8�0��V^2V+ҚS�?K"�:�4��)�~����-9+_�]���.Ny�-yS����d�L��I�۷a�E���Te�8��#Q(|���PL��Q@�{ ��{9�:�)�d��^��S�B�#"R�<i ���]��'��Od�PO�zH�<�u]�A��О����i�;w�)^��d
k������wˮ�X�RU��3���5��㘽����.�/���.��ų������?�4� �Z�P�(�A�3-�<#z4�L��	u��R�D܋�乾騢#�^�<��n�ZR�1��=4����i�h-xf�p ԰>��2׬���R��1�����]mr�'��p5�Y�x(�^�@3��hHw6���	nLAG�����xj�(��o�)�׎h�k���Z`fu]rI��������z#��2�������5ʧ���,`Rd���-������oRP\�ى�U����1���@�I$�J��x�A��|�_~�@:��A�h��XrK,Z��~�m���k�e8�n�D@�:
y�X'���+8U�Z2ϯ��K.�9��A�Q��,�6���6^
��G�*�IWKN����o��/^-�����{{{H-ȵ��H��O�K��xN�Ν^�U�S�������7�trk�h��G_
�Hjݕ�n��:�𼈑��2�X�	�����VȢ"���^$������&	Ӑk^7�Lm���;��r����4�����ܜy�`����cb�&��N`�,ے�6֤���� )�0$\ ���2�X���ڠ�H�x�y���5O�����~��h��Z���P�{�|��F��\:�6�fGX�(�t8~�c�n� �S�舽��A옸^�ۧr�ۏ��dFh�)T�����+Ԃ�-�0сBz=�Ū����U��Vi�@P�aP.?p��-��BnŘ����\��y�:`��<�m|��9���Um4LjΒ�)�-{��� ��v��z�`�sK,�"�����S�A�&��lj�p0ތO,���M`��L�
�{�.`�0�N,���ڭx�`]�Էө�x49�a\O��zyR'2�:].9�h����ڙ��_@�t�8;�fAqA�dd���A5�j-��,0���`gD�?�O͆�q��cH�Ci$�s���+X"�y�VJ�(���?c�G�N��C����N �(�閞={A/B�gj"��3\��9�	9M�`���K�Q�����{`+ɩ6�b$,2=�;�d�b��L���N�Sܽ{�ŋ��#��L#�n�VvB[�?k�r�b��J���$"�`�'R3G����������ڦ���PT_|���[o��ah�X��L9�c���K�m��8eq6t�2�Y��%�5[zsZ���&´�^NJ�����9J��*21�i�A�7ɟ����N��? -�'O���>�̒��t*+��n�^��E;88�w���9:���ń���l�)F��4���a;��;�
�h�i>�Q���W�%j��F_9=�t�5�@�p>��w��=��1;e]=}�����+�9�h�x��9<
�Zh`>�3��+^�t;�V̰��ցlG��qZ�W�(�Ԟ��E�opI4U��:N+���a�꣪����s��F�Y�Y�N�[0�-�!����"Sf�Cҡ��]���:V�	V�
��>�Va��ߠ*sp
h�Z��_��{4?4'���J��b����ъ45ugfG2Sc�E9t:$ڲNSՖX�a4�m��*���Z��	������HCA{nn���St�`@�PQ��1�"������4���}{T����t�:�w� ��(#[_(��(8g7`��W�'�)(-e���jG7�`v%Q,�سH�j�`|:A��r�ֵ�1�%�9��=�y�Io�	
�.Xũ�¯��+��꟩��>k$��%1ci�#$�3��G=�>�N��܂�YWA�u��v2dM�b��������u"�C�޸��%��˗/,I��i����$5� �� ����C��`�	4�����DTB���\�0+�{`��P�|K�Q4-�M�HK@�SD�:ؚ�juU�,dX�=)����*Z���1yL�U���K<���31`���>�1�1�p�i"*��c���dF!#>I���j�-�ʍ��\ZbBf�ā�Y�?~����'|�ȩO��ˉy���b��L����4�uS�L�.f������z��l)(�N��{����aq��:�y~9$~C�s[�-{��JnR��c�|��A�-����'�|��ç��ٔYZN��B_\rN0�UARM���Ky��
h����ZV����ȶ����C�����d�W�5C[Og��1�"�|8�J���D,u���՗��B/�d��7�|C�G��|D��'ֻ�]^L�M�I��Lo�q�����t��r�ӽ�}�M���9C�m2��a��\;e�YZ�~<��h 5[2結�$[[7o�ѣ�������ef�m��o�dXU*u����H�r:[�Rb���f���-+��Ў��F�<��Zr�DRZ�,�W��p��$�����#d)��A��������[O�*:�(�;�u��j[�f˘���#򵮮&<6s:ŨP �%�fEG�9��(��<'8f�b4��_U��J��o�3%���D��J�E�l88ږ.�I%U�H���,�\$�G��J��M����h���9ހ̓�[�8�E��5-G�]���F����%��H+�d���n�;[&���n�DC�H�N��	P�<�� :=�pH�<���he�xAhp��� ��<r���hA$���B�%}rfď�Őf�V�M�{��
��6�� b����8V�C�HY�E5��_�vN˕XV���@4hy+��B��-qcI�+zY6� �I��/iS&��{�c�*�D����5G�퍪hd�����!9i%	{���+�4�	�o^����/���OHE�5PB��AD �	P�N��yOR!�LQ�nx�U��#,&<��MM��*�A�#�T�r,<f��"����&�dΦԊ2�7B�\�|"���jV���F�h�kt�*Er� Cs5;m�7ݥ&·�#����
wҮ��������ϭѡ�҈���y�=��ƞ��)yN����Io�ʷ��]�LN^�.���!HyY�!h�'Ӯe~z��,�⦒:��A�����4��[�"�̖LG�b����=�5� ����(,�23��+d�j\#�|��t#��p����2('m����\���W�D@�5N�d�s����] �6��I�π�ˉ�Y��Ύ73a�MiA��*�������$�K/.�h��6$̿��M7[2x�lӊvT��
!SI7B�&U(���,���6��W��}��[�d	Z%������D�7�R'''��@� �hZ�֮mz'}�ŋ�
}� ���94���i�#���oܠ���fϼ\��Oߝ2���������/�F�����cc#���gtN������kZ�9O�lI�0,0$L���#����Z�7��A� %ڻ�b�݄~��ބxˢ5����(����-4	�*$V��h�V��{Ol_,Q�i�կ]��#`v�<o1|NAhs��9�`�_jۇ���Z�W�ϟ��fy��{�\�g�G:(�;w���E�*��ŝV�L�b�X� �Mp�<��Hiك���|$K�9�t��<#ߛ��j� �~��u�������m��;��|A�����z:�����1^�22?���J�66W*G����I:f���9�=A�~d�!F�_U�!�qy���I�G�y�'I�O�*���Q)f,S����J����2��=Ҳ�R��6�6|� � ��I�%��䷹r�P���Q���#���\	���x:��x3[0FN�LѠ�툰`�Mb�D��i8���b��]��6=��%���]�58)H X6w�j=�Ӻ�e$E�#w�Y��u���tt*D�Oϙt�ie������
�%�e�SbEM���A��-�,��J��42��8EH��Y��h�RQ����B�.2�
���4�J r/���e�IiY�iQ�b(z�zz��ܖ����'���-��.B����e� ָ&l�ylN�ĵ�؜��ؒ�����ʯ@�W�,��P6�odȤAϰ5X��9�*b��4j�$�Kܼ R""9��(�AP�-u�������6���b<88�J��_}xxhyz����f�5P�u�s�H�)�5�V�[�ݴ���T{{��)`�
c �!�HZ��������R\��6���.�8��};���P��V �K?�=r�P���	0�HB��M�O��j�j���Q�%/��TtWd�N�������:v"�2�oƬ+&���Qs.⳸��F�0�Hػ�>����']쫊sxxe�3+���t={Լr��U��>�F��p,<���a�Zx~�'���������Ӌ�kN�ĊP*��޹���O�ͦy&g]˚�Q��d����%}d��²PH�2�p��gM�PA�П�?�tf�t�p��F���t��P�Sdү����՘�*+Uo�$�=L��s8f�c!4:��'�=�c��V�i H����F��(]ГHր���|i@m�;�ҡ��\o0 yx���;�J�l��#�p���NF����J��O_E�S�F�H�-�m���XT�`��!ȵAb��1\ �)ry.f������Q;���y|D��(�/�)aDw�Ŕ�:���$0����U�84�s�hU(��F�Ƹ$��>E- <�z�4��h=��1�݊�HJ������I����N�.-$���drEQ��D�#&.��r�U�8�8�D"�N�6��/Q�s������Փ�Z�ɳԀ�5��hn����oܸA~ş�*��÷К���:���ζ���{}�I���H�ֿn%�@�L�e��ْ}I�g��SBk�(���n���~��#�4w��w{m�N�xI+svv�� ����A����K�p�R��w�,�7RD���L~�����g�}&��Vlt-X�g_}��7�|C�9L���ܽ{�>rzv�
.�`�p��<+l��`M�݅��tvJY+�Q���m^+�>X� �ӵ1�ô��h[fkb*"�g�W��y7�%���6tE~2E�B�ż� $Z���L*��qg��ay�s�6:C��LG�J���3u=�^��C��ey��0�����'O6��߸<?>::�p\�Od!F�}Xp5�n�R^]��k�q�(�jʈ��Z�Q����㤡��k�K�~#�O�r@�C���b�h9"���jf�!��� C:mp���~m���p����sq]l��nb2�N��O3*���ӣ��_��K��+ʰ��I$u�f�/u�>ftȀ���!6( �9j�DZ|�~�w�<?o�50-遠>�������#!�5$!��q`M��k"�,VrL*Y�fC�LK���^!-�
:�+@�j�{(�=�g�D��靧�GX� ==xҟ���#d�p�pl�m�����|uD7vttrzz��Eh�%M��.֋P��)��7��xm�8 ��!{�.l��,{�"�(XЭ����e`>��	��A-T�Ak����
UFR���� 3��Ng�#�I�b�ۊ���r�A\!]���^$}��M8x���^�|I��c�db���Fە�H5"��V�h9A%$1#ĸ�ݴ ��:��N%mTr䈚̃�o޺u�X�\;	���:-��bٕ�2dgقhE�i˼۳`�x�,K`�.�`P�]��%/��)������d
 �
ఠ;9_'�,�s���ҋ�ra>�`����=���k�,/��^�� �n����cD�����_���:{m���yXd$��II#nNr�Ļ�S��
ڲ�o�d�}�#��X�~��<y��r��%���e�2?�|f�)�O׭���QI�0C���)yz�p
{ssU�J]73������Eߓ�[$nc��-(R�`�-/����$�c�ܭ�5rgVa�0A�љ��ۃ=���Sk��i����`@m���T��aN$ީz-޿%1��u=���U|J�Hk`F[C�X M���T��,%l�o9͠X<�{4�&,%�浂�vY�(~+�(�F�����~���rV֙DM�N��3��L��S7,2'��#qz�d.�Ӻ��Q�u�%'E���[d���Y��W0����4���;)������b�Q�� ��@|����W�"�ċ���&�k����j"�x,)X
R�0#)'Y[`fѧ)�+�~qA��e�t�����ɴ,V���a0 ���1���3CE�m�Vy)V01 m�p�XZ�f�w�������Γ�������j�m���ﯚ�u�QJV��'[�쐉ȇR�\�,��!�:�c�hS2��#�W˺� ���#dyw��� c�o:��L�t��oj�ç���c,ĳ/t����
fܷ�Z*�k�x��(����x��F7��oc���w�{rzNNƲ����j�}�����L8Z�~��=8}����$$�1�k�%v"���b.�u��t[۲VM��8��#�C�8�6�F�9�u"@y3W��N3�	VMK�#�me�`0$=�t��y�c�E.+�:�u[�Ko�oR׹G�5[t�ϖ�0KVM�]\u.�,d*q�P¡sS��Vt ���8LV���HEE����R�m>ъ�����I�,�t<�]+���m%����20N�5v�M�J�l���%>�m�,��%�v�@�*]Q�2���$C�^�d�t�H�bk<���]\��Vqdhx&���rZ��ݽ���f��{Ǔ↡�5UY�I4L�ҳ)�z�h��x?y����p�0w��C`�������
���)2��2=E����V�a�t��-�@V�QH�s1r�.����ʚ>I�q��K�U4dҮ�|���΍�Ch��D��{m JyFG�E�	Г�B�N���[o�s��:Z8Kxy=q:����q���K�l�������\���"%��0�;�t�Ӥjgu��Hz��r��E�.��p�׻D;�����^�`�׼�L�Q��g+f�G�������>�_b ��%�ԭ-$�
8[i$L!>r�R�Y4�&:�2�<��^�x�fd����g?��){�&˒�L,�lwɥ2�����W �VE�@��h����_d���M?�/��A&���q �4����训k����.g����~#��HJY7�=���Ϸ��s3�,�<�t>gO�޽RZґؓͅ\W̷{�w�#�qv��j�5�Z�Đ�:��#Wr ��Xf�လ�q����Ѻg^ZB�<0ڧ��4�b7�2t.r�_Z�Dg)�։�����ZZUK��,N�O���_jS3\�����S��vl��U�5g�-&���#\�w��vJMnH�Q�b%N�6J)�O�L��" �r�Bi׹.-�Ϟ<����]��]��ǯG���My*��Ӈ|
q�&z�	�q��e�/���U���#rW�H��8n��a�_Y���H�T:-���� 2�Y�O>Veb_I[,Z����q�R;�S���'R���J;�W�Z6�������&ƥ/ -���A ~�_V������sRh�����d���pokL[�U-]`$ڔŢ\��3�N�-��G��t����g����.����%4�����Er|o���VC�]v���Y��]�{D�HW�Hz�b@Ա���:j )�gϞ]�|n/B3>+�7ju��-@۲D\����O����x��T&��_��[;��O��`�`�j���	�G�u�ʥӓ3A5���05գ�%H����gu�=����u�nG�^��S��],�BZ5�zw�,"��8� f�!M!�@"�`*�p�2��R����7�+�[�ĠE����m��.�f.N��}�q�:�������O�>}����_ޕ`q�^r��4���飇_a/�r�7 "F�H0�^�v��
w����9�X���!&f៵Ώ2�i�N���E!���L��\��_�p���r�գ����w�>ʵ���<vbPK���v�v�I��!��Vk�eSNd�0 ��8 Q�� 8�81#4(�x�M�.6�S�gr��E� q(�=����]:�8n��H�-C�T��Naϩ�IPQˏ��&S;�WXT@ngkn{�},5��8 �(��-�d��7)�cyq��wCJ��YLE�`��6y5|1k�7�j�ilP�b��� OWj���0X�2Z���Q���VU:�����F�z�2L�Ӕ|�@��I�t�Ç��+�"{�إ0_�g�P��Y:z�n����1:��"h(���[�)����N	�h�5G�h�޶\��ePF���!��k�-$2<�ݪ���F��̛dP;��İ$�mL��Nc��l�#�˞��4�b�1�>n�w��)�6���8��Ng�'������ZD�'���4i�4�W��8�u'�m���^�r��Ch]��P(v��4�,��t�f���+�R�8!#����ÜG͜srA�G����Q	�`��� �P.�!1�'�܆Y~��@H��-��hx��*$��@##�k�R;Y�-z:p���H�, m��,�X���WQ� m$�Vh�����ݬ:%����t+hS��)F�g*� �CBONnJ�0:��a>C�K����`e|c�d	�D�(t��w"属��vi�L� ��hf����/H#C��� ������'auj�q��@ɟ�"�b1�f��0�Ma�4�����N����?޾�&*��4��e%u�kj.eT�P�L_ֈ<j�7�Fcfw_��h'��֢�����P���F���C�Uñk:�����4"�6t+��[X���Ϲ�n�"��tS��>5�E��d��&����"-LY��?�B�Ow���m��
���E���|$��G���Q=h����͞聂������a/���^,�"*�ONN9\X�ql8,��f�R5�U� �Yj��٠���~�D�Ù� �E�`�/����)���t{/^� ���B�[V�棋���~�<$w��u�ϒCf[�Ήcu�xW|��5�J���G/Ϩ\r*%�x�!8^3�	 ��=�բ��J]�W���CL
ʌ2$�i��\8�RF6��w�"Wf��ڂ4�&�F�S�HߘزR�l =�����p���V��:�ʌ��o�EM/b��b"=n8��Sf�s��M�R�g���-��ņ�!�)ɓ�!`�-�V�,�i,��A��`�!�xSJ���� ۊ��cV)Hm�)�@ĳ��˚j����͠|؆S�V�c�
�\r�c.���E:����������>::Ɏpϳ�C�D��䍎	��(假���"]���8[,��GЦ��	��]_Ʉ��y�{���|I�S��>�J2e���	_�H��9e��+�����̢���0��(q�9'��bF�a��'������Zy���m�3����w�2��il1f��^Ç���� H|-��deN����`:���D���\�b��=��6v%�%܏���kTƕ%�<'�:5{�ٔU*����  �.�Lz���L���<sR8-ؠ��r��Z��98^�SZH�^|6���i2�/^�h��u*�!��+:��0w�M���^S/"N� �2U̓��c:ӆ���<͐Jԡ^��NXz�K�4)ӛ�4Đi�c���M�
������.��@W@� '�?���$E��M�0�d�*Ho�9��4aD��v�.��� ��@MV�h.	l�j�x��������~���nb�(A2�b��[�
>��JX#�]��yt�R�����)s$���2���m��_� ��Α���x��e�����x��i�$Jxg\�p۶�J���G�0��-O�!�z���9�Y�]��'�W8�����N��t&�������7�C�Wrpp #��L���i���0%"ϩ�٬'P.� �Ѵd���1@H�ǎ�f����#�o�y��m��_|�8=�����p\@0L�Z��q�W'~G���Z85&~�T<�?YY���*èl)t����Q�����.EK�捪:��QJ�q�g�ɇ�fO�[Aᰙ*�Z��W,��-�Y@�V�@�pn0W
�x�@���u�����5�m��>"�کQ+��*�0�I��A��J)��7q��-$?p� ��nv��FN�X%���FB��W:�z7�!�_�&�MwK�|�0�ڞ%ON7�L$<&��(U�&��4��J�B#�V���ɍpvq�~���W�EC���&R\�J�p-�����ϛB'1�:ώ����Dp���8�!.4Ț�%f�rU�$
O=�́t���ൕW��d���$7"K 2Q�\�I�d�y3�BKSW�����x.�i��{N�9+�S&�dz-��<�o�lD�0�����ʅ�If	
QE{dK��ǟ�]��X�^��cM�����3�rĕ�U��$�� �@6���h��-'mB�|Ɔ�^}�:�e��ts&�!�2�)�	���<��c��ĭ.I�P��!TO8e!5��
l4>�/퀔�#1ŵWd�N�M�J�,F���� ��_H�Ю�^���`���$��DBJ)�����g''�@K�u$Q8���4|z��$��)eV�K&�g�f�.;��BL��D�6.ΖE��X�����>LJ�P�W�0�����oC��!eF'��
�� �Q��z�~U^]ZE���$�.t�̦��7H-+��3ޮ�s����/Vˤ�a(wq���3���t�1���Cˁ��[c�MDM�V~��O�z}��]^=�B��;�J�P�7�*1�>[.~,x���sM��o����䐍-K>�_.�_}��iQ9)��\��f��Ч��R�����iK�����d'�RӉTF�ℇ]�U3�ma���9�cC+�-�-:r5n��|�u��u�˾��+��;䭉ɵC��c£����km�l����lqVh�ݗ�_��'g��A��]GM�*C��3���R^��(%,I���C�K�=&b���m��R�"=#8�[E�E�'"��>���J20
��r�A;����Vr�"֩Ԅ����J�(�+&B>9�PiQV�-�B̠?��2��B�:�h���]�t������0,�
�	����h1-a�w�9���x��� ����� �b���;7Q{(�0�o���UB�e���)�6��|Tf�A�-��F`��a�1/K������l��*V�4m6�ò��煞"%o���PI���0��<W9����'�r,���P�̭�dp��&Mm�2��TY&�$d�iI0�?>љ�|�-"����&)�ub��LkR�d���׮L�\�-~��1�73�O>������Dţ{+�n-y7c�5����2�����L��ԁ��k��B�5Ȭ3�WR���^$S�h3$2�y�U�cbu�}�
�%��&���bqJZ�W���W��n���CΎ̘"#�z��
��×�O�Bcfj"w��_�z-�u�s�@�'�z|J�j7#���M6�Q�T��fk�`�b�`>$:_���� ,	�YV��&��NU�A���D,ȘZt�,7��k_�![�����J�E����\�Tw���*�A��<��r ���O�/��K�r�m�[���,z�t�rE��.�N�*��U�<�h�7� 3J�#��2+��F��յ,Z)t)䌅�A.�C��Ԥ<�s��:+IÅ<�R�6Z
s"����X
�Ĥ�J��)���kߜ�љ�R��rѺ3W7Y
%q���#F�h`�%t��^��� �$?R@�Vu#���w\�ھC�
s�2�e���(X�E&.���՘�m�ۋ����+Wmw||���O.�6zDn����0$D!]�v����)g��^7���J5�ȴ�,޴��!:`�"
�-�6�I`t�؃E�N�^�t��իW��Zf���ģP�
��^h"	u��0��n������}˵��	QB�}6%���u�/_���y�Z��E�~cҺ��] ��+\���2��)����Ѳ���;�b�&M%�z��0 K�Y�2����xt|�0)�Uw$���5s/��0V��l��rM�q	S�����i�·��τ�o�`�׮[2Ut�ϟ?��
�b��������@G0$R�hF��99�׮]���j��!�ҕR4\Ef���f��dtW`�	B�H��z��������6�%l����T��B�8�v�Qt��L&:ټ�@����5��.�·&�ZMM@e���v�[_w�l����q�PI'Y X�	T	�b:�2a(;߱���R(vxd��x�� ��^�	��#�t��!+_h�a#���2j��d��fM����@����*3�b����CBX�nk���	�R��bjx�׭���!O��i��M3s����lj�U�I�z�zv�Zb��G*�V���=�XjQ}����[k�$�����Ի�oڀME�26���@�X��l��X�
���d�-�T�0���C���c/�]��X�Ko��$��O�i�� �)]z����#a����h^��A�ɵ6�G�)��oԎQg3�ԝHR�� ��э[Gt�=���~c��_�C]�YVDs�
t�	��{��!��"%�Y]���lop��8�Q�e`�[�(�)`�Rx5эf�|�����lצ�e���4�b�4Ӥ�\���7;5_4�\J�)_+-���	�4�[h�k��k��Шtf�,��T:z������a�=Xz���f�Ō	V�932���?�����e�v|w:�<^	�6��Q�r.f�u��	��x��%F��M���,��
'�L���դ��35R(���]b�D�r!)Qa�$wK�+5��v	�<�j�ߞ�������Ф�p �ڌ)m�a���$��LytID�h�Gn��֑�����k3p|�ڈ�ե�ʩ�\��� ��t�+V���Q��kS~��I`�p��Z��k�c.�q������W��_�<�{��j�_b�FnN�	+�¬d/�Ѧs�F٬��
Dp���M�E!-y�ԋ*����W"� ��N9˽Ҫ�:% �PŹ+|r-�_�P/��dƸ�u���h�|�ŋi�?���"��!��k�6;��2�=�0�FT�k�`"���ie�����$�!��
�吪Q`ȑ]����d��I���L+��Q�eFm#2��n���^+� ��Q!��L���jh>w��5;-���W�^��?�3R�?��G�[��V��k�=�'씜�Υ�ˆ>o�D��O�1�fbr��e��Q��:Ak'c�>=�Ɨzi4�X-�K���d/��Kc�{��^�$������.�&0^GR�p� �!��3�k���E+�I��ǾME4	R���>	�Dz:z4�8=�DPm�V�n�e�_8�:�i�����`�Y�
Z R�����aTʞ���"��+��à4�� ��J��F���ݬN;!J��O!&�
�L��^'�Yj�N4�-�t�R ږ����4���n�8[�J��n$W�P
=J����c�������׃��W�I��jD0�N�>XeM0>�>�U-�Չ/���zK��Z��g윶����H^�#i����B�MD�W|ݠ���s��	�r����!o����6`;	m�ȑ=f�O3�|�����'��ħ�U�����˧����/`c+W�`{�Emp/����|����|ct��A2�[�@�S_HG[k��X��l��t}�QVY��\	Ӳ񟀮�]Xs�|�/^ �D_M61{�86Qg��PVJcD��O�_��2��y9���(�Y.��d�E P)���f*f����	����w�����Ȋ-��A���q�u��!�ܡ�����`!N4¡�da��#' �Cn�������'�������# m�\WJ�n-\tZ���^��� Q�#�۝��W�˶��Aק͢o�1�;;�_�Ii��(n���?��LŮ%�M�u�V�<�(�[,VVo1���H;\��AI��hZv ]*+KS��� k���Q�:r����,󣁈�R#� �6��B�
�N�H�^j��0���Bb��ԧ�~�+������紀�hL؍�-m<Gw��'��ѱP/��qgυ�����º�zj;�x(�P��r�,��Ʊ����7qCL��O��4�\��̦\�E����DE��A���BFM�i�R�E:=���w��ר�9p=ꌆ�k�Ô������T��4I�m��sY��'z��uZ̺��z���PY�� ���������:
)j�uP�G�C�p�*�X(5=���cㆰ�����#�u��?[��͑U6�$*��Z�s�9-bf��cB��A�Vj`�-m~D]ML�`��Qk�.Bw�+��n"P������۷-�$%��_��x���/�H�S]ȢB�!#����'g� �l�����}��$ȌS·;�_]��.qF~-!�Y����S�	������ze��`��G�t����d��`�ʂ2J3�]U����W�a:����g�1 Gk��V6A� ��q2EER���ri���+��A��D�U�����_gf���}l&J $���kθvI"M3�Ύ�K�͢�`�5jYd,�A�u,:�J)�N=��v�v�&���ʫ�p9]`z	��	L��V��><ܸ��ha6�L'l*�u;y��+��/�k��)�
(���S����ږI^L'r�>�X�4 �2��Е����OgzFz����:Řʠh�fS�:��*��6.PH{h@$I�,ݛ�����~���x3�k.2-.�臶k���X�pJv��z[<%���H.r���
��bYmz�d[�8	����3%��`�8��ѧd��Z<e�I%�C���pC��'x�?�5K�N���A���u�ۑ�[P�����Q�T�(p�����ل�}��DZo�\��t�xD��ێ��b-��U������=����(Oq�v|�kLM�2�)�'�^�C�'��0����N�T�`�C�Sy1r���GG�RI��N(@_� �%0�1kg�G�
2��+��>�U��dٮۗ/�n���]��z<
��].*嬍d�0��4���ڞ�,K�p����f���Dщ	X���ȣo�ˊ���|�E����5��2��""�Q����iา��	��J�%I��&yD/��I�RP�B�(s�\ =2�T"N��@$�f��{���m�t��"8�Rֆ�;j�ޡKH������d*&��`�Fj�x$������ϧO���?��emŀ��G�.�Q6������&s���S =�5�p	v�:�e�������Q���V��iz�g9{R�w�O�5��S�"z�[D�����K����"0�*���C|9�3�����pB!1ɇ�`���HOŔG9�k��^+��6��u���ѪO_z��X�q�2p��&$�(�B�U�Ao\��KL�Hf��pc����f�f�m�Z��9)�®&��32�0)��|5�DT.�}��	1X(��
�Π!��ةJ�����̱Iu��Ͳ4������KQASJEo1\s���ҘtSH��U�o��\� e���88�%�p�|���g���D��_��k�#�F�ܿ���?���Qp)�`3�UM"�D�iU��Z�t�����5j�p�ش�d(I2%�¡(���dRfJ"�����k���!+
�p�s߾�i�Q�K-�[e��A�ք~6�j���Eәfs]�e�a��$���\zv�3�S�G��q��L�D^W'g��6��c@iFJfp\���c�>�cIj�_��wsH��<�*�����	*z���g�Ke�'`0�	��<{�vp�x��Q��
��s�A������ڊ�#�#ꇠH]����S� �>�`;���|{+
��������'�;�s��1<)�!�XOf�x\>��lh��"m�TC�E�M��;�>p�X�Қ��)l��-�8�f���ݻpp�{�]�6';�9w�W�����]�;��{��0V�z�7Ѫ�#Mށ���,Ϡ� ��$B�S���lqt$o����[�H$��0U�VT��]�{BW�5�_��`B1��S��� �BP�t��7oҥ�_�&� �s��u2߁���ً�[;�\�W�l$�:�]`�!����ׯZ�S�%*�1B�B.�z��",���
��V�rx�sJ�J��R�r�S.x��~����Nf-���Ś����Z�����;�KK�f���y筛� A�q��ҍݻws�r3W�hf9�Ӝ%�		�UZ�����:����'�<x�����������;Ykb5�i3A�.}��C�/��u�t?�����2�'��a�
� hA\�g���S����`(:��Ԡ�3Eӵ`|�Z���`7L^?&M����1�r�#!��u��YS��݀��-4:��.g� j�l���5[$�@2D�e�=�Q
.��H��v	<9�"��1x���BY�)R���lG�M�/�i����KE��������*h�6ԢkCϋP,b���j�&��1"WRNo�϶�&�E�^IuQ���jd��-���*WqD�1�_k���!��峜1����\�f��qk b����]���V3��k*��to�և��A�z�<����H�܄M���:}lZoZ�j�I3�&U" Am�����cG��9<jaX0�WtZ�� ��4��J��=�Wr5��m'ĸ�{ό��J���������z0��4�8h�T����f��I\�惙��zr�_�K� `b����G;�F
��L�,o���(��y������z͙[!I�@�ӱ��c��R@��2�`�K� US��&=Rh>$��u=�Z,\H�J�L&�cz�%��� QKb��Z{�W�p�顙��M&������R�(;�
���R�q��N劘
�8 "��a�#��F�ŝ��xaq��2�~Wh77���-u�'��C�P�F�׶[Sq%>cړ�Q 2oM�9I4��y�����:g�I9�Fi��	x����?�EhR�����N�0R��Q���m���~;w!�Y��t�qx���H���a�I�:�$4�� mAb{��j�����ꂹ��*�7ѓ�\f�}aG�8�/g�L����ET�p�T�/Յ�O,�c��W^�t��;���KϠ��a�c���2����W)�$�� ��n&��!Ba�7���\���Å���ح7+���s;}8h�&�Qh��m��6+��
�n�3�90�����XR�o,l�<!l�L:�T��ȓ6�;A�ǎ��l-�Nڦ���m^Զ�Q�~���9��	�No��/��̙�+���]��o���w�����G�}���mħ�>|��������m*t�P&�V����5TB
-j���2;\^���)��T�C��?<<�\��˻,*QRY �굅ܠ�Io�� Q� ��O7�>gS8}"|�#�F��l��FK�X���o@W�HJ���6ў���_�6���qFMH������N��	��q�qe�"�NU6gk�%�h��qTVi��`N�n�N��ǝ�2B:%�����'��n#��@���Ӹy���M�(��YH���Y��h�8�"W�L�"MQ��2�p�!������_�
L*�|����E��c�ra�^�7��Y^��b���SٹbL�R��Fm�Zxk�����	N�z��7�5O�
[o�b�q�� ��G�8A;!:%�,��"j��DE0�+�.W���5���ך� ̳��ߓ}Y_��q-q��Um�2��&R��!��sB�*Ȁ��$����O?�t{k�����V�T'ѐT�4�9-���i��R�7D�0���'״R�1'p��	x���hE�M�'+���-����=�x~
�����<��m*H��-Z���=`@-��l:&4ƨ�n���ꅄ�6�J� �K&2��^�06�'�N�0���%��7n\�|y���|W+ڒ^g��#N�nɏ���5@'L�)ީ/f�����Y)��9Aht@��Щ Q�J(�~�:]��
ކ�X�� F�4M$�'��3�$x^��P�p�pP�COL;~�޽���x���K�92^��M-s$��5��R�ة'��$��0�!�B^ћ1M�/��,њ��*�K�2[a�a�y�x�B�)�����k(���t�to��-����͛V>L�}r��q�2��1�ZJ��,���h$3�#W�\��{�������?|���G}����?��Oq<�Iz_>��Z�T��CېЋ�^�jt�tjhS�S���APWa��5����赫,w�a��nb�,Qjl�=�¡�i�k�SԹ�
�G}%�� ���{5~$�[�JIsң���묫2J��R��� 6 4�!N�0h����F�5�:�kIt|�Os>[��}4;"_��f��A{%�4!��i��N�(VV�)������cpU� �A	"���]�p�N�q��
���2��A]6R"j�Ƭ��n����ۇ���>��9P,�.�Cg�.���%��l`ma�R�k�z��}��3�7�f��Y�h�Y�ֹ�СC*jK�G��6���I��t`��Z{i%��ll��*��Ͱ8�9"�w�l?�J���۲��M`�;��A;���l�!��%��k���Y�7f��&����t��xS��0�G���=���,c��.�,���l�a2��A�����:�,�m�S�F-�J�A��ͅ
�.
F�ʊU�$�����I�z�orp�d<��Eaa#��씮K��֕��/ �,�±�a��!����d`z~Q�,F s<��;�x��Eg<�f��l��&��5��n�ϲM��F�z��9�~��%VN=Q���3�`M���n⃤������:Y��U;iJz��^��
��R�L^za�$�Z����}�UPId��7sx�h4	��%})d������F�E�>���I�Ac7��IPI����"{��f�B�������mߥڟ��?���ס��b�[�gzw����z�����5d��x�ѐ:~��9��˗8�Ұ���fN�Œ�����@�����dͅ�>��D�~%��tS��.ܗ^Z�թ]�W.\�G�-��_��@��B*��8�ic�ҧ���4I�v�����Y�?�<yb�QS����+m���o�~�u���7��護�y��9&b��π45$�����j��c�@۠Ul|/�_�"b>�%���p:��II�'0�Ѵ� �%����lMjgL�0(�+|8Z��ܐ���V)a^�*����հ�6���@N���Ж���`�)B�h��0���7�1�U�.\,#:� .��/�3��W_jwٜu�E�,4OS�z�@�sP�A^b!}��' %t�C4{�E��YX�R2 KK��$��d��H�rQ��~��SW������o���X'�(6EB�#	���>���_~��:��O�@���U���D��^k严Д�ućl2��֜f��tr-�5�d�7i����}ǒfPNǋ��N�<��S�Yљ�����TՄ[J��XU��\�be����C�W+p��q@���#�����qH���U�A�F��?��&e%s�;i��ݛԩ��ɐR�Ζ���zXM�� �Q��6Bޏ�30U���-+>H� �Y��\,��-��Y�MQǦ$Ў���3Ԉ9C�����b94��E6�:8��1��^��rI���}���LO�� F+_��Z;�V��͘4��5�����c6��a%�ᳱ�Q���hM�� 9i�]�Y�G�j�^��E�^I!}�YHלj�xI�#�HK�-���J��ʕ+�9/\�p��}�����ַ���'��:9����/޼y��aZ.F&.����>'HFW&MNWCȣ�������l��,i�!�]D�c�3�Ki�.%�J�ٝM�d@�	-����%y��9��������W��S�����{���'�	f,V�f:���gJ좚o����w@![++v��Hg*�Ԭ�xy���6�V�`I-)�6��ʃ9$j��6�8<䑯���ׯcV=Θ�=�I4=I�H���>���.H��o����f!���=�"sv'��x�"y3Pk�������Z���r?lgWݺR���3I2���׍��+�j���a� �̶͠�˺�'�tk�Գ�\�Dв�q��صh�"?�������L&ǀ@��!c�r8�A[ ��p����<x��g;;W�V�W��������ϋ�8�� R`f�����-�HBK+I{��1ǀ�VU��g:�Eq���<w������Q�Y��a���=��Յ�����[�#`��Q��Ȱ�y��q���P��	)GX)�����X�k�� ��CE��4ցM�S�h�7H9j�&�ӠN8�r��C��;�*�j�2��D�#M���a,��t��qL3��� 7}3"���9V�B[�z��3��0���>���i�C���]� *9�?��1��5�*m_�Ē�Zyu֓�8(K��5��� m`qDQ��Z�t):d�|�}?���礩�%���->�d���N���d�f@��K����2!X�GӢn�)3(iP�4�R��2+f��"��[
�`�UI��v�QHU�U�C�pDk^Wm<����?��B�^���A�0mԌ_ԑ�P"��d0"Z?�6h���cn	l׭�aP&�Q���^�ץ��^�j��U(B��Z���J�hr)�.�,h�a~���QzM@v͵���mkL���F/%o1B��).|v֞��^FI�F[�	3�9����G?\��+ͷ�Qom�n���֧7k=3��f,p2QwjWn�A���Ơ�
,tf.�H�/�4n6-Fq	H��{xv�Ɇ�lly�z~#*�%dӓvj��~�*i���X(��%��v�^�������o]��e!I#y tH�j"�h[�et	\"_G��	19&�X;���O����/���-�J�I6"uf"��]��Lյ���_���1m�My����D�B�9:1��R�B��CJxnH͛]��H�?|�&���ޝӳ߹s����K�S$1��l)u|�{X;��-����O�۽�A��l�RNk+��Ax�"o���Y����K>��V�4S�B�|���������7����:�qJ�Z{�ǌ}�L���l��+����m�n�~�CoJ�� ��z&(���tJ�HJ���xp]*B$�P��cA�*#؂������k2 ?�����"�uX_gi!0@C�6�H�Y*Ȟ�e����.j"��r3�uQ���Ə�t�1 ����� ×I<t|�9�O:�B���t`7���D��u�����63R�J���A��F�{�9,�=��(��A��d���1��J"��`#]W��u�����cb�OQT* G$=���gbVt ��)����ARs�!��C�v��1��h^���! o����<)e���,C�L����"�J'6�Bzed����#��Sʰ2k�5���bj�D?��e��J{|��hL�^��7��u���f�Z�u�+����
ʉf� ��[#C�
!�C��%E���H���3�K��8�c^�i�@��A>��o�R�+�l|0�,-�6D�Zܶ렭'��{�A�{�!�Ѧ��e�6��׼,I�u}��n���I�A#fQ3.�ߠmB��O���t����QS�9l6Ցۣ�q1>>+�曬6A7���|+�?�	��޽{'��CV�BV�C̅�O3�Y�M�u�mϼc��{8S�g��tB鳰���ٴ�"���)|��pj�c�"7���7n6���*E,_e��������zR(�=��/%C#�<ܺu�����������g���˿���_����]����}��ݻ�����^ �F�@/A� k�+�!��a]S����������8���*����:��n�>��U��a���ӧ_|�})Y�;w����vt.<:B�ԯ�ʒ�@�PM�$+������@�?z�S�����_~	(�k8V��Y��ҷ���D���B�|@#!�E1���_��sl��M-���ُ�<a8:a������_�>���r�%�0��Db�Ü�4N��Ы��wk�]�v\5e�2=�$���r6���=S�d�p�lƢ2�� ���o���#���$�!��!��T�,tm�hi�a�I�:V F����7��D~�T��'�|����$��aÊ ��Tb�V-�D_D�B1j-aC�w�$�ϟ[@Î�A�Jy����A���f�����h���7�q��f��@`��옷C&�8)I�b���m���z�.�%�߄�a@1*���^T*R&D�J�̸C�,@�V���:��pr�H���G��(�^	�k���� �$�WBO�y�|o ��7G�l��I,ս���"���	�`|ny�XOܟ)����6����K-�1���R�!��Q3*t���j��`8j���TU�ހ팱�� �b:l����r2)j�s�����RP�mz�M�
%�w��У.	;A�4��<7;T.�
&(_��_��ۅ��9u`�a�0�
Ŝ��$�Vj��׆ݰ��`�s�^_g9h�0�"k�65�w��W$���XRX,�R+�.u�l�9'`�b"��Bg��t�==S��-�	Yߘe�Gm�ɇa���؂Fg2zm 7H�5��4�셩�􈣑f��N_��\�7�v�*��a��"����mOJiYmW=FW�.�S���`ލE��<t =���Ï��t"A"uL�gҙ���a|$� �-	���}���Yr݅����S��ha:�@��J�\����!B�]�d�
FB��h��,���o���pk���{~���^�a����V0�^A�2�����×/_�2	޲�'RpD�ĄM�M��!���4��͢��[S�8.���ۻt,���ߧG&hH��w<LM-	s͵�����yh�/J89a�#�jp�Z�[��B��A��-��Hso�B��?��A ��vq�ڵ;�ߤ��U���Mj�H�_L�]�>�'2�ҋZ(*�k-R#�U+�8�y�d���ZI���u;z����������`�zuD��(�'�>��SZ��g��K5��8$$�4�3hM�1`��4]FFT�t��[��AX��َ�B3t)غ��f��Z�!��cII˃�<�H��d��	!l��^�0ى���J��\V�mNf�3�,\�5kqF["s�P�Fo�Y�e���t�K�PŨ�J�Թ[�O-�����<�g�C�fd!��u��={������������X
��v���X��]k�UQǠ؍G�V�t;�h��܉�&��a2:�g ��3��ܢQXg[�R+�RA]m�Z��H/�>=e/7YЉ	~�J��7��pZ�`T�&q���CN����������Y?���`�6z����I�I��`�a+����n8�tX��>�&4��jq��c��L� 豜ԓ"�W+Y5�Z+c�'3s����6�Pk�A.���'���6���iQ�b�'�r�n���=����*?~v�ؖ\v��x�|���垹ě�7�����j>���ByL_�P����As��\E�0i�p���?��R�U���i�<D5JU"�2.�F�Vv���ɢ%�~�R,Ka����t����u�h�5�l�&!.�v��|68����e��1���G8L@�9��Qc�&�Q�|v0�L���K�$�p I1];
�vP����Z���	Qli5�LB�ٌC����2�C�a�?*\���yf�D�p�����K�-%l�������3��xT��`!�TEmDe�����x�0g�e����3�XC����ղ5�rQx�/�_��+=�G�r��w�Y�:����˟���ً����;:9�/��7$����;wH;��DWZZ @(�P������ɣGO�S<����(��%K�
�-����C$sie��Z�o�4��U�bya8��O�H���|ZO/���;t\{~�����o!����1�e���������)�����pv��J�������'�L�a"?m�*3������}]��h7F�` ;J�Ȳ8}֓���.�o�q�ƍA��am��`P�o�o@��|[�,\���3?�-�ij�纼�N�?"��%P��w��W\�L:5��^mfS<��FE%j`��ܳa�h�a�����-����ִ
�0 Ӛ����  p7�/_�L;@�D�}��9LqE�G��`��~��ds�޽�����~��_��%Rr��ܚ����7�6l7���۷�>I0�	�Q��zE6��g ��a^����Qi���f��?���׉��yv6-Y·nW�SL�Jחb�m��wg�J��a��3��z�f�-<�4�Q�\���ISeO��:�s�ܒ%��C䉣�F|ȲM��w��:�`P	�ByB0*�������3�A����"k�,��>r>�[�5���g�!���2�O�8#���d�E��@M*�hs]2S�Q,d!�z�f0Y/&�!��Ec�����'a$M�ڷ4h��($�m��eR�G"�1�7CAquu�|j���u��a�*�¦T���|;Am��$sVa�`��A�!��<W4�*b�֕���-�O�H��o�������-��џeG1e��O�l����0z^21�UI谴��@C�(�y�Q���� ��F��@"m@���~cg0_zN��0_��]���;=�M`�`HFm)5�4�nx���y�Pl��0��JP�i��R� �(�,��b��р��H�1].1j�8�$����G���&����
Ћ'G/ql
b�׮]#ӂ��bQXs�����0�t�ر�(����Co�4��u�De��a���t���ַp��j (atճ��ۿ�ۇ�"
��?d�T�ATI��a�������iׅ�7/���?�u��!��!'���ei��R�z�����;� %���[~x��B�A����:x��fY�42��V�1���l�E����H>y��������{ JJ;)Nfr���������1E6+�k\[���d�._~�������/��C[���V��@o�a�T�E���J���Bc!>�����i��4
�F'�cLu�h�kp�a�̾2ql��>����i�R�]�}����������t�i����<rb�5��ˢ&kt�J�f���B�cF�5jͯ����x����6X�8�υK��99�_��O��7�n� E^f��6P����om��)�We�j��	�ZcOS�؏��3Ԃ����(U�)i�g�p�N����H1*Y���B�fg�K��8MН�=���l�����G�x�W�pJ��� ���?&���5�G�"pP����^)�qkiu�};BZ�ޚ4����$<I2�tY��t��ڃB%��l�v�wgԜ*?~��
�9������FW��r��n��KK�q����6pqQ�nP N:F�Nm���Z�.�]���7"��G"��}���n��^;G��씘�^$@����H��|�L����:&��He�a%�ExXU���K��$�������*�0.e� ���]l�F'$\�bx@�H�4�6�����-@�h�~�!��&	,t���q�c`���p��t����'����"�-����Ծ��k��|П����#��P��\`r2�D�l����B����Ӫ�8Y;^�h�^2^��u��28#h.��E7�m���%�!�M��8g�b6�&�K�/��5ةFI��,MϓTTJ�]���fT:m�2'@3�Q����o�R��F�5�+k.0���f�����>� ���j���իW	�q���%��NE�xfS�������=J"�����ܔ6��rNKJs�5��"^�}����	�ܿ��E���	1���~��<}��ѣG�e����7�XƇ~Hw����D��s�*zp�&t��>|$�=V�7o����3����Q*<oǲ]Ia;[�fZ#��53u��^Jc8e�X�Is��毥�*�(S��y@����G�Sг ��rq�d2�Sw��(q��J��ć��PD�E�/]���¤������<S� m��B�2�F`�i#`H_�Jb����!����R%�L����iumH��c4B��BF�\Jfg�S��ٻ<K��lI�Fy>c�^��k�
7��f�J�� #��J��fQ�~ʺ7�D8��ʘF$;�� ��W%s��^JQ	�p�(�e$	�=y��!� 9#�pE@�m��@�W�l6.�����w�x��O�ݻ��/�'���$��z�F(e��i��@%~�����NKM�J�\H�9៨=.0[p�K-Zʽu��M����D-T%�.�
��r�R)1�M���' ��gl�?�Oi9 �)�� Ϥ� ���8P��sL����c2����:L*pV�k_*.O�I]8��E�2�lP��c�i0�Q���P�}�OK�u�����m(q:����u�/E�H���8d�RQU`�!c�ơv��O ����4Mn�	�V�FL,�a ��Je6�X+�B�6�gӟm1}��x�w4NR���)ю�F��j䲮D�2[��<'�C��W��#�/�:�����U=�Ŵmm������O"�Vҳ\�?}�M��)2�LH�K�)��8�Ԙ�8`1��2�W�*.��[�9],�&�Z*��\5�d��qz��"G����y�X�cH!]�%	$�(���56�g�V�mqF��LVFk��i����J���+9oky[���xC�L�^	�A�C�F->2�d�7j�:H��&y�1�5�+��yz�P�n1Y�s�6��h�_�N��:�ܴ.�^�L����o~��X�������ׯ_߿�''͓,�hҲ�y��i�(8<�E�췦s+������^���s�J{d;))��e͞	��1�у�\u�s��{_�-~N+XQv�w#��o�<���������^;�����������?	�������1ջ�ex�p>'R�O�ϓ^����S��@�Y.W����O������������-Rܜ��82(󚡣�n����LJ��@�Gr>���F�a{�m�i+]X_Xbq/��y�%-vC)�"ۻ��aܞN��шݰ%~2٬�;�S�L���q�ʥ�؈�w�=}�
�L�]G'���%!P��(?�B�4G�c�

�Lg�]�{���o~�G��	F�9f�0�I�Ij�ī���4u�~��o[�y���UB�':�f&H�AR���8�C/�/��q��;�+��%{ƭ��}c_H i�1�S�p98٫�ƶ[�>L��;�mB{��?�����y=t�k�	�8�gR�B:;ڡ��>�O:i����:[r�)��>*��΅��o3��eS�;'���:R�а�p�y G�*pp�g�4����r>O2�'+�mp��y�(���8�'�D��!�;�ņ�1�2f�X���@!Vh`�hW  F�$�G�S��B^I/����A��_��+��]]�ۡ��ݽHȕ�����I�	c����D�|��ݻw�0�)(�w<�$
>/Lf��n�m!B�[��e�"!�wd�}��8�An��������8�&�����Bx��6�;������:2�&�|=:[.�u !$q��4.�z�H��C:��8�I���D|Q�=�tP���,N�e�9�����B�z��m�}��EE¾x�7.^$р�����sS��l�Dx��|	XCz��p{gvڲ�5s5;�+KD�N�Kz����;���!u��C��� s!�V����<�dq(��V��=8=�g�8n��1TB�	#h�a*�*-��d�l!M¡��!i�>=/]\0Z6�ax@�2 �n��zy�i��N=`�|0��;�	@�܅Д��M�{[;��-)��*t�:������ĕ߬�	���E� ^�#�K)&~S����B�8�I����8��u[X�[Jǹ�SKQ"o�N;bc6�痰���
�l�K	ވ�߶M5촇���S*�B��frA)	e6�4�a��-6�dđ�OU1��bq��HN�L�裓�حv�j~vƕh����CY�]�)�_T��{�
��q�&ܲv�9^,��x��rg~�.�H���	;Q+-�q\���P`�H3�� X�쪐w�J�����r����e\J]E��O�,!,>��c��z6�z�����	����n��Ɲ��'-�����w.��᷿#g�c�Rtq���g���O�Q�q��/?��sQ�b��>{��=#�t�ֵ/�\u/�e=z�p�t�b�
F����'o=�}�6��^$�F���L��U�쫇�o$lI����g��%�������W�	�]�z���^j�?1�]����e�fW�|Ƃ9OOφ0�*����t#a<z����	u��Ѡ�~�34Ȱ`��J���,���!J�2;;�Z�X�t}��t��8\�r�.e.^�+�V�W[�����B+�!��h/N�18M���������f�&���{Ƒt?\�p����I�6������/����Uɢu:�4�Wp�i��w��*�^X�*���}�YmR���z�|�l������]��F�������i�5�E@�Hw���K2�@�\�7��tWg+�<H\��6��]:��zN��q��B?vQ��5ui~��_���};����߃=���F�A��a� 2���2Z�9A)$	$:��`���[�,*�(6��ў@NP%%,�=�S�6��'��Zjúɻ��	�L������H�q�l	|K+3r�
>{!�1ʃ�fB�v��&���z����U���h�P��(�����D�CY��;"����rA�TE�yk�6��9W�F7�i��$.N��TnZܚo�y��x ��tiS��P��!�^X�YՎ�����	�1���J£R6�UoNJ��pa{g�'炖����:;A5y�8_����[d&���$�4�������%�pْLh]n�m�`�H�a�s�:zO+��B��!�t���w�^WI�X?ȋs���}��n�c<Iٓ�"K>��^��5i'��d���!KI��Y�[�[o�I��VR7��3�=1� `��C�Ya�
�M
��q��4B��?e�v zN+Hi4�~���3pYK�-T���4��U�|5DmН1ל�5|^j��0A�V�"vZ�	t�j�R�t�2j -�(Ʃ��o��y��uHGټ��I`|��,�noC\��*�j-��r�_P>�Y(���.�@.���Q�Ҥoɇ!��ƿ��^�v͕��5\p�=ߒ��O��|H|���)�D7�/O����c�� �'� M�����>�Y���|�:�?�&���q
3�X���Y���n�_�N�c�4&�����~�/��/����z�n�tP��(zYFVm�����%�	m&)vϜA�w����������7�Ď�J|�6�ep���L:��Q �R��@Ƭ� ��Cs��K����1Q�rVmg��s,�.�R�tF6�^�=2�~��o?�-:�;���ɓ��YS�ɓ ����SD�NpZ7xYtz��z�-�c=`²�R��J�s+�1�G$���v�đɆ����r!:�����DV!��P�tD����;K�'釵�3�*�d�,���C}��?��O�˞�!f�܁sGv>kήE��9�GKf �A#Y��ӷ��ڴ��岰�	S$��;DR�AL�f��lV[$���F�m֖�4�=&�`��ɠT8_S\����&� �y`/d�q@ w �h땓������@�zm4�C�Zp���d����n��A�Bk0QZ�0O���u�x.�L�{H�n��T�3H��6;�NK6J�Ń��菐=,Ty�?�
�J�%��3�����K��S0X���P���NY`´7*)pq§fm#�vV��$�&<���2�s�Zn9�t�$f�zl�n�v�>H�B�n�%��2���p�h�CHT:h��֪Ym��d��!k��m�#�C6�/h5�2,�^�T&l�fnБb7� Yj��}1ᱥ����DMG�5�2x��:������&-:5^!�,R��5��c�AC��*`2�me~���X(л�4�Π�z�&�k��h��9�v��3j�K�կڡ�LH7�w�-?QCx�V.���%�<���_�?^�B  �`� ��vL��s}��^��A���R�@@ȡ��
��zL�,����~�؇����/_��~�H���7#W!�����u��5A렭� R�&����UZã�@�kbSi9��ݖ���k�~���Y���wSx����~�;�9H���rC�'Y���ӧ��@��gϞ�N�{��p a�RvY	��CaE�#��Ha��O\�G_A�<=#SȜ����ѧ�F��矓J�kC7 ����y���0�v��ZF�ǖ�2�����H���sv©��a�,�{���[I/	c�d��f�ҰR*�Z'�W2�K�Rtrk�i\j��g��"�.�l"����uӜ�Ni��huv�t�[d6f�>����F��	g�#faKoi�~�q���1r��1���d��A��kVI�Hς���A���҇J�c�`1_�z�e����𰗜��۷�s�?9=� �Ȟ��(�A��{�ۈtZ)YF@/��mg��)-28��V��M��Ii�t��sto ��2�æ�)�N��ҥK��`�)%��[S�Ac��3V3��b��Q�^b�l��	�Ζ5���4 �P2MgPr���:�4`��+y��|;�*�]�$���6�֗>%�[Y��!�E�LJ�v���.h�h�F����@�t�� ]�z�20qy��ȜwT�¾�$�uT)�3�#��/���B|���8���L:b��$B��JKFL�6Mm���c�$�(�/�-^���$iS���4��,���
<�+�D��%|���Lm(cF���)bN��6<j:�ݖ��P�<;H��3W�� �3@�q�7o�b�똺�@̨;���&�ҲO:%5Gd�a⃃�ׯ�N9<<$}d��R��D�8t�C@I���݈�*� T2�[��q�vĴY�vC�SSO��B\	��֭L���^KC�0<AG��&�a�y͖���4]ԉENI+`M5�J:e�*4m����I7CM�V��We�J�����Y��$�kE�(�����{�w�Ν+W�l_�ѥ2��.�2����A�{]*��=ժi�G����L�A}v��c��H�H���_��M' Z���D�ji��<������w(�c�ɿ�s�g�-lt��޸ti:������w�������gx%~S��"�J�Pވ�nGXa E�{���?���o���>�Z�M�S<���t�<I��鱡
�[�!�Q�"���m�q�as��Jۿ�y��r�A�$���HE� �8����;�����Ӛ���2���l6��<y��jjĞV�n*_d��8_f�d���1k2�"�-J��L9y����˗�vvo^�~p���fl�+nJd�!��bA8Fr�H�Bl�Nu�+�Jp����hG�S�?���.�r9�7l������K]*�u�E���s��c����Zw�j�'3�t��N����7o�|뭷=zD�]����z�1@�p��AqX}��M?� �Ӣ�Ri�W���,�	� o��M^��Iˋ�$*f|�Wr:\�V������NF�,ME��߄UrO8��ˁ�C��!?A*0&5\ jp�ֶ�^��4u��7��Tak,�9���VsOe0JE-�M�EЪ	4��97�K�5�T�R3�W� �В޹�l�d�\s� �sm�H�����6�3����J�C[�"�wܑ9��"�:������V��E@Fɠ�N⛣�����47�@�����o��p�u�3�!h��jEu<
���ׇ��9��X��,BY�z�Q�/�8�Je���T�Q6��G��Y�>lߠ�8\���A�����WZ�`�%��-�����:J�4?B3�I� ��N[�q:%'t��P�uJ��3V|j��.  cO؅O���o1���'��̗E�ZA�<x���ޗ;���G�k�cR�?c�����Ӳ�!�
*u�Xq��А�-;�^���<N&)�jx�g�O�%h3�~���}�Tq�M`��抢�W���d�@yHINS�=��$�� )O��c�����\_���7�j���%|و��4�62Y*�-�5�Y1��=)Tߨs
�� ��#��S�%�[� ����
ͣΎ�5��*ѹ�<!��駟���i��$ׄ�C����G'�r�(࣏>�
cZ.���	�u�(/ƾ�<�̱��.֥'y�����K���!����3՟S2x��"PkSx7�Nʳ�� �볣�S�\%�`��� ;��\��<:��J����y���U-NN_�x�e�^"�k>�y�ּ��1�n�2L�h�oܸ!�]�fѥ��,i)E�+"����R)���˙AD�'E��T�";��@��;�Fh����%��ĝOi@�3Py}L�9�'NKƨ�)"�lt-����.���jY9;C(�!>1�v/�R9}����p)�7�p���g}���ێ�{u�K+N� ���"��/�jq*~4s���5� -�����>�TwM���I=O�Ӝ�x���Ec�Y�Ϭ�sHӇW�$�gݢ���1��:��0��M��%5]j]�E6��#�2��,2 F����ܦ���������"���J�������*j������w�W(A��aM�Y�H��-�Z��ZkT�"�R -Je��OH�C�-��P�E�{��I�I�,V�^�u�v�
�#l=��/��W< ���D;H�T��N���읷߻r�
����w����'����#�����X7=R�>�~}P�uc,�q���bvT�k����]b#�M�C�y��r.2y��b	�(��R�^Ew�z�������g��,�3��03�Xʢ�gym%i]jK.k��3Ή���U�%�����f��ݗ�&A�۶��Fe�����!+��S"���{��[��4�Ti"ݞ�)q	��:-5G���z�	(� ����,p@���	�R9f��4m_�R����J���XG��A7(�	��QJ�YHA
�.���R'��^1�h�x7(��S1Υ�?��9���4h��f���a��o��z�Rj��W��2͇MgX�C��4�hW���œT
<�1߱��͟m��<=D4,;�C���G�S��+#-,��I��n�lD+�A0����z��e#�|U]��� �e�)*�t�JkĪ���e�,:�8�ԭ�E�&e��4���#�N�v�ڵ>����?5��k�>�)'΀���H�j��u�~������ۇ~���)��)� ~��]h�i��"9|���N����ǎ;�	�^R�ӗ�i_0�;H7�@��'O���˸Zv�=]�I�Shm��(��h��k4��p}��-�CuL����CBH�"�$��;;[
�8`��f|\��K���t�&�G8�����w߽u���L#2�NOx8<��O�>�;D��
�0(��n&�d��\� �����,S�",�eqrX�t��!9�xCQp�T<�=N6��-�H��ړ?�N4ۼw�y�<������'?���v���M�Sau �&4��j����N�ʵT|`�4T���]����:C�P��%��j�Ak[��9�\�eq�`��T��xå�Zs�l&wp.p��bgg+:���\$ �	w�f��A��� ��Sբ6iV�2��q%!$1c��[I�O����>i?�%��fm�Y-���Н���#�3��4��+s�|Q��AF���eIt���hQw>eh?�rڎZL-��	9XːћI���Y%]�%T���rR1관�$�C�*�ҍy-nB�pTz&(�<
���9�Z��#N֜����ѣG`��7���8{�˲�N𜻽�ݟ�[FDFFV$Y��TAQ�E5P�4�h�O|�C�/-!S#1 4��jMU.��Y��z����.g��w���g�
y��w߽�ر�g?�ͅ.���1�[|#y]�;�C�(��B�Vko^��r-A;�������'��\-h�*S�p�p�ZDa7 �;ӑk>T�k���u:VȄ$�>X^s� �.��i��"�V!���~ �f�pMd�J�z�+ �)�ӷ�K�����W�?�� �K_����|1o`UE��֑��5i��gʙ��aЂ��h,��zx9Y��U�tv�SP�����t��$t���02�|�r�5�-��,��jZ�q�4�5�l�м�ViF����dzuP�S�F�����0Aۻ�K��������������C }��rs�)���p�O'�d�8K(1[��4��R�8�*�C�[%�OA?�\&4�e���Ej��q��H�6���޾�����/��4F�l0g�_��/_>���k�f/.�,�&����X�`%RK����5���Nr�ۋ٣G�6䅩�&�-u1��İ�����W��Ź"d���K]�nF��)r5�<y�.`���uO=��F��P,d}��=���]��!6�����W�\Y��K����+���m�H�Lǆ��#�-���ӊ�1��bI�($��I����� cvN!$��~�ϔj	'wG�Բ9i�j�(��vKY�[M����H0h�1����������Yg2��i_@�F&��l�VM�m���V�{���fھNƃ��|��/�rs�z}�u�?^�z|a,�?���D�C�1@ψ���X�_,�{���]
#�0₶�'�l�K�$;�6�agm�=" <>�J�F�bF�Tq�5K�Ped?q�x�f,��+s�K"Pӷs br�5n�w�*v�����2��I���zED"5�}�t�v�H�,)�Z��z2/��:-�Z�Q+y���후��k�����:�}���5(�a`4�&i������bA�o��]��6����+\��⁓�#}���A#����M�U�����.X������P��x9ђ�f�Xm6��8����v�Rf�M#���8ݎLPlS�̛��`��aV`���Tʤ��q�܁Ş��WO��'[뻴�[���4�q�	��{u��T8~}tK����ݒ��9/�i���69M�I6Ь��\R@�[t����Q�>���s(��<)X�f�Ѕw�̷���/��1�f@�(�|>܏����JLD�'$5�������=�,A�La� �ۺ�1et��,������A���[�g�-	dZH4���K�.�l��~�ZȒ��J�S#���.�e"�fr�H7d��dj+W�� �Z���ى�7��#NB�R�,��tp@�%]2��?�̺�)}d��9]LO9"ʊ��[�ۆ�l:O.#�]�8�8�9�߮�Q��u
��;Y"+qc]���p����]V����2fH\[Y�Oia�xܧ�/w�z�l8\�׮_�s��'�|�+�4��*�E�\I���my�"�����{�������׷�Gt����Q#���TbȪ8:/��+\�Bz�&"������=ŭ[�H���3�J,e��t�?a��C�29\ ���y)���,=���G�茭�e�	�6)�7x��Ň��z�����)���˗G�j"n+�a.-'���	1�]Y�'�Ō$�nܠ_�����[�D�Uڣ��}��W���~X �O/��k�$h}���J��dk{n��rY�����n�l�����)Z���L���:bG��Nj!����D�&S�X��g�{~�b�s
MK�ܐL[$��������7�uy���_�ݼy�n��;�s�4(��4GX:�)h�`}���N��O9Mz����k9!h끹Pep[�j>���2cA��p�q[���i0��i�:!�yO��!��dZ�$w����;��	|�&���{+���(A�ȵT#����'���3���u: ���D"W�ψȟ��\���d�C��/ո���y,S�m�M�]nf�zJY����yj ��f�����uj���,�t˔�S��4s�^m�K��[0�	 ̥̂gM48���`�@��SLH�a���Q�Y��&�BGA�����ӎ=?3��ѭ��"�G8�Z���%t�6:�wȧ&��Z�k>�Κ����������v�rm����m� �	�e���iQ��f���6 ���c,��,�_8�|:���ZI����"�d��������C����Bb�0>�<>$s>8��͠�;_\�q��U����h�4�/�y>>�F�ͩHZ���w��n����E%����聲.�������9t�bI6���NҐؔ���vxmO�_�p��ԩ�(Q�S�
K��d�����"��������ޞ ��ׯ�m�ݼ�����������'�e�TG�.fSK�A���5� NC��D�t�)@z� +<���a�>�Y�%zE�;��R�<��7Z�(��g��?�=п�͑�-���V�����Oy�0� E���-䮐�&����>E��1����`���k�clPZl[B�ʡq��p���A	Z����i<�T/-�Qr3����덍�|��/�����Ç�s޼NwBa�/~񋇿�����W�������l\��W�r���p�Ӳ���)ӂ�bS��TdM0��nJeB��.S0��\��A6��������6҈³݀I80�JZՀ(�"$& Z�1�H���^�;��	9,��K<�ڌa(E.}�q.�k�f�������%�N�v�#_�o��J.-��8=<;yE?�?����R�  �B��cV�ne���f�$��)�Wg�	nu�U��8�3dQ��}����tb�Z��lM^1�g��4:Z�KU�҉jX��)W���&���� )�_*�/��p�������?����先 �.�v�S�A"<����{��X����M۴JfG�k��5��
}�Fڊ�ʐ7�R_�f��aS���c�C��Z4���x�y���\��d�=,�=�Q�a��$�s��7�4�[�
�TQuF����w��*��t.���iOv��l�x�&O�N�oݻ����`���6O��s��/�����T�7��_Z�y �1���ٔ���u�c!�1_�"�:�����CW�cF"���NB
�1��..S�����9���.�3x
�:�9:7R���`�����m _�2�|��w����ӛ���K�	�������dg��1�b�ݓ'�}�0x�8��������3�)�x��b�>����y��oh���p?z?�}#�Z�TX��4�=/�C�I3�T�j����Ii�J)�,Y�tYz���0,�Ӕy�-a�-��ȵ�͎�IV�P!���9sq,��Ch D���R��x���&�8$w0�o��&�a�3b�u��Z�Ua���F�/���3��d�+-�5���%�A�~p���2Ე��-���a�b���1rv%}�������,�@G��g��U����5ra{�Z7�b��u�_oܸ!�~&s6#�e��x��;zV�������o���lӟ~�쿂Y����)F�v|rhY�VG�a  �������@�PY�m
���U�=�����m_,�����VWy���8g"�.�����7�={����$���?�!�^��>��?�������3� �	��f����Iq���~�������=Z���z�'3��O{�����2 ��KY�04�Prc����d.3
�9\���z���|6�A�Bk-�����8�X��7z�*\D���ѹ�aA�9��JC����a;>z-�$f�����k�.m�I������#�#8�]�S/!õr�@9��i>��F���pL "եe���;M
xm8���dt�/�>V-��`*��FF�A�����x2/�唱���ܕ=��HHu�x� �Y;nPe�� �~:("ϤR�����h?��C������ �ȕ�˖�:[�Z'CKC�C	�x9��d
otT\�62�Tv�/.Ȼu�8���KxF�C��3�a���huǱ5�`Fͮ�Ԙ�3��ϸU8�Tʪ6)�ӦcB���>�UAK�����J�ݛK����B91�q��fgqK��)�$B��l��m�S��`��ݻw�^�zU(�k�6+�v)��+VΌ)�}j����+z(h��f� �|�o"BMK�!�&�+��~���A��:��[�r���k�D�)i��(�eh�V�4�J.�8/�'�BK������k�B-���&�l�\t��شN�������H0��0��o|�v��`��:�`/:&��G���$��Ma��EVK����t�m+�N�PH��k��H�p��mz:�Pz
��)�����tI^�.[&mJ�rU�J���c1�a�˘���G#��p?�eOk�"�>Fq"��~���=�7cG#S"K�3���GU���C"����l�*�^�-�a�1�qϹ6-��M����^�f��f`�5m;C/�%H	�;�!�t���.�8��-y�y����i	�Љ���������&:��=Pz6Q��z(^�)Sҭ�ZE�xɨ���_�m���[;���E�������w��N�D�W�W�/�~t�����������fs�y2e;B[T�2�t��$�����β��A���������������b�p����� ��N��=9~N��i�T�2Sw����X4�u%�e�Y�Y�j��?��N8����k�r��%�(=ou#8���3ţdB� �T����[X��L¦�L�J������&��bl9D��V����$�8V�������Foq�x��d�v�M6Z������'�N\ݲ(>5]�y�ffm����Gm^�K
3������rHáhA�.u�	�3��#8ץ��7�Pa�ܼD�1��%�}��;��UM�����$0�^y��#�C�,��^�\���φil^�Xpl4���X1s�� �R{"�d�3.�K���e��Q���G��~�駠��9lk���:�xs4���k-"�Bf��ׯOI���ir�IF���^�ON��/�)\Y����ْe>t��ʙ��8��[����F'��h����e7	�
��'7󱉊�D�=ҹG �=�(y<i�bY�Jɝ�W���/3���$��f^�c�����	¶�D��b�\�R8�+g9پj��	Q�J봢îi2/?��qfH�=Q�Rv��nEx�2���t�l�0ۡ��2s�ʠ
�%Dx�>!�:::��/ޘн9|ck{�$o�Jfb�z��E>E�xcs.�O�8��i.�mCmF�,�/o�;$�d���`�/�;ɓFc��K��S����4m��Zǰ=5Ֆ)�κ}Ql��%��6ӆ���=48x-/g����!9.��ry6����$h�rvhZ_ߤ�����z���L@/�B	��׮�h�܍�<���tZ�k9��{!Z)H)�ggk�ϼ�s�ʮp�d}k3s�/�X<����ѣ��%��7n�T�z����
;��9Or��y�M�sFtlӽ�ulr�\�`y&���Z�g�����{��{w޼}�Ν7��e����d���D�ǲ��Հ"	�fc�6Q
<H���I�S��tLhQ��N^�>s��iv�� ]�5���S�4�v����L%� ��M)OѝM�������>}9�pj�]l�l������߽�&})}]�浟�x�urS��y'��SU���Lq�T`U��e�ȼ�Q*����~�[ߺw���[7�̍F���e�,���~�SZ�۷oq9�rl���~]���������F=ă&�
r?������7�D�P;a���f.5�r��ZKO2V��3�mr��lƗ�8�2�N�����ڿ~�ק��m<xp��흝�j�BVܿ{�������_^�/$a��֡�PDYȉ2�땝�i:�V��eppp����B3d��	�=\�B�^ᨕʣ쵝f֨�z�鐾��C�5���vU{��7�bf9tsY�xE�e�gD2{]+�*L|��t(`�}Y�Z������˿�2�3�t�={kF��e�/�(s�jL))u>CO'Y��!����@lQ:B��r%#���}�18i(��R$�15%������B�[:�g�����K`Y �o��H��.��EB�߁ĝЎ���S�lBi~�A���}�t�q�Xj�8��(�A۱*/���L���^�|-@��j0S��r��(ym _$�6��_�a���o]��[^x�3���*�|�"���vT�dF��U�H�V'�ؾx���IK�Y��<�Pb^i!3�!�p��WDΚ�T)��)�@�4��A�4�k��@�O��Ȇ�gH��&���r�t�_����</���ȇ�/-����	,�B��{z��NS�_;2�B�S�X�w<fVl���C8��ܨ�B5\�Ztv	��S���[�e����J�j��yy��3�(�r�����OsL#q�P��
σK�d����%sm����+d�p���ӊ;�u��l� ���2R݋v{k����?��ã��6OУl#��|U%3��E^/`Q+��>P�q���u.y$�ǉ�"��{˒w�m�fE�LI3�ҼZ�*�&4B.�rtzb��������+��$�O>��^���c�6m�%=)d�<@��d*B����>�ZftZ�eG>3 ��|�#�h	}����ngg�֭[(v�yY��w����[���я~���W_~�E(hЖ��Ϟ������Ջ�A��sѿȻ����HƏ�����Z�=OK��������\AГ"���	����&!j�;[ᖡǧ���U}i��b3�"ކ�d�=����9˂v�E����X՗�<�WO��v8�9_I������v��-;e�yA�p��E��c3�P�\}��P/f�(O4�b�\==�3ɻXܾy�M^݀L����񠰕bi�V'�`f%��I�)B,&5��t���W�^s�[@:�,�� ���-S��b�!39�|����x��ne|#2q�E���������+��2SA�KdJ c9�.I�[to�<
a�̀߄�i������m����m�R˥Xf�զT(�6� oN,T��b=���kN�F�4�-(`HN���>57�d��
��߭"�0�49�,o�.�\~��^���_V���:�b��σ)��i�:��3oe
�u��ˣ�P�3q����ꍛ{�3�/n�سj4W/���m�0���J��wX"�aˆmMR�.x��;�c�R��a1�2ڀ���Z�֜s˿�������[
27(���L�df��e�ći�
��4`�{�_��!Eg3��EӖ/�൦��S҉���I"1�+�2�s�7�И�B���.�d�)y�LHۮ����d)͙��Bh2�U��i��u7o����E(RQY.}�:���LJ(�I"�n�'Լ6��m������ۻ�W�ã'�#��X�7VCPtUT�,>��BUњ�4Wf`z���0[�TS�IF@�jm�[(�w�L=��ŬZgG�e�P(�ї,]7����r֭%���C(v���̈́��|���W_�'�Cy����\g/�������7t�넑���x����k�bW�t�8K��	-}l7�����'O��͖���_p�o�!}ɩ�1K�&O��һ�>x��,����������u�&hh���!˜��%&��į��*I�Vŝ%J��-I�~�[�"�����k��nΕ��k��T��(�5�:�!��I�k%��N[ƵY�ݠ)�NĖ>6�����ʄ�҂��l�AZ^!fF��*\.�5�-;m45��_��_��_��;w��^cr.�J���ɟ��˗� ��4�YX?'��l=��?��?���1�*}������7�ӓ^ 	%�T,�u��p�q�pUH$ ����\g���I��G���W��<6lO���Lf�^�8���)�7&/��qvzA��΀�&����%¡��w�T����_Z\T�Dr�C$	�٬�iz��)�ctsmk2�4�՚uZ���N���y23�AU�)"�d	9�N�f۠�_E���i�2+�)7�˅�+������X�=R2�� ��01�ٛ7�����,ݽwosss*/�L��j��NY�ΞԞ���ly��6m�ZEEA��V-���G����ri�n����<�V�,X���Z�3k������=E��'`@��K&�;��
Q��;n��~�\�o8N�w,�eL�`C�[�<��Nk��zqg&f�]¾��&��S���_EGQ�6���А�� ��8�X�xK�u�ji�"i�i��(��ܒ5���IHPD�A9L	�:��l��:f���=,�� KfV:��V'g��A3�p���ܨy�N;��[v��v3��\;$ڄo�T\�7�p��2���/�~�jz˧����@#�E�kN��ѣ�tK����X��H�j��G�`7�)�ζ�f�CR�/�����jWIm\���/210�(�R�x�Bh��F��^Rd��.A�� i�e.s*���N\���ظRfV�SQV���(u�O<�)dl���%��i�j�Ś�j�.ai�T@h���tM̟5s�H��N���X7<]�i�=��_$��r&�  �x;O���Zr봆gx����?��~���o�@fhk��ҁ���SuMЬ%֨`�W''%𪊘P������#bƾ��{L	Y+�ڧw޺uK��*�l��R����A?���ۿ������A��nv��ӧ�q�y�"9�v�crAs�&�93���\�Q�&��J"�oR��x�������3	Dp�r3kwZ�G�W��¹]�=� �6�7�T`�Q-Ո�kOy�������̩h�RB7�2Z_39���e��M`9;Mӛq�S)�/��(�!����܀�`�^蘦9�AG�Ӧ�ߘ�V���uz��S��JC�5��������Ro#r"B7pd��=���
���Uї�������t��H�Z��svk�[)_�ǥ�T[E��ZO�.�$�ͼBW�}��
Z��ӂ�CO�b��%Q%�
G�}�E$6kbIpļpu���%f�GSD�v��Jk��8̕����kb�D���%5*�_�y}}�J��htQT	����lYT�.�9�lw��-������<<|��#�-�5ЗtN�Ϲ�<�=2�D��a�`s�m��tI��}�[K� �4I��ގ�#�i�#qLN�0�h��LǪX��)�Fq���2u�筊�,� �U�~����\)�p��X��z������]6�֑F��,m�B����Gl$�\[Ü��5��b�U��m_���LN��4�\��?1��z6�t�Ur盛����K��ڏ^K�ͼ]P%8��Ez8f��d:ECwȌo�_�^_��<K$��:��eG릫W��&K��7����م��L9����A��_���.r��7�[��N�7b����I���2��@����/7�����!�� 0���)�~���\�Se��P$��}̜���q����f������� ��ُ����SV7�|�I��n��x3}�����5��}�k���W�����#�P���=zT�Z������`F�K�b��/��ǟ�'��©�o�����=z蕵��hprv��Q�ŷ�[���w��'�+YQ������w~z����>n�~��y�JJ��������o:ߺ<s�+�nH�ө�V�Q�T�˞__[Y�ݻ������߫HF��MzXruB�tGMLvH��&�������AM��;�x�x2�N&�����g#�XH&��.�l1'�	�3�<�"cƁK�Ăd��-����bL�~v�ڒ�ްY4pUITv�w胤�1x���ۣ��x������ON.G��Q�<��3׌����G��U���?��IS?x�`{����u�)���P��f�zΜ��f>tæm@�tvyh}W�*W��_^��G*~0\������˧�=9C=ZgPL׮��p4c��D� ����Ǒ8���v�;AOkҜܸO��-#�����W_���?���u�������˪� �������J^�`���e�EO���^�V+U�u�%�4�u�),T�����g
� yv��psiB/��f�$FM�)	4B2(� �1��E��R�l)m|m�)A���Ok#�A�K������[o���	9��"�	h���w�w��o��!%���IӐwvL��XT<�p9{�%3�2���YE�+�5Q[��Z���[� �k?T�d:��q5�s��`+�Oa���āeߐ����RZ��X(n�J3{��~�.S(�WpXrm�@���/o�m��9��q  ǲT�y�m��t�1�����bظ�L�� W$$t}2%�����G?������!�LPR�-��d|A'��K�r�%���^4��}��g��|9on��Q�A@����Y�º�Rk;[�h����Zv��0w L���)� +	��,�,��u�O&�x��4��"�0��C^0V)Z�Օ��R�Ң��Ha��)���GH���?�А����e�FG�dlFՈ־�$
fv�V܍�'�Ȭ�bZ�!�gXv �y�P$\�bE���\8(HN�����${���-����H K��[�I}G'����.P �SR2		9�9�1|�5��-B*�r��dP�w9��ܕ�	�!Bf�1�AA��L	ɸ���k8����P�y:qϟ?��6(��d��<y�M�ֵ�\Ӫ:%K�L�fI<N
UӷcĤ�#�9W����S��`'{��+��O��oZ��N[2����P�{V'Ɖ@9$�(��?�7�D9�YAV�SH���ڗ�yQ�h%7z���lo\�,����6`�v� 龖��q�x�ZҐ�%�e|K]8��<-��r�����{��>�裏�W��$X��a���.�_��)�'�@��Ǹ�m&?�XțW��0��D�8n��2-�tD��t�/�s�z�Pz(� ����\Te�Bq���*��K�N�iU��I&�S����fw��g5�+õ����Nܴ��>��(Zq�_v5��^1��t>A0�U��rɀ�X��w�1�f��A���Z��P�(�}'#��wt}o��l�{�����,��r����n���fP��,[!N~	n��ׯ[�\i�"�{Γ��3���B�5��$�����o�G���XX���(�K�͎ �R  ��+��\2�(x�%ٺ��m�����q2X.Z�4CR
/���]w�ܙͦ�S��Z�XBԑ���z%��d:>iL�dJ�C���k��&��=��Gm��jA%�yg���>\\��gNT#%X,2B~�*zԠQ��	��0�L��sTG ���E�P��;�w��-Fe~g{��@`��̢P!�.�t�b>}��щ�KSuPz��Y9.����@l��9�9Z�ym���Pr%�={v��;�Y �qP
�An�4�b:��)ֵê�_Nģ�9Spt�ι��)�H YX�q~缵B8�l�Vrm���:��ڦ-/�~�����:"���C�-2��ie2$�"C�i���ie���]���s�W�����2��ǒ���@���7�UI��͠P
�I���!_��Hi��ԋv�l�.EX��M�r-�"i](����u�M(�*׺$��q�p�chk�����>�+�S
s(B᜖��؁_��)Z�Y1����%�����Q(���,~��3LQ�8s�&���R��*�6hR�at�l�FD��[e®��K+���vPy�.�+SCM�q�9�di����7����6���*'����5}�W_}�Lm��Qq-O���Ɍ�U&bl����[�V��c���1��!��]����x����FO$�|��Ka�"�W��ͻ���J#��˙,�)G�4h�V ��.�߿G��n�x'A��fރ����*�-���'�Q������#����;�@���poH��^�Ny/e��<*�ier:�x��a�ɥ{����+4F2 �q�隧����3�8����++���?�я�ǃV�)�����W=�uq��U��:��ӧO�G��zl׻����%VF����\6����t�sr��J��jv�fS�!�� �ܷ^���g1�c*:���b."�>��������> �}���_��_z��XIo�������Cg������W�)��M���	�S:'��!��R;k�BN���t�621�Q�P/��
x�Á��π��_N/�#(j� 0�Q����p8,~k����wX>x3P���t0�qIR�@��
��C�@D���Q�$E_|�mb+�'�y��١����\��Y�(���]�'<�N�-=�ȃ��k���Ȏam��LͶ+Kf�.#CE/v	�̲(]:%�

!�
�3�VA��sa4����L���۞��\�%�jXpdi���@�1g��o��A��2�����������9�nD��)���r��vHz���t�7��M�ӏ�c�i�O�5ϔ�j��m���95�)Ke	��0e)q��U��u?YV"W�d�3����4a]+�ש8�`w�����q?�(�`=�8�W�-S|�SƜLY���	�-xdK��G��(Y��W��n��f��E§��=]�`D�0����T�â'9�?�p2�V�6N�y�R,�:R	V�s�`�`, �����*��+ytf#�B4��o�=X�%l�v�Q��e�k�]� �Rg>h2=SxT�ཹ�x�L�N^ё���2��`�p�Q_�-����a�D�I�T��v^�|Ia�LƎ�l)�]��L�C-��|��A��K��-}ir�:�����~\�<p���ۺeZ}�&�La�@��U|���H��^��6�x���P}^�Yu�0h�4��i$;���E����f
�zaP���v�Z9�d�<D%Q��g13-�Ŗa�uBoc_�{N��̸2%,�K��L�9�,t2U�#�h�T(�[�,.���a�@�ҷ�]I~�i"Wn'
T�2[���,sP:xz�p0z���H�BR��rH�#%�V�)���֊Ԃ�nb�|�<������GW��S���
52 �!�R�ڟ��Q,�]�G"�,� �H����N�:?��؈��4l��"��N�G��5k��B�ܰ�8,E����̕u�@����֐{�Ǒ�'��|C����!m^A��-E 	������O۴���c�X'C���0� =;�����B5�������F1\��qX�r�E�^���3N4N���J�P��t��q�B�k�;��GC�W�B���j;�xX��
C�����
`�:����t�V#���x�@^\�A����0d�x��d,hW�~	�m";�҂�����
,��2���o�\(C���B���W�T��[��ںy���˃Ǐ7��J/$����b|NC�
�ә�X���*SAH �MBYIj�Y�4��uA�Y$�����hS�d-\(��$]e$1��x;OZ{DM��/����R�+�p�$�CR��N����<.�bZz �聙�,,f�{;�:�9���,�mM��2��E��\n�-P��c�g=�s�/��yMm�ݰ8�t�x�|2�ѭv
ec��m3��5��]�z���t(�P��Ky�e��wBv�#ȹR`3&F���� 1��onu�5<!Ĵh݅@VZevw	�F�7A��f�b��_lIL�	=�?�B:��@�yn�e�������}���g�'��K�?�"�e8C$�XY!�_
Q^Z���6��%��tvyr|pcw3���Xr�����R��[c?U��l!��=��ܷ�~Q���s;����ְtڷv�9�:��)����n+�ݽ��������+��z����xүbZ��!k�^Q�˪�s�~'ՏzOPI����i� 郦޺�Sn<���R�����E��R�2��P�&=Lz�K�=׼6�����ڵk�������X��߅0�����7n�F� K��:(�"R�9��Wϛd��kk�bsW3�	�����ӵ��hm��DKJR�駟�~�B�S..�*�B�2W:��՝�͍��z1�U�6��lGf��M�c��#�ա�7^Nƞ��;�:���[����_�ꕴ�Y�7p<�1����|H�\������H�Y��|�T�7�y��ݻw�^���&[��[�ͦ���e¥XN��I�
ߑ �W�_Ջ�$����Z��2�tr���w��m�g�U���rcs��������[�`;پҺ5@�OZX����2��M�wJ�c�4��k�� j)�A!i �kZ�/W��'��œ��(�� J3�{�Ү���MZ��V����D��ny�|����MH�A�q|�� ���l���/>����܏?���?�9x3Ÿ��^˶��h/�u+e��Z���E�Y58u[�o��o���PZ��c�N�lK�-�qp��O-��{�\&���yX,�*�I�xR�n���.���o�����N��X֩Pp���;j?^{|L}�u��^��%�JZ�͊�A)�Ҵ)�T(�5<$�h��
Z6�sG�y��9jH�=g�o�T��,VV�����h���/ǐ1�W�&�Rzg�/�$�Q��4f*$�^Sov���#4�E;�p~,η����l���������,�͵���*�<qs�t�ծ-��pG�?^hW5�#A!��.C��b�K��'�+9����r�9Tߢ^x�?��{!H���x��_���+�p�d:�ǜ֣��N��`z���]RX
8-�
v�Z�u:�r�E�d���h�ڒE���g�C�7ڦFb��+�U�bd,8�6�����y��1HV��~dמc^�YJ!�>�7����˳�ZN����V�	�%l�o0߾�A7�3�KI��� ���D�
�˞aaE_��sN�|��G��9U���ߣ줣�IR�cz^�E��!�vppW����h*hJvGψ�&�vв�A_�Z�ʖ�:;A.�%��6�'�\���"��8s���1y�hD��n���A��"���w�S1O�S���%�K� ��h�P�7G��	�z�j��3��7��xrqv���4���GGGO�>}���'OX������F$!}З)M<���>��tڱ͌�D�����L1�<�bJe�ɴN+���2�'C��Rj�r��F#qO��҃~C��o���ܘh�]�%D�rt%����t,����@��v��1���]��f:�P���%9��['�8��f�˂㋒�g~�r��e�*3pA!H�!q�*�}&�zc7#m��db�qU��{||\���<���^�tG��H{}Y�N(wQ�΄hh(/l�UM��I�^�ˠ�O��V-�|��󫯾���_%������ZX�aM��r��i��%�a�>!��P�QJطm���j+��q'�
��;w�|��N�ČMkkF�N؁�H�Pw�<phc$"�a�¡RMe��*�L����7͒D�n�>���2��.Y���ӱ��*P���B(�fS�Of
��#�H�I�z���m�b�6"����a�<������b>���D�ސmdQ��V��_UD
�Y�`A�I�S�n�{Η;^�|��4��������x��>xz:"�sM�=­$s�H䚠U%�����f�k��J2.���&i(���[=)�������<�"�B�KO��� �N�(3���\2�#S>)����c�o�:��X\�����Y����6��F	��1��Y$`�K��x��;��7�|���������BH0�\�i�b�Q�xn���ü*���O��*ceB�)�W#CY�
L��U`/����ޥ���}���� NOO�g�7���G���u���n�.!��t�/Ni)�>�&����!"](��Ә��E?8WrzTÀw�x��Z(`q6�K�2ѓ��u�t�����=#���K$(=z�vAv��@�b�u�|���J:��
�Z>.�H^���o���=�sz�e8�C��o���u��EA��U̅D1yZ�#f
kC��!��[���;�2��,�$���۷n��b�q���p���*K$~��3e�UKZv6�6c.�ԋ��b��6��,n��(�����������rˠ���ဦF�4�(t�����*������ˇ��-���S�nbK~���f�TK#�����ȹ��Y��V�V��͛�I�^�~$�(���7��G��'��޽{���U�X��C%T*���d �8V �^�'&�m���f��>�Yx�z26�(Q����m�����L�N�Thk$�ߧ����=2�(�ѥ������1��Ԭ:67��?��Y��-9��3��w
�&m����Q-#J!�lce�� ����'W���:쒾

aT(6�]�fqy�8�g{�6�ϕ/5h=�i^�Q�RQ�N�mh|.r*'�/n�v��`�;��p�ߢ[ɠ��P����T=D�A9鼏e9��y���!��X�/�����M׵� υ�i����g�!d�!��Ο��� ���iI
����FG``�m����Br�im;M���:U0(@�\jsѐ�Yf�t$���d��Ӛ�%��h�,B�\'c+-�c��
�W�ʒ�iQ��K�mH�gZ�ku.�<͙��ɪH�e	�Y��7������C�s�f.�dD��Z�5�%Hq�pxD:�jI�T;,(Y��x��>���+w	H�	�L������0/���f2�DZb�S��K�.e2����q�,u:
6Sڇ��K��4�p�l���$N$�<��6?�+%��Fys,�C	�_�U���--�{N"���%�G6�ɿ7h���w�4]X��1G�y�̮ɫ��Y �$h��|����6�Iј(bŎ��i5���R�j~l��
���pF��#�-�/ʛ�x��u�3��B�:uI��%�`��kJ]w�8��l:�7KH�택���tH�});���P&7VBN,>���C�fuu{Dv�ؚ�8�
���B'�
8����!�����'�<�H�%��g˫��A�g�'S���`_�{�/rJ��� �!�{2��!�O������&N�T�0�d���,ٸwq�,�ȒAލ6u��[�=Z��c�@c�t�x5�`s� -�S]2���O�tx|�8���Y�Yg
�k%���R3xR�J2�a���аB�P���	����\2h�n�~���f��8��x)�P�3}S$U���mb:og������jmj����J���d��?�+�|��FgL쬏)x+<�ZK3������)�V�e����SV�@�W���"���6�]r[+���&�Z%H��K���NЂC��uZW)�`u�Ąp��`��t|�lt}�;@ �5n�9} ��\'�B�vZ���JS�%��VK�0
.��YQ/�3˓��3�,��{>���rO��9��c��A�`�@@i:��|0�Ѯ��?S�m�`�BAZeB1�>�mV��
ؠ�tfe�\B$CWY�� �d#\)M�8����2�Ҁih�\�Q؊lt)��54��	]����]&�"� �+F��HP��@n�]�6y��쯲��ie�7��-_�^����CH]���6ff��M����s���{�Lʈ���W=�	�q�)ZtfdZ���P�`�-��T*���+�͠��\���T
��Ǹ)=���*BN#���ͳ���B<$f��S�j*05��x&�8<��g��Oy5�߸F^��
��zQ�������(��sQ���	%yV��	���X���!'A�xl�D�L�����H����Z(e�B[�`P\A�}@.H����VE�����~�W�׵<{��LA�8��ot6Y��뀀DZ,
�B���r�|V�[�|�t��Y,C��K�Bb��i������~�[p�੼�֑+|zv�g�3�?�+�Hĺh����S� Y㭭����wa<a1识��{o��7�	�Y�P�B�;�*���n�{�����޵������j���+�th��G�!/9ȹO�rP�Ww���֘������������A����h�NQ���oll�%��g?�)��J�JJ�ʶk�r�>A���f��fr9�P	)�|e��c��)?2f�~�)v�ƍ�>}��>H��l1}��G���͛���	_
@�L�m���Ϣw��p��Ξa4�씑I!΄9ɳ�,�RrR+k�h�䬷ta+�԰R'�\�)h��g�`r.�� Gkl֒M���s�}�6[��(Ii�d2�;o�����j8�����ŋ��>�=/�dt���M�.::>+������+yѯz�Ŵ,���J����FY�X	�iۿ�o���+Z���$ϦЁD$�'&��AX�`�̱_�3$�b�ھյu�ΐp!��R����޾so{�Z�z��y��
 }����nm}�ķe�CR��(�]Xq�8�Y��4������EMgD��Ţ�����5�5���[�nQ�zpp�.�\���"H������B']x�(�㈐�2�� ��YZ�\�n>����7o�$|���h��U�8�r�P�R��7
�(�$���+^3��ԇ��(~�٧/�?���-��%I���%�l����ʚ��gQ�h�S� ���jm�0���0�=«�Z>n�KjlE��(�%�<c�ȴ��%�=Ms-�g:ޜB�_��\eI��2(_��{4�e?[B��nA�ߍ"O�ә\R�� ���а�D� +ѩmyK$��mR���&L:B���c����������d}�]�Nҷ��w&L��O ̈0���H�ʘ|��U�db��J��V'̪��挙O�":�nY8-p�}��3�'<іi�|��!��c���e>,�'�)�"X�R�c�M&Օ�$�6�ϛ�h�zp�ҷԡ��-�5'g
��0�� �ش<.��f��˻8�"�bGL� _�,�t�Փ��@n��c��R�+��̜9T%�#�sv�� �=yJ��-�<�^
~F-4���|�Kp������� ��H� �_hW�5�� �9���mO0�\�Ǌ�͕��t��Y���{�k��k�(���r�OU�� {u3�u�a�y�%+@l	��~�N�*�[a���%N���u��fn���(�SnYn�{�o#7m��i�M��=iz�V�ڵ��BE���6r�N>�]��+K���{e������Ç�6��A�sw{A��֬ � �S$�o�-��h���Ķ����`��U����4�5��,i(��n��A�g�O�[^�|	�f~|��r2&=C��d�H��5چH��s�[P������o�@�@l�v����K@�s�.Eg3�)�"&<��Dp����g�2�(�*��'�,�g4�ׁ|�7�x�V ���z���k�����I`t-@;H�.�/f��]H��#��Y��Pd�B};z��W+Q���Y��=�i`�zXa3.v��&���f���a;����%�#��<rRYq}�q���ͅ;�j ��E!��aݬ�����
�qP^����~P�%H!�r0���Q��V��,�(���l���فM��c�:�/���ߘ騽:d���u%T�"�g\2fбMV6�	�
k�2�OA�e�!�C��@��
:�e��V�qZNδ�BOl�C���h%2V"o�������d&O�^�3i'���Z,��f>��L���1"M���6{}��?k"�gKA��C]�x�D�p�+�4'ٶ5$eu!{k����,gg`c�����v�jGƴ�ej�q;[��[�q�+ߢ�����)y�53�/f�ƚy�Ge՟�5
nr9�tM;��)��Kc=���ߏ���v�%+���l�K7��t�D��9��VF��$�/Z�k6�j��'dAci����T�3�Gϒ��i���z8l-t�%��u����G�}��{�w��uI���K�q^#�e���}H�$f����������V��tX��\�L���!�ő�T�E,.�	�twO¹���)L�r<����$F_{�,=�Գ������sj���4�t[	�w(��z�� .AG�i_(��@F2��"�a��<2�`��t��hm��y0`�	Lgh_e��~����7ر<Y��DhaA�p
(��·b?��/t����|B:t�cF� s���;i����X���OZVY�=���k�"zcX
�-��]���^�:88~�����ʗl�zP1��x�z�����e�H�
/�9�;����do���[�H�AzYM8fr=<<$׊��սϠ�(��w�1t�<2�Eɞ�J$�	�#BbZK�%�GG�쯼>�Åi�O�@�k����t������>D�[��c��S�
�Ь0��� Z�J��u_|�Ž�owCw��u+�)NI~��##\(��N����=��Q�������>��s��Z�ꤎ;�U&s�h�$�&�"�������W:�2'�4�{������<ϖ�����&����ӳ�������ݝ4#�h�Q3��倲؍��>������?��?ŨK�`A�U3�������9r^fς�OqB[-�Z��T_йF�Mޤ;�˒ha�P�6��.��ش����d:2���U&�w�������M"��h�<��қ�Ԑ�tZb]#F��|
I0k$Y�2��X
Mj&}@�o&���l�`�kɪ��)p暄�� �^K+[�N��:}e:�#Kx���*$'h;0�Ͳ ��FGخ�:�6S̈Y�F)3��Y2��'M��XJ��w(�LI��fN XT�*e����8��-��u|�SH2��T8<�N�L}�eI%3�2�"R�7��>�#2�xF�$�B!�MK����� \�Nf)� >�P�'��v9h;h:�Љo���r:����L���	m�o�A:��]��!��BY������.���)R_ �����q��t	ʹO�Թ@N��8�v��	������L3��s%ߋ�
����JY��p�v_C��^��I�؆/)3���O�p?2!íd<%�L# ��A���dm ����$�ЦK��R��J�]���l}On�Ä돺/=��򐄐.K������EJ�t�]�|���i+I�8��v���ڍ��Z]@�+>��~��`�&@�
x��e�Mp@N:�W��(7x0p�VGkGX.�V\m.a~�c�QC2��B�l&�N)���H���!B�.��5$Q����g�4^A�"���e�0ݞ&�*Ŧ�#�6}���>{��	`��7�c$.��"Gf�)���.f��B�b[�{X�$ׁ�됅E�,���f�n���#�]����R���077	69��':�z1�Y�8��� �,�B���55i��+f�R��hgn�����%g��I�G�^�����n[i��wnoo�A�l�/�j�ģѿ�Y��K
lGP0/#m��r�����`[aj2_bpb��е_%�����"��+�=&r��O3W�^O
�a�JC݈�(		 #<̺Hΰ�hwM�]��a�z�~����$�V���B�]����d�7�;�
y3��`�+W���)��إ$YN�,��z�.�F��V�e멤��,Է��m ���e��!�_]�f�A���,;n��pAg:��n�hD�ZK��njJ���F"�	*Zz+���Z�u���S�A��M2kؒԍ6s�罝ݠ�ftv!���v�//�d�T�J�%q����p�1�M"�1V�"Tl#��(L���C:e���ҵ\��O�,�te���#���LjK,�S��'x@�L;��Z)�c<����n��]�_�hS��n�~���h�Ev)��y�|�������v.�?_�>N}i+����B�Z�����ZI�m�9	#J���G:�ȵ
M�SwhNW�z�/55$��N�Lʑ��̗\ �
%�̋(�V�����ږ�������7��7o�����W��RJ���9g�؃)2�B�c}7�sc�#�!|2��g�pQ��](�ȃY���H,$	�ꮕ\Ʃ�G%(���Z�¡k5�-Ǳ!��A�oo�gϞ�FcP	��U)�H�ʺ��I$�j%�2��P�6�kټjs��>`�_��vh��j�L��4�N=rK#�J3���oL�Zx�aM�����R���Ե�V��c��x���YQ�\�m�Q��%I�N�|�P�m�0=G��ۛ��߽{�ß����WU�W��s#�>x�Y�BMK�9���]y����pn�^�#'Z,/J����32r��,t��ƈ9l|~xpD�|z~��˧���^�>9����-�B����c��G���2����=M!�\�oP���g"P������`6f�o[�)���x��7Iþ���V�F )0ֺ�[F�0	��RР�(9���+olmr�]�s���M'��������v�������ɋ��&\L�����8�����Nuq�X,S!p��N����tu���g?y|��:�^������^�`�IM7]{~yA��E��.�b6�L&,Z�q4�\���F�]�I�7Ho֨L��olln��I��fE��8}��'�x��l*]���>�l�P�
�U\�i�l^�0u�<r���
L{R��m޵n��F���X�����g�T~CJ�OG�� �dE�ïH�{�ؕ�H>4��M>(����t�Η��xͻ�tԳy����1~uX3A��5I�J��p�HA␚G��+";�;]�=T_�<O�?4I�ɥ���/n�b kN�K{2�J<�cur����|�2�Bq��������I�  0(E ScF˂ ��9�,�����L�S��T��ʥ�>�C�+9����)��B:5P�������n�fA�)�S�G�.�H��̹i�m�Yu{p3��NY�n���Zem��n9�V����1�Q_�`��E^�1�vf!����|����ڄ�'���C2L	�n�k�)<���@���:�<�]^�ҼZt�]�E���W:��"m�
c%�0=�˗/I�nݸy��}�%�kZAN-��� ���Ř~���l56��-K���3#nN��E��wZ��4{k��5��u�X����#��`�#\�%�X��,Ģ�F�$d�]�
��i�o3z�L[����� ��/˃��'5�Eߗ�e{�f����=/�wBB�Vc<g<ȉ��xDۓ'H�$[v�����N�K�%Y^�z���$BK�\Z�N�3m����7�78~�9�8���ׇ���V$h��	
����aJ���\DI��h���-62�F�:xG�F��{*�+�J;��^+}��֖Sp�BHf��
�Z��_�{D!��؉ ҁ,I2��&tƁ�E��.�:��;)a���BF�Vc�6x5	���^�jG�e)���V��>�F]h�m��љ�f	�&zB���EL�����_fo0f#";��/�r��	�SǇG�Gde@ܺ�	�2`gh6q0X��7�H����&P��K��i>��� a��2)3h�6��y|�X<ri�mg�dLٝ&���'��e��0&`6�r_��gA��\�7�z5�Ѳ���##r���X[��RGp��c��
[��T@�X���P� y�-T��`y�ymsr��v	!�|"�d�/��H��/."�kR7ȭQ��H��m�����3d�I/����QD���B?�@�y�xG��
nu��Md�K����2�+�S�/��֧}�CGz"(DN?���%�Iw_�2�p��� ZR��w�lS�X�����JۜY�R6�m����w��~��!Uo����1�$��,����n�	sլ��]�y��S���p�ZY�!'�"ʭsN%�F�ݾ�[�Rd�ݙ�4���{�6���Qץ��ڨ���ܟ�V�FK��"E�*A��L�����Ji���̳ʴ@�
_&`�*2�G�a�r�veuuccC��=�`����F����W�ٸ�w��v��-��r�9�ON��CO �R�΢G�g�3��Y��t��8���E�n�8?=�h���h��Hz�E����7�~�?����A2��==i�ˏeS��C��D%��ՋEl�­�R�l���ȑ�,��ۜd�M����=0m`��p��듟3E���,g$�ڙ/qri{��ɯ��c���ū^+B�6��Xz�Ν����QW�v���m�)c�rδ�Ρ�{\|.�N|��ܖ��Uך��<FDv�lɈd������Fa�
!X	�#8�{{{�O�"1E���̃J)~�f"	���D�L��V��b+u��S��{G�킛�6V;�b�t�S����L!�[��ۏ�8g�(�ѭ�J�K���U�j�B}��6�ئ�g���y��rҔ�8���g�&鋶w�
f3�~��t���w����h{{=�x�F�ekr�M��_�N���^ѐq[w�?�e��s�w�����z��%[��2'Ͼ�����������}�{��ގ�_9œ �P9Va���;�@Ļs(8�I锅�Xa�j2>��sU0*��ك9�?��O��ɳ�>����� �f�� -9.��0K� �1��e���7�\����kX���7O�G4VM��8��VY<45,��ʒE{!��d��m�S�a�F��R�&LM�I:H&��fo	N��wM��p�F �'`��Ç�V}���7o����9t�xq�N|�\YD�E�ţut��TU�w����`��uH��w<πE�"��g�m��z��v�D�Й�(���4-�(��!��Lae�\�2�(���lP��9jq;N��R�e;��������>G+jȣZ�� ���w	N0.d�`�᮵R<�Xp��7��MN��6��<v
�L�C��˗��w��F��' K�)�<�++"����V ��Y^J�ܻ-Z�a�	�|H��-?崸�$Q���a��̢#���:�BĽ���V�R[HYh����頷L'K,jsۗL��p5�U��P" "]�ۍ;/�1�%�UV��:��� C�wX�D�4Ke�0,2�:�l�$S�k@�������=@g8� �'���(A�JwN���:JC"��~�:�RzL�0�}�嗘օ���&a�l�xP�v�JXv� ;��l"�	TQ���ڎ���b[^��T�9<V	aU��& �M�u��:S����>�Gh#"�:R9>I�*^ �i6Ԇ}�mPv`�*^(������H�
U�[^aK�	¿�ŇB���`�盗Aù@�Q���S����D�����4_�rqI*.�l�&D��ޙe�O(;=cT)���fo�H��~:�VP�dy�I͕�N����>pW� �m积���S�b('3ْ@�	�B���c��A��b}����7�1C��̂��n*C�������Ļ�������v�HO�}�:'V�ly�@���TJq@��}E��坲�a�)�z,�U�Q�DK,,�T,]�Xn�LA�6G�H�W�AҌR�à���T2V�ӗ�XW(Ĳ��@JO^� 0�e}�	�V�Tv�h'�u(���#��H�մ!X� Yi'�' (�
c�6#OOk���𚵑܆�:�|j��*  V(����l��rq]D��>MD(pKJmij���?�A�@�Z�)^�N-��ES�L� U�0*$9S^3�w[��"ʊHS�h_�*ŗ��ɂ�	�N�姜r�.�3c�)�v�#b�s`a��tx�K�rl'g��I��f��Tc�PR<SX15�T��t9y�P��k׮џh�i�&�}U���i��k�q�DP�K��'+0C;��ȴE�Sz�N����#eV�����u��&i������;����?y�<=�LQ3��`Z��T�jK�� ��Ҵ�a�S�L3�3^s_+%p��N���'̮�{�.�	E.��׋V	w� A�"F}2�&o�D�Z����pQ�N3�p?�"��1��	ŅU��� ;?_��%��V�VF�mā<"~�����{gĸPp�蠍%��P���6�@枊�flr���$�O��57#�=�K6�6���I??���j��u)p5��DH�p4�Τ绻�(�|��+:���P$�����X��\#����(W�3=P�����i��U�`���(; ����U4�(m�9��ߎa�㹜�x�_�AE���@'�U���=���#Mf͜�<�D��O|A���a��M7Sl������9���dA�o���U�����ݻ����	f�^�IHۼnQGf��յ��h�e�?���"�I.ˋF\Y�[�KZ��`Ę��c�s:ȼ`�s�I�1g{w�K�����i�;��5���+�҂�M]__���<"�/��x��[2���x��F���9�U۴Y�t��6h�!10r�bs`,;EdZ+������0?�=�AA�l-!� $�-��Qgϯ�ʔ7Ň��;�nlm���P���v���i��H�dE��`��v^:i���EߟM):ʆ���˜G���Z!�"�����U�O�Q�y3X)�Z�Ρ.2R��'E�w��I�E=g�gc�z�x������J٬m��Y����X{�K��\l�әO�SW�P=wsR�%RER�'�a$�f@��/6���GH�@����E���H�t�HYMR��C�C�u��Ny�z���6i$Ƚ�@���y��������h��{��p4>ܟ�&���/����>��	4iQ,hl�M ǣ24�v���G�l<�L��?��v�ݨ���<<�S��X�N���`f~����<6���Yä��;����������k�:Af�D���5��������A���v�%R��3&H�������f���Ն#;VR�YJw�//2яӴQ��BqҚ�FV��W�ՙ�2���C���o����1�����`4���}����NP�c��͆����`2�)�YX��X����+I��壽���lf&9o�=M�8A��ֿ��wϜ�����ki��Gì��Mo޾���K�Rb_�ܽ'���0`sŭ�f��"���8��җ�c*�~���3=$��{��2vu�#Hh���BW�y�G�ۂ~+����!���vb%�8�B�u�ͨ�̣d�7(3����dw E�@[�ˉ��w��|0מ�6���p�I
S�+���c�V�^�l{Ѹ�33�
�D��"ڎ�x� �w���oݼ#���J�y��q�aA�őv����䔥���qx�8�J7�̸�M,��><�i�/_>w�^|��=ĺB�)���&2j3�����X<e���	el��B^�i�i���������|(�7⯅fT�2KI��H��V70�%�0qg�a:ͦywv�A�x���M�X�\��p�/����:8�4���3�aY��I\�݀_�7/O��'ȸ��4��p4��h7���	|֕U�0WKQ�z�a1u�7��X�-�R)�Є�?���Dc*��b�ٷ��Tp�#h�z�~�YX�����C�rX�.ViZV�:��k��j^(�>+"
L��9(sC�e�-݂���xd�5S0B���������j�.�J�T�xɾOS�������vvw線�����f���{�ķ�AօŬ˦�m��^�{P������Μ9s��c�V��`�o��Ad����H�p0,�#z̩"��i:%I����t*�r��c��M���Y�0A�Vg�M!D[P�"9�&���;E.�'�v�#Keh��Ӽ��+�j�'�8T�be�+`xd��b�L�P�f#�LG��^¾�d�N���qa��:�Fm�r��bo�ыLM��wgg����?�5[��!$���}ה����ja�8rw��Y>El�h֖�W%h��@�SY����"�|��L]$�L8�������ɠ'e�~���6�R�:�)��Mi�
�SΣz�Y!L}ya��L,���CKa��t�]����8z�
4n�	���*#����*�`p�f;y�ޭ�cX�L�^�Ua�3�?�J&�$N�AQhqǲȦdS*���U���R�Hnmᐵ�v88���er��ʘJ��x�2(4������sK7t��^�7v�>3s����������:焰~P�Y^���B(�5x:\���q\g�I���.ʜ���ƴK�"�1�Y�dv����y�s��y a�LA26��y>t��tDa�NA��Z=O��';���L~��p<�?���̴ƚMC$�X?�W��q���a`)�TM�=�VX����5�fO�i(�DX}`����0������4��K�p�&#m��&U��t*�Kk.��v���xr��Қ���1T����c�I*��V�#5��x�tZ��x<�����b&pc'�&$wV����I�� �>��n.-��b)�BH���Zl�*m���d#��.���D�`{N�:ժ�7�����]�8���`Xf֚��k�#
ґKp�q�z�i�?!��3k ��{��l:�BqD�\(�<(B���?����"�e>�����)���  ��IDATW(Awj���3�{2�]���C2�t�.�膙�9|���.��Vө�Ӝ\��!$L�$EY�;�$7:�P|dnz�q�!��4;���Ά(l�ۦ����nx���[B1�y睗^z	;37�h��7��;��Ȯ)9 d���$��E��ʴH�D����i��K�v��;8H�5���ᨮg���{%�P��	��m�{/d1eksX�幥��U��_|Q����|�2kmU���0O�`�iw!�R>_�d�VC�I�D�!p3m�+�2�,���!#�z�mh9Vz��a����펂�$*th}��P�x�eKi��ב,BR|�F`8��������h&�O�9����ֽA_��u�Ju-o�hmmEb%!;Ρ�&�a�ӄS8i�ɔ�s�C����pFzC�j�d��M��y?6��u����&	��C���]�ݰijE`�?LZ�B\8�7f������BKku����!��J��l�^������Ѹ'��M1Ђ=D�%��C�1�2���a���=)��J��@\�u�0O$�4	�����=���b�"o�q$���Qc��]�!T]��WYi�?���?��s����`#�����ѣd�ް���"��pJ�\u�)��D�SK+��O��8�LE?	 N饈ǖ�qCkh� *��`N��X��G�����q�*5�},+����G�:peXM�qRB������㐏�'O�A��}�S�����ʽ�*\����x]H�Z\2��ʸd!�3��o��(B�t����'D?�/���?���"��<�}���X=��J��6J��X\���!�!'�اԒ��w� ��Q��eT��k�/]��_1�
��P��
	hY�}�"���RZ�O�������FJ����237{��yiȕ�8��ڂQa74���Y���'�����p��e �4+�̥������.^��ؒ��'�\c��K��L܁w�����	�2�����P���s�+K��<�F��S��	�$S�V&;�C���s���X�wOd�}�溪�)�8Xh/��Xo<���F��Q��loo$�1���(���U���
PQ�v����Ξ=K����
z��-��[[��$��G�δ��p��)�ʧ�2�泸�Rf	d���QTăS��f�J�aY��.8c�CY�)g�/EN�ʫ]���a��"�Fᨤ'�\Y^�Z�TA��k��2��ĉ�t�>j}^myyOt����)����[��Z+ܸj�$=j����Dg�x�T&{�9�g3<�dE�5:<��D�����J�Z� /l(L�����W2�޽�u���'���d3m�䍑"�����@Z�#�a �{�lJ���Ƹ;�~�-ךG���;8���k�_�Xg�S*��T(���^N&S�rqBEfI�b_�3�8�5�i��/����/�{���T6:�2�7A�N�H�$+�����ʔ�a! ǣ�m+k�G3nJ�ex�©M����WM��Y6��2�B�[FP�����fE��3vmL��˥�e��`8�6(Ga�f�BS��j%�)}�X9—�X^	u����텢�if1��(�7������Ĺf?Ay�΃VC����C��M���u���CR��:�-L�BH��-��'����%��q�[
k�0��.�S��8��/�P#ZKY��ɕ9���j+i�5�o[V�)�'�r�`[��[_����<R��.�w_<N�y�p�Ν�@Vն�7�7��}��-���.�~X���j'�����?��cD+x�����o*$��>�4�Tx�`�~<`�>����Z�-~?��G��HB�2�ͯ�������[��s��	����1äy��|����Xn��R��JG�$SCJ{�lH#A�d!�i�12:x:��O���Q7U�h�p�O�
 -��56�?�x��(����8��4ˡ�FjApr:m�V&�DͶ�&>=�2߳�m���RvuE������<h���t�L��P1��@5��D���ù�r@PL�x�����R��QVãq�GD:�c����#YZ��cb*�e�8';k��L`&R.�	�oO���v�\�7���NRv��&{~ـEG%�?�PuET�"pؠҩ�C�������Y,0m��7d���Kѫ���ሧn�TQ�ktI���)s���c�	\�?r,�\Rt��e�/�ܣL�R�3���& ��e�y�As7"��S��Aۣ�p�Cx85��������C;=xp>�Վ���J�,U�e�جߦ[��Rba9����:F�չ�̸��g�z�_��$��	����2�N�J�Ɛ�;B�6��Z��R �I	�ڍ��o�=��pa�I�Ff=f�A�S7@�$̓HC�Mo�}Z:�� ���e6�a�"r�JCL_~�%�x:�}�6�E.�[N 9���X�|M+����]��VI��0Ƴ��9����Cv(����J8/=��p���S'O��^�p������\��փm-uK�
cm��{���`�U��
d��)���h}�,ͪz�Fv|��AY#G;ç������&���">&��h ȸ��RC�-k	SG�H��\ۙ�9�c;�4���e�8�bjJ�'~˱5&�#C4�Z�<��T���<��������5�e����BC�g��
k����{��lc���<����	�.w�5�RWe��3�(�R��ϋ�d�ba��p�M���VWWü���+^<��x.��>�P}3M��d�+͎�a�=-��/���x+���бԢ�g�6	2Q�&j�$V��"�ot:�n��}]Z]*M��F�F�-%_<����5��Fcv~��U�����+�E�̼�ͫ��)
u��q���H��_A��2�ȃ�$��2��<E27׬����r:1z҄���O?�#�'u�,�{c�Jc{<�'�=��,]�+p8^zE<6��~�!;|YMu���A�s3q㥌C5{�:�m.K�a�����AofA&�����&���r��Q%��X��q�:Z� �Rl�ʲ�����N.!27:��H5[�X^���?�D�%�a+ʌ6�pVY0ui�h5el^���di��f�:3s���co>x�w��O��k���牰���Fڌ�/M'Nv]�ʂ�ejJ�8�����;>$�4/���<���N&3��[oH,t��1<ּ���K�E��5�L��'b�jF�b36+$y��h^P���57ɚ��,�_�3�z#
�T�:�$��B���s�:�zsiy�^LXJD�K�n�QƤ�b�X�)���݅�`M�/rlc�I�䦠{J��V)����C�tX!M��vLO�N5"!�f����5�R�hI�2>*�c:$yZW,����Ya��)o�f4l�"Wd|�$WF-�+ꍚ`?&���\i�����vg�P�#��X�'N�ݔ�(K3�xם/o����?o޸!U~��g3�m�Z5�$]����(���:ǲv�6��i��s5�C�Rx����{���#L�<�N�Q	�]*p8e�,]���F5��8�r�޽{��%� +w�h4fFO�P��lLc�����4�CP�qh��:(��ƌ#����d�����ϯ3ӝ�����8Z�aq�	�Xd!��y7���c�zظI���`�I��{���hZ���p���NUY��ʀ�N�o;w�!���*u �E,���zr�F<��**H�٪8�/R��8�]stX�$���
S��#�X��ȡoX�7A�l�ð��d̫R	ˡN�G���3�n�.������k��<N�bcC��Cl��xqy����e�����8�<��}O��ة�0��i?{
�G2�L��\(��r�@ ����Us
�p������|����z@ �P:�k��roI�L��\����|�,�E�יnh�[�粂M�����F����� �wmu����&~�����e`�����y��7�i���ZW���p�;3�x�=svzf^ݪ�`bzLm�m��e ��ڵ��'y*���P���HJM8/���鳛PP˫�����>a��	���׮}�DR��Q\a��\��
��˜eLxI��M�s5�Tqp�	kSIxE�$.�*��/]|EA���w��
�@z��B��ta��h��w�Ҫ���oIu�Ʌ�Y�n����䚗��!����k������)Пh�gF�\ݧ$�JpydA�M*˶)�0Ppkm<Q.�x �e�8� �v�;�̴g�f�i�~�^o�N�������֦��u8C�5l�G8��Ț��So��m�(�.5qC���(�W��±g��8=g*.��EŎ�ˉ��)!tK��H@����J���L3;�@?�2M��-�"�����F���1ҧ���O�U?�;�a�r�ӹ�Y&]��-��H�M�����;W�_� �pi�T:o�h'8-l��E-��t��!}h�z����z�֮D]�����2ǒ�C�±p4�;��i�F�
�׋h�&޴�6�Z�	�#ZR�V���`�#�e�"�|Z�?�'��N���O�$lD��;;,��/l}F
�q��%�(���۷��Ё��0C��	��h"��q:�]�s#����u)ǩ���0�$L'=x��-��=��;E8��c76-s�ғʤ�c���P�c�Ç��h��� �!���7���Y�2��fk�����փ��F� ��Nm뤦-\a�t(E�)ƃLG��&�)�'�!�5�|v�v�W�(Ayð����op���L������>�k7.	]����X�B;'k�3.�u
A�$[�N YP�"�{�Y�˦�
�^�¹�򬘌��HK��#�+��_���Kal�}p?������#5�BU���y����M�1��Ԛ��"�V&xj�j6�[U��.C�yeF�#�4���C�9	^p��a:�B��&ntI�M�It�#�������.���}�k��P�P�Y�ٸUx]�Q[U>�'5�;��R�D.3d�=U��ğ��ʇ�&k�JguF�������`4� ����/\8��?����7o&��zC�ĵ:�xeN(�9ł_���B\�E��+�6�6��8vR���N�����)I�T��� |�R}X��Iæz� �to>:���u�=$���� ��?�i�Y��И�]:'<��c���ȓ8�y���8j�sB��t�R�A���ϖ��o�Oߘ�%J�_~����h �˼���0�����D����^3?/$z�s+Z�c^-F�+�8�9�Ԇ>����~e>,�#����5s.^�h�G:P��h�2�7����8����P����Y��
�F�4,���n�(]L��o/����u5�:�zN�e�dH�<ro����Q_�rP�����k�}�3�g���O���n߿���5���CV0�j �FV�WCEg�и�?�6���-`^r�l�D!�I���;�&o����Pz�R.��˕���Dk�ŧ�� �d�&�ςw�9�
	���~B?��b$}5��t[��F��<-����c�=�W�a���ի������73��)d�L-S��/��� �Ŀ _J�2�1q<n,g���=�ڙL��L�{��j�jj�Q���R��LG�-O7��|�yfK.
]�#���Sڢ%�^շ�*w�W�(�ӹ��`���B����^3�$�"��EB-�Y�dmI���M��R��-O�P���3ӫ�g��%�\X^�$��8���1��T�g���";��_�t#��Oj��2���1�q���ׯCl����'4w��ʶ6�Bu�X�.\�t���_�7x�"G���K����z�رc���|��1�г�z�&����l�ZF9��-3JK�Μ���Æ��5qersJh'L���+��f��J}�ҫ�fk��{͈M��tȔ�b9sFkr�4�w�6T�h���W��o�g�wF�t�2��{a`�8��X�Y�Bn3G\͈�\�Gl���>�3K5K/U�C옏�}�nv��w��3<h�Z��sd��/^d�:pD���n/W��ؠ4;;;׮]{��`��r?��s�/_�{oܸ���/?|��Q�T�c���X�lmC�q;/��⅋���o��ą{=)���J��O>��������ۤ��2�ېO_y��;��[�N�(,Y7:qrC����xj �"WS)>�]	�̹����?�ؙ3g�ڞI${b9�����,�����Q���º)������g��gϝF(K4�tl��b6�*~)B����~���N�&۲$Y�y�+W�\�t�Н�g$):$��|��8���_޺qOJ�$r3v\����D���`��?���f&t0"��Y:&D������\Q��Ru��K�������������QN�y�5�O�"�MP*H<pm��ᴞ�d��?��ga�$Tl��F��G����Go�4����1������}�1���A�����q<>|8��Mx��Q=Â����^�T�>bԫ��w�H�]�����B��Rᦴ{J�z_h����;�?������d3:����ާ�h}�,p���u�x��OF!G�^l��:\�q=_�������$�o�p��?r"*��Q%@���w�|���O!��)���J��E):��@�s�����>����Ǯq1�q�^݃�a��m�d��dE{�t"��ёj��b"2�g>� 'wS¼�ek�(�n�S�����Na��q�wFwR��AD�}����dZ�Uwn8(n��M5��>s$�]�_�gj��r�`{{;�\c�c�ay~�B�vsA�{F��]{�W�Ee^6�K�rΫ�l/7B��BLF�'N�666�ݻ�+�R"	L;�8p\��q�VeV�-V��"��`ʫ��<���:���B�K��<��$B��9K׈�Ŗ�G4��Igf���s��Q�+G�CӘ����G�!n�3#zfqyY,�`�D�8Zy���I���Q�D�*���'���sR8ʛ7o6ZuB��q�h��i��T�w�}"��2��Tc*C�-�3:K<PE�^�p�����Gc��
1v�ң���`h�B"r���?�y����^3Ď���������,w݊8���|�Z\���y�_�����i�'y*�2�y]*�X_�6��"���(y����I�z(����k2�Z[_���&K]�e<qj�H��f�B��Td��{44� բlZ+|���嬮,
|���>�/�G�9y��vM��6
��TPI"����k:�T�K�!w�-���v<bẁX��r�}����(����uo5�I�	Nl�hK� /F�d�� ��[MƲ�Tը���\3�O!;X�MV�ۘf�#[R�#��Wܸj�dW� i_��]y���\Ll��!����:d9h5!@��%-$���3I<x�-�t[��^ i�Jɏ`�N���0��w<�y�c�8s��$���y�%b6!q]�L�����}��S����Bdk� �(���\L�ΣBz�����v�0��7�)�����u��[��������%��,0�8���z�cj��G�x�7�SҩI}��j�Ãx���&�f�\�QkJ��Ē�C���{�^��}���~��d~a%�
SQu�U;���Mi�s�r��>	N��Z���E�wx�7�\D������{w��ǝ��Dl���/�(��i%<Wxi'�d�����Qa���>#|�u:��	�y֥J��߃�?�&�q��H��ْ�U)���ōj��Pȳ�ֶ3Wo6%+�peem}�X�7|���dwo�N�:D6je,AU<�dVp?�[�a=֝ɵ�.��f^�^�Bw�m>U��+�6U�^!�~:e��� �f�A��N_Y�,�z��J��8� 9P�c"
:���DI7���)+�AƌNbi�nkfqn����$�˴�`av�g�}�w��ȎOF�tX,U���S&�]����i5��q�|g.��D�#}��%4}DA�2psi����"��¸��wD��#����g�����aޅ�It� Ń�@�"ɵ��f::g2=q���3g��Ή��{�����@[��4�8׳��������L޾}[t��z�;-��1<�s#����������#Y�1b0.���D���FCl�4��Y�:��z�F��T#Lbqb 'k�S�#;g�&b���;�w��]��G�]7�����.��=ߪ6O�bI�F�0�� �J��kl�"h*<��(G����w
���z4�*���\dQ��6��
;
+`+H�83��g���S�*it&�7�u��ի�?��2��9�i����#���s�]^��޺�٭[��V�^����&��.]L'�����I��������a8W���⃾���[Y[��O�:������ބ&8<�a�~ϟ?�� :��,P�?t��o�֒��?���;�ӱ�j�c�i�;'�`8гs]}
a��������\Kw�����)�h����,�����_ ���.�<~���_���O�������(�?.�9s��ٳ'O'	�o̦"]��D��a_+%JA����n���y����_Xx��g�����f�\�i�>i�'n�b�;�z��i�^������ho?ȧ(t���2��}&�Cf[L�6��`BY�XlSդ�$�s ������/r�T�l��%�%͋�qC~�#��(�`�`��\�Q�8�m2)tn�{�j���Ay(��qn�����q:e6аl��O�$���ɓ�nݲ���$V�9�7��p�+���������.4[$�FO����3'{����ǹJajw�E�ky����2�)��db����)c;�%�������6�vduH(Zx_
�t�3��T�qp�}��e|�@��0�/5�X�?�i������1��AϘ#o6w��|6����\A�p�M"G�!Q>5�eG��P��5�g�*,Ƶ��j"���iǱp���)~O��U����}ែQ��ٖ]F�R��"����²y�a_�v$���#DB�,�oCoL�?(q��(\9���ޚM��*G���q��t�Ȣ���]��GF%>���T�ȵIZ(e�u�۳s���1���`����HC/iU|�jQ�ͨG޼��L�@�
/��79uG�U�p�=�mo��G�~��}>lA����,ν�=�N��@����ּT�<c��H�˼	���SZ�����$�q�IL+��^_J,*����3W���\�Y�p|e캰�Ax�f��C��I.I��~���������E!OǑ���5T����]��=f�P+$�Q�QI�7��݋C�wO����k���e'm�S��}>���R6�J�1�+�S��LځiFJO)��<��>�ش�'��"O��]'2��5f�tg'�1ӑ�h�5,�E�|�#+�&D��O>�Nz�l��:-UC��&#v1�/>������{��+���}m�p$]�c�bj5u\yd�������Wz�.�	�6����G�2e��J%���q��ؙ�3K��5�,-���enH#��,�4��u,>>N����Y��e�$��GB�Rs��!�L%i�PXF~qT������K�w*G�n��{Ԧ��HIp�S��cO֒ƛ��	���T{IUJq)<^v��[�{à̚�xIQ�U�#Ɣ���z<ͥ�.fܔjA>���fY�p�33��}�`-C���0vq��?��7z��ą�fֈތs,r��|m���˧ޔ�U�})	�J�7D��I�9�Q�W�Ǝ�P�4p��*﮹�"��q���q�ޒ�T���!tD3��Q�V�?��/|M9���(|��@�D_�����C~K�*K8~.�qYI�z��?x�K��,�]��jP#7��(e�xb.|�!�4S��U���TxID
Ki��^ B�:��"_��)�o��rzE�+{EQ���ɕ|#�S��ɕ�� K�6�b���j*]�K�XZS�I�Ҭx��l���8�v,���dI�~��W_}u������v0_I(�a� Y�QZ׼v�\�6�O��XT��a!��JSy�-�W��^(�5���#m�Z?�� j:u#�p���v�\�-�X�*�e?�t�6�*�2���	�'NXG�.;6]��\*�@��T*rm78H���-..��7o|A��,6�bV���NM MuM�YSij��!��m^������tF��=��nll@��(�hDG��J���(����}��t�v0]�X��]d��0�����5g��<���2A��O��5-
�S��%�Q)3[&IAJ^��o������@�e��(�J3�ꩌ��+���ar���
n�Z�A�a���ze9"�s�������Ѝ����?��,1��L���ċ�j��� �~�1޵�~��7�:^�YYY���o�&�[Ƴ�����>�_��
����:3��!�hu�U�nq%q�F�I�=��q����&2�n{}}򶹹	k��@��x���7onmmmoo߹�P���0'��/	]�����2���[e���ԆN�]�i�[caΈ��{����a*��*�f�&$�mH$/!�5O7��p��b�/��B֐E/�E�%4���$r#]`�X"�ܤ�8��M;-]n�i8�8MQ�#�8uey�ߺz��Y����2�"7:���A����8t*L\�̙3w�>��὏?�8!?������k~�$��.B�	��� �p���E>��K���7ue��[���;wN熗d��1��{Fz�J�<�O�ӏ>��}�B��������8��4sPn��p#���8v���O?}��i�?dRs�5�b^�#�˔�<c�M�s����W^y��0����!�O<�Vfqy?�<<�Z�@+4��u���Q�'>��ׯ_��X����������HFu~kH0K�&�|��X���NIo�F�~��ͱ�5H8w��K[���Δa�wyy�����YcVX�8��dm_q��eÛ?�R�Ŏw���ދ�N]�Wtn�� ��nJ�8��7�ϐ�K�����h�.����_�*�t̼yeT7V������ܑǆ��W�\��|����?�;��/��h���ݻ��&����W�Ɂ�*Y�$T���th9d���>���o��o����ü�TT��m�q����Χ`�/'E�N�f+��`�q��qܯص�2qũ!�,���]*!���T\�w
�q���Ŧhy�Ʒ$nj$])KɒYbqU�������ݞ�<�<�Kg����:������=<��~�3r�N��S� ������[��+�zXՄg�yy�۝&�yIc5��=�qW��.��W/��#[����f"<*[��b��s=3���A�E+\�1� LP2��w��k�h�$6q�d��p��p�@W�Ɨ.]����/�.~���}� '
G��/��ཏ�]��s��}ہ.�-Aeb��3L'�����RT��C����,���S�(N�!|���?��8
�M#���͚�~��5��+s�7q����,�e�.�}h�& ��d:��Lة�t��	���0a4� x%��!s��D<����uX֚�"r��nC�S��e�z�a"��ڌ2]*xMM�O*�/=vv�ƚ �����Gr��T�Y��LNϐƔ�R��*�TgZ��2�4�W�L*y�^&�7��P�����?)ʞm(Id��:4�\J5���A^��8�{�^Th�����8A�3-��l�|�g�g6L�h�8�C�h��yH9֯�x�b���Y8���ف|��<�	gI{��ե(+�=�G}��k��t�9y�_���N���e��a�\�<�e�x�8c:����4UO����4D����\��_����lI���N��,x��G�x�i8���Nh�( ��z��<)~�1�ep�@J��7H7{��˭5�ȻW�u�9/�\�zb�E�B�MQ"�ᜟ�YYYlԄa�6��ms����C�'��h4�K�X�Do�߱b�n��K�36�(u��5�{��<�����G�(�e6\i��V���T�ӐO�eq�x�G�d*�����t��Ls\����!�AJ�rp�q-���a(<��?�4u~千sF��@z�U]��vN8a��Tw_�9=����~��J��=r�"�S��Cq���؈C�j��,�i��X`2��%�S���l�CHH�T�a�B�â�ެ�|<Ǣ�3	�7����U�f[�Iml�`0R��I���:>��#���f#��XZ�Ǔ�a��7>���f�~^z-�J�)�jL+�V�QVR���.~��t1�+�Ŵ+ҎS���Qa걁ea���!��5��.���N����d�CCby�Ӏ29<�=|��U�G��E��*�V�H^�>JNY���ė�T�������q>A�!�w�Ղ⃢ݭ���m�H�m�`���i�iKb=�꠩%W!�\�v�aY}�/�����D�Bh�t>��3��>��O~^O�8�W`2e�;���T���f��J�jI��8�F'�!�H�>�� �B"�s6R�2_ݶF6I]",MT�N�:���g$5:���4�:�F���1D�|q��o����o��[>M��ϟꩧN�8����l��N�}����b�����L�*�	lc������8����A�͛�� ]+�?Y��W�.E⚋����ޯ�Y�0���|����:73;��޺uϐ����'��gΜ�H|�,ݸq�%)���VVI��4��������������C6G�3(#������w�����-ɿ�TV3�0s����|�;�E��±m�ln�>��z��n��H�N���b�4Ò���o�*.�ڍ��A��|)(�.<��)ּ�4'*J/����
���'��Z��s��L,{lQ�&�`ҌLW�M�:�7���)�&�:v�S&�g�D��3�US�L3IO&J�	/Se��I�L�z-G:�Z@����%��Û�����9��M��'O��ɟ�	�P�ƅF����{G�_)z�.Lf�m<t0sàsVV>9sfsfn6��Z�6�����_�������+7��z�F��v����K��ӧ6%ب��tyeIz1�\��j5p��N{uiq��$/|���mu5}	=�o���v�Ν�p��\F����������{@�7�P��O<���3��77���:��s8д������Po�.�wâ�o���:�S�N]�pgjv~F�#� �2�Uf[9ՙ?����"p����}�;�=��cX�f��,��\���2�.�~��r�^DhڭF���p��/�����Ç}t=��;wB P�1�B�����v�|�8�"�q�\z���[Y^���z�ߗ���o���0w��4X	���R�<F�-���f�8"8:���F�{���~	Nu���
��F3�#���?�k���(q��������.H�d���D9�I�
l�~i=u�j4&\�I���XZX�z��?�X<�l�kM�al���Ϝ=u��1�v�>B�Q�_�7����[���d�+b�2>�O�^\�[;���[�����筭��t�5�L��[#��Qȕ��.��ZŏC��)hGa����}9��7���$"�4O�l V �.�m�X�aVJ��SĈUJ,]�\�4�:}�J��R�NmV���!�19�.JQ�i�
MP�D^T�ޓW�M�������
�
�(��*jڄ�5���ș"1(D�����>�h4�b 
8r&5I��C��2��9p�(�����1�jO+Cx`�q3�.>&�Fcemmo�@!��7+་�Q1
HtUn�C�.�]��>��`������(<8d�:t1V��;��X K0;"�����.E�v���h<��%�	���ŋ�|�I|�`�P��DS0�/�9K���}���?T6a����'�||N+I7o�����oݽs���ý��L�p"�Uό��ı�S�O����T��k?�T��X��(�|΄���ւZ���F	�B�Y��c�~
�U>�Jd1��Q�d���ފb�&�w
L�Gp�K�&�)�{w��}�������mE��ߑjr�<�6��0Uȋ�D�~?�<f�H6Rʐc��&�`�fmy�yJFR>ʦT)ۻ:���4��3P%��-�͉��J�,���T�5�hB-`��2��͍�kN�`��=�ъ��MX0�}!מ�����Ӂı�
��Jb��ۧ2�����{�W�m~����6�s��b׶���8��)7�B�u��YB�y��A7�@���?���Pk6�i�ˇJx_g�9�w4�iA�Zm�S�/&�>�\'O�\]]!��3N[�R1"|G=y�~U�~f�?(��Sz���#�������k�Zw�|�_p�F�ƉS���@C"t;�Bn��ٖE���ʝt�(fRvg� �hСNl�pp�0ku�+�;�X�)�{>J�ۄ����.�V�&6G�-�}կ�Wy����)�}�!&8��J����V�WiJW�1�F�F9lmZK"��J%�6	��?��@�eګ��ȴB���'�}��E���Ǳ�����/e%7l*/��U�Ū��2J��+T�f���PL�4Z#�j�y��o�U%�pa)�����������/�!3l��>?Hؑ's�*�����.�i+�B���S#��.).K�W��'���Ǵ�Xþ?~q��=& lh{��/i5��U���pޛ�Ռ�kJzZ�4P����,6��BP��y��c�Rr�`���"�%s{}�(��,m�&��~����KQ���x0�xc8�jKy �Gd/)u��>�}\L��o?(����F��,�-����0����b*=���ʵ�apv�"�����j�lۨ�ċ�Lg��KW�扦�1�3
�ovq����1�<�>��_~�%>����߾{�����p�|�,���[��b��Ѧ׎�x_���1��`(���E_|�Żw�~��Ě��oI��x�׹rRoTN��B�?֬�):7S4��)Ɏ�v����S8��ؘ��1r�q��q�/:.tȘoeIG0V�V�R�xZ��P��կ~���}��p�LX��!V��.//�$�:
K����/�Vh�0X;�WUGU�Do;�P�>p2��J�&p3^r7�#/����<zY:Ps�2D��xG#��Ɗ���w������._�,�=]O��詧�����ƺ�/���}��/~���Q�-�<�_�<����p��Yh]I�`-I�w"#�p鄍v%���/Y��Ξ=�߯�X?w�ܳ�>�[Ҙ��u�ĉ�j(�ӧO���ry��`��R��*�`��"��TUn�O$�'&�V�8�4�ſ������'׮]�e)�o���T�m�>�[<!�D�)�IiP8�o���O27��l�0�$����G�y9�W#�|cC8�>��у�䅦�vŦ��0�AI��N5k\a����6S�Wx���?�6A�fckD�^^</��U3?ZTA"
���v�|T��^���������p/v��TJ�k�z�V��1�����/��ҕ+W ��������;�^Q�:uZ���h������w44�����q���܄���=^	����OC��2�O"	��v�pl(c!������G<���"�)>em}�CA?;pO���J��|�ݻ�#G�}�.]�C����������Pj�[�Z�J ��6��B���=���ׯ_�d�X��㗎� ����?��Ї��Ϯ!�4߻w/t8q�p�:m�������-@a���k�Y��������x�s�R7���S�Rh\$���g�'���W�2��!��{��Lr�/D3�:KzjK����}���ѝ��<����L��e�F$���%�fa�G�bԉ� ,���&�c��C|%'��y�T2'N@�j:q��[W�@��"|���\�1+
���n�����G?����Pu����R���Ƚ��Qo�h�rA�6E4n1���M7���� ����G��#��ᲂСm筞Ыdj�V�����:P�đ����64��>L�]�Rk��p����7Z������E�#CoP&� �}%B���P��f+�ѫ5�,��������)lY:���̞��M#�k	����4��"l�8R�v+>�8VV�wf�]�#>�H-,V J���ET�����z��?č������jC5��
Ij�]!Cޖ�(0���*�kD��':�MùZ�7�j�"����å����^���W_}���?���\T��D��u`�p��������/���+�`�D)���Nd%�5��}�a��쿞�F�JP	���C�TD3�����S�lI�����,�.n��)R��Sf{\uރ��"['�/�:�T'� �g����{)-{��92ek�� Ď���-At<2���kH��EQ���4����cD[�j�V���%W��m˼�8PD���Ĳ5ZM�f��v|���!#W;5�A�H]Qz\�ںy��������J*w�:��6]�d����E�4lR�;���<�Y�I�8�.��wE����&���2��s.6�B)]��G���	��V�@3p���p��x��t�V��G��y4!��Q��LQLS_��g�O�R�}��+%�tR}m�����<�-��(E�E�M�<]��,�b2�d�0�9�!�lsItaKeɣ�Ԛ��J�v[�a 'qwW����v�r�`
x͏�xtq�R�i�U���[��#�g�6�Ŏ�[��P�T3k�Z!�0R��tH�Bo�j�iO.^<���4�i%vZ��7�7 L^��xjJ�LAm�9'J�љ��4�j���
mO7D��5%�2'��mV���wP�v�B�˧��O'�8VV
�ae�HP��at��
K`�f|i��H�
Y[[�_��	��(YYYԉ��T �ׯi��\�h�}��T����W�>?����Q�q�gyd�f~�(]���!�a���P�~Ms�gʦ/�yT��z�<>�� 밅�,������>���?���g�*���Q���T�4�f���.h�L�y+a�����g�0��\s�B�C�!���ԝ�ٵ�
pn݋l:���q����&� ���2�Ņ>]�@�>q�%�]�n|N�9͆�+-��^c-u}��w	�f[�����ow���Vs�N�@�Ã'�~��G�+�����6A`���C%�d�i��I�F�B3ujm*��LM͒l��+~h����ln2��$�7�q}&��'Kk��f֏oQ}�G�lmm�:x����k���g�_��c���Lwi~��t\��1ڑ�����l%&�OUG�n�e��M�}z�� B�� ����$H�&�1Q���[�|;���$8k��ʣvS4u��K�3P�ݱ��2��1i
�R+�O6�e$����͐9��V�iJ���r��!P�w���m)����^?4%D��ˋ��l�U�g�w�p�[�����IW���0�0+�(g��_��Z%iB��C�2ׯ�7��t=��Cuy�㵄/�P~2Gs��$��~~~nؗ��Q���ǉ�L�B��8�մ�c���i;̱�U9~E O������n@a"�|ꩧ�olc��p��i:a8VE�^�b�
��P���|2~~��W^y�����.]F|����O2�+�:�������3�n�u;��o|����_}�mɉ�
�y/�b,`�[��u�p˺ݦ�є�>��իW�I�>8���E����T���m��O�Se��S��ڵ��~����#w�s0��N��#2r~{�HW����P��YZ�B^���y���o���/���c��
����Oa	{�a�!x�I�Ѥ#(O�Z{ׅ�ۋ�/Q�O b�9gΜ��0�d�%_�}4�d<��#c�cT�l�
l�� �)�3ݕc��LG�V30��4�gt��e�����/����o4����� �:#��C��]H�̙͓'����8OO)u�(���e�L�Җ��9����?�����78�Y:���ЖJ|9��>�Dj����jq.^�x���K�#�ҤS%�0�M�VL%��#H��D��2�aiy��m��KAI,./�4a�a��ḏII������r��dB�i>Mu,`���ٓ�Nm�8��&.0G@�&<����p���5K�/��Vuؠ�G��u��˗�>������dq �#U�<�쳗ϟ�<uJ����O�e�~�y�{8�Hp�L����sDO=y�%����Z��o����'�~mn���������$�����Eq��_�I���o��`^�PB))a�!�XLͯ�C��DG�����2��u�&�}����w�KI�-	`P<Wq��_�Ӻx؅�C�@S��k���jF)����׌����Ǩj�WWW�����d4�;�����`P/���S7n�/�(}?U�"�䓏�=�󸱴��n7ww����O�O�:	�H����R�Ք	Ua��!k4fW�N�U�	WX__;s����������TO��D�<����Z�2N��i��f��7�2;�(�ۄ�P8��h��p�+�:-͂e�'��ȕ"�ܱe!g�nIo�P4n�xByc��0��IC��=M	mk��>/��k�t;y�p/SK�S��7��@��jZ��h��3�#�&u�Y����3�� ��c������`^~(ʤ�c|(Ƹ�!3P�sz��P3�(1�h4`����[��/�U:k�z��-r�.2M<�]�p�*t-���:�}7��N��&$�p����K�[k/�����:�m�̤B;~b��c����փ��f�Y�eT��q���=ĦpH.]� Fgiyqvnuq	'pxؓ�!`��T�D~��l��`���>{����0��K�x��'���:������sgᮼ��oC��G�N��N��C��`�;���L���w���<��7o��/�q�@�}�<w���?2wV��Ԣ!ˬӪ�ث�uB�	b���+��~M��6?�`�E:�==n����]�(;nQbϑ��u�4�9���AO��HG��6�#�`#N�a�T�F��_E�C���"
�ߓ��+�ڬ,���"������+���Nd��hWsa�)������ܸO?�w���5�X�'X:�T(�$�9u��� ��{�.$��X;?����g ^bgF�z0�1qÐ\R���(|��u�{��&U�ȊȌQ^�$<u����.�I�(A*D���$t�q�O,�Pt�����r�v�8�Aب�=�t�l�ؐK�����O���aZ�(�R]`���EJ�&�F%��o�v����}�YX]�t��L�ah��&�����(3�l*�w��T��ה�Gb�B;�#�?�����壃>|V��޽LS��MU�6��|��S^�@���Cs���d։_U^B� �����N���n|�^.���|E�������밵PPY*�x�T�FJ)�q�B��~�����<Χ���[�ng<��X�L�z������}��/�*|��џ����1\�6^l���2F�Yi�"|ȕ�-`�^d<���	��h�<��9}Zȼ�^KຌU�4 �\�=eT�5:m��<ʆ��z�&����n����e�Պq��!e�{/.��Y8���0�Go������'%T�(z�X%�R�竟�}ƥ/yz�n�j��SǑ,u/��8P:-����������Z*�*#ͦ��	тQȀL\^�M2�u��lߩS�>���0���tP��8�_|���i��2�M���BU�/z �C��$TjՀ�_���D��X�l�˘��;p<b��GrJZ��s-���K7��q��!�\I�,�pr+�z�a�#h�OqF����Y��Vvf[���XX��{�W���6l���v{���6D�D�@��4#��@1Z�����N'�~,�� l�M�_ç�q�`�x��q������\{FV6�[#�[���>��	n��}�~?`}^�=��qpP������T�o1H��@���z�����,�]�e��H�4\�(�ĸ8j�=򈂊R���vkn'�t^'u��"�$T���	�R#S���K�y9���$y��ԫ:pum�IM��PG.���z���|��04�����֠"��q��d��փ�C���@���ٱ�G&����?�R��Q��~a�!��1��ė�J/+��H=x���_7�%p|���j�mk/���G��
ZX��1y���S0��z���H8�t����7𛧞z꥗^:{����J����ť8��.�2++��d0���g�"N�8=��3/��"\�F;!څ
��"rCSmrD@KZ�ǟ|�����_������nR�5�n�������F���T�>}��S����]�L��hH�@����p�����wN>r>���˗/��8ƌ0��Hl\X�Pn����HQ�Q�L�p�·��-���5��:��*�<�e6��'��R����_��<��Z��Y��	Pnb�Ma��lP��6{B�]�x����#�g���(�$���+4�iª	�y�؍;ch�B�6>�LW�0��3�9����n'��ހ~�/���(���������؝����B'gY�n<*P���I�g;o���1��{{��}�;�,-��q�xX��s���S�ݶ��
�w���z���i�5��������4����z*L0ב�k��~QY���+җ�h��"p�������K��Ϗ��X���"����x��;7	��[�ݻ�͗���>��Y�ե9�v�8|�xA�KW��+�m|����&Z������'?���|l�D��96�I~��f_��d2{�	$AH�W�q?��O?NRe��ey���+3|����Q�
�aqց8;3�U�ȵ2��3���qp*�fu���A �����}�ŗzB%'G!�LݵW��5�@l�lX�H��x���xK\���~}�{�{�W&2Ʒ���tX��A���e�12$z�L��影"�~&���C�"�|=MT,�D��,��܈U.�qCd5�X3�lb`f߃�}�a�H��b%f����Q[Ӏ[�t�`A��̵�؄ M%����1_��u��ݻw�n셜�l�c�)� �1���7�6ũ��O"�U�ی՛mv�	���]��.��bp����Ķ��F���2�ڸղ�X�cy<���J#gↁx\3oFP�]����7�.��w��t�[YY�B�=L���.Ĺ�g�c`r�w�Ѥ�j��Ђ�����;�f�(<�������S�?�����z��IT 5<N�&Q@�0Ͻ݃�і/냕���ƍx(F.`����lIQ�P2�G���'��$L�)�,~��x��ќ�}�ĉ��\�^oPs�L��#���ʑ�/E��Z;;{=�c4��Q8R���-�	q�:�W��P����C����'&�J�wz�i�z���hqh�#���#�'�|~��g�|�M����tr�޴�;5�|(xP�n����>�~������7ޔ���c����{�'�\�rlcMT�2 Pi�Ky�[����{���/0Xqe�����W�yEu����<���r���O*��͓��/����و���_���\�@�d���V��ø�����E�]�T��m�'���*Du������ۑ�<\(,o�'�tK�`dOi�'��I��M�__�����U��ee:�yth����Ϗ�&�(�� H'���8���2�D��bY�B�h�?�p0�|�����&J��^�!�$3���ͳ#��S�m�ֺg��;�ǌ����̝qt��r23[lT�g���_��2S�I�_�0���aL!��Z�j�ۭY�~���t`Ma��39�����	��{��ݻ�A�N�[�_���Zy6�~e�� E;�^|T����壐Q�v��|�@W��jGC�`���[�b�+�����敝
���T��Tz���A�߀-o��(\��$���h�&��A� ,������s0_:��ߓf��2p�)bd"�2ל�4KG38^jvB�ĸ��	Rý�+��J�܀p}������d��o���
����̨텎����Q�8��aFSXX�Bs����(��i/g/��%^x�s����d1UZ���<Mxn�V��L,��gف�(ş��z�}ۘ;�_�ج��^Y�q��"U�0�h��\����8LWI�N���fٜ�Y`x�����;O^y�Qk�Z� �;����K�߻�ޭ[[i�^��|t<1��v��w�Ǚ�9۝���o��h
��g�ᕟ|�	��t�*�T6:���q�!|Ƈ�9��&��G7�� �)�奥n��Sv��{��}��H�0�ٽ{��h0�ͻw�Ψ7h5곝��L���&���*M�� x
8�^T`��E�&�b�vq��$uW�-�K�Г�Pƞ�'#�[o��Iޡ��~�=�G�PO����Z*+gef��{����i�
O�b� �Ѽ����ݘ�t��텙�&��w�����[*����e���Qxc�Oǽ�������n��>��z6M��$������:�0;ͧ&���}�{����N�Hg;
�lXT�L�r�eo��f�7��µ����po
�
FE����To��Q�N{��
X ��@ٻ�4���4��{��΃����%^������O�|�����yl���̹3g����._�( ����f,�X ؂���PXؘ��W����1����3g�����|�B��6�1SrXm\s<�N�j�Fzumyiy�֝O}㉗_~�޽�F#>��#/c%#8�P�zd	���3�P�s����o�(T%��s;VX6�8������pp��Wa�,��w��O�oW����1E����O��nvg������o~�vR��C��W�~��ųs2O'�b�5��x��ѐ��ei~��4&��o^}��jሁ�7F��LB'&ӎ{�/��C1��DI/-i��Vgq"���֍��G��/��N��(�>��G�#��#�����R���$]�􊔙�X�n�y�k:�1�RIi���݄�iy��8�Y��.L	���F�#��[�S�=��Q�|e
�����~e���{��}9xdm�fI@���U�� 5�e�S��tB�N��*tAW�~�dg��cu�b������Y�mIg(�O���b��2�i�V]�!y�Qjε�٪��rI�	�owgw~��m�ŵk�pĴ��2��F;�F-K�(5�Z���ڂv�J�%N�c(QAv�R�7�$\Ԭ	`��>O����X�n��l:�����F�؅�./�,-���HoC��ׯ_�9̧�^����J^��|�gF��z��v:¯?7������Ϝ�d3 >�� �+�\�������nH�x0a�g线��/n�z��������Xg�u�z���@������8~\��+��A��fs,3;8--�s� ��m";�(����vZ�c���/尿`�(�H{�"�y�6\lx�E.s����)�X6��mK�>���:~��4i{�,�K�Li�,���+=MAT�L���������=�@U�8F�,J�F�),4:%*�  ��� �r��
q\y�!۱eͶ|�D�P�R�}�ܱ�{ G��2�]������c)
�x��ԍ��G08Z�N���~+��й�k��$�u]��-�ڛ���3�0$�m�"%RR��݋���RH�"#$��( @ $�xoۗ��J���+����/�[������<y̶k�]�~%T���V�b�yg9�a`��F:hR��g`b�w妗T���RT�)q伆���9�!�?���0|v(���ý��´K"�C��R>TN�I�� �v�Q4�ò�)��`������6�\�Bk�X��{9?M�(�KMr�	E�J�LS���zv&��܌�c�|/^��p��oz�̙�S�:�V��YX^b�J&�$���M� %��D:��jͰ�a3`V�X��h+��[QL�w��N_�+O�Y��?�s��P;�^�������9·�����`����v������B�UӒ^�FM� �"��g�e�A�^�t�$HZj(��8oԿ�a�M~�������B���o{gg�����?�~��ދ]l��PJy`����ɒ8�L����W��y~���'�|B�ѝU}��aO%����V�ɧU�_��CH�%�������1��h'f�C���ӗaȌ����H�Wz��0�3���8�x����#��x.d�<�Q������9�u�^p4� Yju~��_M��tRoծ�r���s��sgOC����d&����	e�676 u�?��;��)KJ�gLE����W��z���9�l��q��?��?�<S�}��cA��Gs�l㚶�e�D��<���0.ޑ��n)�P(��8l�~`�*�~�aGs��$�GE壄N�J� >z� ��hc}�HؖbDD#���\�
���3�c�����%
�=ax�T;�Y\�D�_���2��3a����//���P����]�/����G�9D؜��gx�͍��x�O���H�c��������$�FQ<3X�L�R�Ú��ǰ�����ϱB9/����Z�BeQq��EI�`�����ࠕ�Xt[t��;U�Q"�*lw��%�/7�Z�	�h:�1Ho%1n�\�L;Ng��ޱ�M���>�5����I�μ���[��g��&��[�%{4Q��8v\���0KJ�)�*�C���$M��}_��Cj5�P)��<�a�i�嚏���_Ӏt
-2�� �j؈�Z���;�� 0���LjڙQDJG��6���3�ZƢ2����p���T*=x�@($&cr�0�Ȁ�
�Ҭ�آ�r��R��Qn�ջSU<z�d���9eUWS�\�0j~���g��S�,�g廻{{{�F9�e�K�� 0!�_\�����A��n��C��EW�yso�y�����Z\%�G���z��?��?;R8���kdʓ܂�J������E�	��\XX�&z�
��ݼy��뿄=Z���![��'pk�mLR��w\�}��T
�'O��	�+<{�BP�LK<�t� �Vr	-������a�#`��Pĸ3k�9�J�d��#aS����a[%{!x����c��W՞������^��O����3��������ŞV�&�%�Ow�߻w�d(�L���gLVcn쪒vW �|���u^X>_aє�J���E���C���ĭ`0lR�P<R&x����ÇXJ���+KK�~`�r��j�5D6K_�%9r�Kǆ�i����v¨��>�1����/g���uL�D~]�����3�w����+�NKP+���i
�C�}z�<t�(aW`����r�ج�7�j�R��rdeo
�WX���Ȫ_9>�W�p"�/���\*��%g`��%�`<_����|�Me'H}S��+�Y=��_
�+ҹ*�G��t���$�4ϕ�h4�EU��X������'Ϸ�7�����k$�d��5�4V��tMU>���4������ )~��@
a*$��2\��⺻ސG|�K�Æ�����ޓ�X�l�)c�yC��70�]�����|�7���,���������;GX'/X�q'�+�	�Y%/L����W�Il��N�h��0!x)O�:�� YXŅ֑5ū�kj�x$�>w���g�M�
^�/�#ǐ��aӨ\�]���D�SC���p��]�� ���籐��)�U��`A�<y�H.�aP;�N�E�	x���Y�!3�?�~Vㇼ���Ջ�Y�"�}�r�ҥ�$"R'e��ޣG��l�z�P�)y�	�Nsv��~�A�=ZC��_��#�a�e;����gϞ�OE�+*_�ky
|SsG��z����z̉j�GZ�\�}�/ⶆ��XuA��A�J�W��&6jN���eb��������z(
Q9q��<0Pyf����s���C{U[c;��%Zk�P��aqZ�BH���.�	ٻ��nPC�͕��*��y�>�X_�}~��_޹sOʢ�7B	�$������<���F�U<�6
�����f�Rt�%�H�F�m1 uD��9#?0-�pBW����	)ۼ��8>�c)��ԆilgD=B�V_:����$U�k��Q8%#AY
�
E�:&>n*12;`*m�R�E&Ꚑ�%О�6Íķ�'Qn�)��K�/dU�B���C5�8�m3h�oK�c(�7gw��k錙F��)������/+����u���S�F8	I�B�\�#9�0K_�9���KEl ��a;�̧���_	L?1k�0�4�
���L�=���ʥ����i޹s��O?!h�6'�7�)�hb�)�P�*����H��(Vq��a���*@��Ů\�ܐ-B�hF"�]��l���J����'��;%��3�F�F}6�D���R�"+K�pf18��fKx���/am���W�?Y�����a���-���ϐؿ������[lý���<f����������&U/Ϟ���'��
��x��
l�/��/1��+�h����]�X���?��G}������)Rmݬs3S\�1K*�Բ��3�̼V��m$�$����e�)X�	�vOܱk׮Ѵ�
$Oh(������Wf���f�I�#�!����ɠVR4����{�'b �r7�A�Y|E�\�-5<������ש���'JY&��)Ld��� �?��5�=���#�O9!D�Q�Sr~*A����"�W4hb>$r!y���wơ({m�I=)XZ��#�i�0�H�l��es ��?�a;�a�h.���r��\(p���%��5�呿�*U�,�Cy�I��yqFip%���� ?�Z)"�S����g���K r��+���<���r�YJ��Qy�7c�a���a���$.	kU�F��ð��U�˼p�ɲƱ'�L�U��i ���C���^�ݬ��fU*�C�9��8��{~$	�h8�,��^�xqs�T�\�ߔl��KE{j��監h�7�OZ����um�r��c|v�ؾ��ʁ��7/}f�?\��%���J���K�{���ߋ"g������'�i"��r�R��63���g���j�@yX �� ��Z�EBiĐN��a��x��i�p�ZZb�p�8AA�H�c!7��!�wNmY��䳨�ퟘ��Mv�F�KX`X��SN �$iB>!0P�J�C��bG�����H�Lz2VIR�i��U��zE+�4�'j�U����Sl:�U�\�$�q`��ֵ��W�凰5Hփɠ��9�Ta�ˍ����S(��j^�煾=�+u��r��N��I�0����+�L���pҽ�P	jZy����-�-87n=}g8ݺs�D�� 1��7�b�&�h4Nfi�%5PO�>�&pƠS��m�VB�&�ͬ��L�Lq���Y������������%�O<����m�
����@���+���d4Ƽ�?6K�n���,,/l�=}�����j����
21m���lu'����.^�4ɫ�w�tH\Ë=*,-++�E������_����zv`E���S�x�����>f��/�H��ĉ@GM!�������D"Pe%���?)2:6��@4>�"rP�µ+Z�����mRE7�����GS���$6?���P y3T|~�@�W�EG���@��z�?�p�u^��0�z��j+�l���F� �����J=h�L���1
�xl�<�VlZRk�hc/Ϻ�q-��(�M%R��>�� &����f��GL9���,JVc�6���O>=�߇����$�o$$P�x�BH��ג�UE��
A7�Lh�!m��N��]o�5���ndX�^o�64�!�)�5�J����o~��O?�w�!s$�a����0Y%����a���i�_�HuLm�5�!�Ӱ�Ü67�6�<%{������_������؅yݨ�Ku��uq�%A+mP%i�i֡hDy��fkkk��?�>��N�>S�7:�.�4y�`;���.���
|����R���߼+_���xR�^����j���WqsZ4�����3���*�5`2��8ݷnܸwOJ@B~���쿁+7wN-v{b�+�B��	ݻ��<����ԉ��
8��,�t�2+�D�E1��c1:��rH�P{��������H�=���46�EX{�Z?췺R;��P���f�vjc}4�����3~e2�Yb�<@hX�=A�����U",{���y�������ϟg���9�C�-����|o�IS�Z��q;���7�~4<z�3�T��8�*�Nscm-�ͪ��c��4���F�&N���+$�N�*L�w$b]xF��?��;��D��	\�߽����~JlW��)8h��< y<�Ԫ���^<?{�K�_�'��ۭn�t�)����.��wޑ�z.]ZZYi���f��hc�6��w���߿���E]-"f�OĞ���+H�ב��4�CfA�V��Bq�r��VB��3g��{U�ɲ4�J,�Q��J�̕�6�����AH{?��Vľ~�����O�a̙v�s�*8AR���J����҉g16���3�O��.���&��)tD����~�wn~��F��5��m�p�c�W�Y�%���E�(v�&��pZ�-Ƀ�S��+Ν;�kw {�\��T��'7�˒�o��w��hj�$��ڊ�x��T��
�� ?�;fŉX�کӛcY�<t�=�����$��5��TQgi{{7�[��a{f
�K2W��Gĩ"�$3�@K�0O�>�D�(�u!a��5l��a�-�i'0�S��UdYf��5.Y���ɴޥ�V�7�Y�~���b �l��j�I��h�18e���@1 2�����H�\�����:=��t��F.�U/������I��$�j��Z�MgJ�N��bC��\�(�+��K:�GM�(!�! y�Ԑ�ʅ�&6m�;w��+Wq�h2��i��+�����8 �
���Yp�ծnN�@�ԧYycc&_��h	�)�:{��#�(��Am<bPRw�p�i	мa,�Q������¢8�9�k'�1\���cu�׮]����&�pR nY�-!�j�]�tF2YJ�
�,k�+»������W�
���'��7�_�=t�ʕ׮]�����4�m��?BR�(�Ug�k��Fwa���,,�l���I�#�z�
m-�e3��_��_~����柤uU�G�W���c�k��0����s��\����d�� !�m���L-�r� 	�#�ۇ�%�?�seiYڞdp�H�\�r s&Ӊ�ޖU(�2����L��T�>���-t���6s�X^Y��&}c+���j�jAnK@#������@e�5�����d7Ia���4a��!Q����.�1a��S0lf�d�4�P�<0��r`�:���^+�B*�Q��gp�4A�K=F4�Q�;j��4���>�%��n<c&F�9��w>0rWs��x�Q���Aλ8`�7�	#a1;��1Aιv��9L�(�9���ګ�ƃ>�Y��P&���jҚ`��x�Ǆ@;�	��͓���@�`y楆�>f�zP���D�LF�!znj��3�_���Η��H��(�����% N6_~�DRS�Q�r��`��ĩI�	��K���U2:���9�D���ƣ��e��Θ��M��I�Bq���4ԛy_�S��{����j�+�]oSue�e�*�韠���v�V�1�U(�Ꜵ&�杈�2�No���<0�����s=�c�O�9�Դm��h��?�K�m���Z��0AJ�?{g��,k��(�M�[q�&)3554xOJ�V�U+��)J���|��)�![�d����S�/�Ŝ::R[*>����Q� ��D��\����H]������E�4jcI넁b�]e+�r2٘
&�J�FE@"�P�̹�@���h�Uʹb���Z� }����U��Pv���t�ݘ���(���ַ����ޣqI6E�%��n|zSΠ#~�C����J �D���k4C�*�T��+���͑G8�֍����Gs����id��$��dj�;���p"��v �J�/Sz����mhJN;�e�.a��G�)�x�Z�d��݊-0GA�/�ӛ����Y�@2�,f}�j}}���^��_��x�ե�|����*4,oN3ߒ�8̓٨hV��=,��q!t�b�x�@�3{r�j�c�������w��^8�lD�{��Jal�ѣG���̻w�*��T�A�����p���he�ߊ
�	��*������{M��[eOqa�U��۬rn薬$���bL회�����#�n�Ut�lw����WSF�#�u�� �o�U\f h��zvb�)U�-�9���M�y�.����^�������*w�i�;Wk�^>�Yqq&��d�,
�i�t��>C����]J�S���Neh�����,�d>�-U��ټ���+	%�W#�ۛ2�Z� �G������\��p�?��?��3����j+.;�y�{�O���L/u>�<��ƿ��Z�21T�(�� �����
oO�s�,G2�Uٜ�1�!��pE���G���&5!��M�{�?�����鷿�-^�]����^9}�tY#��M,$05=�h�b#�� WXe�榤Φ���Kx(E"�E��� J���w�����<��E7��˖`��`��Uy�edA��SY �-A����������~Y
i�}˘śo��� �ouu93r��b�EB������Li�B����N�I�b̌e�\���THU��09�M�c)����~'x@]5�<ps���� �c��������	-� ��B�16���7oj��t%��hmoo˴�����߹��>}f��ŀ/B�ܾ}�����ɧLH>��8"l���η�kUù�[1�)#3cCb!{� }�)�h<�`�WW�(�$�K��Ւ��^��ͻӘ)���ϴ�M
��p7��]rw�ȫB�ج�?~��U�����>¼}��$,�@H���-��>FY�P�}���̂����3st�����!] ҄\�2�ޱ���ReQI����*�~J��y��>��Xw�K�6�ŷ`|-w�+W^q��INO���{��_.]��%ú��w�޿q�&w#<Y��L�U�	~�������ˈ� ��w�������/��``{P���+�Z�����������r��	�؁`4�l�/4�AQ�hu�e��b�o��0�	�!s�
CJNŰ?�sN�G�(��<C�kQ0�-���3�'��#�K9�Ne<� ���+;�\@v�����$ �(�m�k�7�N��� �RA@��t����~&y�BrZ[[[�ST��\���P�X#ʍ2¨:���Њ	��Ĵ[Z^�hTE{U�[�TSY�<�k{���՗\G��"��O���B���|���v�-v��Y�,/�u80U=~���h+��]�y#�5$켛%�p�:I�6Ҧb��12�c�5�Ӎ;@J��4'����lcR}|�"��N"��g��ى>��}˸9�h\�����?�/�z��ޑM��HcBK�AI��:�P�%�Lz���$�իW?��㧏s�K��!HL�����*2j(;r�'�av�Թ�8��U�֣ �!_t�_��_H#�F�PP�qq��4&wv�`����kl�,����:�@�0]RL���S��+�ʥ_�4s�ɇ8�D�Kt��o,<��(7�D���
�����3�vX__�J%\͐�V*�f��Ŗ��y���	m���cE6d��r���y~R��;/͡D�Z�)Ϟ<��?R)�+��o���8e&����g�z�.ϒ�5����DNA�t������3��#�7�;�Sˬ=祿9*9G<R��1^wr#A�y/��:s���}*�y�����Ŏzvﯼ�'4f��'���SM����t��U^o������E��z7�[c�07D~j���(ف�tJf���_��j:DffIY�%�hױ��.�8�S�_8�C�xG'��pC�X����e�[(W��^��j���(<_�IY��~Tޙ)j�e��B����Ho�[3�S�%KL�֏ :&H��[���-0��$�0��Ò*ڤڨ��Q�桅!�e�UWh��;�.�3��s�IjƟI��{�f]�'�)�=������O��U�p�D��3^���D��� 6X�E.�������R�w��h��b��^��i�N%�Y��wk������F�/�u����j��I�WY��(��bO�'�9�hAO��Dx�e`,�x�<�����ސ*�T�%G����,���9{j�ٳ��d��ON�ބ��t�2��LR+�CєT���CY6��I���d��x��En#;�3�gݞB����,;�}�~�h5�G��֢��ob�HZ$�E�7G�ܹ#*đ�'aP	����潞&�]��'��Ÿ4nrS��,�!7����1Z��s��cv9�C�1K��֯o߽#���.�/�s��4Ձ�s2�y�=�WW[J3�n�����2v�rUv!�O����H986�R�"�C���ZX2����tIŘF���ž,b���5��̕�*����/
���40da!Agl�����=���cju6�ћJL�:�i�)����Z���32�n{���e��b�O���yK���:[�x>����h��ŋ� ��~M���j2+�0IlH���4��Onܸ��iF;�� �����*M��jdL�u���5m�P���r�*�>ß�{�.&�	&	���|Q���A�f�F�2�Z�O����$TG�f:K�Y16�����D���W�g�|���""/��.���= ��<>��y�ޚ~��.{]����I��>�#������i�����g�g��nwk�� �H��oo;8};;;�x1ЏC盖\�д�����}��!Q�j�j�\��e��CH$���|��Ah���Q��h��)g�� _���z��/�]��'����&ӊB�]}ů�^Y��{7���d�D0�Ǎ`7l�0�k���ce51�$đXR�K��S�F(\Zj �#M[�Ɯ0�e�4�Q�c�M!�߀y��ɓi\����H���fQgr8��H+*K�d �BgE���;p��t��Ȅ�X��eA�)1��E�F2�6���%�-�J�R��9�)DU�BP	n]�5����JP���r..	�K���h*�Px)x5ә��ܴ2�>3��ﰽ�ə1��>%ଶ�٢Y�Y���:}f2;m��GO�$BF���cF��Gڬ�~�˗/��K`�	L��`��
��Q��i��bk�[8-g	��<>8���&���9�ՕP��z��f��R�!}�{�Oo�x��	>�gS~J�9���U������{�VP9� o�$�<z|w88�ҸZ�<zx���3E�Z���\��O�^���-����k��4˳�L�t+=���ۇ������YT77�L��1����=)�����QM�ێ�W�M���nªke�٭����b��@d�{�V�F�hxݑ��ds~��g���{�@c�O����5��Xq��p�^}��{�������t�֨�s��:_�����υ������g?�u�ֽ{��5�:~6��hPBZ�g���/^�x��9蹩~`�=�����G}���O�cX�'^O�>S%O"��8w��`�#t���X
��d*�<�z�A:�'��� ��3�b콩�͝]��W <���k� `�Mk�gaXRmP�ahJ�QD6���N�v� K��F��C��OU�5�f/6�H�k��6�l�$�$aX��&r,dϪ{�}�P%�	��ź�2�EZ�W B��4��M	AÒ�w�+��E~*���}��6�ދ��Z�h ����tT���Vz�1�7�r���G�z��/�Y1U��d���hwa��$'T ���)�� +�`+b�Q�Ҭ��i2�"�K�g��_�u|�B_G�&i�bJz4�1�P��P>dV�H#�9����V�=m�h��ywg���3D[��)�X�(���Ãp"`�a�`���-���[��;�Q?�@�|�����w����!+�5�]҃0�ǳ��TJ�js�Ġd�()3�9�9^���j�PR����u�R���;|�K_z����Bbi*����3,Pn=���8�
~r��G
l1��)��t��^))�v�Q��It�|J�r����k׮�o��������&��=V�z��y�՞���%����<�ᕁi��|��=���hc
��]��s��ֈ����L����Q\�~�rF��j(@��k�&0!����@�d�wN�c�����)^���3�dNԮ�mj;,y���9����F;�B�eM�O�oeeI@-�!�$[ݑ4����q���śN��S?G&���>��s��Mc]K�f�%o �X����[�<�s�/n��"�5��6:�ei}:f��iQo���p�/��f��&�9Gx�6/ȡ�)w8�����?v�:Lf�k<iC�e~��]�y,�c�_��כ������P��_���]R(�n������x �a����w�(�)W-�t�J[��|Sݷ��]�b�W����G�{�9��±h�Q!�qpJ�Z�QJ�B�C��u���Qn�Hvfh����Ӽß���5��n�J0�!�L�h��Kh@�j��h �Pv��L�c�o3E)G	��N�zM:����d�	=tV(~QJj�T�����n޼��[��<:��ˉV7�y_���Q�ʽ���Hps1��(7���7��б�� _c+�x�L����-ɊT�<xG(6�MS�&E���q	,��	��|W���*���n��aKA�8�}�����bĉ��Jn�8f�y��e!���[b쾋C��05g�V�u��^TB�&��g�τ�'�D��$S�������Y]ї���L��[�K�a�?z����k��4+�`N��*��Q7����94"�W�
�,(���X�}>��C���w4��*3�c���Z.�pL��r��t�J�L�b�%�z"2i��1�U*EF��a����%b��Q��E3e���c���P�XIӒ�����˝��o�i�S����G?�t��M[�XʭI�kl-��5�U�eRC�R���:sY#�'�0��'p��|�jz��<�S��#b44�"�և�N� ���G���2%��a�Öe䅙+R�~p���c�L��K7�F ���X{���J��ꬨ��$���*F�(�?�ax��=��^X����E����,�j��XH�X�VC%���L)�6��0���zb�V_�x٘�P:0��0lR���h���l��\�كt�ӱ�=�|9���͙x�S�msL�N���FEfZ��Y���\�����ᇇΩ<��q�_Z���r��`l��E��`~WX}�C����,�]�BS$���,+�r�����ΒIKpza >4[m���(0�i�b8-3��(3^,~�V���bX�޽��+�jYw�CyXZl���<�C����E�2�II(y�7VB������;wnٳ�l�Le��H��L[^���[���ޑti։�#��o,Z�j�qx�,�M�F�j4�_#e!��U�E�%��?��
'F!��:K�4N���?�i�`��hu����b_܇����fS(�\3�-�1�L	h�S�eo��&C�Į��Ro!�`
j��f��/��s@��p������0�)�k�u��L�B�s�1���������;>[�6���5|wgGb�����ncc�7�y�%Ը���x�j:�5�V�r�������
/��5�3�s�63�|����VJSq��r ��}0y��7sd����+߹s�!#��a�,�<}x���ZD��8hXG�<<��	�V�b��8�E�����z�ǔ�h��Z�N�W����aq�'3���Y8
d��i6��d��wP=ex���檉	:������k��^����������'4?(�|-�\��������|m�@���R̬���<��W.]�������g,��::�T+ތ��ʚ�	!f��_ۂ�~�����g��ʵE�������LS�ۆ�R\a���(N�5Η��;����qX^ZՀK��p��о��ob��q��X�=t��� �����M�����sm�q�N�� wr��G�/�6����[�L�i�@��e)������I�`Y�D#�b|V̉�wq�b���g�1��~�)Cų�!p^~��ߟ�|�ҥK�/�}mm�3��(<c�|�#�M�j�k1���^�d�&�]��~Zg�1ŞtI00�"�<-L��u��ef@��L:/�)���-�\��I0�J��B�{���3C������塆��/Y{��IoFE���2�96p�G
�N~f�Y�g�@?3`J�JЊ��4��1�w��B=G��	p6�[�b�J�1h�.��.�/�v��Y��W]��o���/����������)�+�#�:�kҞ���(�f�0A�%��a�)S]r��)�M���Qu.�Ł�8%'[	�e�[Ĉ4�*K�h�Y�}<��9��X�l�x$%'g��W�t�hZ6�`)$�Pkk��[��3��4��w�I}g����s�nw��?&�_�Cվ6˕��
����?t�@�%����8W�����Ъ8%*I�z��i�(D��	Ŭ�۳��4)�8(~踦����ock�\N��fo.�K����f>�	˖�i�A[���qJ'�"B�a���_ms����.���u��>�4���^u�����f�Q�K��ˌs�������ǂp�&��^��[�ک5%��SN��U�FQ���k#0��chOD�r;k=�/�Y���̅�Jh$�<��`E*|a�c�
�v:�˘�� 3��J-w��;�&& Q��W�B��_��� ��h�W�7�}��3�,U��i�U�U���m�GeY�\�7�/�`�UiҭV{{�b�{�Œ2>��U��$��L+���	K�h�F�����ͺݠp�A%M�Y^�7=?���A(�r���<d_��g<v;�\a᪙RC%�)ll�
�\�/�?'���G�j��C�Lƴ���t-r:G�gOZҚ���t��Q,���$&���bލ��*lV
�"�EI�`��_�i�.x�i�̆�d�j��*�o��Y\$��V)�q�}	��s�}A�'���h�;>{E�u�v�wqAp�^�����������r=l�n��1�kO*�����_<9������Q���H�H}0�
��"r>r<�؊�I�c�_b�Q�P�
��f٬�`*�*eo��sv��d��,������I��۲�W����?����]/m��D�p��~�G��=�,����	DI?��������-R�����GO�޹��ً��}F%�������i?�����l��=�;���Vws,�L��J�����=�--Đ���2��K%!�1�����T�)8R8��T��q2�+:3�>?r7i�nx�n'()Z�����4�l�q!4�]"���.cCz�Ĥ�f�h�gO�₝�������p�݁�X�\[\^����t'�������%b���\aM� =��{:�,�b��`_Aa��)R*�ӂ����hb��+Ywe*`SK��D�C�9�v�C|O-H9��Ł��(��J=3�~�i�-����O����6�g(+&a��ª���+����Y4����k��<s^<�33}�lo2��ۏ�^�)լ�;��E��Ju�f���EY��<�?x��"�`I������i�ުV�A5�fҡ�^����F8���|qڕ6e>E�Ϟ=�~�3�l�
����),eS��ax�w��ɭ�;Y�j�:<5�hU� �a-�$������x���˟�+�﫯�ڭ7��Z�V3�ݩ�_<|������ބg?dkkK:�B��n�R/�)�b���!f�x� c��t~d��L�f�g�~j��Y��Q��УG�0���!��fk�pee����nB���A=���bWBy-/���tg&qE��	�fJ�)�
l3���6q���X�p�4�5�p�ت5�:���I�y,`�Y*v��*^V�n�Y
���t&�D+Jڠ���p��e*�j�wE0f{��8~.ټ��F���{)���ZNo�^�>{���������)��x���Q�(~y��͋�/��/�AH#�"f�~���jՊ�͔&�~�V�.v���p}uV#v����I���F+V�h��񭻷��D{c�K��a.�����x���O��h�z���JW��bw�����Z��|=;><rgE6I8���U+��h}y����wnu;x����.,@�;�0��B ����%�9��a�ٜF���;jgp�au`E�XҪ�3v6�봡uO囁S;���U�yۧ6D�cQ��j/�z�
��y�w�]<��-%_��ǃ��{�G�=6��N8�)���~O0����ߔ}ϕ�*�J�r��?����(�ptp�s�x���y�|�ɭ���o}�[�jO��k�a�&������j,0V|��8@�v����z�'��{��g'��J����;I���<���'39t�iJ����L2�5"}�h,h݁��"��6df�*K�M���ڻ��9�Ѡ���I<L��cȞ�����Jf�����;��TwVV�6O�?y�gM)���:_�1�@܎�Bse}���;^�ׅ^�S��'M��z5Q޺(�Vr��͕z��}ngi}���QJ��l�d8Q��Ҕ�Y��� Y���D~�˷���DXYr]�q<�&�U��/--J�ew�S1�ϣ���:��4���������Z�\�6Zj����~���ef���Z//-1�RWԶRW��N����������xK=7�i��t�a#�V��׈��cg���',�0��z�$��Y��Ϟ;w���f�C��_��h� 6�Ѳ�,�X�P����+���wW+	&�ѯ����@�!5����`[*��0�Ci��K�Q=<T��*t�ʺ ��8���B}�歷oݺ[4�N��B_�*�ܕ7V�|Yf�C����N��gµ�Bb���ZC*KԽ"�@g,`�H�*P��E�P��
u�s2�y9�&�4Y2�􎥛���q8��V׮��l�ڂ<��B.�wIIk�`�BG������������{��!ԁ���b	�N��k5�A���h��#���F���Z��˿r��)o���/,=8�Ps�Q�{�-:Ȍ�(��k;��ի�\�tga�0�]���#�`2�r�'����N�i�y�L��/m	�b���"��"ц�vi�5p*X���D��fL��,Kd`{�J�8\��Ǎf7���F-_�joiYj/j:�,g?w��n���S�#k�	���l\�xb���L�h,�u�V=:��v
�d2R�T�K>����������r���0�Qg�Y���t<iԛ�,����{|x0�ǭ��e��|�w��S(���|�����8ӧ��$��0�~#��t���0�߽���w�y$��?����+�wj���iv�m��D�82,�;M��?�s�i�U��������ۣ#�3�͖�&�1,�T�"��Ĉ����f�i���0B�ʇ�e�s��˜+�$��F �{Ž�0�	�~%ԁ��zW�g��y&�Ƞ!4����n�����MMZ�]��8<:r��R���o����P�8%��{2�(��]�p|�cc[�@y�>_�+U�2p����0���I��MH����eq����3W���`GK#W|ٸ��d�׶6�������W��D:��/O�aө�N��w���da�8���Zҁ��%��l�48�Q�%Q�Tj��J�jN�zc�4�N�~�yg6��t��Gd��q����ў�|[MG��xґ�rLѵ�G�{>S�r��f�f��T�ϥ�%�f\u$d~�/TPaZE��Y&��k׮A͒d>_�L�7���R������c�u����H������5�w�\�L�ag���KQ繻��6LkA���m"�����i}DPшob��k���?UL;3F�
�9uW�iˑ[��[Alݿb��t1�jY;�8��D�Zn@�3Aj~I#sB��$DSvʕ���C��ε
���gT7v�wK|����HA���"��	їZ㉃Y��JtŴ��A^I�����Fǀ�f��?���'C\�<�R'��L� ��T?�;֘�n��q���ngA�H�v�z�]���+P~ϟ�����h�)a����bu��	x͉��1�@�n��^�x,a�
4K�!tx���8���/��Nz���t�}�T�M�ݕ
�pڐ����vv��={��8�@�~ɉ�{&�3�=5����7�|}�]������[�$���.ƚm~�n�� lɧ 3�����\lB�m��.�犺���]��`H��-�1AG��N�ċ=_=Ry���%�;�s�(�r�f�iJj�V�IE�0�.�f�R	�dG�DL�Z��kg�"² �H��&��ㇱ���#l��������J�Q�jpY�)1]�� ���2�<���[�XX��S,4�)��S����Lb\%K���j-36��-�o��a�
HV�p�0��,���3�_������_��7��ɣJDO$ַt����U�͘}��������J������[��+���)�(�`����B?,��,֕+W�k��<X�t5�={�m�3'{�4J�G�T�Ȋ,%7_6��@�Ԯբ�,Bm͞<y�[8��������`��p<���;w�ѪK�����L�.��No�e�]X����#�h��HM+�!o޼�����;�Oܐ�׬7�^��Ɨ��#��O�;<Ĩ�,S�^��D�ʨ0�SQF)w���"�����ڤ�w{N�2�n�OrM�H���rE�g��\�J�1�.��N�/5}=���l�d̴|���Ѭ\�̠�Sii*x�쨰	a�1�G=�+� �-�>�l��)��������R��{�O�[&��l*Ԅ��N";�"\�r��礱Kư:`k�a2�����d[V�g��6Lĭ^���$��/V�C!I���(�r]�����ۿ������ڄ�۵k�A���3,�Ix*D�.K����!�	.g*�ٍa���݁��}�'D�UrV8�(#�{���<�E����j ���`8���(���������,c@� �xxH��hP��N>WiH�<�����.����IV)u5���d �\P�f�~��i*�MK���9s-\)xiF��p˃�%Y-���ŋ�U
�w;����R�e��]�4GY2���u�V��@z��]�R�3���VL�L�?њ���]�G-���
�F�����wNA�6R%4J��ā�0Ou��?�XS#Zj6����~cc�p�Q��R�c�{�r=�;��O~*H^������&�at�.=���9�U�b�x.=��{��MKFFeMLMh1���Ť�Y�+J�O!-��H�.���g�
o���ކ�GV�nGb
�1��ٙs���/�ٖ�;��yt������@$^}�2~^X�|�`E+��K}�[�7_?�)����	���В�.\|��7>�����P1����Q@��(f����TLF� ���M1�/Iɐ�둦�K�\����چ��y_�"#-I��K�/Y�����DsK�E���p�D��"n5G� �)�L|��T�X�ɽk�F��U���	�n�O�*�'�h}���t���u�:X^���t��iN��R T�u�C���xb칔BZ�����j�0d)O�Uَ���x7�������o�M�;�L$O_�p=s�����Д�N'JcZv��K]��U�V?'!!�+�Řm"���H jI���� �	�Lv$�{K��>�w��پ�.4�K�����-Au�-���G	�n6Ĵ�_���n�u~��);�v�,���w|����Teq]e��t.�)��Յ�XI_���'����w�jI�-B�w4YX4��Z��"d}�;�!/��]��|�G ��R\���y�2CM�Z��#�?����J`M>��ƞ�>!5[���D�R�7�����w�{��B1������_�������s���d�ck�m���)�@��d%fS�V�E�"*aSI`��[t�CwhME}�ѡ2���@E^>�5L����a(�֣�Gp2h�J&�G���V�=�B����2*繁���Ӷ;� �S,]�$Ő��*�9y�艌��N<���x��p-3Ul֋(�ȝ�ɵ�`�����>�L��3l��?�U!���01a���@w��>�s͇�*�9f�5���D��d&��D�|�`���ۚ�Ԯ�~JM�u��uN|Z���cB����Ծ`h��e����=�t�a]�<YZ�&i̾�L�e�,�f�ᨯp��_w��	,�26H0�Q/�>�%N^��z�pB��:{�6	��HMО��O�zX��1���X���o���I4�n��|��0v��[V�JǏ҄Ri�Cr�_y���h�%R���u��y氋B��ap�ᄊ&)-c��_	�*@�|�ۅ��>>8|�d�ۆ��VjR;��J�N��ڵk�K:h.`p�x��261&��V�}�_��ކ:a��&�%���b�>�ڭ�~����Uu ����~�o���W��e<Ŵ�a��T����Ĭ\�� ?��f�bP�Xo|��O�V#���!H�>�X�G��~�)~���=J�a��L.k����,+l/�H�TO�3�$�,���,����d[=���{��/5/��KRR/�,���:N�z�K4ʵrS��n��
bMƘ�V�fɼq�i�Z*�Z��U�g�?//,*-�D�#�z1V����0�d<~��1&�I������/���M����i!Q 䌜h�X�s�y��`h�^��ƣ
�"׊rWU�ȕ<u��d8a�M�@	���/~Ί�K\e4�ڕ><$�yǵQ_�t,"|�s[;�+��!NQ����w��rym���R2L�\@�~���\4Jr���D!7IYx[�Ͳ2�,�����Ç���4~>����j����|Gc��n�'�Q@"K�(?૑�C
�&NR��e��߹s[�s%�s��Cl��r��KY�k�>�~G�
�KM}�J\S�(>�,#76��d�$��xv��78<zp�n4A(N/Rvq��L�z���os�T���	�-\�ŕ��t�.4�R�3���"O�6�n��|4�������j��bN<����g�k�OB�;�5�"CKW!è�1Z�\V������wp��y����3���L5�U�ߟ��4��Q��������9!�xEIM��$��t\x�� ���G�	�=զ�6���6_\\k�Y����Ԕ$�}\�(A��n�ES�_k֙o���J�W����g�N&ݮGQ��MgiB���p'2e4+�+����0(F/���@�z�}r�ܲ]��[��i��������M֬{�:&�3k2����Iu�����_~F�X;̖&la:�U4N����>�|�2�.�(�n�BY���T�'F��43������B$��ǈ���ٚA�l��zꬬ�t��b�2�A&@���?�^y-B�������J�KQ���n��ZK5�WfG�2�����C�Q�K�1�bK�|U�<J]�#��x�$~i�U���{1�;�.��xR���LJE�-����g����M��r�U�*�Xfr�pQ�2qΓ�jG���m�UȢ����B�ؔ�uݍ�!5V2�C	�͒7�x��믭�����0�ᙲJ&����C'9`AX%!?ɜ�W_�T`�Hw�������W_��qJxW�j����v��/}���<�dU%��%S����?�#�����_����WVV�`}�<
%S������j��X��իW���������>p��c��֤�Y�#�R;��P�hv���/�/}A9�6X��v����Xz���ik��i��/�_T�sq���f4߿
���������
W�]*ڮ�*�@°��h�W�j��Z�7�(rie��w?ƪ���w�R	�B�Ub��Ri�rt�oЏ�-Sd%S�F�!�3q0����z�gK�jc:D��7L��[�y�C�n��K�Q	�(��Ȉ+]�:��"^�4j�{�  �5�#����K�.a3�����*��p��P���F[�"�gaY��S<Y&MFǚ�cFv��5<���R�����T�53x���0L]/��2����{�n�˪j	���n����=aҗS���9<�_�p�����~��&��^���+!9��\�������U��2��q����َ�|�f����Ͳ0�JiFS_4ݬ������f65-PIt|qKq:q!�ܱ�,%x��l�1B�>~���3�Fu%X��u9 &�QW��n[k��zo���5q�G��p$#{��MX�!�O+�/�8s'���H�up4_O?U����^y�gՆ�*�N�
=���^�6Mψ�Թ����P_�8�����d憯ƌ	XlАc��雖5�v�J�MwY~�V�t$5|��8A�^��b��N'a��"������~�,�|@�3������(�W��;/S�sQ��@��<b	;	͇�lܬ�Fg�D�(퐡Ns��x�i$�H���o}�!|!N��&�O�5�dc���ņ����n�KM^bj��Sap7�5��`�9~�Ʀ��M�t�.��b24����8?�e�O��,�����$�Y�����}*!9li�Im䚻�W�Y˔�\y�!�]�Yh�5�'A �0��Y$�sa�l�a[#u>�7�!�9��n������N�98���9���s��IH����/��9F�V��d,���`�:L\z�!'��Xnz�)sD
p��Jv�R�X#>��k��?'�zq6�h��]ϟc���9S�I|�=�����W�288���O����LG���!�Ar�[�i"�wx���xJ�6�2�p�y�$s�u��Mc'Կ�%�n�Y���/e�{p4���Qz���	�#!'!�Q��(�I/Y��A�.d��VГVf����Å�i�^��J�F�i�q�	槻b#2Ђ8�$���;l����3��MH�;���Ϝ9�W�W�g�Ѧ��HD_8�1���p=|u��G�#.�������sa��$� TD�%0�a�@��O9�"V�J�� ��^��\H) %��s]hV��ۛ[[��V�`+H��Z���ī�7�ܾ~������O_�$����"�#(i���1~x� >T3Tit$��j�)�a��`�Z�5��׾ƛkxeF,��)��n|���¥�f2S�$}�Cn�Ͷ���+³�� �Nx:7?�)t�!�cmE'v����/��\�x�|E��A(Ϊ��T#�9���O>������h��(��#�6����"v~����.�:�YS6�p}��	u��l��`�$�����5���d�q\hOm
G�N1/�x
R�4�[c�����խr��-����..-^�vf%�g��seʨ,*�<��3x2%�&I�X��g[��9g|E�7�C7+#ˡi��
ZA�&���0P����������/g�]'�>p
�tE�=(����R����j!�.K�s��b��h؊KD�X'n�TD����(h�0� ��1`��Ɛ0�<Q|��B{pۋ�\ �� ��Ō��׷4�t�`@�`>�R����������{��T���x�]�)&4�J��B��(!�pu�ϟſ8Dd='{�;G,E���aX���~,@B�މ�7x����p������Fx�*:-�_q�WB\%`�>d,���m2`�@�\Sc�hޓ�P���*�\�g�Hپ��U�@k!YC���� *~��$�vc�sh�;�c0�sW�?5��ի%)87�oJ8���bb�D������Eo*d�c7�>7'�+6C!7n޾q�N�N�A5[��%�Ȇ㡆��ݻW}.=|�V�4�%�=B�%^���q���
DҪ�R���Ν��Q�D9\V?���yS'S�v4 �֝�LXn����@����3`��Z�����n�j�fy��C~��zǕ�0��.(�A����W ����@3�Ę�eL�M;�|�m�J�����v;�aH���g��)�,q��۪l�u�wO� O9F�sf���aj��'�`�,��l�i�V�``�9��IMA1��'x����0p���Х���ad��?�96<���_��K�:MVϰ��qJl�Q�)�&��|��7��V;��w�D0���m髶��%m���`b�ų�M!�ߟ?���ƣ'���"�ۃrR��K.���.�uXr�=�t0K8,�3�A�`�o߄ �mPm��FjKdH��g��M,�U@V�.�	�Tė{�� Ğ�.�Y-�#��L�ݝ{wa�Z�u"g�oA�d#p�SCn^����jP��{�!r��J�c-I+X�L�~�����.P���Ef���Jj&ڜ�H^H<G�ƍ~�!�Zc�`G	@ogK:k���X	���G�ٴu�mP)�ZM�!A���(�c�@Og+������4����7�x��Xt��Y��=)�$�'���"�0v�z�L�Z,E���\�ufS#Z��]�!�}�*,�37 ��Uӯ�0��ϟ?|��|s���5e����,����?u�^A�ƽRb�D'�J�8����e��F)�*J-�䙭����<z예0�c�͕�&L%�#�/���M�4
�7�*F��o�ն�B��mC�@>=���0�Y��<���h<�z�-*R�Q%��\�KKKO?�'���=i��`]aR5���gc�i�`0k�9&�a�f�s� 7���Rf`�e��)v!����\@��фn��$Q�����������9T��r��g.>S(��G>�����B��o���_<�)^F�ّ/G��_���>U[��.O��b�X���W�TfK���%|����F��;6�͠g��)V�.�U�*\�l��A�nɱ0��!�d���}�$ue�(� ,�2��f)y��s�Z�sT&u�4�A�aE�0f��Pj�)��pM�%�$<x�8ͽ���|���6�������i'�1d�K���Cɞxs-5�9�^1GI=�X�d�(�Ǚ��'o����Ƹ�<�{�&䦄�Է+�'p$pڕK�Z#��y<�h�{�%���Lq@-�{�}M*�Ԑ����OY�G�FZ����ГOׅ>a��L�1N����c�RJ"�'�:���*a������Y�"W�ז�Y��܁����X��N�0�KbD5}f0�S%��N�`I��|�� ٱq�N����Kk?��%��
�̍3|ka�[oxDy�6ȤK`�Ꞁb�c�O�tZ�jx�1�+�k_�җ��Ƶ.@.;s��3����vIVEkU�$�5�F��G]�^G��n/��������Z���k�������U�.��j���-���u]&	�j�I���$�+ȬQo��	5�T�>�X��Skg.��V���_]kJ �V�9{&Mrb~i�u�؁�{`ie��S�x\���O>&6�)�~�[��y��F ��)M�l�
S������O�0�$�Ӓb1l ��m����ո�c�S�wJ%'�<bRT�|�����XX�T��$��V���Յ<�����e����Ɲ�m��h�z=���r���2s�%�!a��� t�P��|������l�<�:��ƋT��>�n,V���^�V�`!0[�vׅ�Y��@�`~�����q�J6q/WV��+�\��x�Հ��Xa�a�h���s��}Ld�jX� ����K4v�c�1s֯�>�S�����k׶Ϟ��W�������Z2 �Qe��h�h4<{����'w�ޓH�0��{�2a�I��i'�jS3�B�)N�t���Cq�RB>%nZ��8c�;�m�nT�6!����/�d�
�Ӏ�DK5ӥ��Ko޸�3&���O�Vg�էv�S�9¨�*VZQJf�����A��i��*�e�1#7/�Y�a'`� �,^��[y%�u��̊c~0�K��V�`C>����w����fL�RW�X�yWS�y��iq	�{��DKF�n��	i'���eقU�?(�2������������!�F(EI�㰟��#6֡�U̵ز��>7-3g����M�/_���a�7u]�T��
�pQ���|��ÿ�C�QЊ�,s����uW���c��磖z�o�|)�$�����wTe����eB�I����й���#
dܟM�����W)�"O��-ۯ%�:;R�U8M�ŅV�]�[���Py������q=v��p�J�*�=Sc��M�����Lѷ�R8�ɏ~���O�7�_�Z���w>5�/��kI{������\})|��.�EpH�dh���ۥ��p*�_Ș5��
���[�p4^��۔�E=��`<8j�ք�x�I��b�ْZZu�\S�e��JpRNN�E�5��Eq��P�D��fSJ3Z݌.qA%�l��gr�Ν�����Ţ_�x6�]�3b����=�y�OH`�n!)�si��WI�j��6�z���[�)<tbD�j@CW\tn�y�[�f�F�/䥃F�E�
1M������(�E�)O���[�X^^�rh�k�K�$	a��HS5���j���V[�Kk�3�[�H�)�����Ro�_���{���3g�
 ��f�:i�8U�`�si�jȮX�X-�bE����/�gϞ�Մ�Cb��Ts���W{�MgZa]vϬ��,9r��\��
^he_�nqBEoKgh��8��[�y�M�5w�'����4:��B.��f��ߞi���H�(�/���y)���/��I�4(Ic�X�i�n����%\@b���mUϟ�"��E��d����}�(H�͒��E�*�ӡ���P����VA�b�3�)S\-�T���8i�˚�;���p�Z	m��ų�0q����ߺuK�h�:C��e�>yz��`�-����^�ق�����j�76677O����.4_O̔VH\L=N��P�-�����j����Mo�WuuW{��!���F3��J�z���?���O7&�2��I�	��Ѿ��˛���ͷַ���Jso��P�y��^�[߂S�j�K PcG
��D_�.]b�vِTt��f�If�nǖC�YE'K�d�X>�HW�#���R�*���-nՅ>8P�{���ω�Vz�����`8?��t[�&�MCV*S�Gxw�a1�o v$���w����^T��S@%Q�H�n&g�_IO�HOt�΅_�^�d=U~PPl:�r]��u��j4�8�h�pZExF}H] |�u�m&�X��&@5p{�09���|{�,e
N8􀜩"�����\�.N�B}����8�f'�������h�?�ǈn�D�T���Y@O�����<�ty6�eBf;�6��!(��$,��ؕߘ�dU��K�R�"�	˨�5��\�K�$]J�n�{m�g8&���EzVhyI9�=մ��dR8�^���+��$�����O�����ԞK���eߧZ�`v+S�����w�(_�3)��=B5餶;����3�)��V׷Wv7.^�D&��#�0^�[�B���`��	�@+�3᷅��N��AH�v܎g��]6.����ȪV�h�f���^�vOE�	�]��,�^̞ҁЪ�G_6pa�jOc���Xs��P[�E7
(�����{U�x9&]u��'��+��
3-�6_���yd����D�DX�Qy^���˾p3�=|ѿ,l�[g�&���䛼^��Ļ0'rpN�D|)������i+���%A���dpb5x��*��`�|f�uI��äX�hP'n������E�\�RC��TZ�}1�m���wx�o��&�e�
�#�WC�NN�S�SE��E������=���� ޥL!�B�;�q�&�\�7�x����_<}��oY?wNpv������{�J����>WIY�RȞC�p�~�$��=ڧz�y����W.���(���b;�U�TxA�?5K���ཊ�4�����;��QM-6�KN�:ҡP��g
��2V�!d��`iڌ����\�,�Ho8_�r!�$@;:#�"�]kJ�$��� d'Nn���_��S�mm��&Q�)�<��6��ཱ�G���������z��b�<f���PȼK41�e��c�B�8�wGg��9{�,6���3=-/�j*�7_�DU���5/R76�+�p�@5�Z5Us�;<;q�m�q0�sfJx%ȣ���;����Ц��05i
,Љ"A�`v���_a�
|`���a���f��ꫯ޸v�:�܈��?�d죏>��o~3��v��z�.��u�b$��R��)��Z��0�F:����w@�Ԓy/L�"�8���"b���4���~��+������Y]]=sn�;�o$��{��>}:�8��N�.:��(ճ�}��\�W��������v�zà�*�E�)�!��·�$�SX���9Ͷ��Xg��l|��L�z�&�،!���O?�����Ar���B�jaw>���X�@l�.o.��u�4O���ҙh�Wda�y�ۚ��+��������F@�C{��湢���_Wr�GM*ᚇ��Х�j��-ɘ��~�����lKbe��_�b*5LA!��_h� \������X2�Zq��>T�S�h4D8����A"������E���[�Ss��E<לjB.���~Q�	���C�(d���I��墰y�D�R���e/�٫�zRg��"
�:�´�ҙ�"JL�B=L���c?~��<���k�b���BkN-��"l��*��n8�N��&)*v 2�r�*�̍O-ƚ��՘����$��d�!�Fh,�M�C\f������/�$cd�r�)�xF|��fF��"�m^�2�+C���$lJ���Y��m�J�������s�Ӂ��{���˔]!"�\��}dS�+����H���(hVTwI�κ?�gJ�XIҘD#.��\֜�9������� p<ubeڥA2,���;݆���,v/��#�v#��,� &4�;�D��S8��(uV�n�ǹ��!�g���(��G�@�9ŊJ��M��I�]N  �͵���0���O�N#�Ù��(Κ'h}<�~ՙ���t���zaP��#;��y���/]9��ٻ�aF��V�N�3�*�2�g�;oߞ�(C�:��yR⤨Z�2�U'�}���X���Vl��d�g����z�"�t��=����v�3��d�,-�(�l.�a_�h����͛��@�?���+�x*��e��+�S��i΄�p˪uY��ۧL��9A�����Ģ��߫��m�ӓ��z�ڮC��Y@ef�f@P�/�?�F{�Y�Fx	��<[}}��F]H6ZMV�Y&����Lg�>'���30Ff� ��Md���A�]��R��Of&a���H(��c��d��)w�[I.B�|���X�b�\�Asq�������:�
��N#n�ɣ-�z������d��nF�h��&��^Qx>X���G��կ��ss}���>O,?�o��.���t}�y�tgC�:��]T�b�ǢB�Q��Ɍ)�\p�S����&1�J��y����,Ӭ�򮚖�T�3R=2�rO���;�I��)�λ,�'�U���*>�>����� N&O=y���(�n>�W��H��7Tbpr�S��G�ҋX�&F�.Rs�'1��Z�(|�Hf��(!��P�=�f�ن?�h>�-���bKj�J!�2�/2T��)�j�4Ϡ�$xi6�b�m�)'U\���3���ӿ���璃�1�)_�!X�������1�[���/M*Ӿѝ�@���xݞ��j�����,5�~KM7��"Ȯ�b�������fR��`b�u�2=_���<g����|������6�<���0v-|�-�L�ZJ@,��|�a��w���
h���#/���UotW76�իq���$s���ͭ�=M�ƑnD�H�{������I��eqq�B������0(�?����D�W󞧴�K���,^�9O�:��<��Nw~qie:K�5ۭ����h�%���ut{d\"��w��H�g��t\��	e���_n ��L!�E\11���92��:�h�L�)BX8	��C��2`��>)�@#��g����t.������.�S�,�O���/U���Ÿv�ttRe��/�����x��Ҕ6�+݅3K�\��;ɝU������-,���ÂёR�#��L�	rr���d���vC��.�/Ԫ���$倲�'C��"I�R�$`��t��?�뵆j�D35jY��{��n�Ȅ���!�dnqN�k:����\��+�j������w�J���:(M��g3;Z��|�MRH���bJ�,*�V�&���l�e&�9�YLd&�eFR�iv�.I�>n@p[�����q#���gOb�$����P��q`� yt��y�$`Ox�h�i/a\�)�x��[�q�M�.�����l	+CY%��"�m�ҹ璹�DL��|!t�C�M��Ğ��Ί�D��`��R�!���+��xtP�<*��6�Dj�y!@���z��F� ڠ���D\w����y�sD�2��oܺ���o���y�HK��u�!|Rh}��ǣ1�X,�c��������7�XX�����, ��Ś��V.//"z���qpG�IH'���gj�#;ߜg�DS�`�&�tV̄�����o�y��%��t���&�|8zp��㇛��Ic���2,����B�cK6G�!�9�[����FKY�yP��`��0a�Y�c�qe��m����2e�Ѹ�,HD�΃����6������d�g��&��/Ũi�W(јd�F"ur��n��rD:�*8e�K%����Fѓ����r�5L=Q�O��~3,�P�cC}I&������2��sM'��Ǉ!������D}��gW���-N�8ʢ'c�������f�c�<Bc]�*�QX�T(�g��?���ݻ'�J�H8Ծ��;��2�[�inq����' ��h���6c�9�bU}���ϲ�>��w�鋩�1;�D�	N`�ˀ��w��)�x�l�{���&�>��%��N0(��n��M���\+�9�U�J,Ƃ}Ѕ5��Q6ju7�B򘕚�O��Vt�$��Jc&�8¦�5����#H�N���Y�6���@3ƳO?�#�W����ޠ�h��8A6S#_�����qص��L}�_���Zd$Krb�d��*�ӑ�Jh��\��
,>'Ix�D�� ӫ"u2CK4A��/4Ӕ�LaO3��UPc�T-N�ɋ�ԝ��`�V�C�{���qG�Ҩ�@��P��$�l�t@g��e3@v��'K]��]����g�p��$�͚nb�ju�\����&��Q$��H�̛w~��L��#
�r�#8�
DN1�	�Vh�'=�1O�J&�C��������Ep-��X�},^�.���;x���lnn!���b�;��<����~ef�-D2�8Ѯɘ�#�G?H���mo>|�� �_����!��I�x�r%�jMɷ�Y9#���#|��j��veae��h7�jM2,?����pl�(���ɥ]._�L�d���W�Oɴe��?ޑAN�Jv��o_������s���ƤǭT���@G�Ac�g��D�%�Kc��축��[->�[��mNhe�j5�a�/]���_��-�2H�3e�|7�M*+���t�LGS�Ń��Pz�ҏ�b�Zi.|q��Q0���i˂��S%���<�	�5_�P�l�����O0"a�l�C~٨P�
��6j*8����0���7o4ug�q�dtx�#V���s���K�n\�x�i#�������Vp�Ҥ�����-;�I���b����*^b�4A���C�b��K+7��P*i����^.�d �i̯U�y��G��h=>R63q�b~ʌ<��|����T��f薄����cNe��n%�:�����B��^���Օ���/��z���ʲԹ����*�u�,�x�fI�or(X�p'��Z��heq�¹�çۻ�Ƞ�+��xJH�=[.�?����
RX���]�D��{��N���ݹ6�;\�Tz�܎O|a6kL��9�IG=
���Qŗ�Xq�oX&߲���H/�y:�6�����Qx|pt�ν��N*���ng~�I#��:�c���_���"���n��7���2�B��W�|d���l����gG��V'��	�E���ܵ_W����v��K���2�� 󵦲��!]�����B����/d{�I3�6>���P�{>h_�0,�1<MҼ�~.�s������%4��L���7 �'��fi�K�P"B��FUU��i;�x*H�~�Z�k�����L�3��}���2Aţ�e�J�L�L��F�����Y�P�Os>c9OH�4�+�B��/.�Np}�t̐K���ǹ���-�"O7oބ+̰���K2�R�p���g�߷�;��"_�(_�+�e�^����󇠄yJ��l���,��w��R^��������4̾}���v������8�J��M�o/A����!�x\�&���rŏd�� ��E��%�����(,ܗ�@��H��/���v�������FvLoC�}� "�)q���<NZ���U�r�2�ԙ�qZ	a�&�i~ۧz�ī���:5�YW�M�n�:7�Ѩ�/#Z�0ڎ�.�Zĥ��y�eUW�Rض�-��NY��a=������ ��n���%�.�D�F&{���N����K�N�������Ѱ�@��٘��)(�8yg��>�>�W�c�H�b��3U�N�>n��Ht�!�|v�ff=K�BAz���o~�?~�	|�[o���+�H�X�:�������ӟ������ك|���7�x��T5FBŚ<1ˑ��h�#�u�����k�L���2���u���+qM��95��^�9b��y��u.>���-���	7"�R)2\*9�<���VO�Bpx|�եU\d{[&xNF�w�"Ɛ�n���k����WVV8�oN��v����H�*IdX$������Rs�������۷o"B@��yҙJ�$�̠R�T�p�?��?��f��Q�h�B��ᆏ�h��N*�GSA���d<�0c������u���1�:B�|��'8��m��N��b���d�6�Q��C�W4h ĺ������yib��C�@���~I�f*�&k�qȴ�̓�U��\wQ����M9�S&a��$�A�B�'~���^GySw�FS�����XĘH��Ү���0����|[��b�"#�x��@�󳩜�3s=���Eڰc��|�m�\x3'��K+1<��VK�u��>�����W��k�wN���B��s]M�̜�������?W�_q)0��8��1Gd4/lu��,�o������.L9U�ӂ 㼌���YUn|Z��ϝK�vW���m�xL�2gJC� � V���I�̌8č�.uR	�<�Xŝ�%���n#�
d^�b���z�2+vD #��i�8�yjFY���NP�}E@,Ð�Z5��)�K$�� �ۭ��w���7�{W��t��U� 7	�U�չ;� �Av��0~��yҡ�ln�������]�&�5�	��z�D)	�z㙎��@�J� Z\g�.'z�:��,���$������� 8.]K�Ó�]���e�>Čajɂ�g�\*%�u�hv#��@�'�*22c�$H�D�Њ$u�l�F!��V3�ۛ��$Q�1���w(� <�<�$�����2œ�&ᢕ3#��44�~��x͌xGJ�jS&D�:88����ݻ�\�|����0(ϒhs����:�L�����A���A�<�b��3qWjrpBms'��·<�z����p��"u�Li�kҕE.f}4�v{-�(#^���n�d���r�����3;|ɳib/<���Y&�}��aŎ��iq"�h�:a���P�zHb������K���.�Ͷ���98�aK��l
~;��d���-#�եf��W����/V��8d�J�a*]�"dϨ5g[h���t�����2�jYs܃�"'b�<Q�l`\1\�TA⃩Y,��:i�sy@�y��~�N����D�Qy������~�+��Uz�+wJʏ���:���ƞM׊���L��$K�#�V�}v��2��<;E!��n3��x$���N_���� 5�R֝)�1�rr��ɪ7�1��:ˊi�9��mWwA+g���D��p��c�F�J �/�}E���f��c�o��܄�bT������d�'�=H�	, !�\U�L�z
�F�*I�΁)�85���ոV�jM_p�>��ZU ƖO��IvG&�$3�#:���.�N5WEa#��
���w<Ypk9h�IX�c�>��S|���oͷ���6P�~�0�a����Q�84�s�(!��dE�KC��qw�*���Т9�xv�+���f��4��4�hS��x��呹"�y/�V��yc�X{���R%�܎g_�l���0�M	X<��R�,�_�Bf�Ͼ�n�[���r�EQt��j(�E�QB�~O��F�΀+�4;�$�;8<2i:i�Rp�ENgLK��m�/�|y?E�K�NU�S��t�4�n���u�0�	넌§U�� �*r���Y���ia�)�n�������ɒ���t�JMY��A�+"Ϗ�sg)��ɹ��WV
[�N�,�LOk^j�-J�9J�g�w��ʹѷ�I�	�`���z���f�)m�s���v�O�9u�OJ�W!�yaq�qT%����T�8q������<��S(���¶ ;-C��ȕk����rn�_�HYk_��p&�s��J*��e�GQ\��#;w\i ���R��:eiQ�Jne:㗵���V�������%>�L���{����g�Z���<.�.�/�=�����}��b�k�\"s�NR�a�<k��'f�0"c˦ҥ%�Ye�`������uC�r��7A����8O��UK����q���d0N�~����Җ�s�B��w��M��3��S�2>d�i8�Ӌؐ{*�)U�4/	�T!)�N�M�&yg:JX:��eb�kM߲\�ʃ��ާo���?��
�bO�x3���ǿ���?�#�;��W���u��-qj}��k6j�������~0�3wFT������T~�eA���k��v�Rv��Bk� /lӓ�Ϲȉ0dAK���p��*�4�<��3!��Oc����VK2z����\U��_T�
����ZЀ�Oz�4���	Ɍ<�2��[Z��V�Q��,������-�p�TqX��2������t&AN��Ϟ<�|����0��N��ҍk����~�]IT�;Lk
v32�8�t��KG�W4Z͸V�4�ƣ����_�[�����_��כMa��h�x82��#�vA�f���ױk��'p��ޭV�5,h:TM�ZXVc<��(��nܸqI	�(0Y!����#C��"Ђؐ�jp��L��ŵ�Q�O�i�a�K��ol�?�@�c�gӨ7k���t��91�aq[D��=x�`{o7-�ŵ���Ͷ���,��I��,|.�d����Ν;�ꫯ���?�`-RcIR<���|d�e��B��gYS�!��E�D!4�,K�ų"LǓT�ɤ�jI��S���	�&#��������;�Ā��-r��-��(Ƅ�f���kr�&fٱ�8�Pbss����/��r4�t�H-�Y� i�Y`w��QS���6�4�Xi�/�2�,�
�1&֨'�D�ՊH��OZ+j��Br	�����2}b\�����Y׳�,������o�����U�����.`v��F�;�SMz��C|���
Ʒ�u�YC�i/pn���*?1�:� �g:bD�d^����b�Ƀ`�����~���!�������lpB�V�=��OFS����,WV�8�´H�x��sg�ml��{|x�������Ϋ���Y�#]���
U|vC"�F%���G��CxtC��V�i̮^�
�ׁ�d��$&"��:�zU��I6��;�校�l�̉b&H���nj�3�P��)��浣��'2IY�I�UnV�s+��2�k.��Q: L&*9`�[�4wq <W��Z[�i	�� &�
m���P>���/���눪���D~R��|m~^���i�K���������S3�lF�H����&S�af� &i� ���s(6k<�~�38��5�J]��F�nR�!9��W�+�+�O����>|�q�T3��r��Y��z�N�
�F��'���z69����;�|2�KT���A�/<'��6�paqneu�`wqa�#C7���>"Ùff�d9�%ٱ����x��Y9�K�f�ş�%K�d<�`z��pWkgV���;��49U¹����\���#�,A�%K�0��)<\��������l2��۩7[{{{,�A~`wܿ?2��"L2N�[����^^	X)��$�U�LRfa<<�t����"_u#�����J�я~�ӟ�����Q�,¡��9C%��@���w����doo���C���m��3�AyI'r����V[z�
?K��i
�[A�$Q1զ������y,/~���U7�r��E.E޶I"jb�O�v�
�U4I͜%���(��٘ �W�:\S\8-*9ĘiM����_��W.\x饗�ϜYX^����k?���F�S��q�Zl��ilc��i\�A"�μ�g�b�gS�k,#���c�+�̌�f&E�VS�� �F ���2a7����S߸F�_a^�|A��,{w�������Y�L�3)�_-�@R�G�Y!��!�,�jpꕵ3gƓɥK䆫��R�"8aC�*�Y��,�r�nO�{&����/���R�7�+:4C�}3n(��RWOѥ0C�5&����/���bVp|����K�W�e�GO|�HM�t:�
�w�(P$#V��i3��g+5�<�q�&ܯГ�5��v��I����PF2��3Y��v��zS�n�����p�!����z]j���0Q��`[��{��P;��q)�TG���kb������³�~[」��س�#���SD�)�KbK��p��N����'!�\�ڍ�Օ@C!��B�ʩ��(,5�K؝�s����\j慬�o?Iğ ��&3��>7#�۩�r8~	vV�%�C�y�[�����Jr�|���������=����c}Ҙ��p��7�A�Ξ=+��#)�[���M��h�H@ ����r����pdq�����-*LD�9��N�P��8H�i�\�p��2���%�v�'�8ab�̋��n3�O�D	_S��c��C����t�"I�`�����l)\YZ�|�2��S��>�|�v��=bA	 Z�ϳɾ�4	�EA�4�쩇����2�碔�v�P���t�ἄ(��������BJ�cȕ�X�ue�?e^p�������<DA	���o�3���7�2��\�103�/�8P�p�&d����sK�Ge�ޔ�G�z��N���
��,���t��B���Ԫ��Y�Uͳ�|(>�$�I�ڌ,���&����
��S,�)�Sm��Xqn�b	^0pe�&N!�)�}���ڏ�c��Xa�y���?����������K3v7ʠ����]8�(��7�_�ڬP���;-o�d}���,i�w��hP���P(_�� ;B�3�PS>�qaa�A��O�X���AT$�FĘ) �/��g��GN�b���v�aJ@|r������7��������7o�e��NSS�������!6_~��ph��#�����D���[oBK P�,�x���;ep 7g��IC��ժ��fɣ8P�̈́�C�n���T�m:ŗ�fRm����������p������89a�+Q��R\o��Xc�B���M&�x�L�s-�j60���ɗ��!�¥�z2�󊾠fm���_ց���vڔ��`�A�\��ꫯ�����_��2CH����
�ڜ�`�J\��������Ç��F�\���R�j6P�a���/C�Cw�]US��gϞ=~��"����������e�2`
_l�����2��M2\:�B^����k�W��J��+�~��J
.ɋ3kc��d:bīa^�Y�F>O+���_�g?�9.G�"�\��}���F���KZ_;��\�Af3��k���bbE�F��q��%p(��;�l�k%������˽���S�f�j��!�'7j��te v!46��@�����������ͽ�:fa���i�R����k%#���r��?p�#�<]�w͂D�q�)#:62�fłGB:9,rg:+�)q9���p�č6Yl��q,4�'��Ipw"	�>*���V����t��O�+xA:3n�q]}��f�i�r��M&�������O>E�G��kWq� ��w�+Z�h`;!h7���.]z����Tg���~�z������
���yA%��|6�q�����g�}F^�^�$��#�j��e�թeu�$�����4���|���kX'�����ʧ�'�Y�F��W�S��v*�J,�3QbD>h91��~P���5f2��%�\�v0�/�D$�������%�`�u���Q�^�S;�+�N��eJ����4Ճ�d�� ❋��Fnb�
��b6p��S�Yӡ�~\�<}�Ԛ&�92;��ŜX��vJІs+�(.՜�X�U��x�!��L�-�]�j����W_}E��v�q����R�Uh���������.�<��ʜ������*�]YZ�?y��޽{��#��!�����P��uA�hF��wޤLJ�V�qƒO%�~��I���G��!��F�#�v�$���Ё��!!�˔�V�������_ܹs�G�7[���B]�����2�Ml�ZZΔ"�n�s�)9Y�)�i��2����b��@g����_�z���Kt���ِJD��$�B�jLe�&�ڦ���W��h:>s��4Oq�Ϭ������y�CG�7"7����M����_�x;HPVc�/����4:υ����U�r���|ۧ�Z6᱾xv�S���I_�Iȕ�C��x�΍ϫ��;$ã�G;ı?�x|��ef�G��|p�c�W�W`ͽP���+�{v&'�$~�s��BD�h�M��S�c��W���ľ����Ze��b�	��,���.]8�)Q`�X�|�N&ɗ�n��j����n:N�"UC]j�aV"�h;;�j�:<\�,�i@\q����������!��<�0���63Q��m�T���eWWV����]Q�Q���+?)���İ�����3��R�/���چ۔<-8���?$���g��Σlk	��rEO�<�e3�Df>*�� ����ޮH������ffB��VCHN�u�LW����V�Ԏ���"˸"tF6��L%ahč6k���-O)CrNq-S.\��~����O�[�p�I����/��7����=�?�r~������<����e��H�<l1ހ��ΆUo$����w�Y��5�rc=E |�N���to �EA�w�r��;Ӈ�t���oU�P*�Zۇ�ýj���h~b�*
[��H��f��+_[ZZD�]:;@��f�;��bh��-2�(l��d&δ �̚�m��B�7�����y�40�}�l�W5�w9����:��ʨ��Z�������={F(�m�2GZ�!�nk<fyҝk'�)����K5f��!��p.�g�5��i�U#�"��tl�o��}��0��� ��{�q��p�P&\��*B�������VOY0�U�7���CΔ�(bf�H���((�j�,�.��M�퍹1>2��֞�@j#Iqr,MͦNu_,7'���^e�7�dU�J��t2����\<�ʢ�ӗU�`m~aI��V9�����_XT��xp����>s�ڵ�*;hٵ5X�C�}�ſ�˿d��׃ޗv	O	��ġw���[o��q��E��gr���͙Ӑ��e#��x$�L�!�S����Mu$I�) ''}Wٓ� ���l�k���@��#�H_�+���f	����<�Z��#����]x���w�}G���EK�%��*���^zI�ϗ����˽��[jn+X���뿆M�z��L7}LEzF�$�H�%�l? �q�/���PO���N��AJ�/����]��۷oCf�y.Oi���J�U����B�\f�C�;�n�p�d��3�Ҧ���s՘$h��J�=M��Gi�N��Jߢ��ÊVbq>*a��� ���זWΟ�87�U+�f:Ӳ�g!�����T�걑�V��0&l����ª..._��|z�
aP�L����Q���sLC*�Q���)ĵ�$����)*"/|f��|aAӱ��kkB�!���H
l���!ȧ�~* �c�����Wu���bY$T�U�/����,�y�a��><>���A���JMࢰ2
��6X>� �g�e n?�Lq%Ӵ���)�f�	���
 �֭��M.,,J�^�a�����}�	}���4��SF|j(�L2��{�!�9ϦI A�ý��v���&����ʌ�����a�d4��5Ce�ٙ9
���T�<�ͦ�!�Y=QD)���q����f���X�o��Ӫ��(�`&=:����������w�}D����s4�<���4�*�-�OgR�'S���]NӤ=�ŗv�_>|8��N���q�	>��Z\|�>�]r͂��;6�X]��ݯ���Z,);E���{��̵�Uv�����	K�G�L)�"X�ahX��j4!�fg�F-�5b,���	J���b�h�������*T"�{��O>ŁBp��iu��F��rAN���'2���@����+W��������+�y�����E&m�z����ܙ��S�Q�׭��!{�G}���K�7�hc�<lMl�N1o"�;�5[u�n޼�d:���zM�Z����NJ�4��T�A^�ڊy�&�`��#F"�w� � ��K�L�p<�ײ�x��˞h�w{�;��6ң���NG��㑑0�W@��
�xô�lf�<��bH�V��U��J�Dѱ��3����J��x�^�&�`���0S��%�e�O{a;Z�6�N,�`�M?W��7hwp�0�%�E�+�&CӬ`3�
�åKW �:5R���|�����ꫯ���6H�LI'ާ��я�@p�Y�a\�lP��*t$b�8�H�H{o�� ����h��h��m�ol��mVj��U����>�7����\�.K�dp�{�����[`msl|o0�;8�����ݯ�IM�+��CQ�5�WW�_�>���X���b'��Of���������Xݕ��[�7�R ;�f��<�Ty�/՗Z�L��³��ߒ'���T/E흠�R�k'vЁ�Z4�1��׮]���/\��EF�4r?�>:��������g;�m@,wwwe����LD�fVkMA��Q�S�����7�ma�Dq@�)�)Ow�=��ۆ���"���PV;<'�#�&�D�
%2I�ϧ^��ٶ�wr���ʊ-�ߡ)1ʺ�^��������>�*���^[^��-�3�-��d
�'5s`!&r�+1� \N�io� ��f٠7�DU�q�L��^�D�ŞM�_x��N"��������1�
�~���{��#�Z�q��a�:���!J���J+>�;}�_�Ln%�_Z���(�+UG2���0`	�m�GEg����恂�p�9��i2Sw���73��*$� � 4���O�j-�uԸ��%�l�0}ᨮ��r\��Y[����㡖�g<Ɲ����)�7Uq�����G�d	�p��p��'��5�Zq��d�p�o�����ҝ���F|����#�ƨ�26��l(�L�5l��=�o0Ś�lޓ�MA"Ԁ�Mt�ca��B;�;*Q���8�����J8d�3��M�������[�k�)%�'s�%B*4���:��t���<M�Z]b(�22�xa�S���y!����OD޷ ����!���8ܼ��ן���T�{O�kR�t�E`�r�#&�Z���Ƴ�]�ŊX��?J�>cIɜ��P}�E���˄���\�@{�
m�Y��DƲ��X�4�U��;���T(껏I�*	D��7�<Ta�r<;�J}�����rl9�t�8sD��T�^��ϳ�%rs9����m/pnq�^	��o���9)]����~�-Q�l�|2+�������=&کd�����4�-~����cC�Z5:��{}˖�,��%�m�v6޳#V�p�E�!�E��6��=��n��Sb:�)�� ��=}���_܀��I�>�z'�3���HF�A�����UE���.�b�cݓ��/��Y�قs�tԬ��#P�����(f["8�����ƽ�;B�5����R��g	-=�K�L�:^_�aCPa�$��)x0�<�./�x��hO97�PtzE�HX�Q�"?���h�'��ɑ�=9`g�_�/���'��-��r���=�P`�^+e�jyF3  ��IDAT�`)�^�?*�n�S#l�� ��T�����5�dB>�W_}9��=jg����?��Ke���Ś-��k:g��<m�c�N7�p�xg��Oϟ?�7�77n\×���L�4T[ζ_α����-=?��}�פ����S)+�4e���Sp,����B|���[fz���8y?DA�Ks9D���]�b�2ń�c=������$��YC�w5�X\��U<�	��Z���R���X~?�_�Iru�s����^x.�ϗ.]b�{
P;XzPR��Y�q��7Xv< {.�g�9�������G�=בY��:=`��@�V}���X�S��?���i,��ɚ��\X"p���1�{��O��<�w�"@aܼy�62�v���w�L��Koi�c�I�����X�������	m�֞�ۍ7Μ;+��t�V;h��>���ݻ�k��Z�����J�3)#�Rq��>��P$�M�e�q���0vA3���G�TE����1��h
r!����V[���-�3�ϥz1T;����T���2Pnv�� ���8t�3�9���+,�ٟ�o!��$��)/^���ٳ[�naw8�#P|�o�G�5�9ֆR�P��.Q6����c��}�]A��E�V�5N����Uo^��1�<²#�J)��_"ע��2P�JM -��PMf=���ˍ��_�����	TV�?��K/���)M	>*��M�L��y�" Qc���L^�6��������N8������w��6~��DÂ*e>˷��"&vEfu.,w��FUy:��z�2n?�J	"۪�).)�16���w���/�&�6�/�<�"�S�E����R;x�
�-K�@l�MAjx�|M�F?���|�9I�|X�)��P�= ��xm�+%;cn�Dz�}cXERsd�3=r@y��e��|���!1���Z��������c�ON��%I�Q�!0�V}�]U�N�8��S��i�/֩�i��N�s6yʄ�S�ׄ�}��9��S����դ��������&*ӈI�2̈1�F2+�op"����*��b#��x�x�+�˗q�?���o��&�S�_~�e�Vg~�PR*�'g^Q1�dEֺ��f��R U�B{��U��y?|:�%�6���-�\��s�]$��mq@{Ǐ=z�t�E��N�s.^�mS��L��X6�܎=�L�c����X�5��0�ඥ��ը^;$l�sl8��+�\�p���p\��W��0+䕀]ljƟpơC�x��3�e����)���L�&>vz\�� &M�����e�����Y���j�ǷL��2�F�
�c`ɩy^��Y'F����f<��N�&��?�\
{#���uǚ�W� �>(��o�N�
z���&��1����	�CasU�݌r�7�ZH�����c2���΅�u`s,�KJ��!� "
i�rM�q~(�ȶ|vf(��h>���'L_�/�t�G�A��'�ڿ@�z���c�2JU@�B��!f���Xl�X�dѪ5�e�*����b�и��uԷ�_a$Q��G�W�� ��|~�����AB�j�5�Υ���w��B!���J��7,��D�q2V�E┆��Δu�Uv��XoܾfhL,�o��	|���DR�㜮��ŮZ6Xҹ�<��������H�I��P9%C���:��Y��&�A�%j���k���-���ES�4�+��fn;�M�:��^���7""P_�aVʍ���j�-'LJ���e�-^Y�_H��ߺhQ��z��\��On�e��R��W<�V���T���'T=��gWV���Ah��=S~�\��d�"�ǗQ�Q�ftH!��q�&�m����l$G���B٩,4FJA��Jˋ�Y͂��V66.�_ŭ�7B1�5ja���c�	�M��Iþ�*� �������:F\C�v���t����F�"Pל���"b
�c|�p�ܒ^ya����^n���+'�[^��yn]
ϙ�0|.�����,���x֏/��O��#���oz)������k��w�U�c���L:�3�P��x w�-/�f�0v�A�~/4�������ũjv�e_�7��A���1�#�;P�{��.]jv7��[�z?���2�h	o����\(��R�I��(n�'�h���Uu"F� �r[�	lZ�V#t��?OF��ݽ�p�a@�������f�	�%�4��v��O�{�W0)�*�t�^>\\%�U�"��-z�x8�?�y�&�R�(�.cR�k��G7���� ��S"�D�?������Ξ;�uS���*w��j�m2s*������F�{j-�p�:���5>�t��W_}���3md;�y�g�?���t$&){m��M���	 60�c�̘��߽�0C2��!.Ѿz��~��W^yee��RM琲l��3�R��j���s�a#� ��p�>��M�Dt�j<���y��\�u	�LƧ�i��tA`g��YSU�23W2��Ɉ��T��t�x���j!os���NO�K;��� ?x���&�����'Ϟ�ɇ��G�=@Ĵ�t`�� �^�<�D=��p ����:GV���\������������f<_����G)��:M�'z|�߹y�lq5��=� ���+q�;Q�gr|(*��><f�W����1�0d�,,���v���]0_z��6˙?b�Gv'�N�J`>|x��]���D��x�����ۿ=sf]\�"�"����~���&b&:��G��$�W.���,ɾ����މ81IV�	�j�ޝ�kuڞ&iđ@��`����7�#4�c�#IMnm>�N�΁߼_W�F�ݕ+WΟ���#eP���a����ɸ���|[�mo�D�ˊ�e�`:��ue���������tZ���\ Ad����������	a<_����V<IQQ�'\�=�V�)��g	�5�����W(��5����x|H5%�'
\rO�9��c��� �0��|���9����X��xе�>��4�k���Xz4y0����/.�Ki��Kl+�����b;nݺ%�5��Cp���y�D�4D8���)�j�]�����Ue\T�t���H 	�p� Ks��5|��w_��2�`�+��ܸ[�]�ҥ� Z,�C�^�j�(|�M��(�t*���s�P��^��#-r:�������U�kl5ª�~�QU�ь��s]Oȝ+��'G=����y����QS�������~�h�̙�.�1�W�i��`�VV�J����Xn
�X8��"�9��Ē�s�Xy"�1>9_Y]ƃ�2NQ�F�K�ߗ*#4�6�8WX*C�/�&�
5
���vW��fZi�C�:�p�W��|��߇U�x�2n����g�o��_�������!}''�����%�.�W�5f|߸��n�l`^�;�O3E�i,�s<�d�w����B��%�i����sq��uIfi��x�}K$i-���QԄf��y��n��������^��u�r��l��54�ˡ��SM�ʒv��^lmmA����>}�;����ƿ���w�m��|W��3]%�U����[��_��?����V��rA��ӳ\��&��ޞ��t���M�"ϓ�,9�� KE TO*�ώ�{����|�u��j�+­�*�XH�K��Q� e�KKG��~efP5�:��B�6���k���c�~�|.��p�g��	�-����D��U��d�R�\�ȓ�,8e2BW|s�9UbE]��s�ν��k�OӪOg��t�f�j�s�`h=�k^\	�<��}|rH�XD�FT��s��W_}��na����Qr�B��-�� �q�I��Uk6�6���VD�%r��̾�o] �ج(4.�[�Up��,'1�%�#��u�K&���'��o@�����Te�)�������8�7UkH�T���
-��u���8��H�;�T������&�~w������~`�)+5����~dSiz:<r����ɛdG[��Jq�L�A����3e�.���� �|�B���\�P�QјE�����`0��� �lS�QI�qi3/��=�z��Aq-ěm�Xy�q�N���c�6-l��D��U9Yu�����B��o���g�W2nRL��-�NEM��Y�&Ҏnn=����;�{��ϬH`�.\��N̐#�dq�G1�!�Ô�2VI�}N����6�#��%�3s4q���v�>��Gap6��R��X�2��mL�-�߷S�ݾS�G3���_�O�Ǣ���I3$��'����D"ꁖ�'1bUd�a�p#���H&�z�����I�\���2N	������L��G���ӳ����-_�/�2�t�0DxU�* tQ�C9���&��.�*M�`k���V�K�ڬ���̗v���~>Φ�����`�U�sl#T��%��qq~�th��(Uw�>�,�5Z&�W��l �  �8?Z��2}�,m�PZ*��OЪ�D����Rka�[�3I�&ޞSZn��N������L�S�eΞ��bG�_��4J����}r<�S�m�r?���ٲ�.o�
�����]��?�<� �u0�����B��u��ꧧ�og���Ņ�Nd��n�U��qW.�%�����,D%���`C�&C�ǡ���}��"T�l��B��/\ؠB'�K���L�N>�;,�k}�i�+.�E��}�{{�j��s�_�ݑĖ'�j5S[��OyO�x�;wr˵I��"�L�L.ꭧBVz!�+��jK�0IGM�8��
�əI�Y��s�p��?y�Kݹs�9v������y�� ���:�0�O�������)&:��e� B��#ۜp���\���|�;�q���k�����-l]���DIjer���,��P��x�[\f�	�t����`�^~���o���K/�gDX�F��&�v��]6/S���׿���=V�)�u��(ꊝ�Hs�)2�]Nʶgkt�1�]���t2�hQ�$�n����UH3��"��+���:��o���+����5۴((z"�t~�����\H�1��<~�T,t,�ju��Z$�L�1]p�5���g�Ra���r���C!�G�J��ŕ�U.��}A��7��H�~x
^�<D�)Ry3.)a�h8vb��S�� 
NU��a����z[p"AM���J���4�6J�"�	j�If�/��/���q����
�A��sMʕ�p U�"��o.u����~��Q�L��5�_*�K��8pJmy��EU�$�d����~��_���*>P�B��	`-��m���ݪ�Z�ް��/��Ҋ>���21y���=�5L�%v���|�D���ۿM�d}}����Zz)_���j/�����m�t֤�i\�xr�o�ƿ�Uf]�sg��a�ن(�vj'nc��*:�JǚO5�ނ4.,�3��{�>��-�v%��Y�D�%��$��3\a62�X]�4Ѩ��m �X
��<�n�R�����H��OGB���qN�4�&�#�7���xd�`�+���G��I�$��}"]�U�����t�O@:� ��#��M������	t:R
9�t��g���:�Ӯ�<q:��g�)P(+F&���>`��_9��:�����3��%�ʹ�v<��_D����f�7K���v�EO�6=��g�6WJ�cg�(M���H��6(�mwtt@;�ɏ�ym2**j�|ZR*訆�|��#��B\��q���<;���S9�٩�
�+��Ym]�:]�_����<�?<y(�W���7����O�ݻW����b��[��^�y��Aa;����t�\�&�M
�ݓ'�.m�i����_��=\�(($�#7l��:Z��5÷�{-m�䀮(SDW�j��+˪����j�:���B�;�<�l4 7Z��_�
z8D�9ŰN<�zd�,u*g6	R�r�/I`�������w�|c w�|��ǅbe�l����8:C�;����a67��;J�3���4�cQ�j~�����؟�Ɇ��H&A��s��r�9Yu��r��h����G��B*ֿ/_��L�����%ã��)�%�3������h���.����\{ݝ��ʷ�]�c�N3�<3Z��^��S}eZ�
����ϯ3O�T���^O�q.����s!.v�R�o�{��[oU���ӝǏ�����p�t�3��k�[8A}����{��5'Q����6[Ͷ �t���u�|ݺuK�f�����ч��X{��)+�K��t;�DK���2	�bZ�s��U:iq�����l�>V�1��;4��u0OW�U�E���Qoy��l,4�Mo��[�m�ݒyOgr�|^�הj#TBpx"�Hi���E��ٙ���H@\a
�Є�����+=|>�҈�đ���I����&���f�T/bvg�^?�l�ݲt�%="���4��G�n
�k�nv�c*Ƒ��e�.��d-2�~`�|��E��Xeq��\~����W��9m��Y�Ҡμ�s�ZfO�������ʍ��b��D��c�b�3�5o�ׁ�+:9��i2�:����.qYN���4�_Bt9���[��i���.X���_>7���{��D�7S>��:;�+/�B'∹A�k�a<���B�5������X�v�`�������G
�S3w�|��q��B�G�q���ɔ�M�)\�-,E1�~�yw<ŔC{|R�#�����Vc��J\Y]]�ﶋ,��:�� �_��2���2Q�A~b�-�'�ɩ!5���4y�[4�w��������	�¶`���3�nk�s6���T��v,K�����u_T�͹W��/
��A�}r*v?�j�
$ ���CQz����|�ӧ�ڐ��[N��K�o�3�թ�a���tYTfd����*,��Ls�<~�)�_(�)9<گ�1����88܇�mo?B1��\�~��օŹ�啎��%{:1-0\�N ˭7/��=�=�*�[i4F�:.vj��tXxi�%�Ig�)|��1 ��P	>:�s�;׮�}����k0̛����5a�ݷ�9�a�NЁ�Q�HD���$M�����n�=ҧ(ĕ2�XQ�_��_����?����?����o���EIƩ)Jg��ɮ���B�1b���ا�e" Sfb�:���PXD!B�Y�K���g(�װ �Xz��yF�%�Ŏ~IKi*��L���E������5��I�P�����o�� ��U�3��[�a?�N1�Xu_ˌX%��>�zư�	Jq��/5Sx��b׶���_;��!��j��$y���n>��Y__k�ۅ�x���t�\�xe��\0���Cc�ym(���X(��*��D|Ĵ''Gz���X�ܜ��8Ñ7���q�D.��<���|�L��@����-����|��z����d:����ZlI�Y�����pOV,#�
���o	Zmr��J"��@��8�C�auԇ��T�;��}��o�3e�.x���H4��=���ɀXH����Kut��߭�	G�N��F��N�e��yd N:������ׯI_y�*~����ſ�A�7��ڪ�够J��k.u�
GA��t��qODw��
���A�CW&�G�������f�e��+W�fS�¨���8J�vM|�g*]@��{�c�j�0�Y��Բ��F:�cYo����ɻ��I-�r�E��5�Å=�s�K���"ȋjhZ�\1PS�~
��aRj{{˵D�ٳg��}N�t��ŋq'���/p�Y��!�����իW	��mW�o�Qᨴ��\�;G�1���MϬk��b1����X�f��[]\^�(���ڇX�]l��,I7�U��,=RC�)<�l֢Es�?���vԖ1�&RJ��p�v�e�x\��f���i��^��qZ�r1pW3��Z���GG'�?V0���h��`+	�N|5R�*�١��W_	1�/�3��܂.x�o�  �lM�����'�E�PP��&�|��l6V�	>/	"ة�x@2)+]��.֦�eSId+kX�T_ܣ��h*B�$�*g�����L�C���1*�;� [�w 	�S��o`�U�j(�r3��R��t�/!!�@�6�B����<��9�b�[&eF�.d&�/[p��p�O��������U����Å3���.E��B�*U�y��/�����[oq�.+-��za����~�p&��l���;�ġ8�x'�ȣ�^:�)�
|Y�NC
�V������t/�h��LX0�4���KV,�3�4��8��g��?wa��\'�³�K����xM0�]�V�^��X�X���<�BYe�*Qj��F`��6�#�H��DQ���E� ��7k��4�i3Sb�,�/���y�D��aU` �.� {^�*�>*�WS;��Yoy��?>a+�T�'������䊆�
¾��Rza�)t�hez�}��W_�G�]m���M\���RG��ZRߖp(��HX�(�K[�X��a6��'�qςC��
�����}�g�{g��+Ѹ/��7��<̥z#2���
���D&�JT��U%)ݨ(����o�2$����ś)�Q��T��ȱV�	���g��-�|�G��ε�}��ͳg������3XY�e>J;P�N������������?�C���z64��Z7��8��w`1�ȫ��2����F��C���0��	���u�}�޽{���}�]X�˗.1#����#�p1���d6���7�]��S��F�#h�>6������tȞ_��1��u)�i�2TJ���	<���	J��8,y���ȷ��^jZ�� ���$}�Ra�3�n64.k9�s�/�hו�K�z�_$U(?�\�B9C9���Igw�tx��;���G�DIگ6<�?��`�ƪ%��g��)*gidk��6j��:B;���Ij@��J)��=�V7@�CF���;wlm̸:~����l�S�z�����=�tX�<8�/L �cn�oK���lb�TZ�49e<��J	,,:$�s�i��� bw�v��a��_n=����N�UW_W�&�T�hp�B�qXB�����l��Z��	eU	�T����ۯ�,����%������}ؤ�J�A��#��S���'�R抙h$���ԛ-6=`�`Ӌ,U���B�&��ǍF��D��@�l�(1�!���Q�C���1��+LBߌ����:��t�(��̣���ey9�=���=~�#� b�E'D���� ��LX���3g�P�(=Պ�ǣŷ,�H@�S���l����~0&�8�'s�8e�si:
N/��p�.w��uNq�S��z�s�`�ǥ��%j�����<���/J`�0�(˛F�e�K*�Fڙl+��l�c�vˠĴ�O�{q�n�/�8��DKɴ�͂�-�-��j�L��aJ�^���a�U
��K;;;�H�zͺ0.�6�I�*H���a��d�s�s�|��N1&��P/V��Q���M���WWW<��D���v��pI�8�N���f(� k��5db��Z�0Ef���w
eFK�i�v[�e2w	\*�����y%Y]��x�(���%����GՎdI�ҋ�U"�Xy�t�%�$���qM�-��β�H��O���+���B��*�&�
S��
)���WLd���*wdGS���s��%� ��7�,��)T���øB���зR�1�����'?���'����Lp'�����_�mTB��4�������#��٨��֤_��Z�P�X���h6�
���k�h���cDy��(w>���E����ں;����^.)|�ݝC����>|֫/���T��Z��.މ�+�>�%8��P��Ł��&��&�*v�R���[�FR�v���`2�B�U�_��}���I�d|b�ZX��ݻs�o��ښF��4)P�tnW�"a*.��S�[[[B��
����f(
e)�a��|�^��ի�6�౑aaE64�50�Q��:��C�,g�D�)ݕ9|�m�HM"ۖ2@.,���c=!Z�����ч�P�����=x� A`���/�v���<3�4��"_���)c)���i��(��oh��%OByD>�vw�Y�\v�+���~��P��`�5'f�jR[?�F�r���J��ʾ��?��_�;	����8z�<A���F�Ig�*�F�R}�X�8=��LM+������3	�u�t]=_-hGs�Ss<e.���eT;!W�=��'�&u&����t�44D�����#1���j���Nv|9��pM��s�ӓ�LEQ�ő���'��ek며���9S�d�~D�
4�%6�jC++Bx99䨥�X�j,qK䇄��
gy9{��{�/ݢ������7;�w��ۨS�s��گ�	��@��x�~���5f�k�"X���?_Z����P�T��=�lA���7�Q��\q���2�U�̍z��\5�~��4$	�.�2�T���c!�U吜�Q>�ݻw!BW�_w�oj���0Qu�j�y�	j`&%P��43�|Q�(R#$!��~d��i|��&v�-�d�K�.AM���/����"G(�a��A�I�I�hd,���v�z���:�#�FL��aT�tM�5�d졲%��If����M�B��x���_�&.��\ �qGPh����}����e���{p���5�&,����'�qfDʠ�i)���O�ޑ| �}9����~��G�������=reٵ��7lzCϢ�"��T�ӥ��F����w�OA��Z��ڕw��Hf2�����9'�,�~Ox�;+3�ƽ����ko,A�����r� ^p���(H��	����Z�ʗ39�Ԩt+�I�I�Y���2;�s�x�$*�v
	��g�˞�.��i��6�~�vD5ަJ�!�[4�vJ�����Pu�}(-˶o������{��N׋���k�#g�BP|���Eߣ�88N�%�+��������uz]{�b�ئ��Ujw���FZgm�Acr�����L��Ie�]� ט�	4���Ү�C>
nzm1��������:��Ei�MԚ�ѓ��B]O����¼���������� lv���]z��֢�oݺŎo�N1��3�r��8s��J[���<�����a@��O����Ga��(eԥ�10$�7� f��,B3 g� ������8tѩ�(c���_:E���'�X���R<�-(Cۛ��\��Z�$�u�,��&Z�RTS�0��5\�YΆC�՛7oT�W��"�Η������J���2����3%ņ�E֯�)�'�z�KY�b�������y�j%�ސ�ս�a�◙f��1998f�X�bmz%T�ut*��e��DL�P�S�𾽽���zzs3���?iqd<������nSl�'��rR��\�۳�4�G��4�I+e�ց�d��g�K��H��)�$�K��g����d�9I�||�9w���x�BC����m,Q�|��<m�+$��ɟ���'X���8D��w��y�w�c��Sg����y�����f㚹�T"E&��b��j~[hib}ȣ�rkKţr��
e��<�5p��0	"����UP���@��H+U)aq�T>�jFL��&�߼b2 ^�4�
������,��&d����(����&�^ڈ#(>iin����u�e/^n�'�b��凞0�7�d�]�ؔ*:|1����.|��)B�݆ڗڴ2����*��rE�a���5.�1Vuɞh��~�/����6쳲W�E	�"	�LS�R��ŖЃ��]��I��irBS׍�P̼��y��-s�'��f�T��p&�p��[a�[�5�E���oŊ�`LxR\��-�gP,�w`PH�&繬e�q�26���#�$���������=�Q� � ���b�%����K�7��YA�Ӻ�Sլ�۫�P�/\XZY�2
Ӥ�����i�||x"=Y�$/�q��XSߓ/MҶPN�:E՜�=Ofej�uډ�7Bh�Qx:8�;`ݵiw����R}j�+Z���M�f\�9�a߰��ޕ�����=���N��6W������#z���4�py/�
.�v鬬�/��1�a-����Q��(�lA�>�*S)���T*�1F-��8���#�����¥�����P[o����FC�[�� ���½am�80�R,�n2�d��.*q����r�=ַ�h	:@\�Th�e�X
/�	��YV��߸�z�敕ͥV?�+�T�4s����Hܚ�%�	Upzt�_LVՔ�IV�������ꅵ~�����I!Sk9�|LI�_��􋯿 �0���h��I�������<z���C|jmm�����dT�S��JR���*��PI�"�㠣�d��Z��JV#,�u1���� ��2mu��_XZ�K���^W�Af��� �8g�џ\�/�=�[_8Gʝ����[_~�U�H�V����V����G�o���v��������!+Q�LtH�	�&;8�K?~�~	}ĭ�7���������GXn�xa�]����'e]���K����`!K�::Ǯ4�[�gE^���������ӳ������o��H�b��.�5�Vh�b��V/�!��ÁȄz�m�l$8r���`}u�����*�IZ�dBmd�Y6>9;.�\�W����IL+	�(Mq��ڎ���;n���R?L��%�:�~��<?>=w���7�{q��cVז���.u-0ěB�$r�m�~tx��0���u	�֚� K?^,,�+���:t�G �CYs����r�׭'E��U��oGp���k�{:�U�Wڝ|�����{�K۷������ʲM��]�,K�ݼ	-4q�@Lk��O��[�KL"��P02(^^k%�����k�L�
��4荓wiE
z^�Og�T0��xb�k��:�L�ћ�]#$2-Ӌ�X&B�>�Ji��x`�F��p<y����� �U�-����4���t@��YFmV\���A��t{���'ig���4MVC�����f�|�v�D������J��8
����j.�����Q_c���ʕ+�����t�\*GBz?��B{�ǳ���G�?|���P�^O����M�g��8��_/������!8T��T�������]&�!�|��^ǉm�^��q������!��?:8898���y�����^�����uV@�#�xг���  γi��R���e6�����������$}A�@K���������9De65�u��L�jb�)�αϟ?��/�LP�[�k�P �L��'�&lW�&\_߄!X^]��n��&�S���z�utt��>xp�4��� O�k��S��`�3������E�����G)x��BE�:̡R�b&� �A���t4tZ	�$I;U��&����b�V�����'�(R;�1iw�^�u2.�g^o�B�;��[=Aa��V��	�7©�f2��W`�G�?^�.��^��Q�Io� 6�a|vQ�g'�3z�p�88:)�����P�g �,�o���2�����Յ�Q6���Z_Y��V�ZrĸN�8Y�w_�dE~t�����Kad%;��'5�$�r���Ӊ� �g���gϞ?~�/�V�hS�:�4)Ǻ<BbF���H%���_X߈e�J I�@rg������o2��~w��Û"��qֲ��Sｺ��G_6��!�^�a���@��u)�@T%�tV(o��!n��޹y���+Z�k*��~��YB���ʡ �YZ)m�j_7N�gEm2�F����G�A7E��$�����o��u֕s�NS���mAR;r�;=Q����Ŭ8>8�� �%�R�(|r�V���Oxߊ���p�Ə=�J�tƹ���5�	��1��� �O	�XY�He�o��Z���իæ
����T��\�V��I�p)v�X�*�Վˬ@����eN�Ir<��i���]���|�ʅ(�ۭdcc]�vϘ�H��p+����F�H��������ͅ��_��@/}���0�p9�-��	*NKw��%�l�"BP[Y#M��Q�l��3���ݣ8j�ְ�Q*NK�M���6!*��--I�7���&�BGN�h�^��Y�q���؉R�qX�18X�X���o�q�a�bd�<��n�έ�[�_ⰜMNk28ΆL��:1�
q���ry8�0ѡx�u��-��j�lgg��&�A�i1�⮐�H+c��b����bZ�IG��777/+���Ϗ>d������fI-��óA6��s���Z�/�a@��dz�cyٲ������tm9��8��p��|���ѡ��~�����=M<����,X��Ǔl)s��r��y������{Y��V������N����������m�����2�t�-��	�\Ԝ;�l�_�̎�}���<���ns�x��@g���p��H�pq���[�	�;
1Ӂ�G��侟�Cb
*B�����0�(�,�2��2�#>Ϊ Q�;�צ}���Z7M�(�f�2E5W/ˌ���ux�����Bc���ݕ���ĳ��@�*��]C��̞&����=�E�i��h��j�E�D�#
C���T֮�;�8=������1;�1�)�03���R��й���c2�����	Q,aC�$���AI��MɗhC��4�&L��ۆ8Þ_�M"�{5��"ޒl�8��AO� B�M�q�Y.� 		Ld2e�MA#�mi�eaE&Y�mi�	3��JyM'��ca���f��B�yO��f�_� pF [>�<�l@�u.i#���b���΋�UP�!*�dii��1?���5����py�
Q3�ث{v��u�1ϳ<U�7_��m��Wi<�]ai�]�ͅt��=T�N�R��}�O�/�$ΰS���K�j�v�(Td�ol����Ĳ�zs]ϾV�ʠ���D��G�(��L�����FdX��C[I@X��q�PY�FJa��a#��3-iG�Z��;[;���4�8z�Vu��UYY[f]�	o�bZ�#3��_�uj�^��m��
�V~@���-�?w�VΫ��tR�&���͌d$;�UJ��;w~�ܺu�[����� Z�JF���X�����v��B&�MX��x�N��2�;�;�8��t�a��83r���-pm;���^�~�p����X�C�޽��L���x@���E֒�N�,��^����W��d8e���2qFb�K�w�l��=�K#�iZ!�t���B��X�"k�!�e���'_+*�m��y^w�h�,in��;��T������'O�P�����/b���A�@Ѡ:Ι8hWdS�a෌xq�`��9�,�$E³{v�1������{ v8������_��_u�������;{}�������SA��!��+a��,�xc1(�����у�3!3����{�)?Y�Ճ$v��mn���zX"�/�S��3��#8s\���S%C,^�|)��ȕ*}��e���T�^��$����>=[m�oOc�-������q�Q�/{u�@�O�6�� 4%o�o�ƍ�[ <��t�q�<�ҥKX$�@Rß��hO������)G+|�3���e0�Imy��9�;I��γ6+XU'Q���_Մ�3w��x�(<��o���}�6�'��|�Վ�B�H��3)n�X{ ���F�� �	�SA��I|6�t�8("$U56���
��\�ʘj�f��7���U�q��n�3��c���5^��̀�����"?[�)':7� ����3�eǩ�|}����?�E666�zd�B�pW��9��GX��z�܎��t��F��p��	a�>�����%��(�Tu)=WW�����HO�N�_~y���	�'�v:͈a�ޜFd���V _���\b�_J���`&z~�F;|��ousCz8�-�<ޙ�B��肘_�"�JCm�:9�j�n�}��?�#.����nrFS����o��Q+����4t$ �N*p!WXj�#�J�k���M�#�h�T�J5�.�($�yw*�@T�N2�H�w�̇�,*�l�q*ǟ�?��Ǎ-���0/�xz\����#Rڋg��+E�wv�pøy�Y��`������C�<C�aZN�bT�@F�>,�����后����L���.����0,�K���|�Ԅ�H����eP� ��9�K�F� ��,�{?��6v�s�!fL
6�tי*���ցm�"�Ր-h�95�@��?"!#1�L��f�ٶ�l�nI�7<��6-,�:W@b	i��ŊXFQQ�����v�<��V����ۀF?�~`�I�L!���� Ne�8::��y�\�B��4�*�?�N�����L����3�i|�Aԟ�e��-�6E�)[��F�ϰ_��oI�R���y4��O�Id���]3f��`���Z����˗/���KJ��g&�I�X�����y;(wZ��L�#�2z�v���Ƃ��n5?��f�ź6���)'rp>?!���d�����w�`��ݻ'Ai�E�(�fCR������ʻ����	���͛���O��E��-)�L�#�d��fW�,�ө�9���Xw���L��y���61_��o�n�����˿,�����o&a�����k�u�"*�J)t�턀�jS36�b�$�O� �ϋ!i�<]>|����eGG>��EX4]���x���7���)�v�~�<	`?(����O �W�m�+4�øC�xH��s���-��}����bs!�p[6�5T>
����##'e��_`t���_�~�i�iMܤ�Ϧ�N_E^0@ �B`���&�m�͓����^[��N	$:ߙg�����l�Y��@5y�����8�+��'.��C!$$�#X�G\X	e���>&f�A��0qy�p�_<���@}j>~,�T�MEY��`���t�vډ���n��4z�㴌����kk~����r�[��d�Eݝ2��Zy�k�#�n�It�D��9p�2����j��6di-�l`�R���^�f�T�:�Q�'n�'�HO�낺(�òp����l�>f�vdT�F�S*Uiƿ��2�O����������Tf�$���wt<�y#}0�+ټ��tɦznx��nLpc��Zg����4CːZ�9��.�F��02����LZS��b���m�:g�t�b>��D���(I����3�STM�Dl�_ZZ����A2��-~
��5;�}���e�莱󃙐u>�5x�[XB\�� '�i�����a\ϝ�K�YsG-�(�8�(B5��i`z�N�ƕV�<z���K��O�.:��=��$�.��J�}��C�ɕ�5LZi��Yڇ_g��UUOT �3!k�"���'��}
��[rx<nX3\���g���6�|b�ܹ�2	�`��_&-І%��)u���� ��U��,]�~u���O�>C�D�Z#�q�aAe����?�kv��5|;�N��lu�*�D�)�*�e�eZ���P<ߙ�ʶ��+G
Fi	�畸ўV��:)V0��huu�ʕ���7���*X������!���M0$��y��A��q6�֖W��n[�R���_&��8}���;�?������޻��g���H`0��}����W���gc�[�5KW�/m]�u,X�vV `�v<�n_I�܆���Xv��֗�4�~�z��(�NO����o~��W����H�5�����뿱�(0�b�WR=�2��M�2G�?�#ƾ��̖�<��Lq0�77�0��lY�S�M%���1���
�T>>|�����5�����[���ᐦ��0 l')S�2�r.8;y��m�C��h�N���b!�j�dwgR�S�FGG'P�0����1N�6DK�:=�x�!I`e�{37����i��
:�@?����:2��Ei��j��3�Ń���HS,���fn� �p:��#���2�ώKփ�Y�Ӗ�ۤ�1ې�auk��WS�3!�>=8As6�B���㙀��4�˂M�.��藮?'{ƖG�	Yխ0y���ƚA/��Z.���)w��a<�'�(5�OjK���첐�PV��z'sM����`�,%���yf�&o����,���?� -�}�ۅ 5�ԴX���#�Ӑ%H81����78ݺ5�zU�N��gϞ�=x�=3M�U�n�P�����5��4����j�'.­d)�Ny�����Ĉ�Y�$���7�r����o޽{��K܂2i���iR��rf��Ov߼kj�*��H��&�;�����Z�/^��AYXZT�������n���
���{����;��pR��F����/!W����X�{}Kn�	W�p�/^�R��X�.�!��	�.����7n@��Y�|xǇ2����6�X&V-/.	NY={��g�q�ۓfu�9	/v�R�^�V��%�;K�GҦ"2M�N�'�M�=}���J���1)~��]�kKW��|}�:���O�<���α_s��W��N��< Cx5\/i���Gl�Lc��p�j%����Ļj\�!��ׯ_�|���4O�s1i�����'��������H8�����p2�($q5�nCF1(�(�=��@���d@�'��Bű�!B< l1�t�v�-���;��xC)�W��*�K�j�ɛ�m$�L��Pi��kkwo�z��)r'�m��,��	�V>G j`"�iغ�,�aQ�b.���0)�Q�m�,~�_�M�;�u��x\됱�db��B�Q���	��]��!K��կ��G(`J$�Qm��M�g_�UO��s�\]<�4ATM�Ϙ�-�@�ƂaEZƓ��[ݶ�b���es&ӇM��/��f�S��fg��7R���!�C����7�=<YX,���A�)�����>|����o�%&�������e�q��e��sz����NV�}�SZq�� _S�)toU��
j��O��H����k��8��	����1<�5��G��J��n��vu:��5����d ���$%?!n&,�7��z�����9�-�ܓ����b����ܬƾ�hc�Kj��Z1n	g�Vck�5���/��u��/T�Ja"�'2��p
|/@@�E�*U��Ŏ]V^�X�?݌,�{h�VRS�d��CJ�vEK������We��r����7Ⱥ)A;(Yae��������=I��~��(�p��[$��G���������yU������������k<YR6��!"�W4��!����߃{��p�<Ud��/� Q[wc��lz�C�U
�4�C�C�ٮ/;C�Md�X��~��b��rC���ٮs
|U��H�f:���p��3a)�re�s�7���j��7=ŪRj��&-�5\7�V��%ԯ��f��m�R��8�Q��A,�uM������.���+�v��ܟ� �&�-��|&���)v�At�Y�_��,zlF%�o.���ѡ���,�C]J��jǧJ_�F:��u@\Ъg�juYsq%�P&��K3`���7Mӧ��	�%Ш���dr�˚�'��e�By����N�Q�L�e�2����7F��hQB�Mm̈��G���hg{�U��P~�˟�	����d(t��;̙���&GPY��a,�o�#���U��2����#����fҊ���xogk;ֽ�;�1��ϟ.�������g��'˟�����s	P�z'����4Z5�-� E��Թt���%�ks�)=u""y}�����)0�PaD��ſ�Ƞ����0�$��Z���U@�./
��]�{{i]�^/���lL̕��{c��d$��$�13�,�8���V�LGw����&4�L&E��,�.��Q�����é�aba�Xm[�J����}�}.���o������]�&��c�cI�ׁɡ�c��Jf(��GIC������!�f�&��ܠ��8��}�ڎ�
ş��k�,9co�m�M��W�F
����$1.,�65׹�x8,�p�-�.����"��g�!��P:mܨ�9����rV��@BE8N6~��-�;����O>��GB�<J�\M��jO5C%?O����Z���H|
V�ypH'D< {��Q�Pi�{Xcr����7�
P��Z��'hS�Xx�B~?��و�C[a�N�q�r:F�!4��0 S;���X��"�
��*F:7�����y�ܡ��׃�3<)N���o�?=Gr؅{�Ա0ZG��H�YYA���آ'���R�"~��Ѓ��sE����ʁ�p����.a��pԟx���*�:��t.@�[�l&�p�6�Aڋ/~����`C�ŊU9���I���X�R��q?��7�|c��nv�ֳ��<��VP��o�Ք5��,�M���Bem�c��i���Ç�}��Q~(���L�ǽ�0-�EhI�y�c�B�'��4.�8~ݾ�/�BGL��S����@��^�~��O���Ukm��N�o�TY�����ڍ%��d�9�8W�^��R�VV�����ң-�YD T:�� 4a�\Y��..�����;�VL �z|���c�P�x�fp$�1ї��W���g�X���.��Wp�8>)%�bo;�KCu$*�<×���XD��'*�u�����P_��T:��4J����.�a�5���cBV]���ʼ�V�믿n�Ÿ���]��S�j+8��D��/�))�0�Cz��=I��|�l;ոZ�8��A�DOP����yr�J;�����<�3���S��x
��Ȣ�e��	�8���A�ѱ$F��ˁ�������Y�c�#٢���L�����4	t�T���7�q���&��Ah֊�Ў�P��K�NOp���;>|����WD��GuŹ�Ke���s`}���Ϟ��O4|�:!�	-/�o!9t\�
��¢aI�/���.CVb<q���b�K'�:����z�0�N�l�k��$� ��:Hd��C�F���CA$�P�hш�#��1�pN�)f�vթ������14��f�-)9=qe)H��văJZ�"��#?�pj �X�K�ϣ��s)�-<���[�hTZ[��|�� ��f��'RK�~������.|��Oo߾�Nҏ>���w�w����j4�P=�l�h�6�����_��<.�l``{����d3��(���6���5��.nİ���i�(lr(g��^W8��1.������զ��?E,�X�4H��E�l�)��E�d:z�V����d
���]U	�	;34�Q��!ԃשb�w�(Y��hHl,M��׿�5�C�vE9�uNې���s�Y`�f�pAݴ�\Y��]8�th}��6:k�qM�U�<��fR��~����ȩ��n��6�%��
Ռ���~�3����������R,�A�[ڡ��
�>�o�L=���#E����[�nU�Z=��ϼs���+���W�N�\��š��1�ՠph\XH�7�m��0�� _}�՗_~�s](��&j=������	����4�{����N�c���p���/�R�M"�����t6JӫTx� j�A����pMF�8d��Xz>|@� D;_��	�&׍�#S�gh�X<�	��S���sώ=�,娦�j���,���x9 y�md�fn,jc�%��p���bbe5��s�/�~OŲ2=%.�oL�c~>ĻI�?�w��X�R����UJm��@r|�Sa���9����W�K�����L*��Κ��+𝗻���x�"�~G2���K�@*p@���g��9c4
���z5�K�=�{Ll�-P_�?�q4
e�:T���\��>�a4�iVk�6K�Tμ��u���>n�������i����h�ħ�g���+l�j�tgw0��aZ�Զ�Ωlu��y	�_Vg=�sy�m���w�mq�%�QVYF�D˦i�����f4vs��c��t���v;}��\=Y�9��;W��l��*���\rP]�^��τ$�i~����y:Y?�F���G���u^|���M�B�$�?7�Օd��K�I��	_��cғC�é���dL�=�y�"$�'e����N#�P;KF7�4V�J�ι����K�_Zp+�F*�-�GM�k�"��*�����d<�c�m���w>�`meU�P�����V��LO�{�T�Y����25]1$��m(�%-�S$�n�6lD�V[*W�8]�'
�tFw��[\8>��2��Pq��A)5�pcm�̋Y.��bm��XHx��*������a���!�#�:��B��޸}'��5�*�@���͟'�ݻ�6�u<���m���&���]l1�q6Ųx�'=ܘ�VR�<_F��I���j&LZ�q�nτ�E������m<�n����E��o��_���Y^^Z�����q��ƅk�j��$�Lbf��!zc�gE�JFqS�A��Fb$��S��a�G�ʦl��'P|"!��Q�,��>�o�e@�}Op]DSw�ޅ�ýƃ�4۶���Y�)��Ɯ&�l�:�J��t{�W��a|.�(��IQkI��?�Dl�Ǒk�`b3{x�'YN�UU��ʥˈ�#G�}��g�Q�X/�3EB�{u^����o�����p��]X`60RFR��Lѥ�2r��B
�M&�4�ݻ�;��g�+�7yUr�N8WHwX<i�*�g�i���?��'���u�٭�,�Ė��*�^�� ��+i�~��W�{o���C1��/
Ų��x6
�K��>/�D�/��ΐ�U�ǭfFz*�w懗Ϸ�_�K��߃7t��Vq^H��Rl�>����΄�l��o�ghxT�;�?�@��|Y��aC����	GHG����FsN�ǟ����d-��_2���w�> �H_
z��$8&.�Ea_�Dt3��_�`ww
�(����k��o�0�A8��ν<��^a����(!�k�j��8����v�9��4>��k�@�+9���\Y���V�6X���En������O�<E<����GX���䑡/V�UdX�0�x2�����L�t�w�����-*zk˻s������|���譭7-�8Ԯ̃�|��t�X���v��JG�P ��Q�0�v�WbM0��j����{G	��˾v:Kϲ0>�Au��8MG:�><;ÿ����"9��z"C� v�>�wj��0�Xg�h��d�'��xR2|B����������eh;Kn�h�
[Z��b�˓2��~����Ϟ�������
Tm�Iw�m���p��j�&�:�w��_bUY0�u��m>��p�ӬZ�{G�'G�Ǹ��_���j�3���č�`N�ō�:�EF��p�5T���y{��1�i�`��-<eXاO��k�^�v5_�z<�;C�YpΏ>��"�F�s!�Y\Z�xq��˗/t����xk�8>��B�$Y��F|���:A�L��U5�]d�r)5K�w�-l���^���G�qK���:;l�mr�2郑�K�O]� N�3�s��8�أ��u�U,��pEYp=�v�����ZlG�5���P�1�mY<�2�J��j����֫ח/^�%I�L�^�~�E��o,k�kc�&IF2�PbL,���dl���nk;H�i3I-S"9����~ii����v�f��K����W��ad*���[ZТi�S�r L�Y�b]y��SUe�B�����/��ǲ�a&�#�׿���K���µkט������%�@�Ze6�>|��ɓ7ovm�O.|ȹ2�x2�t^�Aޑ�`�'��ÃC1=y	��㮠c�j����d�M�9G�xﶚ����Xj�J��ƓkCә�!�
7��7�~� ;4��Z�_D>�{¢� MP��GDb"&���Np�%<�i&�IJ�̞Mڊ�k'���V���/���m+.nb_p��u�I�sc�o���Z܅{���NG`ڍ�C��#�r.�ȗ�� 	�wYpr�)�L�)�$�R<I��%F���l8��o��RF��FQ�����?f��Z�1y���^�{����曓�AҊ��T���2nf�/��/�8Aˈ�

���;�e�<S+2ec���Xe��N)���'j�Ig7�$�$P&.W�gjI�,TNE3�	���c��da:i���t:�Q! �n$Q��\k�#�Q��!j�#_x��	��l` t����h���<;�>�l*-�A$m�jO&c�� l��8�"7�,s��
�ݡү�	�sn7s��O.
��6z?ji��������ܾP#�#t˼��./vڭn�b��B�B����S�R�̑áӦ�!}�����{6i+6T���D����ͪ rH��\�bd��c�͔���F1Ś텥Q�j6Ջ�珠t?$�LEd��~;��>gg�]�!�瀊����zs{�Vܼ�������\gV���2���O���1���c��s:�D�o[�a=X\pc��F�m����}���1Q�7ǎ���0)�*�14����%%�9��`�љ]�4�5�β[���a��9����}�ݦ.��C��Æ�J"�H��)��=&�X(Y�YNXri�΄�S3V�Ņ�tx��%<�t�(�D��NN�V�R[��]b����ռ����o��o�5J�>��Ӻpq�ƍW�

���5s:�2������<�\<�W5�|S;J̳�b`q�qX~���R`�fݾ}��p�B0���3f@�YDF���)J�l�d�>��8[�.q�|v��x|lK��>M�vf4M�C����_�ur��)�m���LV��ܹ�B��m�v�=�f|d-)WH(�E�qT4-�z���<,�%j�@.�\Ys[�dJ�&�\����˿���6�ֱ)�8$�n�n�rNϘ�>�L�����ol۵B�
�4J]O��U�ז;�Qq������ӥ&�g�� ����D�p��}�3e⦱t�?^\Y��EM+CD�A���Na�Z�$���U�\sZ��+��T���vz�ӧx3��C�m��=x�ݻw�������'2�Ҧ��;R�l��m�ךg^0H�j����3���ʍ@[@�g����c_ �D<��4jzƯc�͛7�N�C!C��ʕ��P�$OG�l���p�컄�C �'(��`��6�'�i|�����b3v�ᔅI�9�9ʡf��Ve,��C���d
�bӊW7�ζ�I"`���g�3�f%������J&qg`Q��:��oy9�*���"��4j3N˳����'�����<n���CA��f�v��w�3��NjK�K_����w#o��xO�������̐ώ:��������6������S7:@	�����Db8� ��[��d[#.�F��2���H_�5I6��L�s)0�{�{q��&J-wz:�,����٬c_2o���PH �:i.�a�E�B��zxs�<���T	�/��vuR�6|��J��p��/��˗�_��B������FB�;-��2S�:Լ���{�1_�'��i&[f�Y�8fxt����v��l��4ZZ����o~����'?	T�`1��X|�q��vb���������T�텯ӎB1�����X+K��%�Y�Gp)�_��W{{;���i¥ L�����W��O�b!J(l7��DΰΌ�_=����'�;�䌏G�^���DO�a�-���A��uU��3�΃����e.�3=�;I1&��W�)����d�6Y�
h���~�`>�v��&|�TԚ��+	o�!L�v�D�d���`�n�\���4FP�_�@�%��YL�u}Aa��U��T
��	�Z$�IR���oNT�R�8��G�c4T�)��k�%�7B�\.6���g"�߂�A>!���-e��P�C�x�b��%x�g?���|��|�AM]hC)p���QZ΍�T�)��d�fF�Gs�n%)�����kf�ʎ4:I��Q���RF���ZyѴ����ѡ��ׄ�ous�ڵkdgv"]Y�*XFaF]6^F(�~����v���X.��/>�_ ]�~��W�^ݻw�tq�[��y}No�Je�=|��ᔎo��2�M0]w�򫯾������B��/��I�Q(U���?+�Q|��]*�����L?k�m��z���v��jI���stx����D���kA3UI[]�-B8�6�Z�dx4|C/!m-���B�-���V�����l*᷇�i5�&�K�tPk���+��h����3�����F�a���_��2�dfy�eBt���L�i
($4�bt"h�W��ȓz�v}	H���g� �j���n3KY��i���sT\�c%"�|�7���O(��.�DL4{�gܝ�FJ��[fm~���.���O��,�ᶕ�*�zl*SI��6�ǂ9�OV�F�Q�N\����|&ԙ6-�l��|��}�o(/갞� �4��t�Bh��_���#��}��|����ɳ-nx��hL�}9!�Y��TZ����YWb�,�o�K��������|[���.!��B����H�s<���m�w�:]
&[8:<=���!����0���X���4�*3���D����jhaI��y1���ә��{�y�Y4i`a�<K��</�<>:-�:����_��F����piu��A���o��|Bp>3h������Vd����@F7��`�j�C���eM��
��5�[j��OGc6�@�@wqT�Dש����jи�Ic���X�yqq�f���]1�>`Q�ٶv9(����*ٹ�4Q�(�T���P��u7S�a�������6K��:��u)�V/T����R�D�������N*8޺����m#����	� �W��b8�����J��UK2W6��092)0yP�3B����:a�p�+\X������+�VV��]�����;5B�?il�/�㢅��6�j+��>�XX3�7��O?�w��7�4?>>=:8�X�<;>�1�pKM�����Y]�݅�� �Y���L�*7��J��5��/n�}!8��Iǎ��?��<g��lDoϰw	�:d�+]R�ހӧ�Q�J��pGt؁AԻT{�UB�e	z�L��0�A��Z%��d�s&�^x��������0ɂT���4�rg9 <�B���޽{��-�������s�{]�v&�3�K�V�$ ֶ�v��Y�{��3�*�(�B�9WA�A���h"�i���3�!�̻�k�f��C�rb��V:�t[[[;�;�����X��Q����>;��M�d��s<�"/�N��(hܪ�il���z�9��Cpz:hu�u%T?
_P��QBN+�e"6)���K�Y�*/�?���}w{{T�tK���Ģ�X��=%7.�n�5�X"�8w΋�{q�|���7��i'�������իWz�Y��>=��F펊�v�p~��.�a� �_W!�Z��Դx۽{67�z�WoF0\g:��0p|���>���0KAa���a��u�9ZW�b�Uh 3�#����j6�;K���G'�����A���M{>{��N�u�҅����{�R���`y� V:L��r3��Sr_$9:B���Ct����\��*��|F��d�`������ ���☎�͍����.�AW�;NEQ�j!��6�K=��L��3�������#�ʕ+W�]I�J&���J���3Z���ϑ�v�C�.�q�O�N�"�yY�H#?������*�Dg 2�q �b�IV�LJ�
�����by��a���&�F:�P�م��o6�r�VV'�;�v��k����Z�����q3��"��5��$X=�X�1��8�Y�e�r��[ N2��¥J[�xTK���%�:N����
&w�Y��x\?����q����iH��؋nR*"�1-w/� ���흝�������I�c[�������F,L�5#�M�z{{1��PX �0,�}�y�� X'p��?�	����=R����?�k{��5�S	 ����D�q�|o�l�]�)-�=�;��͜1�lV--�X@r~�|F��u�6�D�{0�f�q�w(�G�=C;�T��������ra�����	�?�py@z&��J�4�{�cdS=�N��.�`�B����B�����Ⱦx�1S����r�
����e-��t3�SqD�T�G(��ɓ;w��C!�"H^���?��X�Bд�x�ӱ|��`�o|!60�fBK�픳(��z�
�vO��%-�˷d�i��Dn2�e4-���Ų���(�^��*=_J������r\Q.i.�U�*�8]j��I����\I����j������ZN���Adm�K4��������O�۷o*���'�u w4��2O���X��Q��:�3�����g/`��}��+�����{K\!o;�L짦�l?���)�lb5>�EA�j�"����o=z�o�xa��S*�&"����4
���(=���8�O�?�)���D�����:�.H|č�k���&m�*���ﾻ����0�rt6l%�4m+2wha��Tj
��7>{��͛7B���NP��r�d�!�T�v�q�P����8TF�.e��K�x?��	����&+������o��0P'a����f!�6Q�dR�K�$�S��^�����ݻ�[��XD�^h�ҨIX{���}��4���ɁnGp�2�u�Q�qA���?:98T�+�ch�����щ0�#����O37T��\V�J!CT�p,a��?��(����bN���;I��Yq��r"�L�3��y0P��^�	k�`���2��y���-�x,/��h0|������������)ϊt�p4��C��A,�>���T�F��K�-J�R�Va�,o`�y�SD�����ȶ��22��l�H`8�}��]Y*��$��B2��.�B��B�T�l�F͉m���1��-�6�|��i�'� �v�J�f8�<r�#*M5@'O��U�E�6��A;&��MHv(4 �z�/.qI ����/�{�"%|��/�MݔU����3�ÉL�e�H�>�A��Mge>���;���l�I��Δ��ڒ({��q��_�k��(�a�4����"?��D�,���C�Bv�:��Ѿ̛���KC�m�G�4^�5ɳ�~c��9Co�̻>�d���m���~��|�ۉ6�G��5��J	��!�(�`0�e�%І9�����Jg�a���$�sK�͸�;o�RR��${�V.0�z�X��:�5qO�����1�(�iγ���;�'�R�i���a���2X��H`P���|�4�w�کo���!*��}��9��zZ3�O�ʱ-ejeM�f��Uv�U�.�d0��Yҍ�w��M�G�w.�')Ko�l9]�E��*e�f��|�)�� )fJ��`l8�T��	�j���j$��7*e��M�?ZY�Ź�e:���+�XÉ��ƛ���>}��
<�|@8G�@�+y��T!
-Ri˳d�x~�r�H�2������47]��eY���7��:}nR�p��85��N��#��B���W`G�ԩ����A���'��D��im��d2��{�@7���Ud�G��G͆��OdX؛�k�X6�K���I0I#�^mOG��"�,���j�L �uHj,����� �&M_[L���O�_BfX�0�_-�oND��(=ӈX��fR� ���:�/�5q}bKFƊ+�~�p*�R�NZ)�*!]��ԓ�֔T_��#�pM���7��'q��c�C�������7 R�	�J��F���O�����kt4�@�4�$t�7�������GRj��8�)�6�t�FZ#y�c|��s�޳�^2�������;���ǉ;�Z}��H�Z�BD%���Mn��g�峧���'>R{�4N	dY�ϕXY#�MLɡ��b��x:1�&�i�m��k��4-��
[�H4(���I�5t�E(䳒�dS-=Z���C�X�𕹒��pE��ԙD��n��%1���p��&���ի����W�?"#�s�@"�FeX+��	�g�i�"�h�R��\�h=�	~��ۑ�!b�]tT٩���p'_[B��r:�w�Ҧ�_�Y�0&��I�SkE��l����Tb��m�e6˨�!���t>��Sr�0�\&�(��1�cHKK�	�7ISÔ4OX�`z�Q�lF���@�!��ɒ���'�/��ዾ#�+�޵��1�DnB�iĖ-�@����H�gC�vhm�����2�w�n�ظn��BW'�Y!-mjEh���eΠ�8�!�+�������Ee�;�e�dO�����ֵ4{5�4'y��z��Ah���݊�L`�,���S�.(3D��L:�Op�*K��j���Ӽ��J����w�\h��Ba�2�$���%%���C�ۘ���"$�2� >��;���@L+�Fo�S�_���*g�(�X��2�a9��s����T�t��֖���^�g���2'#߾}�zUE��
�6T7k~�vW>������EZ@z#n�-��O{|<$�!kH��@{#�2�5\*�G�GZ���XBP<~H��ꖚ�wU�33�'w����h;_�uk�
�ʃ��X7����������2C�e�e���Q;���"A$���Mu)�f�����Q��^O��7+�>�j'S���� M9�ɔ�9UMc[𸒱�P�,��g�";���p��{V�._���{�����-HV�M	u��BUE�PN�SP��S�>O��9&1T�إK�^�xAWWf���H��?��N�%�2�gBm1�~ܭ����B��ڐ@��x�c�U%�p���>�?�ɪl/�h�/�pA�-���i;Ė���ux�)�C�*
΍���Py�^4�NѧOǟ~�i���5f����ل���T'DZ�η�w3;���5w���k�}__�_����)��X����\///~XX��B	=$٭���<�:�Ҿ`�w���]ѳ0W�WW �=3���#r�1��ijKO�γ��YZYYꊮ�Rc��^�&ݤ��L��eZ,<�V&�"���uD+�qԢ��y�^�fp��y�a�A��BU�xJ��MSKЗ���d���*U�3R4X��*6�H�i���HA�r����iVKє�y�dc�?N���W07��+�\YO�ł�Ɔ��9�o�j�m�p�6��Q^ś��y��������7�l��?�
�Ax��$\��kn�y��J-!�J��I������n�ĺt��=����h��LN�	��������Nŷ֚����>��ݚ�h����p:V�YT��Gǒ<
!ڄԉ	�k��E]�`�wl� �γ�-I_=7�طmε��=SӋ�}U]h�WaUG��T��(2/R�o|
Ʀ��v&����HEDϨ#Dd8��LՑA���7�2���%@����;���s�t���P�(��˛��qQG07����L�N&@�OEiJx�#Op�pbkK/X۹�&!�l˂�!fX]^y���LW�	��*�!Q��'v�%�tmee�������V'IV�J�-/�(�x6�lC+Y=yh�f42=y��\�9�h$j�Ѧ����\w� ��l�fd��~'`��$�ƫ��:�.=3�Ŗ]�jH����v�����I{6��vvv76n߾=��Mv��)��!Y�x0�a[{��'J�'��1֢��$ҁd�n܄a���������}�z1B`@�A%��D���YpS$�u��[�7�
��;���\��	U�S������n�[����@�6���oB�h��Q��Y"a�ec�?B�W�^I�Nϼx�L�S��_��P���c�U��qy��\�5��*�$�!k�$�X[�c����p�es�ht6�%�k�x��VE6i5�.�����#I�J�� ! 3?��m)� �n��ݻ?����ܹ�_0�U	W����P��֛=��Ç%H�������ޭ��.���Q0j��vW�����G(ͮ�ZK�UN��xWZ�ƕ�g�g�a�����p�a<%�ٹ�]&�D��{�1�R�K&Z1�,���������E�+ZSM5i,(f�@�&q���� }�={��=���߅�� �� ����(Z�m���8Ý`��|~���Eq�g�����%��i��k����;�yN䡇
����l1c�2�
IfĘ�t)�~iiE �l�4U�)?8I��e��0�me�ڻ*���qǳõg�q��ׯ�������7In��W_��|�tIECƭl��E����x(�ܹ��Ñ2�ͨ�g��>Ҋ3�ȏ3.�s�g8�2�ZS��NU��<��I!�Z������r)	a�&`H��iЌ�a^ޭ@c)>��]C�Q1�k��Ƴ��76�2=Y�m�~P���3�S��G�	�����N+m��h2��ൢ2�m?d�n�	Uae�C4�58(�����&8B*%aP�+"�f�Q2&��y؁�薁}P�:S]h�:z [��#xe����&ô5����ʪ��k���o>���̲8m��^��ef�ΰ��?[,�$gM���6=�����[Y^e��]�BU�^�QTb8��q-C�r.�` Q�88t���"Jb��È�@?Ԗ����I��TZ���(3ض�dfRE���=}''��BG�8T�WRX��i.���U入�>�@�(�;#��^��.���z	z��z��(Ԃ�	7�Op%��t�n�9iH��{@#����FMJź�|�٩h�\<�:oL�r�
v�oh�/�Q���C���Z��ٰi�����e|j�UkY���K'�����!y�ZL�̤�,�E`�K��U�#��XWq�3~�i_z�Ku$|R�il����$^�8o�&܆����M��W2 �ETFv����X"p~;����SQ�^ý����P��T��wwZ-@B����*PLG������)��ʕ+��xqyA�M��k��'��c�J�d���W�ȽŅ�U�L4���ĸ�o�t,�7F��`Hv�@��EhGp�e�����6�L�NN�n������$��]����~a),�!���[����i�,j�/	�N*i��eoܺ)L,����vv$>�kQ��s�~f�����|pI�,����_�v��j�c�C��fȫ0pӒY�`Z����E�s�@H$d��M'��J9��\I�Ifp���h��~#RY�F>�&I���٣����h�S�k�i�{���mm�g"�k[fڎ����bm�.Z�r�N�@>����ϡv��Q����Μ)J1P�嚤1����߁� k��O�$�
���� ���z���6�����<����O�D�����0��²�#�����ڑ��޻v>y�i֙(�$�a��DL������G2+�6eB8��)-&,H�P�D�M!��=���/��I-F��E�uU�py�u�J����<\��R�1��B���*&C��r�X�R��uhGM�ϸ�꼽�����V��E��tz�-�/..��MZ	���0�������W���4#���zKY�%Ѐ����L\�ʖwN�*ԛ4Ɇ&�L�ф	���0�ʟg�s�Ѩ����M��P���(?,� ���iA�[�n�O�L[1�Ŭ�䐀Mo��ػٴ�ͽ&�$����-sE��,�9_�{��H�8o2�8ZZ��T�WW���nOS�͍�"4�n�3��q�}���k��|<��ʳ����Ri�<5��P��r��C�s+Nz�δU�j�i8�UP������i�i�����Db����`���.X4���,�Qc)�i0�40��Eu�s��ޥ��ggZ���Z
e�.e��R��*�L���C��wVm~��B�s9Z'�9�w��������UY�8�ij"�q�/Pp�VW�e4m��ؙ80<\%b$�;7�ƭ����#%�\Y���U5�iWN/�Ic�A.��}i,�7[[�?���t��49�,=�&}�s�\�8f�R���X�`څ�a֜�1-��@#��ۄw� e!!�?˿b|pqa�$��ڎ�#JE[W��-�e�0#|[�*���Zt%CK�J�!��-��N����1��}�&K.8h}Q�Q5�����|���t=kR�x�Q�m�+�����v������1e	a��` ��_���<�new�Ϥ!o��0�[�'��38��?�S��/�`*$�0BN������D2r1�'
�G�t�L�����o�\�%ll����#W��i)ܒ��ګ���@ �[X�[�H��tHC�����z���ɠ�������7��qW�C��hq9�η�v�Grq��xFJԞq:53����/��Rr������J;/xay��:�`�<��B�pOq��RT9��g;�]^�����G]�z���.3�)J�� 3� x��գG��Rr�'D����)�3�
�g�ε�.q�����X��S�pz��:d���6��x����w|p[��p� *h,�&���P�v�2���7(���c�R<��-爜Pߐ�R8�u�`�g������������e����=0i��xN�8������Z���a)��"u�e)b,�+����n>]��M��Ck��X
���m�`ӇL��g�l;��k<o�\fܷ��i�R���_=���4��2ޖ�˪������S@B$VI�i���mJ�U$	�]����u�[2�0�g6�\t��B��(�D���˩<;t����uW
4�=������o[�k;0����\��sK*�VZ��mܙgA���e��P/�{�P�.˜2���s<��|*m���0
u���VL���6���F\͐(�$2#5���K���xv�BU���9����w�>�lM _ZHlh(�K>Ka��|��a~P�[�>�ǋ�˕m��	-�v�QգƱil�:����jm�����[떘D9a�-���)"�Þż�G�Q�\(*:_�ALvܙIkL�s(H�#^jWx����Wc���M<�OH��˗!w�܁�Q(�ţ �\�Z����,�F���mi��t�T�?���S4�G\�1���	���s����?\Κ����Cxx~�+��S�v��)��f��~�R�y�\RrM�{]��� y�\�10�̹
�c۶���E�~��&8��j�*�֕�9Ba������䈔2��믿�xQX��$Q@eNM/�u��8��~�Xؾ�]�Y��uE�c٠���h�����g��$�\��+]vu���{t0�#�H�G���᳐&;�z#�X�~��s
��j-s��]������&���1�����������io)]"�0�/���᧙L��.������g�$>6.l
n.
��c��E<�8;�-u�83V���$��T�=�J�\/��Ä���&�����<z���F�葉��N��Sk��	$Kt���R���&���;��������;dޜ�	�;在|O:v8K�U�� 
``�-�GE^lgPc@=��q(�S�"�\)i8�,��,[<wϼs�t?4a�ʿ��noo�+�����B�:=��$�Y�3_�G��Ry�Y��o��~��zI�U��{��>���e��j��JL����2�;ױ����l��y[Yk��qX�1���T��o�T��H���������e��qqG�^Z.uB�<;ߒ�� ��.�lSm�*�g��\H.+�x�ؔ_��W/_�MR�_�|�_�/	��~�ZB#�2�����)
[$���0�-�@S� �ʂ���]�ƺ�罉t�WVծy�e?̭o��q�{s���)��^�r6����3�����$��R}������t�	��r�̇��Q���Ρ�Cq>ac�z�L�S_�A��4�����M�h��J���T�g3B<״��S���I����,�`�uh�_Ѣ)!�0�uB���_���{�=1�8F��)����F��C;G�+=Ӗ� ZS�$d@HcƬ�$1����М'�|�@����t���!T���1��2aMF$5����i�#�L�ک��GY�`.qv~B(b���*{W���{��!e��T�����	�lv�9$f�7�^LG�>�^�h�p� p��cI3)�zs9l�zGh�C�?��)ִĄd��_���VM|ZX���C��[��(g�9�\�hN�r�R+/>�������S�=Pjׯ_?��g{+�4l�ե�O>�dsm��ٓ'Q'�f�/�x�w��ܪ�^��fyy�t0�Sȯ�m��6�G��~@#+�)�L:�]�>e:(�c�N�a�w�@<��Ps���M1ū��� V�2x���!��+��uBM���l�|���/�,BA../0�A�q���<28�������:#a���l$1�T޴M8���e��P� �J,n�RG?��Tj�]����=�B���զz����<~c��qz�"4��C)�v�� ������iuF����SN�Yj�W���و��n˫	��� X�E�Z �\x��E&�������0
�L<�(��Ӫb��@�͊7��H�-�����i��}��2|����]R!M'g��燍xB���/4Qѧ�ʬ��2T$Iz����mB�psp���p0�����פy�4�ش�߸q�����?�˪�ª������]�
p���Q��|��v����A1�Aa$�����?�cb/NN�ܻ��[�ǋ`�;�9���&��0y��1��}e�-��8�E%	��;�1�����K}��~o2�w�0�bH��b��D�煖hen�X��~�� BQ�}���3i��@K��TA٣Jz�Ҵ���œ¼��ZF�ѹĥ[�=�\�fa���q�5��s}[z�}��1�Y��UMYb^���8\Z:9::�?�d�f�
��WTA(}"�lƥM�UPC�����'a"ԝ�S��J����=�9����'O�PS	�Rl�r�D���+B�j쑛Yw��x��NT�m�v�:�<��\�'׳ܩ4�&����k!�>�l�^�˥z��f�1Ă��ܲ��H��ڐ�! 2Y� &�פ�V�dj�o�Xd�(����7[�캮��Sx���sH�	��D�Ē�Ԫn�hz�o�驟���6+��2�Je"�I@�<g�>�ߩ���쮇v�%��=g��מ�6����u�%���B�cm*Q}
�%Ccy�����&���N�q��2O�� i ��kOq�2��X�@���'EJ�E�W}%_Z�U
.s�EN-kX�Zl��& �i�Ӕ��-N����[�)I����/�����Br�ZXK���6��`sxxt�ZEn����e*y�*U��6�@5!gV���(�:i^Zl��8�݇��B̦��#�	���Wm�-XaY=�SlU�dY�-�_Ȏ�,�E��ǅ������;?��S]|���R��n�Q֊|JJF^��D�Ǣ�7�{O ����m���o��;b?��qY�3�+�+WZ�j��R6��X���q���1 @�Z0^��ܬv�yܳ5R�tK6B0O0�9��\��5�A3�K��^P�MUV8J����� TK���qC�*�d&%U�T�s%�6q����W�L��>���g�[�,;jӬ�Д"U��2P��NRC�>}��m�ѝ;wn}��F�f\< Y*_z�n^d��E=ْY*�U�(��|��c38�X���d��Uu�?�i6YQ�ꫯڰiNPR��r1�k7#�y�b��Çi��?�P�w|$(��#��:�;��V��-��{�"����~��պ2��������m2�� ZU���<�S�8�[ �5�(n޼	�Aޞ��!�ʶx*�oz���3k���)Oe��?��|��,�|c�^-��u�Y����u��3��o���E�,�s���v�N��{C���|��%*��ճ���ۦ��$��8m�kU�(��>��N7�N�ɖ	��}��}#�k:�+g��:��c��JE��b�-�
���c�����}ʠ	(=��tm�]�'�N�!��������?���lv.�=�tf>�֢��={�d9�����1�]|K��Љ����	�Il�p�GhQ��<��ǿ�+�ASs�o�h��[���e��HV�t�Kk�l�X���p,��1�߭[���"�dZ x�_b�:�NgEA��+�L�^� :/��޽{��Y����Pt2�Wu��0�&��[ �O R05�$0����<뱠���&����F�,+�h<| oZ���C�Ccu�Q�X�$��\�Õwv�qPY���<�t��0R�nń���g�Q�0��P���@����H ��+�l�ܓ(,����S0�Cg����&i�f777$f�~s4ע]cP16[F���D����{���Z�3�ߎrS��`ѓF1�����t�r?*�X��3t��jO����jϪ��ޱ���Ǡ�!�D�a���p������>��b9�"��&�6�Dl,����"�d��o#���/�"0�a�e�#%FќºS�ց�BTao,bഒMs�9�@b<k�Z=Z���P�o�<��VŞ
4|K��E�ן'��J�5Y�B�6(P���SH��P)�z{"�hm9K�g
��7��!D'����WJF䈸���R��(�T/
އ���o���G%��P��Uj5�
�U�V��=!��f�Ȗ�=��K����`M5~��r�
t�f�}p?��8����d�,"_��/TF�crJ��݀��;=�f��jB*��lQ�2L���
�V%0�z�D��^l9�HzX�x�u�@�PD��(�ӗP�E��@��)���t��sS&%*�r6�m�	pJ_�[�����=�ۊM	�T����$P�;2��ڳ6d��}�k��C��[���,�]�g�j=4y�ӡun<���@?��8�R��_��֬_P(_i�ȼʕ'�	�zj��U�	�ނ	��ݻ|�r���*�#O�ɱ�D�,x"���j�(b_0���r���p����s�_�W���:�����'O^�y������߫���u��27�:f��%~|��I_�sk���������߿��ǜHk�����O"s�W�����o��5<�ڛo�������`�����
�	+@��3�F��ԷK�ЕvV����������#l�l���s���|�܎��p��n�z�.�^�W��o����l级�d!IБl�:���`�ID�%n|D�y�d����lc��)��P�%+㴊E�t��3}$�챶27�JYY�+��)aS�R$�{�PUEa�㾺N�w��$R4-��Za�e���D'7ԡ������u\�LJ�ƄeV�jDZU�cYp�I,P�����js�'b��r*X��٩� \��H��V��ӧB'���SX$�V8e%`�
���k-y��i�s��,��JyV���&�&b�'��<|��(�s����bO/�]q�Y���t�n��K�ۡ�fi��!Xy���� +�L����w��`{�G_�ԄD��n�#������d�ew*zx��0�=���,K��J<�����]�����ãl
�����qTP򅅄�:t���z�g�/|�c�J�E�B9���AdR��s[�����Bh\U�UGX�U�)}`�>��jϐ%�m=9�n^�[9C�9����o��J�[Ę2���x���k���t��F�J\cP�/^�-.��{N5�Җ:�+�B�����r?ժ�A+���Q���ʀ����}�f+��-��]���_+7��#�x
�h-V(�n	���N&ӊ>pZ[�*�^c'ǋL�J'B�_��k���O�����ބ��WCkAo���	ǹ��C�G�KC�=���l|A1V��'?���Yy�6��v�ԝHq�6�	5[h`?�w�O>��L��w.޸��g*������m�i�\����D�n�W"�z�7�����a���o�Npie�?~̾�g�8���4��!�ڙ�-uj���g��gb�ګ���Zj��B��;�� y΍!�����Y�Zן!q���v����ce�)"����m�Y&
.�68�['�_�_RO�;��;�������$� ����[�]gsF��)ϟ�LP'H�([c� %R�W��`߀�ë�, �T#T(f�wޕ9Ȭ��.�H��[�B4��2B����9J�X�F�&[)�T�w��˕�\[��)E�?�FI)���� �ہ�.]�Ţ�2֍��0���Q$]s��v �
��o��b>�i��=�k`2s��r��m��/��/�-"����7j���o�����r'#��$���ȝT�
쩬�*1�_&G�s3v��ffM�n��	�����'������9���F�g8d����B6���P�7��ظ�v�h\���S���_�%Y��5�x{s�Oh��Z3�&�1�����i�J�I���A�6V��^. ��I_U!",S�̢���^{%�6���
���ڧ�5�t:t<�~������U��e�B�J�����������M�5k�L���1"�mP�i֫��X�2�B�B;�#��g����5n����؇�b���r=��~�'<�~Ya	�W3n��Ybު���χ�0l���h+��Bz,���A7�
_��o`�'����MG�S+ˊ�#p�Vu�ǝ�o����cs�9��S�����|�!�te��
��~������F�ZS�%�>�VB��Xڎ��ڵ�c؀//w"�CN�|��ms��yh_=��q�d)y-�s�]1p�/9::,K��Kڂ�0d2Hd�RX*7n^�����2��*����{]�!�z��ڐ2�RJ<�C�Fা];����VFQ�O�z��(�TL�fI��<���́�ˊ��4\���^ܳ`/5ѝ۷?���|�[�q�J���Z�C'��r -�[|oʂ��"�/���T��M��衬��.�wm�q��"<�5��80v�r��9>>XW�&�"��4�̞��|ƌ�T� �8�Q�a8D�o��Z��y�㜌Y���rI��6�	M��4T�e�*��__�tI�F�I��	��+:��\�4��&��j����/~(��Ƣ��%Ky����������G�m5��͊<M\]jN�����ts�]d�����y!��l5�-`g���,"V5�����l_���$��޾v�zo�߃H�����I�ϟ�������o��>#��j"�|/~�L4b�J�4�|y����4��K�R��f�a%<gyȨ�t��+
[*���zjT[�NjZ��`CǕ<R�c�z���:\X��~��7o^	� �ۍo��A��p�(!f�?���$I0��C �z���m5�����������/����Xԓ��ݻwTw|x�E���Vp��.�WИ
W����΂8a���
O�#�Q�� 4j,Vl���<	u���5��P�;�SN�:�^���}��s�ҷy��d�PG��j���Ck���nƁ�r8l�Gu����I��v!$�n��`}pe�I��++L2K;~8i0d�(�X�渕M�3�w��x��+l�L3!�x|p�t���t<K3��g�?ʻ&{�eZ�8�]���p�0�;�b�= ��d���á2 � /E�Mʱ+!��{j�r�����%NH�?'�!%�HqՈ�2
�En�_e����;	)"���c��]ż���3�?{V,���1�Iȟ�L��D��*��Ǒ!{6� c_k��K�����,�w�x�j�b־��fiX�Z��W��%�i��a]۪Q ��i��%2e�C,R��F~��ag��
NW9(�����5�Ao�����g�\�)�y#0�ES&t��S0gs�����o�$�KZc�����M���BQTZ�6�n2�dD���ytՊԫx2�ך.��)��9݂��m���dR��̚��b���E��[>�tª�4�|��?ul3�]�Z*]3�����ǰ����4V��cH�i�f���M�B����7G�CZ"�x�E�+�σ5� ��0��H�k��g�y���r�'q[��ЕK.�:�����v�E��%#�¾̧��-�
��}R�+����J)��+�,9�|hRp{�]���mq��]�- aI����e@��>a_{ڻ�w@��O?~��o�	o�C�U����~>~0�-�,T- ���O?��ѣ'�bK]xz:VV�L�OO��?+S3ҧ
e(�����ѣ{�\�����ݯ9|���?<$Y-n�k_������7e��Ӛ�jFmː�> 4��N&�?� jϖ��a)�؇���������چF��ĉ�9/�X]5%�"�ͪ^�}�����19^v�mX\u+*.$�Y�4�
�2�$�̪@��>5����L0�s��@I�P4kDUR�N���,G";�� 5�a?���i=:<�u�Ū�{���pS�]��Z8��k�'���p(*&)W��%�0QH��Jj<KbL,xg�l�2T�u	����Ǚ��c끣�k���a�w���x1:�����Z.�UN�ټ�J]m@�zr��_�[���Hv��P��%<�_&��g��c����މ����vT՝�T�|�0nRWw>�����2-��ʖ`��I��\����C�q�rJ��b:�d�����:]Em�1�n|�ى^I�L�޸�M5F���uk��}���(}q�77������t<� �<��͍�nÊ��zU{2���^X|$����%�H3$��/��x2�D��Zr]8�;��U�̒7I�\?���ɨ��9�0Y�- �ьHl}�� s�fI�.]d tam�V�V�[jr�1P��1v\��J�� ���hmn������i8�R;��X��ž3,��{i:u�M��P�h��<�W����t��Z�1L~�j��"���z:�/��cg�@���%�l�f�5n����T��Ȉ��O��ָ���Q���t����I"n�/1A�����Z����H�e�8�JSv�xv�S������.TGE�,�g��N����E�jT u��T�n{�RD�DL�����WFQ.���Ȩ��$
�A:2o�f���Sk�����*\�����6�d�\�)y�\[��fQ�&N{���/���ۘz�҇�����m���r��k���R�*���]Ǫ�67���Q%�ڵH_��u��׺���]�������J�e�	R_�P{��؇_���)m��iA�<���%�,o�g/���2\D����\�s�nl�w`YV@9�$��կ~��/��e��S��%"Q��Z��^.���x~V�ܳ8�Q�=i�j"�AY�>jb�Q�GC���:��v?~�N���r��dU���j�C�� ��F�R[��Ç���o�y�*B���=��/Q��SqT�	���+���{�=|�`|dQ- #p}����Bϫ
&�~ ��g��H]�B��`�$A=�*�u�5	7@��4+`�i�ߛ��.?�mQ�X�QT.�k��tD��mM�
�e���h�ɉ���鬪����a����n���̰���=w��'��%�׿u��u.\�x����\�Kݧ���f^��;v�;G#�g�g}�����2������o�>]�H�˖��]9�Pwr9_�]��0ɍQ\p��)Q�J��d����]�9A���_|��w�}��W/�^�smn��n�A���Ş�*]u0�8į�����(�A<y�H �����t*��8t8�ׯ_������ʕ+����ۿ�h`p��_��W^ISlU�;p��v���S��o��5 ~iǼ���#��.�����۳���d�&&��+F �����%�S�~j�߬R�ri�B��ҷ+?�:����?�QB�����=�S���K%:�Bi>��j�HQ�A��;#�C6Y��b��M���R.��jʧl���:�wg��s���O{W[�Lbd=z��z"�� ���77]A���LB�;Y(2�7q���{�z���ˊ�v����A@�Jz?6�!�E�'��K����P{ħ�� �V�db=2���S�h,��i땪�h�g�*��ڬq�%�7-��{�U.���_��6_W0��za�m�=G��6+��ʭ�-RX�K82,T�'е��L�+�I�[����[���e3d��r�b�ZH�c��*u׷�"�vQ�|UZЪp���@&�y�)�J���h46��|^���D]RRXܩ1�߲�����+cV5��!�zpQj(����L�x�9�L#7Yg�%�<��b���R빶x`�dF��=&~L�K�y�S_Q.o�� ʽ�8$֮UqJ�$k���Ȱ�!�KU"��~�}��?����g|�\��*��Ɠ����k{
��	����?�����]P��ߴ�����*y��3�6=�R 8��k����n��B��x�$�������ʦ	_�|���W{{{*]שW���������W��i�tp��wU��>�����ٱ��c�HXS[�V�=��O�e�q�~��'����/�.TT�W�^�5O�'X���-�j�q)��?x��L���R	����LX.���MC��ԁp}�>²H��Ef�V��T7C�3�_t3��I��^�tEr����iXv�L�%�N�X�x�b�R��V �T��VFҥh����j#JX�u3�-7)�����43 ̺$eݮ]��bV����j��JE!%c@G�!�� ӣ���Zp��{�9!�/��Rc�9PM�ΝϦ�.]¯ԹyP��b�b�z��M��`�;O_�׺�X{�{�uT���̬�0�Ȩ��x�h�<x t7dΘ���̹˟�F����x��x�֐�7�8�p�&���<%g6�L�'�Œ�^z#*[M^��ەdbM��+L.<�z�ҜJ�^�:�$~�R���ƕ��d����)d���dă�lm���p����}���#YND|��]����N��[Z���eўb>�������}u*��`��(G���02>�Q�I4�=$N�ۻĈ�Օ��@��#�F���n��p���
Gx�v�@E�'��x�� �J�`j�4���w���F�'�$���K�4%�/�±�x:��P%���u��=
U�n�\7�zؤ�b)ؗ>^2��g3L�4K����
�ƾ��1�y;E��@�Lb�~�Y�6�+��0�8���e�������ك���LH����M��;ځ]�89YXrh%+��*ܸQ
�� �6cu��Ŀ��'t'ٵk%[�6q��b�H}/�"	[�]v6I��Ʈ,�v#��c �^���rf���;ǡb]n=�m��ѕV�9n�~ ��4��G{�6��XնM�������: ���"��`��:<��^TP����v-\��]��򣸝3G�Zȯ��T�����5Yqlwk~��"0n�\�*�)���N� S�8��[ئ}�E���k� dה��e��u+*�^�+��G_���^*��xv��.!{V��ݽ{��Wa#UUaC���ŕ���N��(��Z�8[-+�w��\�dՖ+<�<p:��ç�?��*Mn����D��0���^f��n�lh*���dfP�j�����N�b6]�����8,)�r�9�r��d�ZP�s2���o��6|�k�вv	��PjW���%uJ�+��������Ww�-Kf#p$��8��Tx�-�.�-]�'ŷ_E&Nb�v#_�$0�OnuAX�e�֕�[q�Qk	��vb�8f磒�0.P���RG"!�$�m����:����W
RB&�gϞY8�≒�؏h�Z��`��Ԇ)�د?�������|z�S�9�����/��r���?�+F������G�8�ی���d�����U���M�Xa/вJ象�+�a���߽�^x�s��y� ǳ*Ux�F��Wte/~����\���ﲑmD�z�xַ��y��c�R��Z�oB8�D�!��hEp�q3����o���J�6�Li	���O�K/���쓊ʫ6hh ��iM�u$&dl2��E<h$a9X;�7�''p� ��/)��t6��֏4���@�U�>����TP*�D�Hs�$'>�ӄ�z*R�h�Re,��Zy���tLC�k��l����K�f���*�<[��eqN4Yڤ<����A4��f�Pu��j�Óӑ؎y����X(U�ʓE�Z`s̱Ԟ}L⧺�g�)$�	�� ���b3L-���,�/���,�D+w�d4���YG�`к��F���e��kW�"�-f��F�ɴ��l�(�mښU"d"s��k�  sQ��Uz\�"�Mߵn[��'�xJ�\�I�Io�	z�m-�[�W[���jK<�p�H#���f��Կ���Ci��C�mJOξ5�Pϊj�J`N�E�ތY�W�ƒ�5Ic�V�(s�����r�?K֙>je����^-�͓�\�s�t���1s�V�TDծ��y�tzVz��]M��%���k40:RP@�?�5blp2��Rh����
m�h�\���?�24��/X����>� ��'uĪ'�6ȭl7JL6,��hpG���W�u��ޒ��l�u�z����]�"t�=?`�:ą��zؠ��.���zN[��5�6U�T֠e��Y��s�b�hy+ٛ3��G�J&�&�)�-��w�q�&oM�Vx�Iɧ£��pOA%F!�=��⋵ՉJi,���~h�
�6W\2^�H���*�~��=���*Ϧ�>|#B�����*SbZ����	\:L]p �o��\%����o}�n;�.��,\�N��Vr0����ܻr�|�)���{|�)l��(��h�����d�ǹq��t4λ�uJ��g`|��Ǐ5K������86B��"8U H]�$J]���ȩ�TZ
�-IY�`�>����>����
�QV3r�1��ƋjPhdyb���۷o� 7ig�I��I[�\��3�5ܕtry�E�D8��U�ij�#����_*Ғ��M��SNjz�!V�2TA��Y�d_�E.\�����^-�jD�@� 	���������K��f�ee_�ќ�?����b"��D}	���q�4Grｵ^�V��*����Ln�]���m��A�߳�S��q������G:Y"����TW��6���1A�r�ÁR6w��5V[q��t.��0�3Q.��ٚ�R?¸+f��E��m���kT.,໒�έ>�`aI�<�ñ#?fBbԕ�G�Z^�|Y�e4����A�R����Kcs~�������+��X�+���iB�E�Ic��C"$V��i^���"3�=��'�E�j��:�7tH�k�rV�o�:�LT��K�[m�fIkzϺn�:k�ee��]@U�d2���ZiH�b�5�+��ةhX�H�AM_7����rdJ$3B�r$���F�#�бU�ڛi7N5�1�@�Bv'�b��r��:��M�v�Z�)��fqf�u㴐��f�/�I�m\�z�/�6�X��a�h�[֡�Ui�KI%����lZd�=.�)��1X�ړ�&�������/6�~��¾��b;�jº������%��@X��l����[��K�Zh�g���Þ�f{�$QI���"��4^!)���Ԡӿ�C��e&X��c�9b'Sd���Y���n���	l�,zkYj�����E�0Z��)�����+��{(^{�/h㛥�rM���w�@W�����,-?�Ep��)����I�C�^�g��s���ٷ���z:4�6^��'&�gl�
j(�g%um� �H*x�u�]� �F^nص܆��>̉�V�F����8�y��SqQ��6o+s�5�x��<���)�Ս�7�K�M�=�
� ��PFj&�ʕ+�,�(�,6?�6$F����	X�L�k�^�M\��ի�-�.wv���C��� �(Uy-��i=��B�<�`�%����ZcMVNRk�ܹrQK�������`\d��D�I�%������0���ᠰ��k���������	��_�H`�ֆǏ &��UN���B�N�8[|���p�[���3��#DNC���X�*��h�U�aK+컵�����G@��pk��R̷�R|�׾��7�|sc�����$�
�,mp��\��	��ǲX�y��{�]�q�W2^Q�7��Ҝ7�*����̰T¯�`�L�ei��j_h��f��MI!��+����(r�`��}��l�xj]� R*�����7o�g�ᠯW!0+pm�"���g쟍J)�`�%��χ{D�_������W�/p���ߦJ̻<�i3���;lnf����M{����[O=x��4	yE(�kmA�̍�HΆո���U������f5	L4����%p,y�h�[푂;	;�R�+?LM�lE#�e�c��ӟ3�P���m=K�"GR��d(ͮ�@����H}���U�@nV�M�[�f»R~/a��UxM�I�G��+R=Ȋ����$nM����Ð=J,E��/;��ҥ�~V8[2��ՎkF�b���]�I�sVt�����Cc,��P3K�&����QlN<>�D�(�D�j��lZ\���J��$�Na���$r��kD-@�<ϙ�O%S���CSAK@Jxp���гc�p��e[�~T�ƹح�(	���W�y	
j1���$�O6ͧ#V�Y�Mx���k�
U�Z�}�g.˞����}�ҧ�hcl�U�jjZ[���󼠤�-%Q6E$��ެفOe� _������=#0���� ��Kj0`�����,K��a�жG֗�h�qM�>�[J=wX�1�	����t��#dsw�Y�$������C�T��1�Q���Qe_�����M�e��?�[5_,���Pn�!�'�(�9��uF�w��rw�����t��>
,#N6��!�n7�6�2��e�=$��E�����OH�*����q/�c��!�|;�l�V�X2׀�Zj|��ݻ
sȦ�k�9�����gә�ɘ��;n,�4aqB�B ����	k�`��<y2��-�U���t�Z�*���H������KZL��&Vāg�2w
�^�+ D�	5={���ӧ�"]�=Pٵk/b��ܹ#�B+�1Kw�L�ٔ��2�$c�t�ZzZ����ʁ���2�p4�A���j�l�������s<��￿C4������?��?㻶��|	�	���+W?��4��4)SJ%éO5�k2�`�S�J�����PF����j��3�>��I{?��={���?�����D��^��j�u���U�g%7�m�C3.���b[I�>.����V�)La�Co�W�?x\H(v\�l��s)��ӕA �5�?3��B�FO��ѣ���g_������t�yn	��.\� ��+�����m�Ӱn ��AH��X��:�0���p���TkN���L��Ա0=�� �#�HǱi�~ ��y�1hs����ؐ���t��||�OH�0?�:m�hEb�*Ik�D�*A�s���*6j?�+y��=Վ@hU=��g�	�	эFs���ͤ&�3����sE���:vkl�[o�E�t6����n'�3�yJ16�ca��P�4�v<>Ղ�
م4p��3EJ[�JC��IC@;��o��T�l<��c[�.�4�"v�xF�v������k��U�$V�����ۯ����j�t��%����Ɋ< sI�H��3�S&�!c��ѩ��X�a��W��{�ټֲa���/�TO��w�B���Pw���M?�(L���o����l�op��1���O�^/������ᡑ.]������o���2VG��e�æ�ї���f���t��� �����.UeUd�ۨ��qrq�&4�+Zꤰt�|6f���_����l��rcI]�PW�O&B �����T�j�匤p���dZ�M8_.��$�Y���s	���o��C�)�Y;籙�l"�I�#��媱F�E���8��NM[2����w'U�.4ɳ��8��U����,�A��/��brʥ�6h��i�ե�(���rH��w;��p�9uyt����L�rc�U���fggkg�|��ʛ+O�BI"q�̶�!��^l��1�i�J��X
�E3㱟-�}M�j3+�̀���lH"��Ӷ���%�PYͧt�9��Ѵ=l=y,�%�L6���X�~��iV�Jo�q��A��l9�gK�;y;�E��ˈS��a:�T��ۇ1M�4�E�(�4����V��ʕ���� �����k׿��o���խ!�4Y�	 �I[�G������0]�Ν�vI��/X��������wT-���/���Ο��d�&�N��y�@����G���x�)'S�u�@yU3�I.�5�wR�A��xs0n�+DH�����cU+XF��=^w4_�w�����"o�
7�ٳ�ѕ4ʊ4�	��p�����m��]`}����������ګo�~������,Dy'#�<=�4e���t���x��y8[�m��o�����/_����ؒ!l<���v���.��x'��w�����=���}|:6{_{E�i'$�ʹ��P���rܭ� ��^w�f�޺�+q�����3k�Hy�����ؘY�]<���;�]^���?�@����d�N��a��d�ҥ�����J�cϷ��N�Ve3�P�V�US6�\N�'튱�6mX�h���4�k�kgӿE���+�0�ʴI��F��X�vj�� ���R�3���\`cZt5���?(ǇO��нF��)pt�/_��]W���d��*�1�>9=}x����G���`�1::��^- ���<s�N�e������ԫ��ݼ[s
U�������|
@3�� �	K!f�l��/_�>��9�e� �vskC�Q�>}�����_����?��(��,���b7͓d��2���Z�@-��!�El<��I�Z�q,��H+���X�"簔�"��[���M��ݢQ��P�t62I���P�y�Xkm�Y��/����!ړ3�5�%93Kk>K����j<�R����r!�K٦��˫��^�Ƌ%T,�*��Z�B�B6�\)|[?1��gG3�������j[s�U��<e>=�XC�g��ϕ�R�z��� .�mT��Z�+*4yaD��y��򢋣<��`�����t����Q�)���Md�k]I�����g�8o��Ⱥ쌝M��P$ �x���[ T�λ��[��Z�'��8�oł�����
h�]��~%N��4 ���}�l���jY���~���[�`>[�gnLM��V�Ų;�6�f��z9��a\�PA��H���u��&���T�ʸ����F�v?�G3MUn۱���а�1�Il)7���m`_Ֆ�1���	�׎p�����.ʅ<dRё/��}�U۬�4r .&�`�{n���UF�ܤ�Π`U&U��5�-x�T��u��z.ۄ�ŖDd��'Z,����u�J�v~D�7eX�oa[����/Q�h�����y�LZ7�]�8��QeW_��a-��֓��ߺ��*k'͏�N�[���ڸuJV�1��j�4�X�N�+��YF%D���ڨ����_����Jc����2T����}k>��`�s<c, πOg�e�8��,ˁ6��G�.�4�6���Њ��<�I��6���\9��i�J�c F�TԕF+�]��)��Y��)12Z0�z8�a�G�����Һz���Ƙ&�.�9a�D��#8�y�g��kc����g���w����ӧ����z} �����7�}%k��j��3>=0�Ʀ	%�)�'b �~���5�r�H�*���M��&h�8ɺ=�(���U5���5�������c��JC�6���C�|�+�!>�X���}��o��O�0}��Z��<.��rL>q�m7�j���ބ�M�T�w���<f^�S�^���E^��'�|2����R�����$:��S{.;�����J�2�Bnʆ�Z�g)|l�S�V����_3B%H�`�ϒ�p����X�=y���_?��� �����q�&Xf�p�&���^�Z�/����b��==�Nxt��o~����!n���}<��8>�dX5�Y
�����!\�Q��(����ɣ���ǿP�'����
����Ws8x�*�	�����X�J��ƙ�m�`�Y�O�� $5�֜g,A������.��)pO����d��~p8�}p�ܶ|:��p}�L��ϯ�2m8%-��$6X'��8�xR9S�c>����6����O����)���+�\�z=�����_�f%��<��h=�NC��t���U�鴖���߇G��ƍ/��".u��m��������D���� RR��Z=�cb
lc-�Y���w�� m�*��H۝N牧�[1�ř]ʯP	,ǌ�GD@�)@��S�<�Mg�^8�P����}��E{������W�_��6립�LY� ͓ɳ�O�ܹ���}eS�-t:�ōf�!���B�bK��i4��$�0HF����*��Y��!I�<|���C�&����4ɬ��lݦ�X͍�U9�0��M��������2��W��?��ܑ�n��aK��d�՗d���`��1L��'e�L�蘳+(�	�۸�*���w��7[�u��&�AhX�&r5@�J:��D)a�R@�4tDх��U>����7�/������V`!���FJ#"�ʪJ+%~p���3�����r5�.7�tP�׮]f�u��mY^0�^@�۔��ς$
�Y���?�a�q��~D���#�sL@"�e��i��/�ܸ��ZߒL�l�l����?�S�g٭[���1_)�0�R^+@n�6��3��o(.WŜ|��l&�"��_�A��(R�<��SY�������g��ƳŔ3�;"
�I\OF07�j��w�<y��v�� ��FוE�T0L_������3b}z]0�6��H��d�!Ը��|��Ci�k�C�BW�B�
cS[MVϞ=3ƙHR�ƞn�"_a�|��U���ݔ^e �M�3�����e����N� ����P��F"����ˑ�6|����Q�R	I�l����*\����YK��kes���R��ݿ�]��~�����/�0掛�I������I����^Ѹ���)�8�Kw����2��͍0�W��gp�2����o�Ԃ�^0����!mel�s��E˛��ѯ�T�m!�F��ڵk��1�����g�F{{�����{o����o�����n��Ӳ�[�� pt��k��^��m��B��^xAC��/�k(�VYl��)�ht���H0�g3F�r�b�6�%j��QP@��:���Z��L=A�
�T�b+�j�(�]l�_ۆ�?�y�����5��%}���˗7�V�[P�R��PGpЕr������u�*��YJ�j�VK����ʳ�j����)�Lm����J	<�狈a�Җ!i]�;!	'K�U�JZ���a�Z��~�vVX�cM�o`��c�&/���=�5t��Wf��&��b堞=�i)�*��8��Fj�%Tr��N.��M�o3G�E�g�Zj`�˄�O�9rP��d~Nh�i�pp2�x�����m1����&`T��b`�6#[%ߓ�Kt��[��*n�_��>z�h��eW��"�g�}�RSL�Y���Z=,�?ln�G_�rbk��^��"���A�p?@lì=�EJ㚗Z��#HK�n�����S�Ǌz��rD~�g�Jc��"n)�:|��jŐɍ~��yd[����@k�`j��^X^�k��nf0����L�n*���@+�9c�o<�j8�0�*
V<��ĎU�6f��c(d,�DY��5e�!�S��c�g27��TV�@*�d���',^P&�u6��W��&hq� ��V�[{�	$���C��76bS�&��W�"d)��l.J�֚a�v��K�y�p��������B��S�E~�r�s�R���h��m�b���GR?��cM aq�
��y㧶)��f�8"]&���ƁE�Y��!Ie��N4%	 �����U��O��6�]�0�J����h��C[�T�	Х�:��1i[?��(+�8�outV�0>�T!\��BT���x�D$nE^Q���B�;�yYx��֏ye����,�j�%�X���Ī7l��ʮ��aR��}2�F%Q����*��n�p����o�L�+��kІf�.Y�N'�1��?��&�C��ڜ4�%!��`�X��\�2�,s�.��߮1ܸ���m�{��OT�lj����=��/�@Wz`C��Ld�w_A�(����~���?�^Tٌ˽�=�'&P����d�����,pNK�`!G�[i	�VT�f�oo�I�R�~����_�����׿�����������7np�tdE��N�#�*m(��Yi���g@9Ü�(�BJbc�JW�%Ց�P��5���Y�eH+����j"RY�9uj1tZC}7�P+-���ĭn9-D��]��}���.^�O痿�e�����@���0�XC�Ӥ�Ç%���B�4�[ �џYeeb��������n{��a�C�d]���5);�6��_ᮌ��_TdT�L~��ѡ�'rNb\�7�����p�r9g�ט򰛟~��d2��CO�s���x{���e��>��]�6"):U��1�L�32��3�jPDf<Nj�����(j�P���V�@_ԶNi������UYǰdG��R-��1d��sZ��56i]�)�A&s�T��ϗS7K/�N�S�F5����7�@2@D�~��o*�����`��_N�S����}�D��a�W;>>�:bGu���hs�+�Dՠ�{#lĹi���.A~uu����>��sJ{?pH������h�R +�7�Fu��]�;8��|��1�leZ�����q�1 ��5��ِ�b<'n
#b�YW��ȡ˙��\�=�����91���ɲtT��OZ�=��*xs��w4;R��jg֓�̇�a9Y6~�p8�yY�7D�q�G���r��ɮo�p�Ղ����yt���w���S�BE���i�=��g�1,�������Ϟ�NY^��<�q}c�]��� b��>v������s�<�ݗ7y���h�[�L�ő�m�k����!.���p�n߾=Ϭ��QZ��k�ǿ�~�o��}�#��Ʃ��^+�N#jWm^��b߾#wL����^Ri-P���
EE'��.`��C�^>�`WK�j��5��T�|?hf�������?���~����p�#����k�k'������ño/]��њ&6�J����#"�Z�7>_L��63�`0�_Z�u�	.wx�.@������;z�?��	7�3 7O�<�"�����*��B{A��>I:�$���~h}8Oq��T����
��v\#+�k-iv��HE�斷�\��
���	�������Tt��f�"z���&�:%�T蝼�=��4����J@`�A�_��<�AS9�o߄���޻x{:�}��'o�������_~����j�u���������v�����z�ݦ�R<Ņ���2��˒AU��l|��o~�ӟ�ތNN�z9�(wLC�����+F�\t;\�~o��u�Q3��;_�-�k��[i���I��'��T4>�B�n��s���F�W�-/�pco��0h�<EW��^с5=>9�s��U�k�j��� vך�FW���Qߺ��狩�>������̋����������}`����m~Wg�zְ�������T�mQl�>��>,�`�a�R]�9�k����֪�!W8�D"V���R��Bf������n���������i��A���D�O�ё�:�=x����<�?�? �*�ʒ�S4�usN&�;H}'Ze����96>��j�e۲����n�L�=n[�����}�ɧ��/�����ă�&k42��MEZ�s-0w����?y���?��Y�(H �Z,���2[V� a\LE-�<ikOAU.m����߿��5�ќO�B"�����LX�š26�h<߿����G�ф�&,Ov���aڥ��$ù����xl�Z��0�>&)�F��VVe���G�?�D������b/l� 0�p0Xm��??��[l�N>�ÿ�����޴��X����%�1�ܘ���=��M�vq���|DN,ͺe!
�O����ݞ�h������t���cE�C"�e�q�6V>��2�ǒ;��p�-c
Wt�;Hn(
���x
㶻��U4�����6�&I�y����JQf���y. 'r�^ew�)��
=B"�����|�[}6_ޙ9�9��x}��5�Xv
g��
ym�㙌�<6BC�vMe�p<s�Foa6a�Ժb��ρ�3%����_<~�8�Y�����?�tpZ����4^tuR�[ms����Mu�ܖ۔���e���:����-]��1.Y|���U� ��C�5�wB�c���Г�O�v5Y���N�z�bE�{E��;��Iפ��x�2K�;����U<ֵ����j�L��ȣ��$HcV��l`N�6�0���ƿ�QS�(k*-�
^�]�K�3���u�urrZ�r?�a�j����~J���o�,��ZʐPȒ`)�5��ր:�"d��!�OOD�ホ�B�3+ʶ��r#����OQ�z�6�מ��^5-���Zٔm���2�Z����4�q���$]���F��3ے��*n�ՙ�g�4ق�p�TU���K, h���P�/������b�w��?�����������t��6%�y����a��;IT������T���O���-���]��VĢ�-JRL&�S.O��jEIii�`#�6.W�ɹ��S��!`uH�"Y(��=�k�k�/��:&�wf��d�lX�7�rXSY���ې�CN����/��7��M��ӧO��������?G�b�H���:d��w:[�0���0�j��{�B�[�$�-P>]D��u�`6�g��&g�����|�^�>VF�Wt~6�#2�(�n6!�VC8;;YI�gʦ��.?����D�j#��`����k�]�vN49��ܹsG?�=gk��ڔ��Tr`M�P>���D�~��5V�`m����~V�C����r��]��Y\�tɳ��D�*OE֩�ɍ�4���3�D�6(�ڷ���u��G��Q?��Q�W�\�u�v�5w?<Z
r�֭o~�[;���-�g$�(�+c+V�V6�vEߥ�Uc�9c�ۥ��9]�o��5_�6���B�*[qs`Y�����+�5�Z���ư�0g}+w�q��s�r�ЫJ�����^�|B������}.����Kq~rB�+Wvq�OO�?���ؠ�b�����3����Q(|o�#Ry��%8Wu�z*�ȴ�6a?c����y?1*�+W����GS���W�%���J0�B��g�vaǁ���
�@2���my�U�7)��:�:�=�h:��+q渚x�b͒l�s����YlC����U�9��7mKKX4<O���ƕڱ�@�4J��A^I
OF>w�y�U�G��qxc_<᳤��!�/uR8;����<i�%>A��09��:��T|V���w{�Es��!6a$��S����1܈��;.�Q�Ϟ=ݳ���")A�zJ4�#w<�n�y���_��O(��s���h�ٰ�����l�LJ-�3;¢���3��zic���sc���0k��Ǫ�Jì@��4V�e��y5�t�ׂM�{��ϗ3��"�!ց8:��_�����Tƶ���"t�w�1Mf��2��H��W�h�c�����~~H�~Q�\L0�g���"�C��*P%ʽW��MoBم�/��uʕh-��3^�Z���d�#���a���j2��?=�5R�O���>���)-�*��*`m�tT�g��H�O-W�gDh5_'�7	��l볜v0Zj~)KW�ę��t�V�+�խ:�z��U��+M�۷oC9����ݛ�'L���}��2��ͮ�w�\Σ/���6����(���f� ͧ����g�}&|��X8H��L�
	%�Xԛd���Ͽr\*>��A?��)�%ш��ǖv^o��ϸ|R��zX����J�|�Ҩj�C�9:=��ܽ{:"r�J�%>�u���b���ez-���h��3�CI#�UzJxdt(�%�b�SR�0�S�ɡ��3P�jM,����������\=~������	�{3��pNT������"v�X��p�%B�ʈ�R�7J,���O�Q����u�+|f'�	%��f��Sbu�k��ᔷ/��݇�Z꒜��A��dN=)q�F&�RM��.��׿>9>������H��F�6�md�_WmP:�E�cU=��XF�VF)S�.�B0��`��=�hN!�D`M�ht����q��>���,��굾F���Y�NP-�
^с��\����~^v�Ʋ�}�3۰g�3]��E1�_U����eb&�SG�J�ַ����2�up���;Jc2?�'���
����- JO�W�>�F!29)])PjŇ�gʏ�I}��z:u�/!�h|1;|]��b�Ʒm����A�+�G�
$v2���a�,�@�T�������[o��#��U���
`�A��e� ���:��C���<x?m�M^d怔!תܡV���g��#[���B���c��|D�z0��O_#>6ߦi�XUJ�&R�(&�7n��:@$�-���\ � ;Xִ}3�6QHZ1 q�@Lͣk���|I�wV�u��"L��9��8y���fp�E~�b8&#���ČX��̏z7i�kH{G�R��;Avix�h��w���?��?��8=�ԟ����!V��\�X�/W&�&�l��;E��R�W2�r%���jj�p�vS)4*�l�n��b���1E�R�S,N��~h*�lO�f2F�_��9TW���آΩ�l,l��R����]v ��t�_q{Xܼ��E�������2�"מ�)Z�\���8���G�Z��F�Af�8,���晕��Ċ�n�Ue�I�����5�������JYavz�N�>[%��#����_��7��ʫ�
�B��_��͛�@<~������������N�"�=�\���M����{�G���J���Ϗ}�t�E�Ίj�AX[%n�l��[��-Nf{�����l���ƕG�&qݴ��1s9Hu���E{�R�^�r��;���uNҥ����+������A^��\#J�����ʲH)��)�	 @eb�1���g��x�;Z׍6ĮޤU!����Q��Vׯc�(��4VM���T�=�[|�y~^�^�����k_�ڟ�ٟ��<��Ծ ��|n/��H"�z�|�L9#�,^�vx#RJ��g~��i]�TJ�Jy���ስj���6N��^�'?��C<QkY@M����7�B�J���
����EU��,Zi��x )�/������:�R��~��_�Rǩ��q'P4�5�/�*�_rx���s���|ߚ&w����»�n�TdS�TR}��y=W�	�+�C�I�Z_<�F�a��\)��1��NX�P���q��:�� �d㷿�-,�j���?���+`�_{�5��Q�j7rm�g�F�4�k0��Q6N�e�L�D<@ԯ��b�I�:�p�U���sX4Q���[������9v��F�D��Y�oQ��jEFZ;�Ы�<fT�\y_��!�\О��ʹ���[ 
���䃃��f2�)[�:���s�������i� ��c�
�.
,����D��X{�'ׇ@A��E�ʋ	���ܫĚY�l�`�r��{���_����z���m���N^K�)خMO]��_������3�j*����T�K�ֹOp��x�&`
�eg��O�T$,�S1e��n�:,���үd�������h/�m��PP(+���
����FuR�nT�c&ȬYjZ��:K!T�ue}9�ڱ���b8��k_U����}u��hq$,lsklҩ��ٜ�$����.��Qja8���6qQb(�.b]��a��̅Q�U�g�;[wqz!�бCQI��m�)U�B�.�.���֭[rJ�R�� h�f��T��kz��jC�C~�`���_8	^b�؜��?4��,�i���R�"�+��#{��8%mԭ�k�3�ʥ�m+>�3Dr������Z]��G(l�m'��
�E�ᲔJ�ݻw����*� �$�IF���op-,7�+��O���o߆9����6��:>8���&ǧG��n��0�~a�s�d���F��������~�����לһ�>�vwH��h�{1�{�!<���_%�R�gK�NO�0h��B�D�)�% -���2,�! #�T�Tҝ;�?~z��÷�~[;��2�*��j�w;9>�0(�MG6削�#�t�W�x<�wﮚ�`��m_Ul����ӖQ��2�Շ���� C����Ƙ�bߐ.��iӦ��tJ^�:9�Z���fX��df��)6]udO?�0S�K'b�h��d��dŤI(NN�ݹ���\��U�S��x6?�
*Ɵ�*m���\ف�ޟM&x���4i���A�D�?�+pw*5��w��x�ݧ|9�X2�mUC�EI*��N�ː��b6������.]��pvv���kɢ�z��ڜ����;��޾����g?�	�z�`l?��׿^�%�g���NNLOV!(�xDո;���>{"��ӓ�� �W��ի����|����ڲ"G'V�ѣG��!������Q��p��;T~Pf�g��HZ�m#u�~(Ȉ��1����pr��ʬ��ڏ�nL����V���S6,�VV$�]�Z�$�B�|��x����wຼp��p�_h��
�9a� Z�Q9�an�UF��z�yz�"gq�[������^O]�l��]ݔ!�k_���O�Z��傽[.�$tP�@�p80V�%�77���Y7G���Nk$������pT�loܸ�w��_�("�K������N�����ʤ	�v4���yny�Xx�EQ��|��0�$Dכ�hE�FCy�+ٰ,wc�����DT����-�VL�6F�u;yk%???"�&�-���b/�7_~��w޺y���'� N�W������:��<�q�ϵ��Hv#�����U1G��7+5"uٗ�e)��3j_s�AS��.b&�9B�
c�B���buS���,gA�'�ư+�>�l?�9��>����&�a�Z���l��η�y��_|�g �0���&��$�0u��OOI���%����+M>�Nl$�a'�1��v��3RBP�F�3���S�$0�� n;�+m�V61��-Zѫs��\�Mɖ�s���MY���"4<7�����T߄E{��/]�$Z7�\�y5.��s;� /^0�[��n�^�2wB>���:m�/ C;�gs�~��k#����'琫����LeSy'����akHB�.Kl`qƝ�0�o>�j:�F�N��s���f�����\߅1�ڬ�&�ͧGǇ��k;�[�.��U��^������_���_�ܽ{���M�3m:�t��-��0�Z��g���&����;��d:/��/B�ܬ����m��n�P�3f��L�];��㣩�	%�&_Q'���1�감GGpBɹĵ���0����y�^�~�����o�:ۻ�?��������鳻��*[4v���v�U/�d2�6N&m�;�Wn���)"�H#�V���Ս���d)�3|���'μ���'>v@r[���H���&�dO6���
��c�7id��5��4
��fKeY��]�%��|~x���?��?��'?���c/�TY�����le�;����ͨ������vc��e����TBh����.��~{�w��MFs��L�"��g.5tH�R@0(4>i���$�����1p���v�n�|�{��^��4�z?������PyF4q���B���9�a�DKRy�
���T��s���l�>&DK�cj���Q�s����+D5ٴJ��s":5p�t xY\�9`,�l+��D��6�c�1�]!Mer�BJ�S[����3dT�b�_����o�!�@�#r��������={}��'uU�,_Ȧ�$n�j0���7�DXUS��xc��'��K���8M�g��B��"8 r�&�23F��?������J�K��E�l�P)��Tl]�L�а�$�3�g%�FjY�D �$б�nn��V��!Y+K��w����Y�	*�Of&�S��!�D��Ccd�Z{&t�B�hȯwF����p���2M���Я����;�(��Ӫ�b,������CL�o(ftb�Ret��8��M�@�t��zmM/�	=ǅ�۳�N��`��lCģ]+�
o�`Yd�Þy.��ߏ�dݴ��������Z^܀S��nl��m�ېE���^�ì���[p%�#��o�B
��cCb�"�Dg�}�æ�ʉ�Ί��XNk)v�o6��TV��2_6Qǚ:��������\�驍����q�:���8B@4Y�i�0]�p����r�dEf�*
��M�P�ʸ�i0ȅQ�R�ВM{V9�1�C�j�Yo����Q]7o0r�Y!����S�Z�7A,|D�+v(�;�tʍkY������`PX�s�\M�qP���:zkֺ�B�.Y�������|�%诬K�G�h_��8l���`�{�\Nb9+,?+	7�A���O]ME^y���{��5��u%����!S��Ė��<y� ʄ/j�Uvq����+�	k�*"�{��������M�]��쥡���JH��J�3�9��O?d��+a�1�1��,��p��¡r6T�h�U������}��S*iL���
XJF���т�q��m9K�W�^5�$��t�����#c1��>��ڌ�tdq�#q���6�!�r�pٝ��+W�0F�!L�0�j�ml6t����ě��"_�uH�y!��h	�H�F�;V�� ���
���}l��o��o��#�J|iv]�p����&�a=Ipt�w$�p�`��~�KEV�����=?��P�C��>yI�L�n�@с��bU��l!J���굧�)�����o��x��%x�2�s5����8_�ΟkCox�_��W/ݼ�G�q���dq")������c���޲����p�+�X�q�v��
�Fީv�=q�.���7�ݠtA�?���
^j���U�I2)����4:��kۄ��h��ܹ�c�s4��Q�M�j��c�s�lv���g�W����
��4R����|�Z
�%�g�X�l�gU
�,���UF'iP��6,���?���ެW��:<s�7�N9�ER�K�T�%�p��`���~�S�?���7�Wt�Ï�n5�hr�.ð��EqJ�ɜ3�|c<c����7H�v�CD*3n�������5Q�7o�d��P�|�F�-���ɂS�R��.�"�/�%�Ru����� ����T��2�k!T�Ě�|+�j��h�-
�a�^��6�����Y��E�1��aŰ��ַ��O�����G �(Z�������OvT*��Ñ6�1U]�i�mjm�x>�S.�U#�rI/��E?0Wz^r�V2��`ɠ]�= �`!�5dG��QP�؞�e�x���.a=�p�|�������W��8�5��꬏C"�.;p\U�c��XpT��l�h"�:�3/�͢H��S�y�#Y���ɠ��r��XB۴Z~^��c_gS��v7�چ�J���j�.A/DX�q�Zm!%�X�����^S�����Y ��wE`=��#cTՄ'���zcvm�vB����U��=�z⧐�t�č�3�)�|*[��|'[,r[d���iG6J�b�SȐy6:Ӂ}m�B�s�~�������%�}l:4���:���Oj1���1�&�F�T�o��ao��w���B�9��.�s�i��J���'�������B���9�.>��m�6���(j�`v?t��t*�k�N2�x��G~O�a��H��Uf�#�������F����[����n�q�b+�~iX�X��c]��D�#�2�=� �*�c@x*�����������+(�9���^�)���Ռz��^s֐b��ᓿ�k��c"l�΂�SI�2����:L9V����FA�B��e�Oun���a_�%��y�-�*�_�|s�f@G��O O�NH@�ס�GP��;^*%#���b�֘5LY��܀��������7�	�M��z�m���5��=_P��Λі+��i�|�}�SS���<�����ٌ�\N͠OmD�������um���]���������)쎜�
}R>gn�M�m�p����k�ٴ1:~�1��_���fb�k�`\�M�e:qh 6?</�)�kS\(�l�N��j��5by��
l���%Ƀ'�taKN,�f^X�OaU�ZQ����E����?#ߴ�(�n�:Ц�(�$�%|*<#.�S��_�~����_��_�w�hdH�BR���wT��(�.6t���0�V��!��OdP�r��FF���
zϞ�������G��{�.އ��L�'xptKخy"b���mƀY�d�r�����~����p'�����vm_J9r�(`��xk�+�B	�A�R}��߿���Ѣk�=d5�llY�W���O����m�gk�lߚ�`V�	�.#��U�M� �y*CJ�3)���\vGE�q������g۴��0�E&$���O�/��>�
W�F�� A<�����qk�m�g�(ܺu�F6�>ͷ�t��~�����{Pџ���W����W�\��G��ğ��e�"�
y����.׎o�Y��o��k�44dF��,%=l��ݕaG�J�$E��e�ɱ2H����k<&g�w�4�9������M���N��a�[B�
\��l����I���TM�	9b��6I����d�X�
Z�v&����v�����B��H:  ��IDATo��g�I?J6@raI/j�\����u쓡1I�93�i58�6�@8�!-���`���� ����n����<�16߸q�ѣ��y�Η1�	b��!I?Z�W�a�D��	Q&�?Z�_� ��7�ɪ\���ϧ�`���������eUP�n�hJǸW�֘
ϸ܁})���3&�n\#�C�\>|���=~�@�W�͉���!�>�����ޫV˽��j�X�X��/��ƾ���۸���� O����	�,mb����#��k8�n\����l��u�<::].֫e� ���kh���h�4����wk�s�w����p�m�TꂺZ/xI�����KaJ�q����!�p���c���8u}��g's�:5�P]����Ϟ@��_!����m�iM���C�uO�<}�����Y�Dpv6}m��{ܔ����t�9���J�H%�{�~0nu_��<f	Q���_�������X#k�5b�����/�?�2��c�37ud:!�ɺ\�J2D�p���򉐓A��6���0gZ;N,Q�%q��!�"?}���S��������Bs�M�z���Ϟ��̲�O�?�bV�i�z�U����q�i�����z~{�`YW���K��|��Ggg��Q Z��
N�NN�B����"��v��~to�^���G#B?�8;;�n��g�g'gg�K-��"��0mv��ݽ�/�˿��/߷��ω����;(d��!bu���]��8a]����޻xp��/�������[BJ�ul�J�qM㹍�����G�*l�oS�bWb!Ad�a���s1�	��umY��h��ռ��
�6b��_���𕄚&��9N�Z��E��Eo�9^�����^BEn���gW�e��X��:�̲�4g��o�mJ?N'���)C� ��Ԫ��� ���յأq7�WuLz��F�^n3mq��^=4AJ�̿X3�m:�E3�y��_�������ޮ���x�ʱ��.�f(ݼ|&j��:<z@���<�rk`d~�Ѩ��5�]p�vd)�˪(�x��'���\���*t�\O�@�ڂ:�#L7��X􄆃t�~�)p�8ػ�h�rlS�I��.9k��s���ʕK����훯��ſ����]��[V�]}��̪��I��F��qd,ʱH豙�t�s� ��������\��첥&]v@���u�&ʞ�d�@�5��w��z�ĺ�J�����aj�V�����`�����Y/8�<��O̹�G�Q������s�V���_����
�w�������0*�*��v
c�[�N���nP�rmHᲉ�^_�.S�2e{������9̑���e
�uL$3M�F�^
�����mCEm�5�d<0v�&�g�b<K�s������۷�����Vf�����O>~���c��x�8����~ SL�T�+�DZa[mY�?��#�lҁ�h����+��p�t԰_�RM5�{ؚ���� �p���Z�c�v+({xvr�L(6��zFL&_Q'�3v��|�NC�oe�^��bFT�rn�=��ˑ%m���~���'�'x��)h�f�ӭ1n	�ztLb��p41ؾ�N+p���Ւ��f��b�Ml�d�o4��|n-!�Wo����z1?QzQs��O�J�HY{l;q0�����]����D=5'�G�/ƣ!�.�ڤ͢*&L���ظ�J%FѰ*�ʬJS[9�@E4���D�1>�(m:OzeG�����4�9�^D�I��ji*5u��\�[@|��������%�O���jM��T�p<���f-W�\���B )��2�b�x���/~��u�"���t���Ů>���b���"�_�!ʿ�����e�=�)�Nc8��P�h�W[-'d��I%ꀙPd�#����3|�
->���-�T�99��h'���h31���ޥK�x.ghZ�	��6c&�C(ס��U���=�nٍ�||z�˫�A���VF��V`���S�?=[`�\�"'V�)�=#KM�4�z�y��ۙ��:� �����h����D��L�6$[��X]k��!��0�/�pr��uU�"��l��g"�����_�V�����c��|��ӣ�z�A�������i��y��4���>��xa~]�h
�
���j</�qo\.K�;�f̹xv����M�^�ǂ��W9W�?���˗��x	�;U!P:F>j����vQ/�H�����!3�Q㆞1y� ��/����Mr��8�p��P� 6��(�o�e��)�5p�������}��l�?��?޿�1l�-~���ëW�V.x��/����ޑ>ԕ�M����#�?=�K�(py�?�:�P~�I�&�oT�N�7��:W�> _k�t���r1���عO�go#�l����f��	 
'!�/��B��G��ˎ�4<�J�Js�����Y�8����	�P�).&��q��@��u��v���W���m�:a�\F(�y��.W	�e�X�Z�Vơ���MWG��@/�Z�RjM�s<˝�#�iҙV�����ހ��Ae�'#g� M���+��F�����C஋oBl�sxz����aQH��I�$$�
GG����u�{�Fj��2'؆�s��)�ƴp�l��2`�
W��$�� �mU����<�d���s�����.��UdN�]I�~EŊ����-�)N(��"+G��j7��B�&HU��_!1�KbJ�tp�]݆}X<8mx��3;$=Z��`�Ԙ���?d�f����smG�X��P���Np�p�o�æ��bvv&	1��&��q�^ę�SW�I��zv����Q���K�z�]rH�t���쑴�t�>�;@�>���S�f��8���y���9�����HUn�c)Pf �T4(Z�m��n�(h7,@%�U�%�Wug��p�0�'�c|;�E<��=zTy�J|7�۶9�����C����Y�J-5ψ�ѓ�%�m���;|�R�X�_���+��26�_�.D�״Y*�F��0ܳ�5(Y�(1F���9ҹp�.��*9�+'��'$��|���5�k�D@�Nl��&Zf��(�}�7_p�m^B��5�N�����QgBA2��]K��JCȼ)�m0�hjmM��:�Xh�������)�¯<~���Ç����~E��E��}9�giU��,��������ݻj��f7�E���>!��̛?{O:�Ӎ����G��e�Cnぅ�:����^pZ�hQ�����?��?��A��j!����3�	ߊp�x��I�-d4��,Q��$�4w�S#Ô��ږ~�3��|��g�Q`���>U&q����2G!M�#)�XN�dFg/�9(:G��l���Q��h�����65�T����؋�P`��7.�+�������Z?�Ր!(2����+����P�%���K��W�0�u*��M7�b�UP�ߣ&%3�G�f�<������h�h��cnݺE�2+^������*��B���HNE/էK�R����>�+v6��9˵w��*bW<�G>|3� � ��d۾��B���O)�j$j֜�cj<#<Gf�E�ںi0�P���W��p�L �״�Q5�y�����)3ٰ�k���H�9_,����"˝���#0^(
%,��lY�~�L����As됢�6�~CMF�I��:���[�S�c�ZwqS�C]|�;߹y󦍄l�ܼ���~W����;�����ÞЩBY��Ԩ��5o�"9`�$ML�:bMV�S^^�	Ri���!�s��Ǿ���<4������N��n)�.z����xH�YO�s90������ ��Y�Z��2a��o}���/�x�W�3��V�P�We{X����5m���N̆���ꄽ(���N�m��lh8G���d,���޻�/Ǘ^z�����G�n��B*}��u~������,Jn[öCm
)�
�'T���O�\ƾ��j4�)�;V^C�F��V�g��I>��+P���[,&�����e��7�ag�&�3\_Ľ�ǀ���ȴ$�֊���Է����c$�c	�J�p���Sb�k���iN�Ŋ�	�Ub$����Q���P��*K���9��"�<�/��?.����sh �n��E���2aq"���Z>]q�oLX���H���p|`��p�R�����A�+�~�cFħ<�6s�G�����.�X
u�`%�ܹC�:���%x�)N<��p���'�޽{���N\���"��g�TH���a�g;UX*U�U'C�u涋���K]#�vl�[���(��1_ 2�`�B,~ׇ���*bu8~]c��8��8���߷��4�z��p�dc�Tl2-��&��p���GOx�SG;(�
�W-�:�*�i�~���/kD����+8�.�#�4~7	�cS�eR���hV��c?P��䲡�JF.�o׆*u�n�Đ\�������P�~j�ܥ͜��(̬*�����/���&s\��(����O��֣)�t��W��)�Se.�CH�V$6&Φ���iEr����}��_�f}�K_�i��R�������e�����ݛXG�ns �cU�����ț�$��6�ӑh��M�;�_s�H��+E���[�X,ae^}�K���[o��C���'�)K�=j�ؼ�P;��/5��=��W�J�'���S��>eE��������:�!�Q�LKN�2,�Hn�V;K)��L��0��:��B-'d���󙜋4��+H]��	Rc2��neȴ �?hX�۷ooM8�Jk��Z��Δ�àGc�@�L�����}Z�W�:�j�C�5\H������Z�~^��;"ZY��8#)r��Ŏ�"���ΘS�i�E��쥰�]f�0`�b�&�,N����Q���!1j��t{g�{~fe�Lc-Qk�<	1��eX�!	��Q�����.F�SZ����(M��3�_�I=Y!��[�/�=�_�AB���FV01qj7R�n��>l��)H�N<hpl�&������ǡؖQZ�!�
$O�q:��Ý~�m$%7�%&k�M,�l���U����۬w�
�;;�Ĝ��p�0H��K�	��g���	��:QF\P[��Ш��[�?B
���$r�����ܟ�5"Q�V�Bf����K�[?�����{�ڳC����逳/��}��a��[���4��b2,��C��*8�If�އϗ���Ir��󓣣���`n^�tywjh��`4�=���u������q#1�D�Fs|�r]>~����щ�o��Gݞ���1�^���k㫝洞s@�9<���;;=~��7����34����jmj�e��ZhbɎ���p��i���xK��zY���G�C�=:'����������;=8��l[E����,�zU�,<|ȼ��'O��ٲNy��£m,�"48�"��l��AOO���㣣	V {m��f�ņ����.A�D������GYf��r<�䪃z����,j�/��y���>~���ԓ���q��q�(��8YDu{)}���{��1�ը�n$�;��r����/PR
�)L��������+A�0��h�G�.m�פlDݲ*��qhr���}zpp��I���1��Idjun��p\{=6>i�fO�ԼH��'�Ӭ��Y-J� >�����|�+d��c��"ū���p��Q�&&��\T�r>[*JTC���/dk�:ܸ[�-�V���t�J�H��&/Y�y;R�R�S!Y�
mc��#�Ң)""iնH��o4y�� ���(��<[#��G�S�Wf� �����?�������!�*{{�p��X���D�:�[�'�S�<��Q���u-�AëT2������=G�W�dt�5f�Ȱ ��{�_!���n��(����L![�\�]Xi�a"dƭE$�?��kH����?{��ݻ;{{�A��_��!�C��U�K�c�*����Xy��j��8;�KF6��5��z�r�ux��ò���n���@]qE�ёV�q!.�dlc苞��V�1�[b�bK�M&C��8��c�p��u�B 7Jm���C\ �������"��Y�ങ/��o��̍<��H�2m�j��a/���n0�E�8=�u�.!7�w���e��.l���Q�����)�Y4.��(O��;j���`�ڲ�I�1)'�{����n��$�1�7��M��bc��͢�}?{6m���ށ�_���ֱ�\����=�y�:B��j�9^#�L��mb�,�Gׯ3�՘��ِ��|�`4ގx�;?k��0P����~$��]�G3=���$5��� '��q�V��c5������<�e�4Ê(�^<��l�(�8>UM�?o]޿Ļ]������Yb�|��B��H��Ӈ�R۠=��+ε\���_ɋ����"u��6�Ҍ&�����;_`e��	D��5�Z��ռ?(��4.�:aͥ+4_fȖ���W_7;ػs�����dg��L�6Uzن�����pr8������+W�!����
�xzrp|����O��ƣ��)�5�I��!0X�c~���ۄ˥�0�W<|���>��}�w^N�~���4T]�6�ټV�y��c��"���i������ф[]�$wdl�
��5kb-�4ì�J�()E'���=Mɤ���3�ȓ�A�����b�������s�����8�>�(�`�G�3�g
4ں���Aԭ���&wnߪ�5k��(�Ek�)w��m"���8_o�n�iv �knu�T7�����,F��˲K�?��zRu�B'�.�����V%OX��z����>�xB"6�|����R�����^�gՑ�o�^��|�D�}���������fSX�Q�FbQ�f#�iU��}��@���|N7h�QO�r&9@&�*&�) �a��X�Lxb�J��X��°������Ze9�nuI�-���_\�"�-W�Q��?�V��Y� -��)���n�{�R�狺�g�(�`hH��O�nѸ�Ʒ��P��%�foǅ�b���Ms��)��?1�M��n����U�vq��Q��(����'�g�e�_�D�C*g�d���d_�f��a��
�/~|ogo>����.�ZϞ=9_��G|�;�����o[j!�"=%��6�G|lMc�|��Y����0�aod ;�mkNu>��;7m�9V��"h�������dI��OF�R>���w����bW�^�??�螅���0��a�a2NO���*&2�!H#�h��8^������g���^bV�}�����}��l�~WVQ8yɀI���l�Y���QT.����z�!XU�9y;OQ�Ϸ�/�7^R <��U�S`�$����!��6�Dlo��+�t�4V�4kk���fR-��N|mC�})����-,�Xwy��8|�NF6�L[79JtE��N�M�}�'�.f�6���?���Jh��ҼՌ#��>I{�uyz|r��`�\)���s`�����	��2ݞ@۔M)F��Ӓ
�2jZ:�(���� E]V����/ۢ��2F��M;�<���3�e�/��=�ēď:şP"ϟ�h��%�8��Be�ȧ�$�te�Tָ���{O�_dh��ڪ�q��i��G�j�i���m��$��*�_���'�^z"a��3@_�YcL�%�Z4���t&�$e�(Q�\¤�e�r]�!���4��{7ß&��9�<���^$@+�!�D���>5;8���J�u�'w����֐��Gv�^�:�V#����yd�DH"�j��64we1�/��#b*�����2$���/z���X��-+�ï�n~� v���4Fj�a�7��:K<���H��)�ޠ�=�@�9�/�=}�T�!{\�.����b�X����������.�Y�G1#����������MZ���q�H��1���X������H�aA��B=z�IuiPP�! �N�ϒ�^[]<��kOK�2�&�J��*�-e�����j"�xo���|�ͭ���D��P�/(x�2�й �H�ىS��.�_��H��hn��yS���+�0������!tRçlh��0�?�l^_�˥0�vל^0]�v�d��Zi��3� `�pJ$�i��&����n����t3^;E	�.���v��� ��^D��VT
6�ڼ۵��u2. ��tJ ��pB�{C�D٫��a��E� wr��U����x`���o��)�^���,a�r?�]�Y���Vۇ�5��4�X�Q2�D/�B����R�g퓑�`�ʿ��ם4a��ew���6$���.T����;OBeI��+q֘-{������$k�,~$ C/驖�x2���\�H��.؏�999���[ �D�Z����s�E�����s8�ʫ6�@�tZ�K��b�Be|/[�a�Z��\�����nd��.�z�'G�T��(��0�
�K�(�+aPĥ{�}z�~��y�F�(c��#|48�:T��m�K7\��;i���fR���U�g��)�����M�MQ���f@Yj!��I1�nI�B*~��_�v���D�����qp��jnlg{O7L�o5H@#��H�S�T${Y��UE���{N��Isu$��W	��;Z�v��� ���Fdi(F�����S�X7�lPTQ����8=��v�/1�d���C���t[��|��1�c)^}�ջw����ElBT��m0$�D��~ppy~��S�.�Cj7����"z(�*�S?ҁ�G�i�K�K�VZ�H��S1�e7YA�}���Y��)D��/��j�n���ݠ ?�&�G�����[oivDm���>��c٪f��i�(�6)ä��S��!�Q	"q���ζ̥�]!<Sep�T�50�qW��c��ԁ� pb�yW�!N�7�zPnV���~Dk���5�����s�f�����>����ClK��u��|������%\w�v�ڵ+����!.��K/_�y�%��A�C*a�V8n8��n���:&W6�h8sr�qba�N��$���R̘^-�^�W�,L������)������{��O�;��M5�IN�S�.|��?��� �pF�@���q�j����}��9��'�B�U�7�?5��I��<C�9GnӘ�E�!�\���OZ��H%�Tc�WY3n@F�:l����V��L�"�esx�X:�_�4�g���Ώ��6��	ɋ�aN�Dgk��vD>��>�x4}�'�5~�<��Ϥ��dA5i�����S,gX~�|�N&9���\%��ҍ�"F%E���K�1����#����Ӛ��R$�;4��q�m�1��lʧP������_n���y9fA���ܻ����>'�;�К��B%;$A�vu%w��j��^�z�u���QW� y~�w�?g�|jqA@:c���t���>���|-���O+�P�.��q��MaVuy�ZB�޼yS��x�2G���q|�}�݃ǎ!��A^�C٘��ơ�!Iˆ��ͳ8�/.cY���{�eV'��!��5�f�2X�;wna��z؜�V|?��a��z��ׯ�e�:?1��w�Ø��b��'_���u]�|��Xt��[���%�D��3�ƕY(e�6C4$ۡ�P^P J�a�Q��EJ�y�r����#�c��V��֞4Җ%@T{9S�8�P�Yy��6С�⋔�˷�[�<er7�k��z��Y�uf��0�]����'�|�q�l~W�;�?�
��_��<߂ֹ4�}�t䇲*G��}���Vk��*�kX�AU��S��jMt�&��w��]����¦�an�@Fʃ��Hc���g5�s�8_d�ŉ3���Ɩ����p_g�g�6��Og�Ykg_�=�瀏;�O����q��W�LmL3��ҀQ�W+?��f�L��Ε�L��B�:㖴��n d�O猍��)�x09mX ���L��7 �.��Ll@�Q�ҳ�ܷ��I�\���E�I��m�#��� �����4��!��ٝ	�C(���1�\X�P��3Ļp��8�$�(*��$�Z��'E�ϔ���
�1K�R���f~0_l6kc=�����Ts>m'\��5��V
}wo��5ݺ���׌Ｆ��\I���;ẓ2�Zd�yU!,�}g��O���Z�;۷oܜ��.��so��~�����o���Ւ�dAb!46����Ɵ4�A����&����*������E�a�$��Mk���>���#�!qY.����h��]�^-�nЋ��1S0�Y嘹ʭ�ԔB�dA�(å����✰��M�"��l��
b+gg�|�@�e1ꏘ'-�w�y��ٹ�o޼��j=�8�DK��5�&�w��
�ҏ��eC�.�$����z23�U�Ъ2jh_��;���e�s<%���AE�T}s>��֤����1�I�	x���޾,b�`�TS9�`����b�9k��:qaF�&����󥱛���G��s@o�脶ֵ�ڄG,���kGy�p��'Ɂ���`�&�4u�,�,HE�j�ee���:�vc�}'Y{Cj*�9��Ys%6�����W��>�<y�����c�kD��#���|�
��ڗ���O�0%z����
����wLa�����l������+ �{��4�f�ԯ�ܵ���ɧL]FQ�ٝ���sC4��ww&ׯ]"�<�s \,��N���W�I�:���|.@���nf|�o���VHT=���G'Ǻ���L͙����5k�Z�y�Yf�[�"���>&N��l�%��m�K�T��ॅ���l�|NM��ӱ�D4�-��?������u'�>gw�r7�H�<��i�Cp"W6�p �r��6Q��+��%T2�Z���Ɯ�[�p�G�A �FKK+�kN&]/�i���e���u�a��B2����{с�pK�ҽ��.�6�tZ�� ��5Xd�}���7�j8*U]�i��F��`�bwO��T��°�����P$�u�����{k�:;������?�4���y1�ߏ��ܻw�T�q+�2�-4��<���BRI�Ӗ��O�� �	�,5EZ��hjj-7��lh�A����3��PȪ@��jL7O��
�Z���4����ġ�����l8��D���𐖘%[����G�p��tp@���^���r6[	��\��61��~�K7�cw�x�O�}J�"���Ҷ2�8�8C��Y�V�WD��t2�1Vٚ�Q)ܢ�c&}4�A`9�F[�8�1=��h����}����e��i�[���z#��z��kk"����C�Ɖa�� ȫJ�p�9G�_���'j�ԑǝ DdE��>�r���٣c������4^�^_Dc��M�J��','xB"�.�~�f�������mP�q���t�������^����p �<�e���
�;���7�����7���vv��'�l<`v�֍�wn�E{��_�._�f��8%L�?xW���ݘC˳E��S�
b;�4��X����E�unpS�<����+f�eE�zh�8a��ڵ���Jc93��<�~"'ܕ�:�UKÝ+N��v�5��j4���O�\�u���EV:*WO�=���<���������)ʊ#��"}��L�O&<�(5H�r7�B�hnѬi~���TT'b3��T]�.}&�l-�M)ud���u^'�=@��Y'm�O\g�~1Utz�g����b���jvsl,F�h/DJ<ֻ�/�[
��.f����h�op}9�p����:������b=�xr,|X�i� ��ɈC]�{�cF<��E)[ĒMg�L'F���A�'�g�=0D�B�{AZy��%�)V φ[���l�~\�)���~��jo��t�L(姱uJ�6���
v����ɤ�e��+y��UU�V��#���nj "�{���c^�|^���9&q��7o�~p�� �����3�D�17��q\�x2�
��"��/Ws�f^]R���\e��b0	��ݿ�55_N)�9�ō�7Ԧ�J��>Z��������_�n<:�\k_;;��-�1$���,
�}�T�O�a�B���f[&��f�gL7���g���T\ǹ�O�E��Z֋��%���y׉�+��t�Sؘx��s��?��q����S�*��򭭑��
�	S�c�4������,�c�G��_��@��x��)�)��X$<����c�R	��*�(U�ۓԥ�pg�w�m�u�d��A����xL.F�3r��������;r�<�,*��WPFU-`G�ݙi0��,�2�r '�Q�VF�շS�RX����">���+����o�B���X�Ʊ��xq���/�-�҈D�46�L1P}BCS������\����-ܲD��+��/�z<�(�-���3^�$�Lq����p�l~:���<�oe�,M�J{�'�|�,�r9�\�ƧR��C�YB-r�iϟ?��
wGᓜ����V�8��U�=�7b듞eWB���&������܀p'��l���;���/P1���w�2#B~�w�A�I����@V+G�&���i�{J�Sv�l�'o�TZ���Q���	w�)n��"-0�	��������8Ş�=�Պ<e* l29��۫��qWQ��m��?����J�m��CjcC �h#	m��!�:=�%{eT�_j��d�����/T�W���͌�0Q�-p����iCU(�jP�t���Y�J�	�$�n���`�����7~�7�O�
�/|��?|���c��Ew���S�nt;v�<���s��L5<�LX��vj0%d��?��p���=�K�phE~B���
7�wɺ6�'&6\�j"��Oj���(%	 �	��TǷ�~�k����������?HlX�Yh�0
YeT�:,�3��j�H͘�:�8����dU��&Zw�� wr��h������g
�6Fƛ�@�hN=���E��X]����咶n���n`!�J
�*U+��L�Fc�g���q���"R������#��ؓ���c�f��)�b~��@"q�,�-Qb��D����ڈ|p��'�z��۷o'S�4�c5������Ո �<4�!�vp�u�b����9�x�M��TF��][�M��Z9��ُ#�Į桢���[w�i�;Km�AP�^+r�UY�2�u�tF�����%�����O2Ȟ�jV^�\4�V,C���+����p��-(/}ȀD�%�Maj��3���9pf-n��-+c�c|������3�D0���Z��=f�.�X�`�!kf�`ݽ{�0e����W�mȡ�Q&'����&ZR5PJ�nDO%��=/i88��̍�Hc
�VLבo�Y�A�IչP�,�a?͍V�޷C-���`�۷]p��,��2�cڞ��'-�%-!������"�9�-��W6M���x�Y�&���Ξ4�@+l��q��Vk6Jk�:'P��2�g�_��0d��ޑ2Y���|��U <#�ԝ�i�W����kⶒWp OÈ���ݽm�5Uhr��Ȝ�l�2��FШ��!��������-u~��F�)EN��K
�;����I}�q�pL��֭[����'����6���&��A�y�c���%g7���ZLaW.<Nm�N㚡���p2����	� 'r��K�n+�0����q���6~7��!N�v�%\A�x�C��r3{5r.�KSDGpp<CsC����W�����T�5�#�~�#����&iF.�s"B V��#'<N���4��!iF.�_��׾����?~�P�e�.Ȼ���|��ɗ��P��)績%6���bXS�&t�/Vo�ƱK��7�8��2�CEd�H�������
�����{�y�_��m"S9lI��*�^���雸�������D��yֵ�#�.ݺ?����/�]��J�_�)%�TT&"��8���)�۷n�{{��6���.����D����/~���~p�.&���믿.q!��d�ٗV���m�V,�9��:@������v�8�<���L�<�PW�ޫ�(S�1��4`��̙C%+@�֐���K�\̛�OD�4(��R~r�R�M맮��,qYf�x;+��l�ў���;�
Y�3�U9$!Oa�	Wʐ�a�ѱr#;C{`�́!=����g	�ˢ�W�Y̖a_�Lt:��n�^�4�{-�c�Ro>Hh,�,#^f�A(Ւ���Z��w(&���SsRH��x�n_~�e�#�I�k�k�riYl���X��!'�A�h�af��q�k�X܅�k}�x�}JԵ �Xȧ�y�&�v�rvr*I�z�K�I�"u��E�P�6��o~x�#�ń_k�J9��Zs#_\We��ܲ�j�����t�e�(��p��Q��G�熎_K�C<�����F�)�J�}B%NR	91�]��C���;;g������W�ܰ���%͐@���W�?	��X@*�Y�$������<7��Z��p��)S�r�&�k��&�U©â�.VF\pi�E�������� bYF�V��}>����>�?ѡ���}�<�>5��S۷�=	�B�v�AB`��~jI�����o��O�q�m����8��lV�j�fp�,}y^5<�g<k��и����&I5BT��?5�Xx�~��kv(�	nwԄ5�|˅i�X��e�[�!�XI�س�BK�-���Ϟ?!_^nVٓ�c9�t�k���	K��s6S@�Z.b5�^�T@�?����]mhLn$�����8��t�@_���a��VV�.~����镸�,IOf'���r5�)�|?ye��?Y/Q��}z6C E}�է^�X�����P��y#���)K'��gs�A�M���Açb?S��y�l���Y�+xx��p�<9��
�=�P��C$���Tv�`!���X4A��DJH��5��8�2��2� �r�#�7�%��������`��ƣ?�I�,׫$K���%�mrD1��2G�@XV�'�G�֕�\����	�ѵk7�߾������?�g��U�?��?��l��K�X�>����2@)�̚8�խJ�@�4���8~c�7���W�[̗����!��qtpH�S���7�_��J�z�&dy;��������p8�$0s;�L����n��8/zY^Ğ�����8n��ñ4�h��}�����!q�z}t|:�������ӧ��m������RCc����W+97!�U�V��
���f�I2���K���Mܭ���l��.�H�TS����
�����6���h2�V�����N��aH��&K�����z<�c�N@��$�_�ړ�����CĠ�-O���yCD��t�R���pRle�46Pń~$�޶����Cp�6�V�'��yZP}��<*�Jp�Xܛ��1�T0_o��ܐ#���w�a�<sd�6�`�I۳��n�t�ƍX��,�Ku=㓧�Y������` B�fvI���'w��%u������,-G�UWW6a*��R�I��gi�zg	M���PH��f5(�ȵ�
�W����ĨAǨ߰lIn]�YT䌜�^۝NG95��7�Z�/l�|bO2�p�^2����ZQ�l6[��ܾ}Omh�J��<�����-<x<O�ލ��3m�`(����	dg���`d]9G�'GM��c(�&>��nb�}��ol|^�b�r冺8�����׮^���w�r��'��69M6]<|x�OFS9vb1k�)���zR�
��u�Y�L��P�	�Rj_��{�)��c}Ҧ�΍Y�nkg��H	8��\��R�l(�[���=5Sq���t8�&)�a��?k��ځn���$]o��K�d�Nh8x
i�u6�������Hs�NOή_k�u������q'ĉ�k�b��t:9R.uf���c|�E�>��6��֠4ČQ��DĲ�:E9���ށD(�����[��k���DAؑ�(n���-�)F�!5�� h$V/$��6����`�p%�}IR/�x����у���|����g/�4��C'�W��͛Ϟ?�Ef�Vj�_,fXm,��.����e�����2ؚ԰�#�Ӛ�O<$0x#�'�ڌdL6Ԃmǐ^�m��'i���'Q�z��1�US�P�[_��74�	^Ų�����L�4�eݳ�KLB�������S�E����;S8Ы��6�lkkj�� ���@�a��̏�j��˴2�hD�'1�B=�!0��L�R�-{�W�Bc���w��@��by)̳,�>��w�}oH��ڱAWco7�:�G�G��}��=�h��q�1�� [�KW�o�X��qn�Š*��Q"md�mfmṰ�7��05���}��`4�oS��I��{8&ƃmg^��!%���٩r�U���:�����,D=(�_��:^�q�&'|�F;;���Z��DY�ڸM�׭8o��@}=a�������(��p���F�^������`ov).���F�n{gBqf�{���#e[�[㰗�����C��x�^O�>�f�6W�SZ�V#��nL��I�|�M��J>.h=+�y�4�y�19ζ�bR���u�!~}�����_��چ䶰'�.M�H/%k����<z�Ն��~��]\��@uW��bīB�T�-VkxbC���)�×�2
�	'X�ԭd������Vɸ�uᐌ������T=��
3[#H1N3�god��j�j0�Æ\	E%�Ň�z0f�a�H��]�v.O��cg F9�ڛf����V�I�Ք Z-�A�,�#g)�T�΢��]�.��E���k���L���<�@<��I��˚V"�,Q�O�@��N�;S�KY��b &ִ���������%:�v���y2�T���S�Xp")��x<���5�*���f�;������%7��u�g�6u>F�D:q�����&��w�:��|Y~���"G ��I;�ۖO����j�
��f��]�CU7�G�dfXWrn+��Z��NV�+N�ωk�CD,�M�O8�9.z�������_��*���L`sK''HÚdӂ@���Zx��^�h�]�h�^.�Op��
�Ӫ������8B]�:Y0�v�JRaya���fd��Κs])UG^o�I���5����Y�M�}��ε<n�����36l�|S���l<�?T��9��E	���@M���4ʔeV���kOR������LYF�6�����X����ߣg�'b�Кs�K�9�D��
+�X�U���6��6.Q���:z��/(]�(�Ŭhl��(�it�it~��Ś�:��nf�B#8�gGKd��^9�=�"�6������:�(��jmS�%����j�M:e�,���3�q��q��5�v�E3쿲%��|�ȧ�"�Q�c�K{Ą�R*�(E<�)��s7�+
N=7�w��C�s,�^K�K��?�6Z�#�=Z|�S�-��幃�n~>�/�o��Tc�ć
俯�씐�j=�@�)~b�
&�;+�*>�*Ź�OG�����V��̀���Erރ���(��m��(z��!�v*G�E�qdMϜRUMH�f9Amպ4�3�h����~��Kw��tG�O��O_�8|��w��w&�|g�2��a����&�� ���F�C����b�T+��Z(��X�rb�Y�2	q���"�'��&ZAm�����QѱA�a�O�\"�r��#�N��P��7���X������}M�h�����O����?��_���ٟ=~r���)���<0m}�4�HO�'d���#�B�R:?=�3���Ӫ�oc(Q��3n�bA�Z�FJ6�31��N��4�C�E������ͳ��u�M#���&:��o߆I�v~��Y�Ky{eŌ'�� G����S������A�_�'��(��f��\����f2�Y�(Y���*��~m�y�u�tE�	�����W�^%�}�@����t$!�at3i�f��i�����n�z���Ǐ�g�:�t�Gc��7Ӱ���~�W�v	����Y*O<����%yZ�y84�Yz�3 ��J�J���k�]j9�(��bj؈�Z�#�_�r������j<�n���Ex�F���t`�<:~	\7N���|v��gy@���JL�e6����MU��p�m?M��#��o��M,�I���}��2�0�Z{��N&4L�k�O[!gN&^�y���׾��h�uJ�`�`�J2��~����9=��t�������������'�[_d"����`��㑥�`��	�e����0,`�Ċ0Y���jȻ�O�4@�U�W|{*	E�1�K#��̫	�>-�Տ��wݛG������k��
�@�_(AK0$W�'��R�ɭܵ�U�Mc���FOҺ�g��]z
-9��<D��]-Ɉ�mD�}���4���Pc�uKB4#�� H�A(��+�yz([g7ݏ��5,�	�v�;E�[凰ie*�A��*ã�P2t�;1o$��t`q�����07�����W�
���4�A]x�=R�t2��&�V�G��D�ťs�rr�Ǆ���B��C[!��_1��q~>�އ�y����e�U�Oln���smř�1���ٹ-X#�̨^Z1ֱ�%�r�TYpMe�.]�����G��v��zv6il	�R6R������N�ْB�پ��7��R�qR%�}��@K䧱l@�XX�)��@ÿx�aD����n{O�z���`�4Z�B�LV	�����80�8Y4}^݂��MR�r�����SK�O�L���*~{�^2�?,��'�;V��aI_ye��6�3Jj�I��+��:?��<y�;)$�Mpe����	R��������}���9�&bo����`��tz���T��O�H�L6�)���}�Ó&Ʌ�&A�E�##����=Z���m��񀋘H8����߄����k��	���^�;4��\���mݚ�k�^mIOg����i9�"Ӵ"�eJ��פ ���,z:���Ui<:omFx�Al���mQ o�h��}�A/!B�yQ��N\�
;i���"!բ��=�~�-H$�[��X�	���vz��7�d��"<99>7�J��󅀇�t�M}��N�_���!	I耢�d$W�u�h�Np�����V*�k`O���Qב��fY���	tʞ�P�g��$V�A�ZG�k��z$s�$*-8�w��och���$��	�Y0�V�Z�/�NJO+�%�=ߺ�KN)����w\9�g؂�h:�a���:������z�����k�O7x�kϫ#噐N$K<՘��R���"\둡�\S]#}�>=9��:O��O�Zr����e_B1M�3��F~'���m�}엒��А<���_�ؼ�s�N�n})��a���(�'���5H����>m�g7K}mV>>{c�V�p3�"���>}
3q�����b�a�
W��2�\S(�T��jMPSp�j�οXpF|l	b����5�l�M���8%1ps#̃rM'4�L��&��Jk�Z22�U��n�z��4�b�Ŷ8��T+���(Uv�,��h��t6v�v�'�%�V�X5�t�%,�6�}[�G�,�j6�����GUg�ȿm�aB�J��P2`�Y�Oi}U��J��m��}��MiXhE��1�DuU~Z �n
w��~Sz.n��k�~`4���e����/|צ��!�>��7u���ϝy� �$z�h#�i5�DPH���P1P�q���qY5ƋO���^2���}�b�F��V��M��֢�l-�кb�ۃ0��,7�	nAcUu�9��o�43�/nV�`E�����嫯���;��k��*���}�{����q v��WC9�"]G>�Q��{��Pe�{ȍN.
�JC�Bh7̕V��$M� ���|ow���+�X�b�̖���L�-h~�7m�״�����YV�Z�p�`��˲������{E�)�Ep�_{����w~��=�ۊUͦn�����7��Βq�P�8��A}�0X��r��@�Cn˭����l��svֻ#/�e�X�3Aۄ_D����Ă7��� �i���˖��<F�f[�G�/�
F����#`�˫�M�1�d���$,D��ߚL�wvGc���*?��#����.+1�biE�,߷3�	�HRή�+6�.G�nCe��ƛZGpE���SFt��^AЬy�T�kj�e������Z ���k�A�2]+��"bW���Š_à���3'�u}��x��8�[�;��I����{[ӝ�}�p��hYlQ��9�=	7mV�r^�Ń�%]�l��Ϳ˓��aa ژ ���D#I����������8R�m%]bCe����ɓL��
#�b�gaY&[�W�^�O�T���9����`>[ΰ�"��ɠ?2�w0����{W�`5�F�$���.wPTt�&��۠eI|�B��7�%���R�<���'�7O�������k�׫�Z��]'2�d[:��4���:�j��`�1��4�9Vbk��QD�@��)N��P��ӆ"v�d"���];�(4�/Ԙ���� ʵ����̅�<q�:S�z��mB]Z�}���n��C�(�-��U5�B��V�-qxm8W"W�S=��Z��\���\VQH9�ڦ�B�Ϟ���Ȳ�3�)wy�GX.�l�6��ַ�utx(ؾ�2ꥮ�O��O��9�F���2��Ó���|�u65zjAKZ+��ش!�. ^W8�.�y�jj�fܔ5�4mA�o߼��|!�	םkNi����O(�����!���U/W1I��S�@:�Mې��s��`0z��w?����T|�(��ɨ��ӳ9�����ؗj,s�g/�3f�Dael`b�k���e�*	��͋~�d<0'������h]�Doo�vu\�a}FyfŬ%��������u3����Sl-�8[.�JLL''�����bŝ�G:�
�Y�V0�;�S1@%��r�ܷ���oݺ'qr�^��O����]���}���g����/�&&�0b���k#ɂ�pz'��5l �o��V�9��.W�u�T��sen�O��l��|���G��d<?xq�ڕj]�����:��{��5%w�e��ڇ�?�F��C�Ck�%N����6��)	|>|��)yZe�i�4�����,��fV5$z�~a�u���&������fW6��%2��9���9)&2<�ۀ!Yݵ4�u<�L��b�ƭ�z�:��w�����x2�q��bu�:_7m�X�	�1ݖ9�7�	׮]��������M=}����/�����'��'?!(����z�d�.�>��z�+���m�t�����Vs�RN�w��q���E#��4JK<���T1BDK	t$C�/'�y����̠\�̸G�z��ً/ʶTu���@Կ�k_����{}�1�UYJ4�<R)�s�7���\���NBh������ S��9۔��r�ukm�S��^�F��M7b\Yb5x��sTuD^�~�|��A��=�ҋR���F)ARiЭr:��,H�2B�@0H�Ϟ�ʸ�ʓ��>1����Aw���7q��/4"̂0nn�i�[�H�Ē0}�ܞ�ᒈ�BP97�l	Ǡ���5�Gg	��r�S�t�t�Zr�u66�l$��Pf��_�:�	��g��
���Km�+����y
����rܴ�v⹦,UR��"b���������W�!N:�\�F{{;Buy����S+D6��Pׅ`��v<��+A�j+F�N�;�d�G�PppJ�2!�sa.zM�ݰl��g)3��KA>��_ ��ۻ$�Q�S	3��NA�=����ƌ��wQ���*?�FgV¿�ԓ�]J��D���L�&�-�>��{�8���"I36�It�j#�"�E�N��-��}^����c�]�c6��mCe��S�=��Z,�ZA�5�F&�m5��~ڲ�[��^�FB�?�����!�u#f���ƺ��.p�v$� y�1�bp���������RY�uVb'vS�:�"饸;܏�T̚�2șXJ�A�42��3)fa����}O�i����z��̆��;
G�6A;�Fw�D���v��p��"h+�h{{Wn�<:f�l'$�bS����d���)q�v��/�Z&Ip�qc
�c��SQ��C�_�q,0����.YO���E��j7��66o&�H����&�r������Ø��:}�	�zc����^$��ƾ��,��Ц� ��L�x[�`j�B�	i���k�`r���q�<[�4�^�W�0,E�J`�}Ȃ/R�:�@0�r�=2c�����/�RP`;UC��ٌ�ڈ�����k�ǻw�Z*�9�j��{}6���7��;w�<x����S�i#_*q�;Fj��]l�����4&đ����en�9$8�򮗫��<��3[�5��,�$0j��/�A���mc:
��X+���$�p�)��+W��O�@��կ~5�WZ7��z�.��W_�~���J�T�8;�'��m�"u��Ca`A����/៫3�@&��ّ��韢؟Np�IG7N}C��0�VM��z���V��B�+�"7`NQ\�G4��˼H&{��M�d��d~=�Z\?����~���8�'ս��6C�@|ļ�|�&+ܐ;�F-)Mc4�S$z��͔Lm��0�j=�g��9���S92Z�J��˅{����K��6�ʹ�Ӓt����菏EZ4O"����;�쐐2�c˕C�ݭ�W��g)�M�ܪ
YF�튱E�Di��`�Dt�)i��=��lz�%,5�̔P�p�1\檌_�Z���B�R�x��oe�-�������q;���Nae�ʶ\[3�B�Ɍ�2�^��T4%���u�y	E��G|7����aZ?�I�Tq��d���F>��!"W��n�,_�����}�	{a��J��F�<9�OY�ӕ���p�:�,�
��|�4[Y'Ez���Uk7�B�i��K*s�Éз �;�8�Ue��u/fyO\l���<��ҤS4��q^E4��R�",S�'��oy��a-'AާZr:߲�h�E��,U곢��a�H���|!��a;Cp`��f�gP�Po�'9�w%�e��󺿿�fC����B6Ya���>ǰ�J���p�ɪ�^}>��XV�*���>
J��8�<o�:�>"%1�t;�=ݗ����~����������=�H1l9e�Sa>ن�x��@z�^�U��0��,%���pXm\���gr+771KQ*�5!����Ґ�������ׯ�ikw�`�͔&H@6�I�!��ۅ�	�x:�:���P�l�#o��Z���U鼰w~1!�o�ROa�5��"�Ո�AC���M����+J�˪]�
𩻊cfj�*Ԍߩk]�r��o���D��Q�67���37��~�腀0-z�>+�[�1�M�B��z���V#�SpH���1���C�Ch�����<|��铇O�>�O^����}����7�q�ML�]�&҇�
�v�DK-�hNy����/��J�E�	sT�ౖ�YF�N8u}H�QI�e~{��ت8��+W��{l�\�K;kyk�Ѓ�10~���'#≨K���7n���;BN�����5��J�YyR��s�E�2t��`�*5cEݟ^�|��!x���m���`Ŋ�K?���x}�O5��Aa<��+��,��ݾ}W�����3T�VK�'�_�r[�O��&me��-���u���f:��1���-������j��ݛ7o*e �,��`J�W!�hTHӲd<��;���`(cD��N�ο�Y����)��k���<vn��J�F��7��,�	[F4P]�U�.�"���ME]1���'�X(��Z̈́<�o_Vnj�nCI$�^�e
�d��}�.�"�Gy���$��1�ʰH�Z�B'{m��G�b��@T��V_�X[D{Ztg_n�Q��L
&d�ZO1��%��4�[�1��^X��ߣ���q��>�FfgJ�*��[�i����xNOA)��vp�,xqz$~n��Z�`�~F6W�s��{T:V�t,�d�I�Cc�x۵k+q=�d]*�,�!���2[�N���;F���H<��XH���z�D�T�p���N�K����7��-�A����޾��ěӄ���{�+ϳ�6���%� ��z��F�����
���T��"ق�ݠ�ʵ���+��܋ǰ��*K�
��e��3�96�|.-�(�b�h `k7�~��oOz�p��y�Yt�C�Lb������>�F,tZ
Y�b|��(��([��=9=���9:��NFn6SJ��A��.�z��=�I��)Jp�&��'�А�ɥK�/^��w��/���l]r�W�'�/���m����'���G�ܿ���_Z~!��D&���N<�O-j�U%��b�q(�؉*���pk<�ϖ�dW���O��#lM_��+Tイ��ޝnMu���g\#�3�g#o��H��]����w�	��x�wu{���b���c��\��]YM�&��5ڭ."�^F�K�a�5��a�:�@*��5p��(��&��'���X-k\���f�ו�Hϫ��eb���]�@���Lq�kfgy�K��>n�b4��je�0P[As�� ^e�ٜO�P�P�������:�Bp��c����[�i^�j��޺;w�2��f��$9ub�EluZ��������c��W�������כ6�v]�ak����kЃI����*;JJ��!�I��+�7;�R9�$+"!�	�x�k���v�9�Xk�������s��{��f;�7~ϦK"�`;$M
[%=��d�v)Y#�BޮGi��n{�30Sga,颊2�7vn1w'��������[�L�q�孹n��A}��w�yt�z��D���'��۱Q���0��9K;�)K��؍����_�t�5������vL�o��~��YZVC�na��������������K�������ef�	����,7_l$�C�H�b��"�ȹ�([�-�ȳ��"su���v��t�g��jf����A��P:����ˆ}ݓӠ���@Bj�Sz]���Qx*I5��8�y���j^T���- �I�Z�k�S��X�YY���>����ӄX�4��v�H���cd,��ɞ����q�b������ޱ�6cyM���f��O��þ[_9Pg�P����K�^>��=hy�Hf�f*�y�i{�w��6Ņ��9�X��%�Pm��7)"F$��ńx�T�EwE�n�)փ\��� ��YU�d��b��>y���ى��W������>����ѣ��|a�_#7���̛��=&�q���������e�����ɩ�,_}�V8:̏t0%hX�``�82JY�~�����h�M��J������E����7�S��u�=��l�	��<���w�<�P��nך�kＶ��c��-�3�[,�L���1%��/̧i���hz�����%�������l9�T�)�̘�{c��'cj6�-�&�bg�At�v���`���!S(I����g��?�����߿��;���E�����a{�'&�&����wʶE8��~Z�9����%�j���6�TX�4}�M�Tc�')��u��[_\�F�߰ߧ�%�=��� ��m4��r7���ٹ����TY��Ilh�O���r��{��}]]�1�*n��ް���#q��y����0v��څ�S3���E��n � �2�2��l�4���}ە�ي�Z���u�X#��p
m�'�0.R��d�ᘦ[2<�����؎j�ՠ@�\�ۘ�89Z������,l���9z:�ls���u@�$��_��y
�hSߑUYie���hLv0sΤj1�5�u���\�!84Ҥ��v�h4�ޒ�ݬ�ј�������z_M��l!�_�bAk��T{&�Qfg��8�}bZ֔x�e�4�b b7.4�tR��G��l��\_�s�6qR�Eh�,��q(��+۟zߚas�_��ߠ^�,S�e+";CPxL��0[8�������� n9sIm)�qf��V��Ms�~f��G�fߺf]߻�Z�X�DP�W�� ;�*���43dI]MD���0�fy�c_��g�8@��zUŉ�cό���ā���aoa��z@q_��4��!��L�!aL0_'�����iu&b���拪�M�<A�m�O}���v�8�so���_���[O�������7��4�=�̗��8SZ|Z"ܵ���55g�tZ;'G��M��nQ|������j��;����.� pS��}f[�fݸo�H�5p����wo^�|��7�l�6(ոޜ���R���Dd���o�s-*%�Fz���,U8�����a���L�fn��/�XB��1�2�j��G�����k��E�)l�252Em���v}���][�yq��㷓�i뾨�d���?:;�ד�d�dbw,L\�)~�����j����|�շ�u�U��t�_������=}rqw}}g�UN�ukаڍ����$k�ܹ�l��F��@m� �Y�f��0��3c}~z��ѩIgӢk����%ͨ�of�<��o�"�t�l:��vǞ���CO�g,L�v2�W��a��)M��&x֙`��M$�؃�w���˗];�J71�0�ծp���U������֜�����|en������ϡ+>
�X��&f�J�x�$̵���,�����ߺ�,���b��''���r1�I��۱�>��ۏk��4�q��L��:��`g��͕�S�rb�h�Y�cQ�vW��X��$��;��Ƥ���ܞnw��X��Z=�8�o�zw���Q�n�n�Z�hXs�ڨy��z�-�Is�R�D�+h�+�ּh��K�2�	�y�4�@�����,Ϟ ��(�ޝ���̭��B�,������ ����g1�ܱ�L�ś>�Kd�����IA��tD�֛1O��3���@4n�19>:���3};[qfR����4�w�6E����kᆲ,TdP��3m!)L���@#�8>E|td1�ёy>�ͽ
��E�0@C�J��;кM�zYL��CǞ�i�%�M*�-

l�/���g0W�\#T�s�o=z�8y�(���)g����|}�)Uf����J'ذGrt�!�It�9I��7�+5&���-���'�~����0�)ڎ5��\=��*-Πvv5еsS��a��>=ø����H�+풓��*'?I�K�bs{��7r�{ZՄꥠfv0�.KB&n�i�'�kp	DO��5y����M�	V�4�7��8���w��YR��e%�Hf�I�4�#Q��O�|��P����'	;h'��N�W�o�}��(���իW0��ߚ�1v�.P7��y��mK�������&��w���7w&HfP�l]UL U!����ۆv�Յ�(rӼ�	`��|�`�m�E|&of�w��7m���x��t�p�ڀ�z��wM˘*@��Ҩ��B9ȱ/��-D�ɶ�<Yaҙ��&=�1�.ñ��>e�����|�z�������[��"���2v}�������7��0�і��G�Bv�<��灃F	�& ��p)��1�B~:�\pK��$�ϦsW��f���KiAm�]�¨V�lM!eH|T�ϋx�[2����6��[���H�f�?��[�<�2��e�������&�)��/�z����d� �@�*SxUL(�?=fº�}�~V;�z�t��#��Tb�r%�ת�$l�.�ȟ�ٟi��]�=�-�c�Ӷ�_����G�[8��yh��µim�Li�g���`�Ș�=��*)`��;?�L�ɴ�(a�MPG���X�=��{C���l������?��Ǥ���2N,�u��*�B�Y���ϟ?�)�Y�����_���������APq�����e��K�����P`�9m;L�������}��SU3b~dt��J�;���%>4�p���ȅ�@'x|����I|:�����
D5Fq*�8i�r2�O��ڷ�^^�j7�����_Q�,�2�'�-�z0&IΕ��]��1�B��\��ɵ���HN���D��8c�%+���J̀Κ'O�`�r�)���86�_g��X�tv4t�=Zz gF5[����>���<E1���_�|Ψ�SW���?����o��6(��VإS-Wi���a�\&A�������
$��3J]��D���������aZ��9p|Ռ�x��f#��>afώ"5U�{j<��X�Nu�A���#k�[��E��^m.ui�~��C-D*�p/M�8 :�i[�xjX��Ve�1� ��:;z���������� i$]d��GL��~��Y���4�*C'rČ0H��2^3"I�	�F<���1�5_��a��O���\Si4��؈�F`CDJ��!��|�����ym{̆L���؏�d08��$8�>ա&�wT-]�K�EN+�E����oz�ⅹ����P����CtYeQ�J*K=�DXo�%�1�
6�}M���đ7����"��YT鲳��#n'8,�����!>ȶo�g~�00.y�p��j�p��Rs��R�%�%�� ��n�3Օen\�Z�P!Y�N���~��@z�?��	�/~���F&֡�K�G*LanL(���ĭȿi�<9T�������K6{��ǁe��=zt~���/���<K�?S�]�%2�P=���vJ��Ȝɹ��e%-EZ>PZ�D�g��{0g�l��#1Y#�gϞm� �9zms�5h����c1�,|���Jζ���$������.�8ns���<�Lj�L�mG4*Tg�B��foB2٥;���K�٩R�i"i�{3!�-3�է��� ������,X�"'U�˗/m�n.�h��Q��&9Ղ�ݥ�v{9�.�hJ$zF1Ϫ�X�	���cGϝ��L�"��g�E����&:���;0�:�G"%1R���#��@������`K��y��fֳ���N���� ���sy
����W�dv �Eu�RO�=�:A��F��^�������ӧ�aI|�1���XB�*�/�H�=�V��E���:��ؓ!s#���?�@�{���<��ݽ�
u�N�C���������L���v�}�GЗ�6 ����T^%xE�䍩�-��}�&���ɂ|<zz{�y�/Vt9�y\y�&�k| �:�g0���xv��nem���L��fp�P��AIҥ)�� �y��!����L�-�V=[��MHt�=0�o���(IЊr'��3�c���
�b��b_��.�Y���J�znܘ�!mh��Ӥ��Ǣ���H�0m�+HRg�J��n���4����
���e".�T��8\*�vu��<0Qk7[�.*��\v�'O.�{������ t2^IDWi<n�@�U����f�~A�� ]#�-�Ⲣ*C��cEa
�S�.�I�u^�1ɑPi�B��	��LM�ꏉqS�����s$z4�"���Y�~f��uX1S��^?�Zߢ�R��?�����ؔ����f�Z�8���������(*γC�,MO�!e�
I a;�����ŭ�����?�J����lt�߼yc6W����w1 ��ws϶�UME�?m���@6"��Aͬ�zL�I�Ho�4aѧ�W$0m/]�Ѓݡ��$�`�2g�t���dk����T�����W7۶ݭ���%��}�4xp��_�k��M+}筷�nn�}�Ā��H�"�̥�i�g���S9:���w~}��W�I}�بc6���|O��ңm":fǀ��	d[�&1��4��� <K�4�I�e���u��t�zS������9������Ǽ�ڗ����!�_l(�v`x�0~��	8a�uW�ǆ�^x�H=f�a2$�O�b���ġ�K'�i>�����p��]�ѓ
s��J�Ő��Cw��Q�]<:N�1� ��D����F�餜L-��̅�Z�U�tY�pT������?��׿�x��W���t���u{���juQ�uSG4��&�2]%���"JKr�8��S~^Y��9�� l���wssɤyurr�5E׳�Ֆ�vXjAb�Ť��_HM�Q��O�Ū� ������$�I*�Y ���TBDd�}�ѣG��m��T�<K.)`}	�L�2G��G��Ѝv~�Ig�'��C3vm��W���O3��65j�X��S�\̉p-�vt���ظM���`��J��2�$'���c�e����~��|����_}������3S�����qj�=Dq�)�4�k�{c�@^chۏ���ԁG,x�I��D�51j�u0��"�1�f�tvr>�?�xR�o��T�Y��#y_� ��A�X- +J3zQ�z+'�w~�C��_|anz�L%P�������n;�}#	H����RjJD1�c��i�G�����8}
9��e�uԀZ�B⪄�ܱǙs�$�[��v�Z)���9;;�1z����H�0)H69�tD^o�$��	�=�|�	G�ţG�^p�J��%��/����I�۵�L��
AJա�3����߫�io�+� �e��y�9��v������i���E����a�C���C!�d~fE�����C{����J��䎑P�'��>5��/P/\H�o�ѫ^��r6U�����C䆚'3˂u�N�B�^&�NE��6�f���ʪ��#p:q
��e��6��m�ż��3Qm_�D�Z-I?�
ǘ��ͱrys�/�%��b�
ُ�ԋ�B�SS�'�gE駔��V��2�'1ͨ�c���~`���,	���N�Jz��\�����#�A6w[[t�f%x.s`6~�����c��O�$v��h)�_�6���^2�$�
j��_��m60h�����Ϻ/�g>��?��M�j6!E]�*��L�ͷ���>ae��b�7�sEfHQ�BW��wan�v�n��s��(X�`'��̮imHƽ���b����&]�ةg8�@t�2�{̿���t��L�v�~� ���1��|�O͟���Y
c�`>������|i���ɛ7W�_�'��޼;dg!e;$ �S̎!�R�ް��]��\�mh5�Y?��=�2��LI�̳X���99;�� q��8�'5������R�+��M�w�nk����dM�1e9 �����rs{o���yB�W�"����5<��Y&ww�E[S���l"�Q���E�K�RM1�3�k��d�]i���t��s���I���n�����zE��OQS�"�$d�%��0v�Yf�Ab��-����Ȑ�Z@���j:?��o~��{~��s�V��꘣5�.L����|g�3=��d��}���@�Ɏq��� ����g S�bQ�Έm��v&��3�ZG=��%�=��!G,�,���w!��k5�dV�] 3��v��r����R�-#�H���s�w�f;.������}���u���7�Y�m�nbOn���1һ��f���3Za�$Ƶ��}�Y
v9�mA�Ċ*�!_n��^�Q���!���Y��g���}��c�.;e%,w���Aǖ2���
gL��9��R��r��5��
���5�h�	����K�V�®cJ�������uGe(��sCGqט�U��$��]؛����#��)G,�Q��\m�T�=e~�����R���
3���HH �a�%{�b"���T%�7��F��f}F$D�t��|,�y���6|�>� ߺ�5(x��\���*�l��06�F�Fuc���$���f�.�2)�ַ���
�N[�;UR��VX�O�����r!���#i�i5�4Q�j��[�T�Z"��J�B��ԥ�7&�0<Gz/֞}�ip�aɃ����>��z:�y�^���ͧ�8��,�9B_}�|��(�� �r�dB��^,����L|1Le:�b\�4��FD�%���(F�>l��&ߝ}̟��w�\�3v��5ZC���׷/_�j�������J'Q�!fNh�|��q��-G��B��f�t�rq��q]Up�,v`�ճv(n�K����Xm�鳑��!%�C���S�Dqov (}��U�S4�6<���-	`=Q�H�٣�����I��<�
���6��7G4���~�z>G���+ ̌���W�`��a���`��@�{=Do;��;I�P��u��g�a���mp�����{2�����7�j�={f��,��y��3��� 5�EQ�-�#��k�x�,~��#I�*[�>��B[��L�@�����3�&�+�7$_�.�-��5Ѵ܇1��PO�=��u����F�}
N(̗��%˸���F��_�>}
A��@��#�YTl�h�)��~�ӟڥ~������3#\��>'�D"�Ӳ,�E�3z��3�0��G�;�d�b�9&�����]NO2��c���D���Cğ2�Z�X�CR��5\.W7j?���W�W?���.����/������'��=�7�/^���ٷ�x�R�P�v�yɃ�S`̸�;��N#F ���a�#@�\��H|Y_P�I����Z���<�2HE<Aca��J	)	��T�>Ř+H�-��o��m���յ�.2��N�Q�67N���E��:�҂ymtГ0rD�X����nL��������t2NK��P����-K�~��S��7��h��:6�T�`�9�b3�x��)��=z'�8��R���a��8d��훲�#t5�i�&���ĥ*�nl{2 �Z�y ��2d]<g��A8�����b�1U�Qk.��Yh���á-���k�-	C6bpS]a��͖�hI��[\{��)�>�ᎎV	m��g"�a�x��ٻ����S���4&�lm���n@Ը�|gN'O��X�|.w\�&�������ڸ"L?��N̴��U�H6Q�H��:5}�FC��Tz{O-d�Cr�mQN4FP5�Ő����X�������_t;�t�?�s�RM��İ��;V_�0�7L���&�{x�M��X�ݞ���� e��̤�Ԥ�}k5���(}h�%�:t�9{.�i��Pw�T�<�4*|����DT�I�]�vӠs4+c�!��{���Öm�d�!���R�P z�x*c/cd�E��v��7%
�Ѓ���y��Ζ?�яn�����1�}1�ޞ�^�@d\+߯�S54D�JFh�YR= �F��M�E_�TѺuvv,����*���r��`#z�'\	~�ڐ�Xk_ʒ8���ߥ���y4ͭ�KO���|A������l��)�ۻ�ԒɈ�^pbp�c��T�m�0�$�����ۍŕ��C����J+���^������ĘH�8)��?� ּ�8�E���z~���hp@x���vv�I�71�H��~���m���o��w¹^�GȢn�F�$L3�'D�t �H��`9J��������0�3�-�>=�����w��C��C_�Ĺ,�Yr"8��cr$��Շ�?c��F�"dgA�G}����Mu��h�����>5�����2�a����� iD៨Åj"�y� i�\}/�,���,�%O�菉R�s��`dV�4�':2.#3n`�?�^˫�q�=#�o�*�Δ��9�ER����fA�{��|a!����'�|���nw.��$�.��_��%�|�^�1+�YlU�$��Y�����P��(H�ؐ#�~L}�O1�j0
Rb|����U����R��μ��r8eǗ˹�����A>�y��݄!p����˗v�KDX�-سe�֨"�w��'���tæϵ�����Dl7܉��>�R��BU�H�Q�ԅ�I��'q�E����=�k����\р�x2d���@�nQ��[�i:�Gȧ�g�U;lp�Iq�)��"~İc/M͊1W�9&�\��D60����w���y �Y:�<s��[�d�]3�tz6y �C�d�5>%�	5��P�"�Ξ����<v�8U�i��O0��Bfw��diuA�Eq}}���_��,Pׯ�b�`P?��2J���@��W��G^�Ah�>���W�,������=C�*E�L���N��s�Hv���f�f��V�Je�r�s�O.�>��#��j�ɀ��W+�c����fb`1ڜ/��Q~sP/6�p2b21��)�������h�
օ��y�I��xr|�,ym'�N�+ӻ�$�0��OB�=�9I�<_��kVAÃ��|+�{!�������-��5fVA8Z�Vu��Xw�*{�_�lĲU<6z%31�u5�Տf���zVc%��_ʡv��+�r��.S���~�����Ee4����1=�b�x��(�3�"}�(�b�M 
�ど*?;	��Y��E4bUK��k�!�EE�G��Փi�X��k&�Ժ���y鸈uB� �jΨn�I'�8y.��|Y�WO:-Ǣz�T�;�pz�����:��Hy�x�����k
���?��?)#g�a=���{�)o���]Z���t��$��#��m2?�Di�[�	�g?�� ��6��	���H����!����ۦY��Xs^�4��� ��c���a��ş������?.,I-�_��L����?>~������k$?�����V�(Q?�/��:]��)w��ӆ�R0�՝��d؃��Ө.ٓ�)�mCOb$��q�fj3����A�s6[�{�@q`r��p~��>�}���{��uM��Q��}�������hҪ<��|�M$�n;<Dt��;Cbх���q��{�h�з�uc22�沩�|h���w�<bh����k�y��-�w�wNME���]��zZ��t�F+�~��O|^����{͞����mw�܍K0�Ǜ;X���k{C�o����Y�s
NX�2��c��{�sn�������K=G�_�GGS#����U������͐($l���Iy��+�B�.fnҤ�N��z�JfH3x� ��¦��KIm�SӰs\E�,��ʶ�3^+N���f{���(����޹���Of�d3���&�689>����6�5��{sv�) K,��0v�_��\!������+� we-KY
��p3UY+�|��<��jվ,�b�Y�kq�#nȅܱ<Ke	Wd����)���*��9���m���m6����BPM�C���=���=儢�*� (����#�I6�Ч��Z���}AA�&W48��ȗ�d�gP�z���jV����U<'j�3�m�V�QJ��^?)�Zw��	�V���J<j����I��s��6	��5�Fz2��{�[��4k&W�[;�[�wĈi�ѾK��1$s�ؼ�V�Y |ZQ��u2���TH��+��h�D����$�/&v�����d�57�����|���E-{9�o������G�������W�
���&�l>YMכ��1m	�g�)Ǵ�ʵI�B��F���B��R��`��1%9v�{s��f'?����>kܭ7c����c2�^�ػ=*��ꕔ�����&ڤlx�S�A����M}�G������I-��n07d��g;R��M�v�A�S0vMe����1-*�d�V��O� Gը�]�ǅv��o֫�eg��ꚷ�Ӓ��d|�98Sqf4LgΦ��6 �W�`�}�L�ӛ�;��f����#d"b��g���0�YZv�65^�:��S�$9����&��k�z�d���op��s�FG�?H��-ū��Ku0���I�<}��$�B͔��7�)Ȣ8F�S�U@��QЬ�^I{;P�V%�`s&�n��6;��(v������G�i9sb��{�T�:�p�:;y������o�j��7�r	��FTz.d�ַ_�r�@b'EY3��×x8C��7	�b_gMrҖP<y����d�i*�C�����U�aѯh��Z����I?K�TY1�$����է�Z�����v"x ���N�f"j����b�MN��V��T�t���d���_��U�PiE`0����_E�����ṟ��A�3�3�0�� #&zn��v2��`OŴ]U�:h^pU���l�4�%�>� �툴����>�C��`ƣ2�o�¼W�����I,��j�ݚ����f�n��"	5�v�S�54<�DKm��H0Q��m`~nL�%²%��Oi:�v�7�5ʐ�`��G���Ӊ�@V2-0��֡����/�뭛�6��ƹiC��r(=��A%Ƒܾ$=����̝3Ix��eC������:[M��I�HP��3<��P_̨���Lǚ��rc]������cǔ�����?d�00@h�[�2v�Sr	d��@�$���C�CA&�-��$Y�h��)$�X�%e"n��nje�ߘ�e�`)O&	�t*��Ľ( �8M������ҊP����2��*��=�G�^]]�SX�|*���<afO�;��x`M�����:�+m��2�g�,��.d�=t5=���
Q8�A��m�N�LU���XJ���~�ŗ�,��W����D�b����3�NY<;9����z=���^	\��<������J�b�7�@_�5�Q�+c� �EZ�Q�ez�Ե_��`<��ej>����9x��vVA7����'��������������\"��o^\>�\���{te��4a䥶ʞ�w�%�r�x��q~0D2nF̲��ɲ=H��ﻘ��y�nws|s�5�z�����O�=h�(e=v�^3%���P���z3��A�i��ow2���M���*��	xx`�#����bFj݃�ru�c�	�GB����(C��.�|r�ھ��}`��j�YHX�ė��R�A~�#�E%��	�8��o�}�'F���A��R�TzJ#J��o��/�����;�� m0S�q<v�/^~�w�w��� xN1_�ի��6�H�4�9�#��{α<lD[�yw�}�g��0�b�������w�1m��B"+��J�:�b1�u�B5Z�2�0"�<::�`,Ef~�b��ODۤl�;(��Pc@�O~���Ej���h9'������H�lؕ
��/_s�U��䕲�9Pvh�R"L�~B�����y�pM�/Nl5��v_8'	��\�ظrrg��-)��%tr�f1�t���8���j�k�֗��N���t��5��r�>�<�o�%�
_�]�������W��J�,. l�*����"�B�.��Υ��i%8*n������М.���Q���D��t0{:�
��ߣ��$��`�;� ��6���f�P� �b�߬_�~���MP��f�zbr����$�R���'����X����N[
 _8?݂�ɇxb`�2�R�k,� Y�,��sf^�Q
��?WZ	�����r,��;�X�Z�����M9ˬ���h1��&	����FD�D�ˇsU"������8f��8�b���V�!�C�,W����Q'�-}�E�Zݤ\��R��	�1�I���򨙓@��d�k�D �k��f�*o7:���{����Ą�X�̯��w��}AW{<@�F����%J���ż�ۍ#����餾d�$$U��lѩ<f�!f�0�j�>z/�����`���b8��j��GY��m������kW7<��eY���Y��Xq�f�:9R�\��L� k\d�8a�¼ˠg���c���X�Z�8H9i0�`U���s��{�7U-T�������TG�qd~���g?��o~�k���Vb������)?��ZU(��I��e�g$JR�5�,Z����و0�N�z��������j �D��_����.�{�bm�dd��l�DM`m&>�a �b��;�F� 0ǔx���0=�L]�&�)Ĝu���ͽ�k�t��vFı�6��b���oѯ�$���f;&&���Hٜm�;]������?ڙ���\%[�G���H#��E�l�Fx���j�vjL;�f-[6���I������W�M&NG����ZF9�:>�����(�I$�M�k07:]HO���4wNz���UAr1�ʜCmo��.x�f�:VP
�y�Q���p5b.�I'ǐ�G{�ؚ��蘧X��a�!�t�������~��` ����lkL3�%��c�)�����f�B$����>9T���"�40����hߋ�  N���i��Oƒ6/|�@k�2RD<%����/�"]Y�:	�3���t����p�'ő2#�nw}�_����k	�rFi�Sk/��l��'�U�H�4j�nf8���S�pQ�1�{DY"�JA�� u�(�3j$��Ԏ9��0�:��&�ƔJpt����kX�`�i�s�u;w�jx��s��*v�U��D"��Bp-��	Ym���;[����O@�I�C�5C�P�=�p�@����h�\8<�8D���b�Ǳ�1���J�[I2����d�XX�\dAeH29�b��+�u=r��^�G7�I�"��5�������9��2]���|-58��������:3�������v�����vt�&b� �0�{3]8�}7Ea�\^���фV�Z76Q� P�}�*Ј:ߑ�'��]r�����Et���Ц����3� ��xJ����4��`�hU2R#�������Y�{i����Ìʡ[��ٕxf|N&�� ���5�W�G������ĤPP�����׿��o?���+<���-Bi��l��Tz������G|I{h�<x�&#.��t&;�="_3�ږ��o�m��v����R���;S8��|=�4���3�*��:pG��f�e�!��駟���-���*sm�N���g^1���T���I�mq���+M��'9^-�eG���ӑ�7h��w��`u�E_�~����7����=��c�	OK�qh"nI�,��?9�3�ўqqr�Qtb�P��u������^60����)J�a�yz {Y��(l�Îa��ytdG� ���u\%�O	8d�<Y/��45���M�*��!9N'�1���]v.s<�C��CgQ��ɣ�ݵ]C$�o���XVR�H�
2S�m�D�1�g7��!N���)$�7JP.Xb�tI6�Vg���������E<��7w����OlA���k��7�W��Ie2�qH2�zj��&���N&(ګ���&h/}P!զ$]��K4�������&B͐��������/E���F��E���-YK� �rds��P�߄T�}��.Bߧ�ٚ�ߖ�U�{���Þ��ϊv�+��~�������c}Ңb��8ϒې��˃��O����a�~Q����j�w��{�?:���M���T�D�*ebP�C��=iKf�d����gtH{$�U�jc:t�����a2�9�nuI�i���ֱ��f������OvM�����h�\<�p,,��P�����0X�i`q�i�œl�hm�����œ'�lw��5�B���<e^ɄK�T	��=��"1������k{u�mfC6��D�N�r\}�I{���ՠ����bړ����G�s5�7�޵�,J�}k®���.��4Z��#r�2K��9���昁nG����Ac�fI�W�Z�	&*���cn:dR�hS�x�4P{wwSL'#M�	}�.!MT3z���e��`��d�N�VI�2�G(���e�L[�iJ��f�天A"c��/��bJ5Ц���#_�}q	��)@v���Ӓ�o��n����|ur��gF
���B#V(��a
	�T�ڃѬgR`fo���8%�ʽ��şՄ���hĔ.�B)�Qa�g������䧺ݚ���=�b#TBV����Պ� � L�&!d�Τ�N��Re�3��O�$��m�k����|RL78۔M�s�`l
��d>[�d���N���G�啞�b芪Ę_n�iڦe'C��:�p�����h%��Y9��\.���̖�|zrd'���hS<c�O,xٰ��0fv�啜�>�����O̶�jR�������$�*�:3����O�>LN)�b
 _NVߔ�I��3b��n�4�Y��*KiB�Z-�����F�۞!"T�n�ѷ��ufA�fu}y�G�Z�����V�X���6:�2׷71��[J������p+\ji�AR���+�r�����E����$���E�d��@'-@s%��~&a�Uo�MCL	Okv��١������èE�0_̩��Q�y %�;�<5��$�,,�kC���}=G�ڐ��q�M�����a�Ch�W������%�(N*s�h]Ѵ����<m��@_�EV}��r�+��D4o�����ݟ�K�E'�V��F6w����
Jk�Y�%�띝���
C3�2�OIzh��ow�bRc�*�2��k����2���w�Q�-�.&S�$;�M���g�G�N'�~�1�d~��"��|�Ñ����ggg*���y���?M���������VVΊj9ڃ&%r�fV�DA9f�g��œ�&����J�ܲ�OR
�ln���Nx��I��o�A�1��Z+���_$I �ȧ]|�c $�`���b9�� �u�n:B�g�����Ť�Q�"�����6H~�����л�i�K����"��{��ʻ�d:��Hx�k�e�n�qw�_~�L̤怡cl[kx�o@�!��i<�J��[%��wC��-�s3�Hyջq6I\n��	-f��lV��0)�d��p�0�>	8�W�0��g���sqd�EzL�A�f4�i`���:p����ݍũ��?~���	7���Z�}Ng��	����	��S?<J�B��b�ɑS��ꡜ�+z�b2���~'.־+��T`��0$A�B��0��֘�����@�bJ��Yѱ��l�IF������كg���C5-�:��5�����M�R��y�1�,3���*���b�������@'Q+0��5w��^w{��SaR0���Q�^ډ�Ds3f���Җt�ؘL�<�Hl��(�M5�h����&M��ݡK���~V!ٞ���Zp=�r�8=���ψ��k%#C�_��DAI���X*��o�{.�p��M;~se��s�vC�?���X���������P�f�⟒��bjίtQz ً/��^���I�_�-*�j�޽b�THT��P�+�������|��Y��{�ϐ��OIms)E#OR���:��P�,A���8LHc�i�����������]��뗛����#�f�G�W���^��
N�H+�AsV-6��ߙ����W$f�\`�3�49k�7��7�}SE�wС���xh�M����}�믿6�����oNNN�j׷�ģ���@*v�bM5�h�����/��R�S-���J���ݍ{����(%���;�_�g�)��$*�x����s��/ևr%/�qm_�xa�fr`n��
���b_�]�y<�"V*0��0u7*5������&P�V���Pp3b�5�x̲���2W��Hc�3��U�l�0�%��TrQ�_B�i*v�Zw�j�h�c��}�2�J�(W��R>����~s�i���^���a���/ ޸���0���c@�Z�x	���ŷ�~�2x�j��bf��}�#m!��/��4W̩@`G���K���H�(��J�сV�J���b��q�y�L����}�]����ӧ�z�px��͛h����+WWIh�K@`a�Ǿ��K��
��6�0��������	���X"��_n�wb���GJdGR����(�y���B�l#	��Q�[����g���
c\ ᫖��M�`g+�y�Ǝ$w�?�x�X�L��I�q'9$�$�J�@d]hן�Rw�i|��՛f�Y��](��e�z��NT��m�`�*��)�_�)B�諕��
>nQ�`a�(�M4�D^ܡ�=�lUG���GSĐ���Ņ���B��i�'J�L&�3.�<�e�G���WF�s;����wȘ�%=ry��{��g��z{&���{�n��*��1�8A�$�1'�Jz�Z0��5{��i@$N�c�
r�곓�
�nX����A�T����v�8E��k^�暞L7�����O�&8�W`ܻ�}���P7�ro���+J�hs�DJ��E�����	Ex��$H�&I�:����i�(���T�R�% w��)8�;���;�EoO���<���6�)v\n�X�����/I��1�մ���)��t���J!�� "	�1����C��toD���yd���.P/ES�8O-���vL�Ͱ���Xe�-Z�N=?�&o�Wk+GO 42� wwd,7�f��	5M~>�.`�:�Ø�7��)��
)7�nM[e���nJ�֣	w9>P��U�!F��<���>��Ow�-�@v��R��}��s`�g��6ߎy��p�R�������@Z�~�8��ڟ^�|):yͨ�E��;��t���v�;\�'�2tp�����(�S��V	�\8i�0�Yh<=v�;�Y`$��Pk�5iG3�m-��-�� �q��&����9���Ls�Zߌ?��gJ�	ٯ�@t������x�	��rU2�ϊ�qX�/=z��{����w�yg{Tx�M���������Ԝ4����u�Y�ѳ�bއf(��b��0�����6����$O��&A�t!�uT��(E$I6W���;��2?WM�5֪�d���t��`�p: B��]���j�<��a�����88Y�@f>��"�)3��s�����s���E&UgP�$|�\���b¦�l�ߎ>��QGMc��u�.�jM�]���R�	-�69��&�E+�OAE��\`�U9_�5{'�ڷa6hDWD]z�0��s"�虠�R�&xD_V�S�Y��(4ɱ�����)#�Y,���L���٫_�t��m�@��jJ[���|ƾHiEi�$�yǿ��G�$zC��\�!8�C�b�6�&�Ж�IS2,��C����� ���j��tJ���Ta��1��u"зC�z��Q�cL�v+���~d�Ȼ��7���$`�b����XV��?�!Vr�g��(y������ou�Pfʉ��g���<P�W�Q�9��z��q0�N�nÀ�!p��:ϴ�I(��o�(''�� 1fB��Z�l��0�;9H�m��$�Mj, 	l)��p����//�K�c�j�����6�^:cP�2Ӈ1W��F��1xaf�~3QW>�$J#(C�Ӥ��K��')�RuŮV�����vor�š��b`�������SyI�Y���30*��6+^3�҈-8t���Ph����e�?�J�8r2�?��'���y}�������?��Aѩ`�7�,���m7�u8r&�k�]Ю��h�o�Ϳ���ema�D�.b� !SVYU�5/�I0�*���sf�g6I���a�����������E�M�}�j̓!�����Lԅ1�lU*���0G߾D�m���?\�+A��/�+B�2����8��.e���3�?��?��(=~u���4ߔ�2�-��2�=�%�C4��
DY�	I�$V{�&�_�A=�{R�=�=N�=S����y]f;�!��YN��s�Nr���j�v*���(G�>�7��43J���J�R�{&���B[�]��4�2v�f�P�<~r���c������5�����XѦ�yl�]h%c�)	��-�iG�r�=�9V�㈉�A�]��g�U͡����`�#��>��������i�,\��|�c��S��>V���?�1#^`O�iRI*W�L�}�J�c�"X��3���ӳ�2wmWn,��8&����� ]Ewz
L��ve�O$��e�Ϫ��&ss�0��1)o�v�k�� :�a���tC�7ww�e�5��}����aC�dO���@sd��}C�O�c|����gD6�I9�[��Aĥ��) ��<ӧ����U�^���c� 夶d�թQ�BǤ*���*�N�LX����M��t�v�gʂN�צi��&����f��<-������IY��P�0v߂*�cT9w���OBD�	�$��x~~{�[�a����������/�K<)�0'��;�� #�EҦ�N���@�XN�&]�9x�-�n׽�.�2Mʦ�sOSQHL��D��{�\*rk27: 5��z����\l�m^�E�*4�Y��ȃ��qi�f��y-y���Fd�����^�&;se��(Q���5�9�_����}���M7��#����]�I`Nwo�q��]ϛZX+�;�Df����<Wj��u���΋2tr���6���˗ׄ-�V���Zᄅ�)љ?�O'l�V��mw[�`9�)�����	p�{����������1�[�6��ZI�Ct!JQ`mSZ��M��"�n]S�m̞�L������qj�~_�.M�1O\۰^������݅�T=y��*�aR� SK�_.f�]��w{`�������tvz~.f��l���Z9�^lAN32�O��z�mM;�	P-p�����s-�ϖg�"Ԃd�ϪDwY.��fr+���e�?y��|����5e��T��Y�M����t�����g��$P���|��V��:�87�]��0���{�:��^��T�|܏�w�¨�<�ڙ��E��yt�T�nz2X���%����T"�I�a��0�vR������nf���������}�Ϧ9��O�4M��]��rߋ#��e)�XLtw�[�}���O?~�λo}���v�7wv�&���5H-%W��е�!Ӂ��n鬥�d�.n�����9�L�����i� KR�^��k��G��2tMM�n�ǚ|���:YQOد������٪�I>Z.SNe�g�CgR��"�%l'ͯonv����D.���h<sIf���(���Y*�nL+�ӭu�S��+���������Y Md���M!�ZU���'�ۓ�:>^��O.�'n-���1�׻5��._�z���n���(�	��f��o����Kk�����v������k�ۛ��I�yt��������@�`Z���������1

�}�����D��-@�d����:izpQ9E����i�����⼢��w�V[TT�f�+ Ξr��H@�kn�k���ۘa�����śW���ҩ��sf�Q{�+�����P?:;�T��?�\�D�)��EzY�H�w�n��<_�(�����Ӫ	�&R$A�	��4�Υ�Y��5-T�Q�o6�1��od�R�et��#B�F��tˤB�M9�>��� Iˉ9fM5�~9��TB��v���h� e'z�Nx�e�UB�/<�����;�p Ix�����%�R;���ܢ0��ݮ�&��1b�J�Z3+,�M_3�	�P���k��1¸l'��a�RJ;!��uʢ7�bi�� %�+=����c�����������׿�=�lH��}UZP�Gk��x��� ��9`��!!*[�7�9I���ד�mq�����n:�c���s5��~@-y�15�q�`�> ^�0�/�W�ay�C`��)GY*���[ڳ�����)R(C±ϲy ���H���[ԅ�D� �޹����sCi�B	Bnra�_TT�,��2���7��<�m& i�Q�X�1Di 8�yLu��}�<����'Um�0b���\�âW�K�6��e����իW�N~�73__�����Y�>9-�}�nXt�Ӏ�N���L�ܪ���ƭ��M8�0�;m=zj�1i{��5��&p�7oP�1���.�¾�39H��a��K�������I|JND���!��jM`cy U>�(��86��yH�a��
���,!����旿�U׎Ϟ}ɬwa^��_~��'�p���:F�y��A��D�f�̥����G�����N�M�J)@�9*�vsz[j������!��$Z0����֮ʭJ�_~yEE��W"K��Xfo��W���g�<9���)_B�HbRO��*��ǠaT��h`a�Ή��32V�Ǔz��^O�w=��vZ7�-���M5�Ï�������8~/���n&Fq	���������3{
;�*�˧9����E/��Wz^'\��fD�kCa��2L��r�I�Z� c�3j�U�,����"�rr��@w��W�E�	��]鶇Ќ�n8���~D\(&���CK�z*��шfC��P��T�/_�|���jͫ�*&NZ+�˔��/o�9�>"?bKi�zs%_�S]�I�tr4wEc"�T�U6�d,�l
�-���6��Xv�uC�U�u��F+%�Ȋ'U(�z�|u}+�8���h)*0�\����O�{�;���L��B꽨��"___�������%���m�~z�J��3%fr��4�R7��@�D�B��n���(	\f�J��Wwt�\#֦�{h���)�$�H��=��YK�흻�s�ƥֶ�d����j��2�A��j�����/�}��_��*.@t�C��!�I(R׍�4��<h��O��O�j�7 _ܤ��Ʒ�ib�����Q���r.����;1>�.2"mr/(?(>�-+�!K)�u+��sz^0�u��z�f�+�0����^�~����R�a�j��Z���H�(>s�vF'�a����rK���9m`�XQU#;��s�23��8x$A�t����7�ڿ�xvޖ�3J��w��S��	���}�qX�<5�xl�L��L��V�ts玎V�pΎ�z�v��f���?��[O�y����\���B��7o���]�B#h�&�c���J��9��tlJ4���S�"��<�-c%�u�ķ/��C�G�^ȧ�`g��T�G`���9���suu͔�w�̛��["D(?����s{��a��F|�U�%w6'C�|:�2���W4#��Q�ĵ�c�#\���ԓ���9.Q�cת#R,�SS���"�B�v�������ki-�����NI=�;���q%��"�Ԯ���o����e��{s���04$F��TN'��cN���T����0�m�G,�4YU�R���3v�,FXY��0iO$�=k����v�?��C37���ܯo���І��Qy��O�&�wdEYЕ�;���ŋ����x�S����ry�68�'E�m�jZ�߀�s�ds��l����7?�ܼ �4�"�=�c�Y�죨T�D�ݱ�Q��ŗ_ړ>~���n���������Xs����R��mR�f�JY�4)	.�=t{��\�N3��ZKm:D3II�Vu"�T���ڶ��d.q�|�ͧ6����孜{�vL�E?��rvq��ɓ<�i�$��E�D���eSblnFT�Û+.8����kOd�V�<8��H�*q����|da0��4at��f�ɂN^�f(�U�EHP�9�X3{F��~�����������0�h��������S*�0�ޜs2�]̠)�<�7k���mϵ-/��Ox`t%PT�]�%��U���3��?��gZ��U,�S�r����hfT(��h�W�=t���4�3>�1@��Kd%l���D:��#�T�M�+�wɻ�rno��?�`3�JfP���E���f�Nh�B!v�̟T�Ä߮GKrQ�rl�������هѨ2�8��M�zi��<��JBNЂ�x��`��"v��f���7!F�������?����?���Ҕ3�0�>�<�Q{ý�˧e�ϱ�Rۮ8l������N�i�%���2�yHB�H�w|������QO�1X���7��} �I�I�@��5�� )	"���t �z�7;b�#��_-��F�8��M��"S�$)�i���D��;!<����� x�T��o(*�QP����0��ӡ�t!�x���8&�n��y9�-�n$lW�+9�����D���~l?��,�+�4�Έ�i��
'���榁L�0�׳$�1ԛ� <��9rc�h/��)^@��k��-�\��qS���R3hJ\��C���"�AB9�b�߅o�{�;&s�w�21������[P�[�ёYt�	��t:WW7�P��F&�����Al�R�ϳ/�_J�w����Lv���Xx�LK}�n���t���O�a�����h'�ke��=�����[3ygϙK.�"w�>�s�� �b6���E/v�f���3���R����~���	��z��jYͦ���ӧ���߄�gy��L'�W1#R��MH ;��_��~o��LT'���B[8�� �w79�8�Z�����a��� L�z��-O���$��{c��]Q�M�v�L<�6O��	��n���n�S���S�l��oTI�R���0e�/h�=� \�j��Ѝ��y^M�}��$�5Rʶ�l�kZ����Э�v\-S�����<G���d>_�$���v���by��{�_W�<*�n
�_C�P�����ۑ�h�۞!2��ؙ�P2������)' ����r���Q��ډEr-C�B���l���0J�`�V#�c�Y�~P�S,��)O�/��Q��13.��,H{&&`�7�ҋ��T�)�OBo�E�B�!?��G�Po�hkN.elt�5�vۮ���E���57]������g>�7r��=_;���&f( �;:Z�����E}�Tؠ&P���cI4�1�LG�QfØ�G���ٹ��0vd^O��{'���w�0��J�)��b��"�J�$�w�U'�8���K�j	��Dqt"�����~Qf��jr�����sJ9���{��X���n�nU� zw/�>�W҃.�	1�+[�̏i_���裷OO��5��LI��hi-v[9A��X�2��w'�Yi�� �A�}J�zme�V'���tJ��=��G�K=>����a�m����-i�=����o�XYM���mn��&�%!$Hp6�6�Eb�����0Qx��$�j۝ڳ4�^���)����(I&̃|k�a��ZUG;��6�Ik�V��βY1��r����ܥ�ԣ.�,����MX�@\�����	�}S~
 ��d2���-�bދ}��;�,�v��-�l5�����_|,F��f�@'wt77��̣S`�i�� ;C#١�d ��3�8%*0�B��bj���f�iH��硧oL|IIƢ��y�"�r����*=,6ɶmS�V���vԻ~i�A��|Zq F(���(�'�u�Zz(~ѕ�2;�榧E���o%#�`Rf�������'��6���jM,u���~\���7��k}3�tq|t*��b�+p,�+v�����#9���M[�Y��Z�[բE:>}$�ұ�&�u�Y�3hn�ݽ)�z���c�dR��r6EV7 6�%��b���DS5���\�I��-{6?`�X���x83��wx�ӟm͋�E��^'4И{���>��f���V+Sd9��mV��1T|���{���Hlw@jt-QSr2v�6����@.:E����/�����z��N'��lzs}WҺJW�SO���0w���%Nd�_�Mhf�`��-WsB����8��[a��صf�`y��_�ZD��b`�E��Q�ەf�MN�3�c��+9!w7o��vj0�'���=�Ob�l����D��*s>�+�����6{q�۝�P�ǋ�٫����////�>~r~v�裏~���2�����db�6�Y�!��4�o^���lq%K����\���8�L�=ד'O�*�g�3�1b.�r�v��	�(����>���j1;]-�>yL�w��Ů_�_>��g��b�Y۱=;:�Z0+f�g�i��I�iZ����D���Vf���x�|�����]���1M�_��݋��=�S��������Tq��A��W#�cz������x������������A�z����]yl]�؃ِ(���&տ���~�a�gf��O��ww����W?��������u��^/N�T0K��13a��`�0=mo���5�ґo�D��8�\*9t:ؗ}m6��S?�d��k+w�:��Or����T���#�)�@�K��"=�#��'`����B����U�<���"I�"Lz���P�i8<6��M�4�o��b��v�2dy�	�f���<3F���� ��E_�x�0G9�6���A�3 	�	�G�'<0}�c�*Bq�|+�����h���,��mS׾a(V
�����(-V�!�p{|�Y��rDf��bq..ӣ5��5�/}��}���������?��}駟�֖�����(R�@�y0MͶPdk�x2OO��d�p���A�N�9*dY���)�����#����0�ǅ��������<[x{|�K�wyW���U0cv��Ϙ�+�Z�^���7��^���ԇ�c��p��l�L�n��,)�Ԝ
s��/��*��74�>�%�X����u:�ئp�Ot���;g��8�g�XD7����c�1��~�� �d�)@���M`II�DM<C `Cڌ�^�B�28x?PJD�0F���S���Ѧ��5�ǅ).r������\��)�].�Y��t��5����n_���}o��H�:�ԍ{ȫ|bŉ��}��x������Ge�1�54�f�F?�z���b��@ ;4=L�U�Hk�xsy��7/�}��뗗�|��w�ɰ����M�z�킧T�7_�r���P�y�<�0ۑqg�ONLR�voN\9�}����J����P,��Ov���3��|�s��^q���*��2Ub���}��:�����!b<�7Oxg��wsG���S��о|���~#�4zZ�O����ɕ9j5IP�����_��9�(�Ljr�{E;�y���K>��R���羛9�����2,�@�Q����$����_��S��#�z�J���?co�lGv���g�p/�* 5�(V�bw�;���MO
��E�N/
�z��n�&�(uSͪ"��*���Ϙsz}߷wރ���E���<�{���o}�5����2�΄���CQj��a?w�m�!�K�t(ʂv{pΞ�@��N4�	=�I/j{�&/;��5�+�|dζX�D@@B��,&���V$^\�$cw	�!|�A@J��aYnT���H@W�k�`�!��/T{W�l���_��{�������b���R!����
E�Z�ug����n�%��y�Ǌ2T�6��nm���W(v���4�1Xu����g���-�vMŽ���9�����a݀���x�z�{4��(��lG�;P�}�˗/�Z�R$��y^���ku��Z� ��Jb=z4�-�+����,�W�v���|"�l@?�Ja8�_»��М;�=n�_�_�v	�)b�6��^ǆG	��1"�	*��-a�mDa��x�x����{^��	�?|�� 5�����NI@��<��q�c�ʧ��g��w�'y��r`�E�^Q�U�C����װ0AđI`ѷ���'@^䚬FYw�b',T���T�5�C��\�W����O>�(n<�t�o66�d+Rh��u^�/��<u�-+�Q�L���F�M�*�T�	t����v�@�D�ดN�t<<w�2��x��#{"�wKL>����lUE:3h��O��}�H�~zҐ�ݩ�b����jԚ!�X���a�#7��&b9ۻ0�lzj��-�'��OT�����,'IB�)���Ps;�v��'��e�x�����T��=�8i���mV�8�R���#5T�P���2�J�p˰��vr�",q�y���f�24o����.o7�XL�ſ�v��/��mTM�?96�4/Ѯp|4�bX����ý�{��ƞ+M�)�G0Θ%��L0�=vD{m����؏La:>��R�J�T�=
�#��x6��X�P��D�M��z�l:�Ѭ�,�s :��I����.�DH�����y�C]�(������.���f�X�$�"�V�&��#�GFhb�B4����P�
�L�V+��R����x �f{<��K,p������r�0�R�K'
.v&f�2aN�4^w��HR��85�AOrG}�Ȅh����*�Zt*R;%�K�=��}V�K�jQ�Z�ּ��8����o��I1:�t���&�,��0ՒkXJ�~��ի9Rc�f��W�z��ٿ����ŋWJ������t�Hxg �88Bp�1���W���B�	|L��߾^݈����v'\�5j�w��tM���|p|l�6d�!s_hA�w�g=�e[VM�Jm��lΩw�r���?����B�=�/�˿���3�|ss�I��}u#evq��(-����	˽71}��c������A�|r���zL���q(�����s���ď�cy�����r9�k6���?���]<􁚑�i����Fp����+����k��־8Gᩕ��;�*0j��X��z<���VC�mm ��c��S�F �(�)�=@:�A�y�1�������W&9�M���R~RMDM8�K�b�"�4� �|y�+t�Ծ0���o	h�(�m&�\��3H�#��\F�y��@z���� �����l�^$� J����s Ǖm�W����������Ɋ�;��m�`/�zL�ܧ��Z�A�IBT��2p�8O���Hn/uٞ�M�r>�AU����	Y�ė޻wĵ`g[+ϡ{3�'Jy�^����2��p�vR��ShkO~yW*�k��d㙩"�
�|���3}r���$���2񯈳�@�.+��<��ro�:D���k>~��Y��s2����WW
%������^K����]��]R�� s��z`�z���L̯;����%��R���YN�����]s;�%����h����Q�:w2U�n��_�~-�7d!�Zm�����b.��ƙ���%�DI�RN��+*������{���)X����S��Ξ?>?8��[�=w������f ��)�p�#�?o�s{�o�������-�`������f�?����|��d��J��\��nݱ���h�qnF��BT:υ"�M�"�t|u�4�c��/~�M%�L��ů�%dF�YC���5p��.�����d/�!�8�/��rS|����*������p�)��~��=��HA��q�ɓrG�?�������u]*{B����Z҅��{8�ՙl-��m�~7/g�����HmpH=���D�~k���"F�np�+�N��F�{��W���v��eɨ��b�}�����z�2*�*Ox�R�ĭo����Ȕ�.����1�)��֛$L��4�mD�稒�è�Ѹ�c��S����l� �O��D@�U�F����r]�'w�@t�9�5��G~��S�����9�˵M����G�He�웧Y��X�4�2�tHN�crb؏g@l��z��C���;GG�����������I���U�VMP���B��E������`J@�2�Ԅ��qm�2sګn������m��+�z8��n!���r|���BeYi����F���m�a�fm�ۨ��y��2�0���F�ŁyZ�ϓȂ��=����m1���Zb/0� X��r|�����^6�����39DY����s�ɥ��ԲW�|V���IZn6��Z���ǟ(u��fo{������4��`GCט�VԤL��u�%�ٶ���tm�1��0RB(>��`@�[)@9�V�� �l��k�s���!ZV�r����ւ�؈��7�G�����m7�����DdCPm��D�K��3t�fɞF�ؿ.���]m�����+���\�A)A����#TD�|�K�+� `�#���M16d#U�yd��[֗V�v?vFNOOU�Dc�+ǭy�N�[�Zko�!4���O>��?������ P5��@��R-7�������N��#�d�%n�w.�t���m�o.1��hʢ2]l�n:�O�C�y:�x��l"F'[��oQ	KP�ТŲ�������ƾ� �zn�He�l����ک��_PT��k;E;�~Ah�BTC���ܥ� ������O�K��s�8l��O+>;;��$�x�P��c���z9�����5[�":����>>^����~�ӟ���W�����_���m�^�iZ��l
�U�:���&�����wOOq��0 �YK�f@$[�,��5�9�zQWˍ�yt�lD�C��JR�g��**�	��~����1�P�E.����/�S���qrs}q���d/��b��aA� �Xgq�O�w�����K�݃O�k�6������]0�͎�9U�]��U�T��w=����d:�O��]�,���'�Y7�0��
8��#��e�b��*��bҮ`�W��s��ĔmI��u�>��1�������V�����2
'����|��¨R�	n՛�4�6a�i��خ��v����||t�����8bЁ����lt/�&-�,1 tm���	@�������]\^oV��$�n���0��v۵Y�4��`���^���'�|��>���`Lǿ��Wor�:������/�G��f�G����O��O������՘��eD
/ϝ�f���`"���y�bh딉���0���vF*Z|E���,S���w��8ڭ6��������|��W�78Qd�����v}]l7�&7o�7�/tF�U:?�E�5?8��i*0�JM��=:9��ᇏ���nח�ga�,�������Y�ސ�("{]p��إGq�Pr}�v@��QӚ�0�t��ã�xJo�BW���υ��]����˗�Ŷ���#.����n�Y[wyq~~�6���hʭY�r��<{}xƆ0F�- ���v���3TR�k .�^A̎�Px�+�$�:PK�]��i��w��"'�+�e�L5�-�(�`��to��z(g7.�sS�Z"	����vX�mxx��bL$�A,.M�u�!��9rLϟ顠3w�s�� J�] R��:�;��N���&��4g�nn���d1�A��N۾��4y���v
8V>���&E�V�����@����=��d:B�u ��y�c�Y�ģ��<7[���U]���Ӵ�wN���7���K�m}gi������������D���a����G�ݚ���О~�Y� 8'�����w��b̶g?A�΃���,?�GW@�(O�.��c��@�:�`	��U�{�ov��fi�~�Y��C����q�GDPڢ����[��~ �Ff�c��{�d���_�Yd�����JB1-��JzW�]��;^6�;mY�KĮ\���f�!��5N'1�W����!��2����Hit��4Y���Ø�,I�;~�*���zS�J�µ��ת<�U�%����(����?���c�E�ڼ�0�Ѧ�bߗ���\n�fv)��p��2��2י�Ճ=9<܀��n�$�2��K�1I�����v׫������Gx���<���~����=x�n�GU��)�;5���*;����f�+��ߡn�����8=�b�u��{�wc�-J�*�󳋗/_���޼z��
v�V+��	�ƫF#�\�3��
���{'rׅ7��U��YI̍�`�
m{*�H7M�Ҝ���[�P�au��Nx,�F$�v�$x7��L�xE�����{�7��|}��Qn�0�#=�C?*,7�+�ӣ��2]�Y���}�����>}��꠮B?
C�i���y;��F��>�,b����龜!I�8�\7��'
�S�u��|��K�~�z�y7�{���_�ߒ2YR
��W�n��,�s*��X��Nu��ڦC��掿t���w4$��@fk��	 \���^�gAJ�A�Jb��!C���S��#G� ��x���1	�_z�m�7B���s�uK����nK=[�Dh�����6�^�:S.R�@�U���Ȏ�/�m�HەHB�܃t��]>y�S������z��{�`�$ ����B�A���db䩽'�7�'�	aITQ�y��9°y�Jb<�Ly(�`~��d��Of���������<W�:�P��I�g2�d�H'bi����W����M�uy~�QsO�1�K��#���P����d�h�z)U]Z	���N
�k{V��2��G�GG'��V+���i25�⛧���΁f�P�ZDj��:Vc]~U�Y���іFa7IIw��T� �C�F"�L���yq��4v�T����cS��k0M��q��$Ac� �l�bS,���(zg�H�Z�H)���g��=�H0Y?�k��g737@���R�S{�_>x�����|B��8P4Q<h�F��$�[W��H�Ɠ��G=&մ��׵ةUJ��烃Ç���?���m�FS���o0�ϓ��G�=��K��%��7��
�۹ށۋ^>��}A|&2G��7�F����XH�3����۷o�4�F��̍�V��nC�ݹs,��J&v�A�A% =L0����!t�q���¹ޱFq]�g�e���2��>bJ�<u}FL�YT�.�<��U�T(�0s3�0�a[(���O�lܮ�h�x�z�?��S{���KZ�k��FS1TT~d��&K�c�R��F�>I$���ҍ�fEu�ԏ������A�$����'s��	"���!J�+*f%h��Z��a�RMl�(�!�șj�{��¾��[�ii>�X5�#8����{�Nu�����)Cz�H;W"2+�Oؠ4����(��6�}܎Q�f{ƛ�C$��|�"�\���r1��w���ŋ�5�\���i�ʊ�D�v~!�����u���v �A�nNi1(�G�)��Q�ؐ9�g�QK�k�UeQ�%T���L��DuAUY>u]�K��gɔ����$d�]�e-��A`�2�ɐGn������cv��u��F&���Ň>6��$d	��yw:w*|�������!���������o�͟ɗ�,���he-�i��+|���=�ח�~%��������~��H��cr�O�\�H���2����ǲ_���Cg��ͫ�Pq���4FA%wO���|��3�D@�3
�J� g]�������h�g�g������Q�V�"�Y���IQ�W��|�< ���v:��1$J�?��{�����Ry|�ىZT�����G����b�'_���?��Ͽ���b-��m<|#�b:�H��)Ǧ/���]2cޞ]s������%u�}2>�kô�ڬz8����YdT�o�Ve\j�������B��x����m���ؐT���MA�ǡ��m=���[�����f՗n]�;�g�Q��5@ɤ��H
�N�Ȧm��T��Ćw��*GYH�N���z\���Fb:�xi��N]�+�8^"AK$r^{U��Gw�9��]�	no������mI�r;V����|�h2��I�F�:$��7v(c�J�MUL��8���mĖ�/>�J��11
Д�f�j��Yr͏r��ۍ(��<���
��#� �hu��c�Q�9�Jw{]���!#���8��zɨ)/w¶
*B��=���Xyz-�=�us#7A.�䵲�Z3��Q�I<N�?ʴ���GEX�(ChKaT���S�@@�P�E�!��:���cf�We<b�\c �kg	:%U�D��+�`D���)s�:��m�o[����vZ-�>�w*%�@��j���#˓Ѿ���J�� ӗpS��͊�Qb	�O�
�9d�!���v�9�!�c�m�Q�/_���f�K���_m2�1FѾ�|�}���G!�p���������7os�{�����W���:yo޼}���W_=��_6>�iC���WI3C�^���B��O�����Ȏ�4R��9�=�,��C�����H+F5�T��5�|Oos�'��h4O���
:�|V�
Q����ٙ���]eʽodr졘�V��m��$�L]���`�3y��\"^��?����._�x��;��V"%#�ԃ����s5�*�����MϾ���S?9�g%l�%�Á���Ae��'�Cq^!t���t
M�ܴ�d�/L���OR�/݀���˷o�-�S�fV�b ����:��O�BN�O�;K�.#�+S�95zb
\ `LA���zG��f�`ɲ�!��� �.���pa
��"o���~6�\
e���5d�d�1���ޙz
����Y饠�j;�,&]�/h��W�Y�G1��:����3L�ڬ�F��h�x>i#%�ի˭���0.�57�/��眹!�;���Q�F�E�%���,�@�����=fߙ��Z
A�l	E�l`��ͽ�>M���;�f��ͬ�n� :fx�fE,���}MS�6BbO�8=�8��ރ\m>��iw�x��`��Ԟ��8���{���1�+uc���K���!/DuK-�<}K�ֿ��I|�~�>�0x%�M[ܲ��9��Kn��MFn�Y	�,��E���t]!�쒶ra�����=[���Ms��l�����&S=���#�a	�F��-�8�����'s����1���}w�X�]���q&/�>��C-�X�8�4qY���0��(f,�3-j���� bv�������θ��ǁ��K�3�g� 3˛�o3R�z��(��dg6o|KԞE�,!�
�jΞv<�a_��B�{4"�:�o�>��H;��v?��-�{��}�=��-Q�]�4
��4 �+���e]�@.��#�n �ě�S�&L�k�q�b{�i��2<l����-�[Qܳ��端��w�)�%��&�W�k�O�붛�(��v����Φ$]N�+�}_��F@7�Ի&>�qH�������E&*�U�c�P�������M-�-/؋�x�=����M 1H�SR�Ȋ;��6��k��[^5�~P�I��٥���:��y��(�b�v�Ϫ4M��<��HV*��1���3k�&��F�%ݘ����r�ظ�XB	5�)�I��l�I"n)��;�tYx�,l�!�,*����Б�Ҷh�����|���<i?Rٯ6V'B!�j�����[�ǘ0���o,>�u���O1�+�71�?�ګ�Z3��8O�z��U�%��H�o�������ۛ����L�?{�
�&�(Y-��p<q�^�6p��f�-��팉ʃ���� V"o�,�h���"��x2W����N�M$��(1��m��#�6�VK���c��f�}��;��\�]�a.>��	��d6��T�E3�K�؞ c+����q�q�T&��&}k@���L�]aҾ[�i=�u�ɏ?����>x��A:գ�CN�./.�"eER�ۃ��
ì˧Ͼ�Y^��|�͓�����o.���r�eG'0�i�Ī�q@���ѣG���&�m�p�%$���8}�i���f��YF����j̉ؗ+�C�w�^_\�;m����z2Őz���x��Ջ�d�l��$ӫ����>���u̷n@π�|�D�w����I$���������go�I�?��?!+b���b�޸���=*<�!�/�XL�.L G1r^ML�?���jM�W�7��l<���HF��l7n�c�������v��HQ�ۼz�\݌�(	�$�/߾�/��?/s�1L���S�ʂ��fyqaJ���8�	���b��vc�!���&0�T��N�X����a�SOT$:��Ms�O�A(��f���)��j�5�|E��q4g,LZ�w8n�SK�TuǨ��r�>UQ�E�3����)�!k{.����o���d	8f-"d$�'��{[>ޕ(j��Q�f�͚��|:
Ď�=��&���h�w�FC�!�&&I*�F/��zf�\1�o�ۘ�>::0�GB�.��]��b:XNRಬ7��j��Tz�"�F���*v"M��@2����@mS���׿*s'y�r�r�+��HP�Q
���R�t���!��kh���M�?�����8 !��K��Wju�s�!Z�Ϭ2���޳6� m)���	I��Ը�HR������fC�����Ә�"ˢ2�M'�@:��a��-�d2���R��O��@�0����?ܰ���C�}��zW��R]���?~l�
k����WBy.x�d��n����QNV�$���o�+a\6��t����o��n6Sc��P����v3d�c��d/A���r,m���j���3�I��p�;�>}*b1��<=�C�x�O%�#e��h?��FҮ���@ei�WC�#�I��rqu��_��br�O'�Tܿ�����|Ի���Z�N9���J��d��LƐxiA��;���v�=9���~Z1���o��$��G"�f_�����t��Z�7�Աu1�7�-;�	�/c�&�<h�uc�� ޡ�'��!���|�$�;w�O���(4L����/i�U�I[�f,�1��u���M��W��� ��l8d��F��&Q�Fя�t�jw�$�������=_i
��1��K�*�[S���$��@L%R�ɟ]�ٳgu�㙏U��<ؐ���x�����i_;i��&���wZ������}wU#��4|P?��G����믿���K�j�F��� �\;Bx��I��t�����ЗO:*1�67v8�0T/@��s<�Eu�����vp
�=����N+S)+��x�P�a�����G�%��&�7�c�F����� ����԰����Q�+4�7R
�;2DG ��O ϣQ��}
o�FUv�Aw�|�R.��`!7�o\U�'����\�ھhH��wӞC
�-w����϶�6ȑe)���N�7���8)㣜,�MG>0�ґ�ʜ��9R�ktlek1�.�(�͍��lH�G�\(�>�!yBg�ob~�O׆M��9
�е�_�~��gV�[H�� pA��%��:R�����K*ߪV�U�!��D�e{ي�//'���_C��vv�����D�W���������s�r�j��a"	O9��"��H�5���{?z�Ͷ�������a{���3JЎ��o��Nu��� �\Q
�9�6W�Ӷ�`�ƈ�A尞��`����s�cNm��xa�D��N&��@�#�C�߃��m��ΤY{?Z.�'�������}p;mF��]EmHt����`��T<o�@^�]�K�'d�wI�nZ��b�i�����_�4���l�>IE�pd���$&d�޶��t"�4��(��˕}ER�7��>���sEB�� }@��&V�ҺS�
��	8׊i1�)�#Stz�W�ވ�e@�)��zz���7��0�B�-�>35�:��/6���ns��S�Z��)9��R}۴Q �^o}X	�"a�z_�g~?zܴY}�՛`t�s��x�,2Dz#���nk�ܬ�}i�kd)�c��>_�n�n߼yC�h���`C%]	G����pj��!�Cdv%�ҮGH���X�Z>>>���l+��mqM���ya4|K��azӌ��`���m[���:$��`���e�"��8�����8��.� �ʼI����d��7<5�*�����z��#O\�@�X���b����97=�Aa�>Q'��&�Z_�^$b�j��bl.A�A�)���I`�_�y�Qڛ�7lS�C //�]zx����2ʊd7�m41�:GK;ޒku̞���X�6baʔ�6�l�y���|�G���#�{��+�[lQ��h��z��N�����O���_��!��t�j2��tiE�2���(/��,�HͩR��18=��g��?���9�M��m��*�W� \���	F�} �[���[�h[L[�������w1�4"!i�����p�y���Of��o���<�$E�d9�&�z���ߘ��OǄ!?�я����%=���W�{��+��m���fP�ȎY�� \�f�!�6��b�|�/~���'�_�1���5a�!�ps\dI�Z�u��m�ׯ_���|e���Wg��Db�����9�W��w6OH���5��A�v=����q�؍��z���rx"y�s��[�@ d�R1#��w���W8�$��:u��l��[�Ǯ%t�,6�����GS
���+9]L��O�6�h���<qÈ;�#[Yme许����-��}0K��d˴KJR����S�9���9�[�f1�!��r=X�W%���RdP�F«�P��� ��>�_��	Y�����A�k�'l��a.k(�e�DE�3&+�C��R?�C%�0�x�Uh@��+�-t��'.l���s)49��5yV��d4�����)oc�{���~��)ϝj`���38���t���X5U��Vx;X��3A�ۿ�4F�?�̧,�I��\��hbI'��,軚4j��G��,fs�S5���[���==�]�
�՝h�N�^c���d��l�M>:�П��Z�0��'?�o�{-#�5\�U��I��V��)8J�}�T�=��m�9�Q�&��V#!p�$�+��:��g"8r�3�����m�{E4�y���A,��+�y��~� :Q�ep� �<��-�V��$P7��m;�t�Wu�v7���Zn@���3w���A��
���a��(��M��D�㸻=bND�y�����_r_�_�Aè]�6]J-Z�቞�����^�ձ�5;�`jD�gMS�0y���Ý�Nu��/_v{(Nf�bQ��������E���sY)��@-�$0%z1tȆE�oW��8M�=�~�lx�n��E�!��G�\]�׍)c�L����@|��m�+9�'�ڞc(M�#OJc��zy�4��������ݟ���o��o�jÎ�,f��]����������*�)2$���lQ� �cb^���7�awy����������A��s��D,�u���7��!����N�Mj=I*���N{�������&��v����������k���a�I������2V��szy��ITbbcK�ڇuH��b֦��d�.tV��;İ&���)�1D~���E<i	�=rJ����5j<�=&��v�2�>��=b5G��=�v��Y�gv�Э�)�;�,�I*��@�4�^�'�Č���H�M�W�ˣ�;2�́黎�m� ��l�.춻���]��zW�&���cd����ڎ�:w�^�6l���u��]l67�f#fW�kԠ�
F�rg�c��GCNM]��`�
V�\�A�m�h�5	f�E㖚���(����(h3;���)�>�L��Ma�ӱ�iv"�lwU]̢1q�d�Eq��5���0�+N)-�ۍ�����]@��6Gc�|�y"�\�GI�AR&�U�4b8�L�4�;�����8�-2�H ش!1�0.�h�V��$z�4�$G�zc:�tH�d�V0gM]�Ao�I7�1�a�M���R��ݶU^��`������i^�hCY�{���_�z���r��f�\����C�F����n}c�K�X\\\1�s;�b�f��Ij:�bb�r<M&�פ��F��d6Og/߾����qޗ�ؓ�1�ؑ������`k�!��Q�MFUS�z	�:�L5���M�mv�f� �~Fȕ��#4sU���d}�7�����;�_�x6#PH��o�ooT��۴nI��&��9���<��g�tK���Lgc�m�w� �W����x5sb��l���0���<+�jS �3'߄�AB�� ������]�w������ݭM���⦫W���[ 'U��x�U���d�Ɏ�ͺ*�����o��ͫ�|��ٛ�2��զ�nL����]_%�3�m��J�"r���w����{�c}\)J��kC��M� �DB �Q:z���L,
��]�@rp3Ǉ��<x0[�_|���Є�g(�va0O
��o�����l<M d�{�'~Xt=N�{w�"z�Z�#H��l}�Y�Ma�(Z`�;��.l���_����e��e��%:Һ�,����X��x�o�(�������xb?Oǳ�����-6e�ǳ&j�hT6�j�1��'�x�W[���P�(�G#���s��������d;��LL%�p���+�t`g0�@��]�m6L3{WTh�jmwe"}~}S�)��$J��K)g����e��X�`�[�f�#�+������=l��$m�`��D���j�mU��,��Qz|p�F����f��>m�c�&�N�� ������ ���:��gD�C��F>���i��ۘ�7ً#��U�:��q�IO�Ĕ9��s��L�As��#2�@�i	ƍ���q�^�\^���#ik���2������WƱ�)4��<�ã�d��We�a����#`�nZT�͛<��/�r7���6�1���|v۲�U�t��b͹@������I/9h��B$s��� ��1�f9M(�?O���DE��l<w�����#�W��(6���W�٨m�0-�d���@� ��#��M��{;=:Z��_?}�Ȝ��W���8i�m�&;K�R����,��À��|�.(j�뛳�/��~]c�N/�Z9os�j�����>{zr�}�i��w��tҴU�%}8�|��Ӟ:	>���+-(�O�-��M�쿓�&���@�P"ˣ��耕���f�*�e�fl�Iɢ��Z���'ׇf���7��b���D}O���`n�'������X��hZ�M�>���Ҏ�Y�#�g���ӻ'e����_n�͗_��f�Ҥ׼�`uU7ˊ�$QHv�F��|�E���\VS�P�¾��-�KRx��{=�`z}�|��i[�"c1�8�A�����7o�0弩��08�A|vmJ����Hwq����ӪXd��E9[�vMؚ/i�x�8}{��R��q���17y�Q���!�`~T߄�Egm�*߶�(����sS� �3�����j�s�~H�d�3�8�ͦ�17��!��)Ѩib�{�}ժ%�l����CL�~��cy�
.L����M�4m�'����y�7�猒c�]av��&8v�)x��g	����Ҋ�I(3���ly�1��\r�@ �hZ2g�ȶ�Vl9��Ҿ)I�WۢFg��������^<cʨ�햻BP��Ɯ(%��Bgb[�H�k�c�B�#��gG�G�ӃC��Bn(�ò�\a��u��M��  ��IDATfGg�w����4��P�ЌM9���*������!9��ǩ����,,�G��6�b�Z܇h�9s���
�l=\k��W/_��M�"��\㊂��.f�6`�^��Ng몶�1?ݼ����lb.�nW�SX�a��(D]�nwi>���jaN]I��\�{S9�H9��$�H�o\�
�`/n*M�#��e
H�~郆�d��Ev��xHF4�����Ԇ���{��(Nͻ��ۙ�rrt��b��ׯ_�y�����#iƎEs�l�� ��\��4iAh�i:9�{ss�ab�-�-!���ɽ��t�;��'YMZ��o�ڑ�8�c��R��*m	�:�#��a��޾=G'�Qjn0�3����N�\�V-4��|�6���C��C&$r̉z}*��)�wp��2�a��(K�a<bS�Rxv�M&Y�a���s��HOT��>� |� ��9h͟)�MfC5TDYf�uT-����3Z�L1 �O�R�٬̓Y���㉉�n�����,�[������9,� W���o�Y_i�C��o�0��i2g��Ef������a#������,���|W[��<��z��7�<{�̴����z����
͐��9ƙ���s�h�����~��B�l���G&x�P���/�x��a܆��N��sL�_��
Ji���E�>�s4S�Fψ��Z����B���3�Ij
v|p�/�F��B����Fe��C�����y�ܼ�LD�ETZ����8sT27�D��`�50D��zi��G}d�͢�h��C�=���F��� Hf�4�������I�"�t��5m�;���3̓Xt�7�{_��r�����Fa��nY�RE9��Î��իW����zG;�߇��-�=�U䆝�V����t�
$=� ��vDi���/������omoFc�
�f^`ABzS(��[\���Z��b'2;�rj��8�� ��0�s�8���Җ�G����O4�ݾP�<�O"v�J�i���fi�]܎����S��!���B9[*�@@��W��~�s�(dn��]��zC�&���:lD�9�0���rp`����M��H�d�嚓ɜ(5�(U��t��rʡ��������;�]X�T)�嬆�z�o���b$�����\9�0�	wp*�F���uxO��X��Ԫ?���
lD���xC�DNǲ��8�7���Cr�0 �&�����`E�J�5�F�9ɔ�o@����4	T��؏VY�.W/�W�Wi*^'���OX��.�w��R�ĹO�c>�B��*���DJ6����f*ww��6d�i9���z���̊�I���u�4*�g��r3a^Ȕ�Đ`�k?ۛIݰ��7���?����TVi�eå�D"
8[I��T�ۀ�3e�
�+�i�F]VBdr*�:f�;߃��T���Լ> �Ƥ�K�IĂ7��:�j�2�Z 6IQ0 L��q?�^�Dx����ŕ�����kA& |{�>�y%�+%���H%��{����ёY�����ѩ��5�W�<
C&@�>"�6��H����m�L� �K\�	���\����B�t�{�6�ߔ��p�����&��T=�r�f�,�]�[�g ����x]Ͱ��c��o�U��ݛ�#� {�.�0pm#����H�~-�� �\&��-�-��?�SSn��v�k���H�mU߻��Q#��%91��~��ln�ux���W��lv��^� B��m5�ڍ-��&�C��[��nS݂絯�k�9:<==�e��~��w�<��U�v�WH\�hsP5Bb��ѳ8�~"�p+���r$��y�Қ����*�2j����^�n�4.�Ý�5<��"M�>X({||x�Z
���h�&
s���S�y�^�CO@� io��ڷ�CI�Ո�������
R�%'a��j	�-ֆ$�|!@�EHǚ�lg���y/ҷ!�_Y`/���*�^�`@!��ց,��x�St���]�+���v0;�&�f��ݻg���̧&�]S�e�Ʈpq��_	���6:�[����I��#����I4(,̳��h�l�W����̗�5�_�@C���u�������"W��t�浭̛7g!YƩ�C�|�$��?�������4gw�#[i[9�� ��zL�'��֟�H	2�	%�a�i@����(q�`>�*}���o�����e&[����xP�f��A��YtT���l�X�BO�"NO!���VD�5��,1g״C�	�&�-���d���V�X��ET�l��$�7�QbN��[�O$5���kj����mhvD��<�\�)9G��Шkk9ñͩ��~����ɠY+ie�;��������K�}�")w$�[(%R��C�y$ls�4/Z�ܖ�'zS����sn8@�7IV�#Ԟ9�Ĵ�k�dL��/��^V�dL�jv���݄���54�0�%��U�=�"�$> 6B?;�.h[���ڮ��a���4��'U6�OdȄ��)����"EÎ�R�@�R�$pUA�!"�y�����7z�Q๳B�b�h�U����V��zn3zS�pz}yekrŜ�|Ժ�t�x'��8�R�MI�7e�v�����%`1iD�;�k�,X(����O���^�o�T�J_��ѥ�z��C5��Gbo�-ק�%�X�$k]��]�3@+�'�9S��۔��P��W|��C�S�P�-��v��}��O��'Oz���Mcg*$@O#z��b1w�:gsa���uS���9��f�)ҿ��&1g>�9~Χ�;Q3�2 jgT�iM�B�D�-���ΰ���
r�Z]c��fXR	ؘ��hC��.��6JZN�� kU�P�ioC�]�F�Ð�qN4j%f��Xm鲹R2R;�e�QBC��Y�0�������� � ���h4!��T����＾������{@�j�>�o���Q받�v�ݹJ{�7o�l�Ҧ���pwԥ.U��@�ͨBS��;Z![���x�D��26k2C����g&�Zm�(�4��~e���PP=� �>���֕z�����8�q�C�@c�z�ރ���b�ԍ�`���X����#0������]u}�=���ъ��~hK�H��	 k�\�IZ���:�+��;n�,�k�&6ە�����1�ΩU;��2�`D�)� R���-���^~�nߟp�U���u t���)?#�{O�������
����]���e�<�!��N۶���9~ك�`#�U�C�R�<i���Up^	������]@���@7�݌}j�Q�r
�#ȩ�3�]�nD,�سbA#�|�Üǝ|;isn\��6P�C9���f�����28�� 3+�C�7o�^�m(N�����b��M��p�-__�M�y�fS�N��������.//�va�ȲqS8���0�a�����
5=��,�=�8˓0j%` Y�c昳��|ʑ$����ve!'I_�s��Ki�|���"���o�F��(Ly@�	JHp���'9����|�3��*�7�8��$Fl���w��YpP�A����y�*���:��"��%-���*=�I%�l�DE�.'Z�d��]A�d���ߩL-?��g��5a���Im;���.��3��3.�l��WD���[�[O�#d��y~�!k��a��lǝ�֔6}�E�4g+��^S��}k�s'
9�;�α�$�y�D"��m���)� ��}{sy��1�,��Q����vW宜O��b�p�P)db����9���N����8bR�3��y�.����*[��RJ��%�
�a�S�.���j�r|�! ���i�2X�6CJKZ��/��e�ى3���b��@��z3�E�&K�ޣG�2��򡁎S5bO�=��� B��L��_���h&�5���E�^�p<_{�).�5�io��P㡯�1���nI��f1
]�.�x���)���<���ǈ�Fv&K���*�#eq���&3X�.�l/˸�{���9��Z���Isʾ]oʾ���	�H��8��0ڦ��'�C �ayfʾ��4�<���8��s8�:2���S�&7�]�o�y�ͭ����<�>�����j�YU�KH;En�!�x:0T�?��N��'�y��"��׫�i]�~;�@���Ȯmq�vSlF
9㸴��������{2��r���U�f���Ę�J��e�|�1�1�r�nd�i��t�cp���۬$�7,l�S����ߵ��{{��M' Owq25�����8:���W$ʚ�;_���ځ)�+�D8����/׫�����e���۴-w��fmw�X�\-�۝�}\��n�nŖ����n�s�1�3��;}@�b�hJ�I.��YM@�����Ŝ&YrvD[�۫3��iȻ�6�>nk��*�Fc{)M�8<�[++�����ݽ��ݶVDG�������_===y���ݛ����-�yS/ޞ۷��8��Вú�W #k8�B��s��q�ȋ�ʗ��ho��\�eM�����ٺ�|n�o�k6���	<F�@�؞��?�����?����>��g�}�Ï>����/ϯ���ʚ�P/l����L�B�0gyjO��ne�=Y/�׶��Do�ߐ��ʲ��%�;�L1)���-�W/A�q�-�-�I�ۮj߮��ۯ��o�fyyA
��(�9��d���)�γ�D���58<'�m�
wȃUi2��)&)����T�3G���B��gH<h �z�o!�Q�Ԡ�a�2�uY��kb���� x��~�r�3Y*J 귻���^nPx90Q��2����t޲��w��H�)��r����q�)#�#9��Ͳ,H$�7���%�̜N��P?P�\p!�tGm�l�5 j2�9Jn6�.w�d��˹qjZtʣ�>}|��x�z���Q	��h"���BcUq
FmpZ�C4P��;���]�\���%3��ߦ�q[=m�������	�\���Ԕ�B�eM���S�zlͰx*����=F����ɶ�;A;^GN.E.dv�#�I��R�
�G"��<h��3�pF�	>���F���U1�L�.�qk�/�ϱ|$�
d�Q^�oB?3ᓉ�(��2a+c�!E���'uN϶�ď����Iz�'ƉJ��5�y]�~of�n�K��fz?�
�µ�8�Ҥ5ۅ<~�j^���7��b��6���\�[L��;�Ё�z��f9����r�IG.T�ϑe��Ge��>!lI�+8"�z�9�ն2U�=�=�C�p�]�h@z\�Ţ����'�s�����b5hȓ�w�"j�򬝀�bf12�m�O��"lG�;���p98���n;Wy�׆��?}P����Q�:!�\��*:��zHуR�-� 
�z"9O8(�o�
��¹kK��)��6�Woj��ݻwOI��C�eq�`ߵ3c��ޤ�w�8ܝ0�n�^{���;�!���,��k� �#�)��n���ǒ~a������#�"9˩��ȣX�����e����ж����gϞ�_�����0��<բ�d4��|�<x ����H�3����
�gEo��A��>�w���|�~�E��!������~��ٙZ#�l��׷廭�jUs�� �˧O��b��/i�o1�W_}e����$&.�3�#�j
��B2�W�Ra����1�������P�#.SпC&(�j_�%+�o~��Iý�bM�i�Z	��U�~�m�^@/7(ʙ+f�d��ݒ�In��w�c�ʳ���ΞL��!�=�J�+����	�$���;O %R�!���(����Q�l�	��]�,�ۥ޼~�d���5�I�-eooK�LP�əNņ�ّ�&#|�wʭr��Ȕ����B���^`\.�ܒ%#$��u����<�4bՎ���BVPU8���K�r?Ӛx�4Y��(�L�4ٮ ��k�8��+Hj1�,���`	�Y�4�\5��̃�P}�P���(�CD�"7��W�b{��7�,�Y,$�P"h*��)��
��g�� '���.��m�S��򠤿<ֺF��4�h��E�$�z� 8��,����/V�\�D�BG���4+`t2Y<1�ͱ�1aM��$S�e������)5�w�w}槤9�����«%B>r�n9,HW�2Y�2�As��y��jPڠk�!ϫ�S�1�$�C�l����(4�k�a��3I�ٻnB7]�,������H@��턘ʹ"
��h�X���m�4�^��):ly�g��H�U��#�(�	#�M��Z�"Q�F��f�x{�t�*�D�{���u$��wCC���6�J:���\�;D�Atl+�zR���s��A!p��S��	�d0�2s�h��c&���(�{q�� ��r�� ���'H�����L�b�:�Ev���р�;���cGX)e2�K�_V���Ǟ��=99�`���)є#�����4U �1�@��(�С@΅��C#C�W_球D�����T�{0�
,;=7�Yvsவh|���e$�i#�Q�G����\�����%j]���l?�k�S\�)��-��\��LSjׅ��\�ȳ�|�P���s�,������RcOW4�~�war����;��y�E�#dRa�*&`�m�)��be���a�y�@�vC1Ϥ6�鶀]`��jr��)B��JD���dk������S�v��Ӣ�Ð<��X�K�M��'�G�H6q�zȰ�Đ���	.�`���x��%*L�Lߋ�m��%��Xh>�p���f��E���9���C���\�~R���g�E}R����w	�������鉅4/^>�P�����R�;��瀩�P�i}�� ~,ǈu�_[[[F�1�r�&7"Y�v*�.��O/X�RT�R<v'8�I���O>��<��_��_�_\�F �%��g��=�lϿ	`a���������}��a`9��.��Ev�ޯ���W��>-)|�QN���*���~��]nK�P���Q���������ze��ᇏMK��_�ߺ���4eI,�kh6��uui/�:�$
Z=t�(��q��[�Ls��Lٚ<��!0k�s�?��&�������5>��<�< ���^��~\��r�|r�.8��X>�؏P˛L�@����HK�N�`5���{�˚Ug�T,�ZH�)����<CS[U#N	Y��<^A�����@p���-����c��m�H5:��i�^ަX��c�����/_���=?S� ^�"��C�c7�H�n�b� Np~:���FG[���y8,i�Vd��g� ��%�4�#��j\k��q;"�d�Ne���b�7���c�N܄=�֝c�FZ�BT;�=��?��U�DJ�V��ۂ�n��j54]���1�����B�X�R���A8����d��R��͖�}#��W쫼�F�F�L�4�7�/3��Q�nj��.J�IS.F�nr��&�	h���W�8:?oʼM;�*/�	ٔ���@�E����/[O@�#co�����,Q>TJ~P�5f���4����K����K�8�؂�B�)�^#�ݴ�����+:ǋ='�®��q�mA�Ȩ��f�>�L��{v�խ��{��7)*��I|/l`��2%�B�K䫘6�K���[SZO�nA��ӧ�
:3$ݤ�U%�DT ��=P����g�}f�\��Bq�|���Z;
/���ݷ~��}���x�p/8���W�d�sHV�_�>}��ŋ�kia��A����$��93�W����I��)���S���:��h�)��o7�"��jz���lS�=jN���g=/ڛ��}�+��(����u1Nk1*�,���iTB���Ճ����������M]������α��P�I���˰�
v�B`{���/1��g?������vq���Ů�R�6[̃P
����		,����R�I��������̓Q⽐����>��̱��<�!�7$C��'؛#��G+8��n:QB^$~�oGJ�О������4��j�.�7�PHV�F
ڕ+��̳���v������A��Ͽ�ke�V�~V@�K���)k2�R���K�j�t��+>�7�;�0��-'6�0|qΠyt}brJ�Jv�p��mk�T����8�lO��>�l���E�T6f��R��S�0g���ƄD�>�KxJ;��$����S�iը��\����r�QB�٥�<ۈ�2r����~5<��C�g�Sl;d�6������狩YF>=8#��&!�����	��.N�J7u�����f��ܕ�WJ[Yk�=�vJ����\E��2�Q�	���4�(���j��#�ad������0P��	��*Ho8Rۅ�Jj������>ifm�Mi�,*e!���ΝD���2������I���ўp��6��p�o��iGL!�[�����5���:>�����4cZ�)�ӄ�؁5�ԍ���@�=�#q�oc�b���B%��z4�1�_p]!U{�8J�\j��	����jE��U���lo^̧������ۮ��ؕd�8��=�.�|}�N�#�c:�͘\�v��7x�M!�EEB�h1] mԷYlX�>��in=��?SD�US7�zF�[���!�=.T? �c��H�noj��M:
���J�?�
d�6����!�,*�v���� s`FR�'J�E�N������:���4Y'B0��:�N���B<���� I����h��wyu��@�I����b�4�����=��C�i���;�c�o6#�^�,�����ٙ��h>2�����X�|�W�w�����slV�u�诸�[�""���r�!�r�\h"Q�7e�\�4��ֲP=���.��mX4�wQ�`Ol%���A�k(�ҝ����۱0}0��z��L���w��`EY��i;7���;�!$����uˉ�5��֜�Л�ڶ(~6ɤ�Y���#�����v�q�`�4��z�"I�a@N�`8���-L��Qm.lQF���x��yC�%I�P��沩�RmA;VA:���Q�F�k�"�5�î�Ewc^��6Ѹ�E�}�Va&��\3G�w�����ERf��/ޞ�_�Y2�󦗢&���f;�U�k��t���?��~�`e��ћ�g1'���Eb���@qZ���,
��r�j�Z�+��	IBa�l7��,�:�[%#:_h��1�	h�Hш�͊��!�C�HU\jsQ�;�J�������mM�M]��5�������V�`$&s!���ޮ7}Ѝ��s�g�ƈ�"W�}3
GM���d���C�>������SF���nqT�U��zUͦ��U�Z"'GY�+��N�H����ޒ�����Z��t/�r�����W%:�l�_>r
�|lV���6�$��@��<'�S�&y�G}�ۯ�b1��]�m0���jC�������0�1��������g�Wc>��&M$�$��ȦH!v�gw�'��{��!������t4>�L��k�r:��k��W_�����3vLБ�$�����D���'�t��vp$��Q�Qj&�N��ӽ��;W)gYt'*sE����u�Xz�Γ��GM8O�`�r���{��h}��ϟ?��������5.k���%�7h��G#{І�}�4c�A�	�y���`1�0^\(��_dj�,f�x~E?->
U����������-���Y�,�eG�ܠ�	�B��$z������ׯw;f���w����U�B��3I�����9���RIy���_]����x��J��B:�S�Dd� �T��78,AL4���)�^�x��--� ��"P�9��W��&vc�n����l$�	��ł�h�9�sJ+@�Zm��c�W�jY,C�������q�oN(o��n�����*���t�۬�.�Q-�L��a��"��d�]�Y5 ۘL�W�Y�6�3Ow�`��a	P0x���XEEŃ��ʴR���zq1��!�r�`��Byv-�%s[�vĮ|8S�^Xo�0Fgn�:�2b�?	�8��x��^"7z[�v
B�&�@M��Vb�"G�����tբ�2;#_PY cK�/�����
��B~ ��U
Z�#��\��,���mm�������Of�r�[�a�Jd��N�ԕA�X�A�魊�g�V�>���+f	�
�ͨ��ҔUs���X�{ΣT��Ɉ�L͹�hl�<Q^0���ws�����U���(HlX��X~wΡ��#?�M5ra�����@=�*�1)	+��NNN���1�-~��dla^���t��N�k
������^�|�������z��ur�Y��7ˇ<F� �R�Us��7��׌�X5$g����Py�!��N*0ڛ�N0{ۊ�1���Dcl����gO��x�B����������C⚨_PW�&g$�ʐ�Ls�N�j��۷�Ϫָ��Y,l�i/u��*?3�K�t�Z���k8d�~�9q�6$���T�_��Y-~"�ݙ�������{����>}[נ:F�&��6oh4�TU�kC�6v4y�q�~3#�ԁ���ؚfϦ#;]�� J`�G|
I$�-���ϲm��t5�����M88��y���<����7>h�o���W�!�7w��$,�\6r����۶�}��I�I� Z���>��w2%̂�p��l8��V�l�2�����W���$�+d�u�oH"�w}o .h;�u�DJU dWB7N��ݠ�D@��Hf���^t��%S<2��X]�n�u��в$U����n
1C���2mY��߿���$V-3��|)��:鸒]Ns�qh����'W�\R	R�]nwU��������䩃�ԩ^��������ԙ�ς��=������G�iDy�+��n'���iƮ�s��qB�8��^��J�*���D�8��F�D3��q;��Ȩ�¾q�U����al���h����]��C�1�0J��u�<�[;�&�p��SoƼ�T�]`d�"���0�<���?fb������T�qer<�j�U��;�v`ľ�߮VR�5����k�BO��Ǥ�����ꖕTk�{�UB�� �L��KB��:��k11:�oZ��!��z��tː�3�Ǟ�������(���Y����i�HׂI[�i�k�`mv�xL%�b'WiPA� �Pd��]�S���,bm1]ﺤ�#�hۨs�'u#;(\�gC�9e>����H�@��W�a���F�<�=���1�;��&�l�"�Jr�8JM�װ�4��0Q��r�C=!Ǎ�V��5Ţ%��.u�t��q3��S�%�3y�D;��j@���"Ǉ���#CH�1ḳ�J���P��qu�\Ȭ�l�vҟ�|fα��Bm�]$�ik
Ӭ0u�	 �ef�}!1����z��%��C�4P	�0�`���dCF�j	��|��l�V��vd�-�	M�"v���q�G�	}Ĉ �u����V`7��\�A,:*%O�e�@Ñ�؛08��T>"�#��N�_���ݚ��*v݊g��&��rZj�6en����Œ�zŐ���
��<-2��;��~,5OG�����M�eǕ�ӡ#eei��@w� �i�O���]��H3�H[3���`��$��Uuu�T�"t<�����e6�aXYYVVf�{���~���q�Ʈ� �x�b�+��Mpk�)��ӧ��P�u[7��N��"o}�u\������������ѧ��Ck�:�?
l&r��ֹ��!Gb{�P�b��4�U�N�`��M�F�<��6�#�Ox'�~\�H�*QD��wDaoG��iά{�����ͱ��^兪�{�,q>e��]�6�TZU5t��q���[H���jNIf��L��H~6rM^N�2��F^0N��)�N���zG�䮴=��˗�����8{��5s�VŴn�G����+;,��������׾[��.�+�f�j�L���\,@�ٚ����w��پ��_������?>~�X]�����nM\N�]U8������?nG�d{{S�>J��[Qso0���haL|��H6h~�IO���^{Uȱ�bk#��Z���m@�������S���^��a��x=n#-����oݸy���ܻw/(�����$ę4���ϳ.�
q�=��U���M8�����̯���;�M.
K7��ȭ�:�E7�Ʊ�/X�**~Ѓ$����d�/�)9b����� ��Ζ�f4Z�o�6��R�Y�b�7�g++�����1�z"����g񄜀ک���A�Oc��}S�(
����Y�#%Y��J)<:J`��*��m��c�`��(�nB ?��������2JU˧[Y%�|:�n�M�Ue��*1��H�_S3�r����:�ς�ڧ��vT1��V����M9ws?sz|��	D�DHR�1ŗsM7�,����?)i������1��6P���LxmlE��A{�:eW���.M���,��u�Xq��)�Gqb��4JqBt�^)�X��;�7h-Z.*�,rJ <���
3�wP��= G���.\Z�*]3�����<8�D��ݣ�̲�u�`΃�U��T�.�WU�������O`,?;��G��ji2�H5��^�T�@ݠ��
����e��
�?�'G5T�M��F��L��Y�'��|U�^ׯ��Wɀ�.����S�[}O�@�w�[��$U̥����f��hd����M�㰶�-�E�I|I]'/q���za7j�R|w�i��|w��Q��?���F�x��Εm��Ǫ�L��j?���g/^���rM�82X���-DI�F(�>v�"�6Tl�|���`����'T<b��^N0�g,�M�+��b�i��W�"г�p7�:��on�?��߻��6h��>�T��k?a���s��O�H��a"���867��<],��	q�K�M��<�P����8�Y�Ah��pf�!3��Ga	�4���r�~�8|��9��ǯsl��Q��L���Q��O�J��?UW���#|�_ו�R�Gp�)�p�ji����k8��˩�������/�yf�-��9tL.#�Þ<y��,�Ģ��|�-c'�K�N/�[���P,_�'`Ԧ� �V��X��B�
)��<iq�kF�,�bK����	�^��GŁ=���-99>ƅl\�+�*P��j�[-Ͳ�=Z�ű��ճ�X���ܝ��[�n)H��1Z[��9V2� \mJj�z���g��3�W�K���h�nӃ�}*y-M3��h�UNy�e�����J�s��h�af�9��$�'E!kUZ�+�4s<�h�I�PiI��J.���t{��I^�bƫ]�.�Ų+29u��u1+XM�KNA��n�&�!y��13��q�&WK��2��<^K6��W��\�)C)n��F������^�_�p�����)"`�rR�h�t�Ɣbp͚]#�i�[`��0���B��OsЉr�3�R2N
,�>4j0;���#v@w{�YH�P�_�����Wq�'�|��~��a�\z=���V�ߥ��'�����^�a�e�	�m�i�1�[/�o��h%�	�Y2T|l�Q�܂�Y�0b���s&�xk�A�����I��4�����4���t�r7:����S3�M�رxj�_����o B�?����e��&�����O���I�����p*���M��5k�n4qQS4-�����(��h���� �dsk���|]�Q(�x�H頦���<���Q�H�b�#	����m)�W���Eua#Uu�z�/s�=��ذ��x�!P+4�~d���c�����>~��Cf�bq��e��4�vl�7��cKf5���Ռ��r�eM'3�#��H2៨P�;;	����@J[��a���D��`P;�xV �[�F�2�M�3M[��Y�!��P��u��%Q�ݲ���g�}��[J�ZY�gM=g�;�nq��`�����̫61��H�Bgg�la��9r�誖��� h"�ӎ�]9�T{:��Ѵ��7��?�������7����f�M�uY4qY�͌L3"�RW��)�x^a�*�i�g���8�kƋ@a�q�kG����*��¡,3Rv���WE-��X��Eq�eXr�q+��u0y����D�l.G�E4���%��p���}�[��}i�\�xg5S�]�+�>�6��}�JŽ<'��t���p����Q��;8Nʹ��rz�Ϻu�ƫ������	����������-�1:�>13�>�u	ʡ��C�w�F�0:뜳��ln[�u�{qO������k�����q"�Lgʽ|�̵�F�]���E�&�
NU����pW�v�^g�0���gc��_�[�z+]�RC��Ţ�z�5���~z||�5&;�hX�>~ζ�U�t���,̦����+W��f�����3�a������ݭ��sM]�Iȍ�јx�``2o��2��\��N2n�[p���ؙ㍭Iܤ��<���&�|r��ǟ޻G�E��5\e�^���n*���~��c�ݼy��������)egC��9���v�$��+�'��E�f�����)��F�Ϲ��,�,W�H�������D��"�eb��q��J��7o�g�&gJb��Pfߴ\k3-�/���ݳ�w�����Gq]Y��r}vz^������4���li?�	�xYb𕥝�^+ �Ä1����xL��U��Y���Aw8�_�F�+ �{�����M^޾�������ٳe�5V1'e�y]��*�R�B�f!wEo��Vh�@�B.�����
n�r5�#k�*�Mȹ���#g������<
�Ŵ�T�MeZ�0k�d�&�FT���U��e6{���+�<]�+w��]�|�����w�÷_���?~ G��ǃ�hC��Ϩ�Z�����a�6��;}R�qjbkS�-$t����2*��I��4��@��2VݱT#�vw�>�*6v�E��|�LQ#uAFZU �e�OQ�9������b����CL�(��
��h��M�y�:���i��'',4�\�{������H9���j
Le�ԭz^.q�&����J$Ѽ�U�~�C�&��.j�s��g�C��s�Yi�3�,ih�U�Jʃ��0���jܻ����D�
��ŸN����V���%�#�dww����7�z����O�nnݺ;�]aB@vœ/�§N�&#�l�~���fÞGjӘ�k7HR�C�l6D~ C�����STHuGacjZA-]ڍ��KF�ilDea����g\�=~�83}me0c���L�Å;�ڦ�̕+;�e%�tu��Ӹ{"�q�2a;Aܰ�767�
��Ӑ -��4����%f+|�&D�kasc�6�e��ݘ;)'v��}��f�|���B)=�XU&��f#��\G=QFX�\���o�1Ӿ���Ԫ�~�^��Е9��1LG�d�Nf���l�"7Gx���fω�Z�srt�/WpCw�܁G Ī�$�q&Iل�2���N���߮��&a3H��A\�2<���c�����}��	k�KJ����6�F��.�7u	N�ϔ�/i/֞�%���%�|]�iyzzj����f�A��ʰ�X��½+{���իW�~��d=��W�B�V�S�K�~E��_��9٣c��PW�lM��B�(�8�g�<~���No���(�#�Sax������[��rpu���U<���wL�%/m��(a������}Sl���hϧS�)��_~I5'=?g&Q	&q�xW�K���p��v5ڜ�Wv��Z^�V�����e��Oe�B�t��U�q�6���D,X��N�U�:�S�b�Δ�K���|�|UK���R�4�&8W��:�����R��ʨ��zE'Ղ�=-r~�%��ÁuZ�1��YS�mM��L��|�\C�D���P�"7�k.MV����z��w���o�����������Ó��Ʋbq|ΡL/�)�gIY�LB���5^}I>��_�1�����*fJ>Z5��� �mR3H���ڤ ��;��5�������u%b�퓵����[��V�X5y�pj %
 rf���: s�bIy C��ٮ���ڟU��|�P�<������	�vg}���Αʉco����������c�@0�M`�텕�/�B��@Ϛ�$
�r�j��8͂�a��:p�bM��*A����I���_��l�P͟�������k�H�/0���BH"�ʷ�G�ץ^�kV��^�G`c!\C��=�
AI�`\�J����WZ�^'Q�M��dA�8�<�����sR)Z*��j?�G�۷o�;���U�~�w�������Ek����r�x��������<��*�a�.i)�O��#�(7�>ߢ8.4/�����2�xqq��6��͋(�FI���Ъ������Ҙ<�t^���dK�f%+*���Mn͜��oX��H.��~��y����:���uG����gM�ϻU��r�R���.iM�6�>����"���Q�c8Nq69@ M���I�[f���}A�����v�ǐ����R�����W>�M��T���i��
����ͩd	.���%�c�x~�e���XY�����?z�o6�q^���R�V�[	��T[��d�A�j=߲�O�u+z �qE"�����������^	�e f�ٍ�%��π@6���Z���?�ͱ������#�����$J���J3;7�/3���!�e���I�v�'*�	9�)���{�8�ե1|�\8h�5!�C	>ZJ�%�Lc�E���Uy���%0�{�5����ub�#�+�+ӄ��f�QN�^:����7����k�|�ݫ;W�?}���ѣ՚?�볳��%5����;�BW��]UDT�IS���t~+S�4Y F8E��:�-��~,��.���`�'{��Y�y�"V(���4��(���������\�Zz%��}v�b��$�
e�`+�z��ϟ����M���~�mĨ����裏NO��go��a�pf!��k ��6�^�����e�c�=��[L�]-=5�
2�Ob���L:7h��}1/,�Wnae����q�A���>}L_��(ʚݾKfvV����\ >����{-�ٳg?�T��3�ll|ʯ~�vn���O�<�Q�g���Ob��a�������1���
2��k�ܢ�	B��2˘0�E.�ʔ���g'�G*OZ����2�6��N�.�z>x��t���n�4[c[�l��섗1�l�S�
K6�ߺ{��/����w��O���3Ϗ����Z56`Ѳx��6JM��G�[�Al1'�C������P���U��(jƩ/'gD8�3�fV�}	q�dFZn���nM'K���Ɠj�ٸ�S�;���VH��03.y�T�V�S�����5��8~7N������ۿ�%y���*(*z1P�NrٖtH��jt�-���8Eߑ�W�
a
p��<8�XLF���}X	+��K������"P*����p(/��M�QXQ��̤����f} R��+W� �Q.|͊��'���ˀ˳��)�:v�{�uzNP,�$��ܽ����{]ί�%��)��>���Жs�-�#���W�Bf���qC�У��P�q�^����涔������õ�rX>,o�pm�]��u�z�u�|iA�0d�[�)lܧ��ŋ��N��_�*d��uZb?9�c3*��$���S���訚P�T"���ĄmS�b��̲�6��i�)�4q���&Y�%�+�-�Q��N�3�Y�o��&9a9�˾����k¥���N�VA�u[��Ű,m1���s~����� @3�z��h̆�d��m�=l��xe�d���WT^%L�(�.��e0��ͪ]�D����d�X�F��Zd~�@웨2��,u��m>��/\pT;/����9��C�OO?��S`����88�0��:��\%b���Գ��+p9��`��J���K|thj�?��~�Gm\���Ћ��x`���� Jw�y!8��P}�r������?~�X�M�V�;�̓��q�ƻ�˄��c�����ovV�}9e{� Yp�(�����z�$�7^�;hDL5��f���aw>��]EI�se�.v����`�sғ�>�5k#~*�*(�m��n�M��B�	̺r�*�� ��ݿ{� ��I^J�#uE�ڵa�M{R�Kg;Ն!���VL�_��h��S�~��̝,�s�,.ot�/q���F�]���	�b��y�)H�f�S���˝>z��_�))����4#�[��"��mS�D�x�OE��0j.�:�г|����ՑV*p���b`�'�k�R՗�Ց����p�~��&-*�o"HsR��8$�ZiZ��������ȥ�e[ӐzcSn��1��Χ��'�Z�=5��1չTs-���������g�9�k��,�Ԅ �K8�����f#�a�x��g��_>=5�t6�%Y������9���wz�AbӚ�:������bU$t��ގ�.�ƚX��^_����oͻ�O�=������]*�n��I��٤t�e5��AO���p���\
��,������Ӣ��&8IdouC�pN=k,�>aԷ\���Yi:�p����t�,Ԩ�GW�RTi0�ˊʵs��0�M�( u8&�7�;s���S|�0H���±����L�!��;p)r��Y����v_;#m�wO�-g�Imһ&iVl�l�����寒n�/O���lQP����wY-�������t	�YeE�ͰV9U#	��1Ϻ��E�f�c���Y/���ir%�V���/e�b��JiQ��MH+�l[�+i�kU�)�����V@j�d77���~���re1�Nj|��ؚq�˗?�/W{-�/^ݖ&jIo�����7�q��Aü�7��s6I��T��!f�MV�dۆ.���];���(��E�3�0��M�[��;�,W�S��ʧr%m</IC*+aG�{-�r�p�����*�vMD�q9?��O�~�����G����BX�r�%Gui�:����At��s�#�ɭY���;�&'GR��v� �tz���g�.�xS�霴 c�&��	,[Zp����>�b��A���$"���	B,���|�\��$�'���OnS��S��?�����k_��6��������<�YC����w���s%!,-���3�yY��y����ܷ:�������i���&���],��D��Y7����=,��hL��ݎή�R�ĥ��=R� �i�a5[�uƙh��<��f� g,t�V�i�d����b�A� ��ʃ1���k�D�}��9~����p:��w��M��e�t'�9;"o����x��]8�$�ÏaU��ƹC�u�L��T�e�����K��1X��q�Т��80�y������X�[ݔl��"X׮���V��r���͋U�`c��O_��?hL�/��QP���o~�?�$ِ��8�'��-�������d:�؝/��`0_�Ǜ;x����W�>�(�D�t��C�K�W��DP0�fxFf<7���K
�/�;u�6 G0_���C�Je��͎�N�:��	$�yy|��F�qrrv~>�2���L�8H��l"8D4��G��׿�k�~�����C�M8`�W���g���!_>z��7ob����X�G���4[��ѕ�����5,�b`����3+�
I���ɚz�kH�Ʀ2V5X�����<s��"(�Dzq4��p��s���˂#/�ۊ�M��:�j[g���([�f���bK�5��GYs��������nm�d�E�ܹsg�\���cMg6Q���>z�^���`sH���ϲ�iH_���/���=y
H	}|x�E���w�vz�����ƾ��'4�v�w{l~�6O�E�re�7�ꪀ�<����9�0	��-H^)�?��9���Iu{��`лvm�� '��}뾬��k��)Է�s(��ݺ*���?7���E�'͜p;Mfsf(�B�+\��e�<MN�fī�c�����Ǫ-DVq9[Y�p���,�Ҧ��K%��L��w�R�Dq죙|%v �:��N�Y�>��M7��
��+S��լR��Z���z�w�:��:a^�|�����<x���YNĈu@��/q��#�tvvY���fЋ�z������$F��5�RG�g�����^�����4~��U���&T��#¬Ӎ�tq��<9�q ���5xSY��?)0�el�����������le��1f����~�������$V�9�v$2b��e@^[��A�!$�Iv��f�3D�[�����W�4ce���a�u���њ���c�j�x�%������ i��JΚ3v�o��֖�ȭ��Q#-kP+�i#��k�[Hh1�q� <��(�i=���a�TK�������)\ݛ����o/N:����/gj�z�& �j��y�N�����}���0��1;�'��5b3��9�P�\����`x�lmS/IéRՙ�U8)B�5��1c���{}�:�q&�3 �ӓi��S?���^R1 �+�H0�umq�"�#��?�n�l�"<�K[H�g{;��wQ�G��˓��T.,����HZO�US����_�7p�v��d^1I�ycD
U['+�ҩx�h-�SOY�G�z!���H�Ъ�2k���I��n�r����I�����#�n�\g��h�B<�����"�+����Of�)�)����,��;��7ษ�2B.�Mk�D-�w��ᇝ��
�*i5�x	_��`�w��sMSH��ɓgJ��_�<U��Ur�������$��X�2��e�\�(L?���㣗�n��^�u� ��mVx�^�_,�o�q����o�6�~3�3~۬]仃۴�2���i�U�T�f�3x���k�Ɇ�8;?�z�T�����͋����3����
�m�U��ʋ�+�	kSxٵ;7���E�x���D�P�Z�-	�d��D�(�f���R��eN� 4�S�bC�V\3@���׷��k㷌~��ş^�ȱ=#'�^$KQk��t����|ڈ1�L2���O1�̢M��Z�ap��g�d�p��Z5�>�v��B7�Z]�b'�~R�=�R��#�y0K��L\(տ����D/����B��t��Rčs@�z��� U޲�u���Ȕ*���lHm{QE��ǭ�4�\u<I��wz�  ��76����Z�Hi�W#��U�F�g���	�pwݬ:�J���8�6��7쐰.Q�npW<v����Rӫ-����}�W�h�v#�WzB2miZ)��tԖ��E��tT��]i��cB�n ���/�[���h+ ��>�BG��[�`�DO�6'7I\��Q�i��52���X"�7r��u��8%�^j:�x�r4I��Km��e )�d�$6��(�"�1��,3O��U���3�8d8$f^�Ȥ1z=��Wx�E)�M�/V��������G��㌅4b����������#��ʦ'�k"<Q��(�����64�͕E��VD$�oY�Ֆ&�;��\gߴ~4��ԍ7�ȡJ4�tXN1~d�5�Sx"�ҋH֗����ES�V� r���{�я~����Y]Q�y $[�->��ӓ�������]JĜ�N$L0d�ϒۓ=TL��]!}>���3�P��Қ��:�%�6�)��f�͡M��Thv��1Q���P�j/��	=��S�����UƔ	���ͼ	�6��p��{ϥ��|kD�ݎS�DU�6g�P�e��k3�3-�T��Z�S`���� �%@) |�Fc�om����I�$Nk�1�.�%��K#�/Y�'�j�n�dy�3W�����S"�gc��}2��G��]Voߢ
�ӧ��&��V����LΎƴ�E�fn�y�緺�"),��mV�׈���e6�۵\̉�S�Y�f$Y���?�~8������D����ʆx$���WSc��nk��]���l}�*^�BW���v��p��Ej|{���������/��B"<k/{8$Ӱ��<s�lE!�\ 3; 2�YsVY��u`%N�.����rulu�_��,��'p��a�Y�V��h���ˆ5��(����F`99�צ�m�n!��pt�)X�������Υ����x����'�Z�Q��h�f�盵��l��ڽ�B�<Y��X����q���t�V�#X%b�Q�Zೄ���4CȦ�����D��/��bb�L|4)r'�b�KC�|Pܞ����~�mqV��z��w&�op�[��c��IwMPSQ�c7d�q�؏?��xta	���]�;<<=�gB��4A�[$�҂���S#
��t��
�,��[�����F��Z����Xލ�m�B��E������?��b!����9���Თ��͛7������1�r���Y{��)@R�G��2l'�+�[�\�	��^}�\����^�hX��@����6���V����R����R�xF{R�P�������zk��)UMm-\6� Ƹ�s��Ů�t�qX���>K�.��[o�e���9�-e
ڄ�����+f�G��#n�-d���.*F��jZo�t�R1)�#),��ˢ3�bk�FTm�{Bts�.�};�[�kI_[�xm�CJSXf�_1�����i�^Q3�&�j	�20�sg0��U��EF����E�u{^ƙe��X��2����H�ڢ�>�/ ��;ݬMsM��%vwǶ���{ lB.���9=�f�g�y��ND�|nT
��3�}ĕ�c�y�٦B5@#�� @
W	3��=��/��l@��wM.^����0�T�pUSӮU��>'c���a�UDqJmĴf��"�̦�`�p�6��t^|�$�i�Xb�D�k㠘�v�?���C4m2�q������Yilc/Y	�X{��-669�nb�35P���+����5�k�l��hQbSGM��U��ɱ�֙k�~��`��.���_g��|��%������ˋ�tK��+be��]���_�w�8�9�fy~�ĩ��^� +��r~��Rz���}�%c{]���N�?~�n& ��YL�-�6��"?�?�7t���A8>Yu���*�Zx�,o���'eӭë�!�\�e h���ږJ�/��h)R�j�Sd*Hиy�k�:�{U�����l 8]dM��><�����{� mB�ѣG�`F�޽�4Q(���%��T�[�A��7�X���]nk��WM��x����c+KP2��B^�'�psu�$+��ޔ�.C�ʶ5P�hH-���>�L�n���8��t{�P�{��7�w�ܫt��������6_I�]�"��1T]p5y��WA�o�X>רG�:3~:fp��Y-U9�dQ��]A�pȆ�u99[�u�(>»��x�Oe�xf�$�pv�HR�j?�G����s�ڕ���Ç?��]	y������FV_^���M�Y(��
7Ʊ,b��g��_>�v�%h'W̦=���={3Ř��&�d+E:԰��/MuE��IM45G�`ӄ���X�zY'�qJ��,Q�b��tx�0��QQ��g'g�N+~�"~k���m�#�b
M-�Q�����)BP"L�~�I�0yg[1"���Q\۝R�m|�*��)����K�4
��#��*J|�B�C��m�m�?)�_l�D,���������k���^{�O��O�,%c�U�vGU��S�!�$U�\�f�$���1`P'������gF}{GVOp��b:A�����,�!3fIL��o}
F��W��o���4�Sw9_�8K@��a�˪�P�șH�Ŕ��&2m%��p�)
��43��Q���8n/�gp$Q�O����Y���H,���^!>8���1��{h{{�ics?3�.��.Yշ�c�������
�^|�|F����F�.hڍg���K�s�-�t�N+6Q�[�%q�u�k��JԪ����U�O�h��N�d;�uU�fl�S:�xb�x�2!Ca�� �8������BK̫�U�j"�%�i�`����N��=�|�@��k5�'~&��!(y�j�j6��6Fl�Lc��%o��6n�"�5��O�a���tvrz��O8E���l����]��v�N�ƽ�"�ƻ[��,���~���6��up>���]���wfc�lln)��t���9r�w@m�:X��M�b���Xa�fp564%�$�,�&� �FDY]��'�1�/�k����h���A�T\��I�[�I�N9�v�*dUL�}��Hq�^g�Qa��xo���O>99��pXQR6A1_Fa{�a}�lJ/�F�nSEUXŝ �J�-k��!��;d��x����b��d�6]ژ���]V#!ꌩ�yk`c�O'sN�֖�m�zkK�em�
�j����sǋ���Y*�q}g��5��]�y���*������~Y�-^��Χ����3}�xw2�	Y��K�l�zQ�銳�Wp�E��v��Bb�ݩr����+PN�Xȩ�"��*c������q6��+�G�`�n�ì9g�Q��}������2�f4ۍ�߀Y�]���Ʊ����_����=��6���Dqo���.���$u� b���ӌ{e��(�ꦫ�qǺF��r_`P�p��-M�`�h2sRWqS;a������EMr^J�' �����H��M�P�`~�{�����v��>�zÊ&Y���Ic�~��u9Q��Q��k�^�Ζ�����W�ek����Mf!��,_�@�<S�X��t��82K{���Ԉ��XF�<��Q��uo^���z^�@YF#��+7ܺ��AF4\�ظ�~-��J �L4X��(y�@F���q��!{C���a����w��k��ʕ�K
��į`�Ȋn���^Y����:;W��X�e5�ܼ J~e�4�_c��d�7�}�4p'�d�SVkp�gg'�ٺ���H�`��;�P��Y�,M�2��nt����XV*c6>���(��:�F0L뢄寛
�n�dF,�8�-M��t:Y�1�iY��?:�H�UiAWp��-��bm�0�Q��c ��`#I{�NS&����C�<����l��F�jU<}�8ɬ�nݑ H�=�U�6`�j�{�6�Q5l�Fx�ꌺu�D�}z�R���~��`^��<Є
����D�� ����;u�t��(���x<8=��'�ճ�O�_�� .r�N'�jX-Hb��`gw��x ?����f�Z=ß(Lp�VRs^�` iD�cf�q�c���:��=k�,H1��T��\�t`�=�aV�6r�y�k%rbS��);���	�Z�[���6�<��]6׋��Z禎<�:=��E�r�
��]S^�@�8觖B5t�κ]�2�_�H��!R3�; ډ�ĺ@رTՊ�J�e$ ĭ�\��嗘|3'�$YZ�Ы����*�ةMI��A�ۯ���I��ƛ�r ��6/�'jΐ�Rng�J���Y�G[i�C4�|��ȑ8dP��?{�N�?�� �9<<�����&�Е�2gn�������c7� �T�~8ЀA NLy:�W��+ML6�	+�y��N3:z�����Je��/v�H���)�a�6M�A$[)KH\a�^��z�%�&��n~��Ұ:H��i�$�{ڙ����&̼ċ/�$�ms���K9l�S2�Ϗ(���!4����v�$.W�j�m�4qr�ͳ�������=�G�+x�(`�{4�B�F�qg�kcl��tWӵ(���#�c�	-���:J^Z���5eS:���D`�H�Ԩ�Y��ԝ���ܹ��a��a-�����)i�8m&ţ�^<����x7�#��b?����,éQ�ѦڕK
=��񝎢�i�pܔ
Tt��#���b���<	������o;�b<���ƍ+׮N�+�M�| �<��/^�@^�v��ۣ'uj�7�+���l���T���o,���9�(&�cZ�ӓ3E��/�(�g�5*�8D��i,�Z��uvx����'{�^b_qqbJR��B�u��0m�Rt�����Y�X�mE��{�9�8xｯ���{6
�'X��G�ﭭĵ����m�r6�D1o�n��A�cy@���)70������ϰ��W���.��w�VE����%�H��՗s��~�ey������8	�czOa�s�������v�����^|�ғ��Y����(����5�����s�/���1���B�T�zK�r��Y�6��;�:�_ӁQUS�@(����X(����^Z�n-����Cm,�d��e����	���Ǵt��L��B1�h��S�)v�L[�׾����"�X�&�����m�o�����Z�9�fU'K�J��'�ՕW�p���E�OOB��ԙ�zl�������'���.n�w�y���F��Z�����_��W�O�sv�uL���<���3N�L�0��B�}����,�X�ۘJ�T��  ��I��������
]d.e�T�ů�:]�o<q\��k��D�����b%Rm�z�Y���J�in��03n��&"[�,p���ȳ6C����gz�����m���ׄ���ڐ�J�s伎�uC\3���ÚKPi �r�������9x7�[V�l3A�ɠl�)�f��	�^)r�@�\<8u|���Lf�ai؅&
l�9����ן>f��pL�)�Ɏf�X����>���g;ƞ����'8u���K����|��J����W�7
y�SGi���rs���Q<k%w��1HM\.0:��������F��5ߊJ�U��"��	�.5�oޤu*�@�O>���k���j�����8�d�ݚ�,�DgPГS-�Y3.B(�'80���22�:P�A��Sm���;9�:��6iP��MM�������u�ܙ��%8I\u-5g8,�O
�aĪ�,�Xa���ǅ��Dp���:x�5���!סh2�1C������W�Z�c�j8mf�!�`���lv�G��Y^�YlfR���5h��m'����]5��m���-[A�@���#�W���5���fs��z4F�6-`��s���q���'�B�,�n�Q�Ƭ_�=D�FQ�Ap��U�S���.y�v��|\�w�Vߔ|���DUI";*��q��h��o�sJ��ʼa�5#�i��_,�y����B؊&=LS��,���=�k�W�W�w.8�Zt��������i�ea����Z����I�"o��hL��!����I�,k�X�+����U<NR!n)��0A�br�������={�L5��7o67���3;�� ~j��`N���\��g��iֻ]0�f��B�Q�=�w�'b�5��H�(�Z]�	�&ttה69V���M��g��4�U?�k '�*^J�2���o-�fzڔ'Zuƥ�C;�w#,$o���W�^���_X�P��;9=��q�F��q��
�(E�E6D�=~D�fP�-�ǒ�%��|����_���M�	��
�#g���1�ĸߘZr6m��$��d 1E~Ĺ
��x���[ׄ#Cb��px�}���;U�s��\|"�7�l�3.-ˤJt�(�+����Wn�;w�l%�2>�|2կ�����\��؟�l����$�⶛��[��l���wr7}5����3��>�5kƗ��˧�8҇F|��qI���oONn�JT���D棈Վ,`�0/�$��vn��orm�̫|
�)�	�Ŧ���QQ���`�p,I;4 _����^W���@O_�a��\ꕣ�6]� �A"�����C��Ђˆ�zL'������I$Y$�����*�Q:?�(�ː���*A�"y���ʓ�Ֆh�	
Mh?��� �Z�&��/�誜`^r)�Kq�s?���cʦ��xS���kW�/�B�x���*� ��vD�k6�y��t�u�y���Rr�ڮ
|"��Ö�QEt�������x���c�?���c��v��ӛs���%�.ۥ����鹻aJ���m7�2RV�XL��Ю���@�*I5��h;�&��HU���"%�3�YZ{m�v˵nN�:5�P�0@��+����7��8P�]�8;������7��O�|���q���>[�t��Jv#���|U�E�n�:ƈߪ&o�\mx@+����\�$�k��	��,!6-�'��b�Rz�&2(r���Q��������Y+j[�r��.}+�ʴ�e�X��p����w�� dE4i��D}Q��c�~�����UlV�����5�
�(�![��j�d�Y:K��<��Е+~�e�D�La��7�d��/I�U^�O�8y7�>���7�_���_ٴ�Ɠ�����6E3Pɿ�3-��ݻ׸Β@���3n~l���I����P�+ڮr�r4���W��LL�$J������sec���T��T�=9���1�Uo.u�j�����n��t<U��j����\�X��6�0����y�ޞ��f%�gHA������'1��k�D�/m���l��'��z�І�i
�św;������d�dc�ޝ�֝+���ON��F\5�_�d�5	���붍��>C7kY���ޢ
0�/�#�'bY���>
�?1Y\��"�D�A����(�}�i���`?M���1*_�j[�U.jЍ�d8�^�b����d�|�,�������`�������
�����46fӺ����q��]���:aN:��l�'��^6_����6���Q���;���:��i�����Å%Q�5e�f�7,rV��r�_�n�����sl���w��o��*�Lڗ]���E�ϯ��ȩ\�{����(!��/�	F����n�������n���ر�nk���r�cff��&���,�^��e*�4	�l�0J"&p�W^\FDa�V�]X\���-�e�b��t;M�w(�zo��u�:�KF��v�3.����ҵd��Q���JF�p?8�=��jo��I1K}~�Qt�GgFa�s	���N�ILMqNC+r6f�Ygc��8����2��fd�PǏ�kؾz��c5�Fۀ\Fq�b]�K���A�*��ܔ%6[ _�`"�j����ի�&��fI�%�5�Z�]E��&UЎú(=�"����-�+˧w{�Ǥ�U��XN(����9��;G�b�RRH֫�+��ʤrb*�Yb�dj��]X��Fؐ�C������*ȗ���r-���[������&J�"��l4�������	MA��~|DA���	���|
�s���a��3Uώ+�P#�h��6Ǜ������WI̞�$��F�)Ǐ�w�z�����m��'Ϟ��g?�ӞN,��E`a�s���]ǖ *��>=?k���ЪGx@gg��9ԕ~�`зj?����h�1B��
�RSeROC���� ��Z/���)=Į�s�e���l�;�aj��H�d�ʧH�ײ�5���87��O5̧�5P���0��u��M���V%.N�J��R�B}
)aa��I���������}��
��_T9�	��Mu�Z������ѷ�Q-VK3��*Y`	c�O�w&������F6i��Ջ�}*�V�����n*PHAhk�eSoп	@���kfP���Y`�5�g	���q���-s�a�٨Mn�qe��u����69"�IJ���Jd��Ǜ0��4��V�m�(N�d�C��T��<�2���Zƣ���"
q�d�W�;��^���`rww�8mr���XV��a�L�;�W��l��:̂�Sq&��i��P�ɰn�����%,v��z�*R��e ]�7���%DN�Ә�We��Mb�u��5�P�l[�Ŵ��V�p>������)����r����O`5y����ͫغ�?�X1����'k*I�/�����W��A<|y�X,���kW�È}�#����-��X���|�4>�nyU�"�϶�N���%e�S�z�����K�Yj�Pv��m��{w�U�+b��,�ސoők��S�魊|���x`�-x�����ߖ[�2_|���������k�����O������t�O�l�����H))�?]����O�@{[[i��aǍ��tN�EʒpM7�Ƀ�y��0����:��=����?�E=g��,.ʨ��l��bE5�rr¨�]EA8�$T�m��5��u��ؓI�c�}>���&1t��I;�ĸ<9�稸����W�ߒ�5�P��|g?�����ⓂyQ&�}X��N��4� � }����'e�1���Y/�Ig�=䬀��Ȱ6�5p�e�ѾN��䆋��Np���{?�

e����Y�=U��ꋜ��,�|5�MN�N��@ 0~�Aw:��,^�x���=�����$,�a��ҋ�ZD+E��G۽ B��V�A�x�P�鷡�g%5�iݝ�9-<��,l7yॽ����=]��v���t&��vS��c��"�.9`�3|bo8�W/�����^�$1�)�lA���
�!g1���J�&d�x��ßj���,��U��x�aذ9�X��h>E;Y휃7|�,���6�0�|_m
*� @n�֍$�N\��r
x�	���Y���7�S�j����j�]��v���E3��]Sx�h
������'�����f@��Nv���k���2��O�hA���Tj���@t�T��[+7[<�Lj\��XJ*z����HAMZ�����'�z�Y%�9�AC��� ĨvrvN�seG+��y�u�\��]ڦ�"�Zw�2��zݩV�˃Ã���������a��|��ϟ���W�n<~��lrk%�`4\�e!Y��ɪH2]����ef:��oVxp�`� F��F�/��l=��*\P'���b3xQ�F+��d���'GS��5e���)#��X��� ���D�՘s�VG&A�,�Zm�X�������1��g�*��g5-,A�V�T-�(s�7�#ѧ� Ke��a&J��
a*�9��;��c+�rz7ȫ�q"�T�5+�'#��^�#�<���̝� ?�.��D�. F55�Ƌ6aI������q\$�Q`�@>�U+OO9�.����+: �WԉZ�ƅ�P�I�����q<bu��`�-U76��&�y�V�W�\����r�nS~���� �?	}c��4�N�1��s��U]ܲ=��c�ء/O�
&e��+�FcMXͷw�8��m�3�d/��/ئ���5^�&����P M[Ɔ��tC/>�?X��ҬX���'��ﭷ�2<�	ə̞�eG����}SX�y�(aP��c�3����y�o^�~�S������I�zsF�ׯ_״PY�d.5�ZͿ��U�PnO�x�;;[
ɬ��F�����0�3�f�9�;W�Tk�u�|4��c]I�G���I�3��ȸ3��J�mή�-��	@T>���m7b/jv15,��W@��y)�ʷ��)�<��R�~�	��=�x,>l,��^` nt�#\��E�����f¥��D��z�.��U�d}T|��j	�x=|���p��u��t5�W5��[�ӱ���|lO$p��L��5��MnQn�ꟕP��v��ޠ��Ꙋ�.��{5��f�]X}I���"`:�ɪ2�S�����T
�M\3����o������=|���>٨���i�Z�a���}%2�	�D�&qʢ�5ZRx�\�e�5�fژ�f�CU���*.?�?e�y8���-@e-䙱�V,����ގ�|���v��!�t=G�@6"#���<��><����܍�3-mW�Y!0G �o�^-��p��x�A�d�8��-��앱Ej"'��1g���w٘�X�G��ǽ����˅Ž�!4�%5��⼘%�Ef
��.ԕ<_�k�1IvVm㮋�J����}sn���� P���x��W�� *���S��9��p� 2=c�u��_�u�ַ���ǊO�v�ڭ[���ts<,9#�Β��������l(�u��@�?_s���۷aJ��//��9��Y}��cʓ87P��vA�ʕ��-�d&��AꚎ�rV��p�R�G21v���������Z4s���=�	Ng+�R���Ք�4���VF�I-���v[�����V�!�ە����_�����g��J,��V��y�ލ��.���z:4%<��Z!9瘌��M|d��Ly
�-���/����{�i�2U�r]����c����cj}
B
��FЉR/ݢ�L#�t�($�D<qkQdc�4N�8�;-��h���*tj�4¦H���"-J��J�\�j}�<�N�9���bd�r�����2���@-~�\�?9.�m�ڠ�t�:�h�}�7ܐ2:j��rS���С�8ۂ�ɂQ[F9��u�����2���b59���N.��	��7]�#�X����&kxu�rv,����7n0���5P����Sq۷I���^��}��'���#2�n[�o��DlA�ݥ=����e�rr�F��i�����s�t+3�B Q�4�C�*!H��Ǽ�����wn�QR�g��@(N幸�<�KVZ�5��Vٯ���_����H!��18&����{ｇ[��?x����R4�/^ ���;쐨#U;�b��JD6ܝR�2)���".�J��ƺ���#œ�x�/�D�,.-��nV
�l32��e�Z����ft����yY�^P����#'����7w�Ј�:����ѣG<ȑIU�b�������$�J6�4��t�6˻�i��j��-��RdfkҵXǦ����P���n���X��1��g7�,4�4�\s
xA���r��V�R^[���7�#��c���Y��µ�ZЯ�c�b��4sYa���[J�����p��U�DqY;��y�������Xp]�F�e���Zl�g��ʕ�'�X�[51	C�ř5�K@(&�|�V��ө�@���)޺�C�nAe4ą�s�N�����ӏS�U��8��!O�zM�.}���]�eH���I���`���Xѫ҂xH~�YW過�ԁ�P��q�\�H����2�Z�N��[�}eR��l.�瓖|�w�:�S��C����]}y�Bk��ǟ��`�nĎ���ݻ>��o�U�E|�J"]{�n�.��Iq�=�m��N�n�k̤M0jժ��B�¤u�_�+�3�ܝR��M;��T1{���8���	o���h��V�Y�w�?.¤�NN?��󳙬�n��7��A�#��w�Dil���@�h쵧�PǬ�,�f��VK�yOdtHM���iby4�)67��-������U\�p��-�Y��}
��'(Gx�֦5G��`q|n�+���J��SU^1Sq`o�y��(�ʼ��b(`�	F�d�t
t�-	�^�Hy�Ɗ��o�i�Q�X�I֩6�����t��"d����u$��2p�Z[5�-)�	B6�#{]%y�(�%0#�*Z�|�L�JDf�税�u=�y'��O��##W��1�_U��Kq�q��i|��s�u��8n�v件�K�Ĳ�G0�����s��d2�c���"'�y�7Ԡ`y[��w�h��L��^N��\�w9��o����'��_�Ej]Ǒxx��(`��l�9��KG���k�X͓Ӝ^1�V��2Y�O�zs���i8T2@�j��2��I,��}�?n}�;��?"��K�n���Yұ4D��O��S� ���F�}�K�H�0=��kDM�V �캱ͤG+8>]�gR�����r.�Ң�6�-O�J���� {��9k6��f(��tN�%t��Al���e���Vc�o(/o��ZHĹ����v~�1&�|�Rif��)�s�t�
>�~UŬ�G�ԸӡsZ���;� �Sy�p�g��-3V��� �&X=�|������$�>��Ns�srr������B���9	����'֗ ��a����F�l�|9yT��,ol�4#%_��I�*�����%�	���Ã��yh��Yf1����Tx�����dؙmŻ뼎Lb,��[l]fe��o	;jc1֤3�g�������
��N~��w�E�a}�o�r=�H����̓ZS+k��ۻ�Un�	L{]�n��t����󊪞��e�N띁gǞ��� �9�/��䢹�2�-�*d��W�#�<n�J(�`�Ze�\�Y+�ymE-�V�w�QΎ���Q���l5��?y�x4�]��͐���pG�����LYf�f��w�̻�IfX��RI��7�;�t�U�fHMt1��~�H{͒5�4.`46�������y�$(���o<��z���3��C�v����F�I���P����=�L�<��Z�A�ﳘM�%q'���|��;k�Ô��,M,�گ0w<ҋ7!�hc#����W_�s���۷��(��p8�r�W{c�
��"g��2�3��$i7͢4ٳ9$1Q�l~.Ke��}���T_�,�q����@���X�k=#�x8�$~���)��%҈a��@n?��� �5X�l���5�=�}x��Mg���UG#l��ͭ�[���b�XޏX��B��f�^㒨'��G�S�s"7aҥ,sa��7�����G}�@H{FXs���u�V;YU�m�k��>׶J�Q��tDZ�M�W{:s�zQM�b���������ً�x"�.���x�/�2.�
�01fnT7���{��W��UV��j���Қ�K���|�(�Y\W|oI�1C�$�v���%)�~�<��m"��Ѝ�2S�݇�]˘��`���adb������Vc�B� ��GY)�˟	"�@�hccl̻S�"l��(��Od������!�שIdf6ݯ;ܸz�����v�����?��l>��&6��M��6��i�
�.sYr	�3�;Յ��XS���%qm[�+�]�e�>bi� M�_O7��.MDa�J�3�{1�n����k��=tLH�9�4B�/��r0||��mDDLW%� �dm���&�EC5K�I��^����1�]����Zs��ȡX��S�
�x���W����}'���u V��+wn�l�&a
絘ў��!"T+a'�\��CI�EI��ٌd����SQ�%��X�kp�ν�ݽ��w���Ћ�X��"w���ϩ�u���vط����7n]���-����	Æ��~���W�:;j�.��iw������/n߾U�XEmd�pzR�}�9⫷5�.a�}�ɫ�t�>���Xr�7�<�T��V��e�N>+V x���_S=e�:6v��Ȳ�U�&'�>�6��e�����d�&Y�w��V�^+��O_�8��|:�g֔�$r����Ӏ�!_���uV�D !۰nV�E�Y�]��6��>���Fߠ����*U�C暱^�'N�M��Y���Q6�:��=���8���XƁ+���s�[μ0�� w\�l��'P�$�y�IQYZ0u����	X��.Gc5�(��	�J��eߺ��6'[�Q��5��E0��mē�A g*t��li���b��4v��ۥ�%�T���w;�ge�d��s&\�(k�0�j�\`ollmo�,4�z\HM���]���������;Xf�����x�8'�,�2y��g���HI���Og6R9���$h����I�����"�D����l����رY�U�B�n������4�Z�<뗝��e��-tBH?�6�(Y�����mS��ID6��e���6�<��Њ�=����gϞ�t��t6���<y"�8���O�n��J~jm
QRF믎�T5���2���R:�0�Ea5|z1�X���;4	��X��i�x�2nmi�N�P�fy�^<G񝅨ܟ����1b��h@*�I�g�<���'���b�u̈���GN@ !�����l�Z�:�6P����q[Q�}n)��qU��4�u�"t:��"h�-�;v#��V:Z+3M$��C���͍�Ղ�V�f�0�Ԓ��
�g؞�,�-du����cM*kL�bi��Ç��)aj���pÔm��g���8pO���9���jzr@U;N��(�nU�Ym2�:���t���'����R�Pe�[t�9%�'W'�m᷼6�R�s9
Xl��rk�)q��
ĥh�4}�������׿�vuoh/�B���MM�g��-��S���>yy�S�jf�%l�����E��_�rf�NL ����g4\0baĆ�$Ma���ϟ�u�ڤ�cϐ|ɡ%)~�a�*��KL�z�9|�5�a�jc������������7n^��&��IF�F�)i���Ohl����}�+�	��4l�_����ds�����r��ry��w{ҝ{��!�f��|1��zKS�v�0��+����.���+�C�����Ǐ�,�z�-q�^}������$�sS����~6��f��'+�B�Y�;�UywmG���F�8J�jz��My�q;c\u� �hwF`ElJed���iV��0����$�����ia��۲��F��t�G+ܯ�p||�8Q�X+� xK{"��R	�CD��:���D����L������b�/�x�nL��B�!�;��*��Z4�xJ�"���\]8Z`[����:8Q��������J�-�3������{7n��k�������2蕤L�ܙ�j�l��b����b��TZL�"S�T8�����,5>N�Z{����9{y<������5uW������~������m����D�2)��|Գh��ʿ�����6��5�`�J�%���hŊ��׉(�����8(k�,}��]����Y�s��@�U���Lb��7�,�����Pm �b���q`"���L���,b�f�EA���=l�8ɰ;k�:?9�>yy:�gǩ`��q$'�<�hkk�6��x:��/|��S�i��\����S+v}��M����e.~E:���s�q�l���H�p��j��H��X8��f�L���Ux��h80��%�[�:[˷�6 �{��hԾ�&��ʯ[>��ш[��o��ǝ�LV^�?�����4i��.�o���7�2�R �n�,I-���;�s�>��ʍ�1a���u�߭�=S�Hx���\�D��#�ɚ��=<��nT��l��9��jk�=�X��h�RP�e�?����َ���n���Iex��\�
E�a�gҘ�~����yiH-+3r�)�`��6R�fbN��׵1q�E�-l܁i�c�[�3pCo��Ж[=z�ʳ�qU{{{�6=�\�gf�Yd�ٻ"�kѾ#�h�ɂ�ڡn�`p�^LO�Jd�ܫ�uh��*�2&��g��2�a)�y.;�˛��Dir�F�Y .�_a���#f����δ5A�gɅn�m4���K�Y����߰&x�է���%;]i�
���$G�?go�kIz]��q�;����X$e��$�v��6�?���G�����%�c͕s��'��Z{ED^h�H���n�'����ǵ��Su��a������x~$>Y�$�[��'v�����+ �З��q&�d��n2�D�{��J�y��R��4̯J�|$Ϙ�`�0Յ�9KӢ�� Z���X�~֡����^���/�*��f���0���6�*UaMF]/�.KE�#�q�c268aL[��Җ:+��� ��	z��%���)��z��R%cdN�#��1c�)4�ax��7�ou�>ziU�����I��~�vmL^b��K� vsn�q��Fu��uK�0��(��7TZƹ�X;�/��{b�P�%t�P�խ̫�:�}��n�)AO�6����zWа]�,��]-E`����i����d���k3l������(i��c��]|���a'nd䆸����X�h��E:�0�Č�vj���;%���^>z�*B?��ɶ���96P�quuM7�a��yO/�o�g�x%��E����<��ӝ<��ϋө�	������z^ߖ$�<v����R��ׅ��8�	,E5f�y�D	�iu)f�9���D�mx RS��F�k����ie���Wy݃�k4��tm�!'�..�_)1��U�C��릎�%tm`����c͇l����f�Q�k��r<�U����#���,4<��';dCSɅ�/_��O�S� &��}sw�
�,2�8�'��@�́�Rz��I2�g�,k����J����p[4�u0R��1����$����B��	��7��lݚÆfI�n�$�VȠ���Æ�����d�|;���rmkI�����/n�o��o8��$�q��ٯ���M��t�#�U��H��Qww\�(!b1Jb�'��򼊳�[6JNc�c&ql��u���S��2Kes,�hh3@���Չ.{P�uE�
��b:|���#��qz2���G�����තRK,��_J82JEL�n( �	�t<�Nv�靲_jq;0��DI��9�u��A��V��u��q�i��⋟���
<�UB^��h�{��r���Ƞu��q\Q���ȗ2�'ՃU��z
=�l�@�k�N��<%n_7��|0E�j��"<=f.�͟>}��������4�2n���H�BKYj����M�R���֪Q�ֆAcM �X
��u!��p{C�U��Br"��^[��*n�JU:l��=�f簾2Ɇ�Hܹo�1q��C�f��:>m�	�����ʪ;�\S�)���'b���D_Rݸy(K�v�8'2q��J;�DV&ʛ�ݺ�|S��<m�ZSȕNi��N&m߽��?>������ɓ �zG�`BV�[�5J�SC�������R|���;]P�{�����;0�c�
�/+5X��6�q0�B3'8�ǹ~1���������ǣ�׿����^���Y;���m���E�P�Çf��h�TE����1�n�wo޾8;?j�2��t<;��T#C[Z��mʺ@��A�[6������Q�0�,M�?���q�~���Ѯ���Q��]a���x�㣓�>��y�������2YP�y�R����5�c�F�g�
,ưn��k�_�Ԯ|c7���F	�����V>�2��B�>�� �[�I�q*V�{����z~��/���qLrh�(���?�2'�j���T����
������4�pƂ(ȳ�
�5.�8|y�ڝK�ƍ��s�0�-�Mm]V�tē�����;D=��}q��:oq6��{��PnB2��7���C�������,�AϠ��Ύ���O?��?���(H��Wo�B�rZ'��=w�ڔ�ԩ4 �������rHTWs�_v̨C��Mӷ�8V�������f1TF�zQQ�a2�?ex�Ȃ�toGݳi��EH��NA4�C݈�w���?��??>9q,��'��Ȁ�p󊲚p0!��j��~���o��&�ņ@��|������������vx89珎�۔,'��}pU�D@e�&���`�lb��6�MIYSR��pFVh='�<���{� �X�D2��k__�,#��R���r}29:��&��b���m�&3�MY^�ۼ�&�ɡ���փ���g�M1��SS��eY��wW�)���h�d��x\����!��aT���?�)�+oY�m<�Nn]\N.��������Vxph��N���q�v��m�q^+���QS�^�~���N#ğ����%�Ly���sklS��Y]Y�>P��]�
�.�_�L�f���̠���z�¥zq ܲ�f\$/�^����WK���$f���j,BPzQ��Q �<}������~vv}�T���0��}����u�������	��������{����j#On<Id�)Ɏ���خQ���MfʼH׆������7/~��#�u�p<�3xk�5��y	[۷�ŀ7W�m�˲4
�C���q%f8	���e��f��oʞ��bq�}��!��j�������~4���>�����L��6��NS�Monc� �%w�/�{�
Ƒ7��)T>�./`�M��o����`'�'w���LR�l�A@���yY����|��)v�m�0�6F?u<VX1�n��#�M�"���"�ю�0yq��IN��b~�X6��rĉ�N��:4 I�p�p'��xX����Ӈ/�#k~�ؤ�d
�>]�
(��&ݯ�*�o����.ۯ5aͷ�����*��?y6���u��>�1�=�K����H�2on��C��t2��������'�YU[�?�`�6���.Z�z�-��}�A�>;�	�2��׏�Ӌs�?��O�;�C��7�@��1����(3�+ #��h�������O>d��hA�ǣVi��n�ˠ-Y�?@��a.W{���yY���[�ۤ��ݝh(�X�[��%0��"/�K�OpL����������xr
�8?�0J&��G���a*�u��f���#����>���Z��,��&����3ػ������_���h<����G�=}v͸�@�0����2���v�K�ș�G�>b�����&�/�ݒ�Y�`#~�}�9��X���7��w���C���"��8| ���!�-�N&���f�X�2o?	��'�[W�U�$����zU7t���%�SC��'�1���ᅂ;����gg'�؞����JJM�F~w{�B������歷���
�e� ��6����e��G�E�P�������6�l}�d���7X�����2����7��c���G?��尣�[5[�'|4�Fr�K���)��$)�=Ԙ��Y�1SQ��M
/��C�VN�3�9���%1*���t6#�>�/�}��;�|�A��-oq�F�I�ßnp�F��d�^��F�Z2:O���Q��1�ق:L.=���O���߾T��K�,ww���z�o��L��ܧU�F>�dm����Lu9�ksW��: I�:��-������T�װ�4
�}B�qzh����!����0��Vi�$��^t��A�(��*��5si���¥�xp�ّ��᳷��v�ĳ��y@o�h�=�����vc��!I���xB�����yP�j��͢�']���A�H�|��������4F��Q�[lz�S�O�c.��!r��n1��Qw�=~@��a ��"^�0�Gz���ft�VpX� � �hΔ��Έ����X��f����_>~��ǁZ�!��=7���mv(�ǳ@%��k]�Lo�⮌y�tw�M�Pb�\���>��ۮ�oq�pBc21�G|`LKq�)�s��<"��yq���nON���J�&=aD����ѴN~ȎO�-Xoi�WV�w�*3�OlZH�ɬ;�l�-���KGqP�$�f��ALZ'���q�.�n�W���?>��ϙ�/��_�X����co4N�!�^L&�n�0�,l�uW2��Ǥ��m��K8߻͎��Cƞ!���!���p*�We�+�g����
\�G�l�X/��6c�hL���b)A�s|�����Gq���
N��h9���XQ�C�ӌ���B���;
Z�xU~u�6���GH�ݸ-�U/��f�QX>�mQ��� �a�/`L˖9�O�+��0����wգ�;w��NƬ2�p�'q㓞��e-�T'�"6q���܉x�n�	(����4Nߢ3�����E!6���s,�3Sp�6֯8���i�],g��j(�q�v2������]]�q��&�����MĹ�ӛ�F���9.�&V#��)���9�������-��( JW���~��[�M�� �uG�U��5�gx�%��Ç��J����/^����/����G� ��]U]��V+�٘MV��������.�5�k��@\q����S�M�����ψ�<&�{gy���}􃏙��l2I�H@;6Ͽ���=�9W����Cs�TW�e�6���Qw
'΍C���6�35�Wƀ�0��S�[63�zrg�/*�K�ܷ�T=�l2l�z���\���B����,�8~<���O�<���Q�X{4b�����hq�:L�иw����OY��_d�p���ނk�L9�,̃��I'M���)��em�)H���2��?�_�N��o1�g����KJ�/�m�6&�s�b�^I���XwAlp5� L���⣏>B�w~�ۯ��J����3� HjWR*/�D��yu�6������ B�\�\)�n%��S�4+��X��E����uT=��3�����PZq��0u���P♑�1��(�wCl���K4���=��o�L��F��uf���r<�������o~���������t\�&�ė�;ƇX�@��8�:�1��L�P�[�ج1:KI����RGй�?
y���k/ �
SÞ�G�@S|��7:�ֹ@6_ԍ�?<���O?�tN`V�,EVO���Z�8��3�`�o߾��R��zf>��n�:�u~�fq�ӱ��xL/M���Q7ɮ���B�5�h�rd��`���t/� N���0 �[E#�������_	kHrW�P9���3H���$x��D�������콂yןbࣚ~��}	*iW��h���B������<��)�d^�z�_�ǧ��mt�Rs�*FJ��#��X4ΉTmC��ᴛ����"r�e�߷Y[Qk+Tѯ��ƚuN���}l�&6��	�6���+��q��Ʈ����onoX	�@Q�4W�֌���H�;��n8W���W}S��@��ݗ����"��|3*�R��Ֆ��C��Y���L ���\�=�`�����e�mǩ7����ՠ�!Z�׊���)��X�����Zcy�z),�F$uF���:MD7z4|[��@30e`�R�t�2z3���7=���Э^ͺQ^w����)I��0V&ہ4����������'C�A�y������3�%��^U�������!Qt��.77KJ�ڠ�*��g"��{6_|��א��d�f�.MfZŦʻZ�G�Ϥd��Ll� �a3�~>c��+�s��ծ���&�)�T6D�"O�̓&�g�.����8_3{����e4ٮEM�7�̻7o�w�>�J�I+QԒŴC�X�;�[cޱ�:����{�p����b=�W�Q(`&�/��p9}cHm.R��Z5�t���G�o�0��׼��e�+���n�XH�3�.68:���K76x�(G��P��S���Ko`cwyǤL�i��p�d|�I��q�>�Z�M����.����l�qd�{L�T��ᢸ��*����íJ8l�{;��j��?�o����S 7+VA��zm7�����
t���WW��;UT����������:w�$��i��w�
�7x�����-'Q>�<�$"�s��0Cķʺ:���<6c"�/0�rD<�_82X[<�-k��R��숺G�+9�Q�\�0,p�4��4O
��peQЪ�W!�p͸����N�����wƗ�M��ֲh���#%���Pԭ?Fޠ��}(A�O�d���j�aOO�!�eUHpRD��bX���Γ)��on������'�Wu���[��tB�[g�gs-צ��\��)�AR{ḱΝ�IE��[�m��+���ԻJ��yP�Oj�jju�uЇ�'�A�d�[]�#�� Q���o�����u�Sf`I���hltf&o�1�
W�o���Zx2�\����W]�?8�V��:�f}�� o	���z�GkO��Ԓ��7��>��3!�$��A�rm��yU�k>�8� ���S��aS�G�Z��-Ϯ�呰����	C��9���lr�T|���ȹL�b �N�C��X	�C�C���F;i[e�^$�e�n�?�9�P�&�\\m����~��#>��ztB��T���"�5i]O�{�0_�ԝ�m{*̶�lF���5�;F=��	@�7��5�I�Ӫʛj�./IT�%M4Mˎ��{aoq�[�Aj��nV+ʌb�0<;u��V�-\��,�ؐ^h^�m�#	m3\�!�� ^?[���������g?����qO<c�o�2)�.�g�q��fMhs�k��{�V�<_��⃂2.B�*�Tyѡ��s�f�/�),-Q@hMKDt,%uU��2�k��b���2���z��5C�
	a\����MStT �f��ǆ&��F
���9��-������
Ǆ���~���7�7�[)K3����?����(<y�0*0|
� �ӱy}��B�쩠�1��E�M�<85�zC�vL�iऔ��y� w�(vD�2L�F��
��&��]ֱN�	�U��0j��A���xv�����W�q�9����˒�sz��26C<���7<T����}���X[G��ΰZa���Fۑn*���a;���26��+��s���%+i+�{��(1��(`���2�Z.�����{�K���r�A �
������e�*��dv||�62Krwn�g'�I�����q��]i�JG<�N��y��X��VF	�c���O��1�+kUC�@@��9	n�������Oy��樑�>� 5�W��j����il�b����݈ho="���\~�jO�KX����M��
q+��V�)�J�`��ȴJ]���e���F�p��*d¡�B<�{�n�jG��&sAwL#�A���$�7WO0CyEZ
B�f3X��� VO����g˜<~�ñ3��
k,�ZQ"d&�޺̬�A*�̴]S��Sd�������uK�b�^W��Z���t�R�5�O��'?!t��b�����?���l��9�l>om@�0���G�>�6;Ǟ&��$�-�Ȧ$P�}���ό$EHc�p��D�#������\���{������y�O�3y ��� ��T�m3UI���({<$~??.4�IH�����7��f!D���Gdv-G��x4H�>f`!�2/#kKd�z���x��u�g�R��Kwy�qC�Ye�p�D���qz�>H`gA=�N1�R`��Η�g_|��n�2��������8J�j�Q�"����<+3�c._�9�8A�Dׁ5�&��
(~K�����fA�XY��j�z�������#M�Z�)�Ɯ�����O�>V*pN�3r�r��3��ߧ�t��K���nx����"0���z?K��^� �#KC	qi�<��I�Y}�
?���\:/��j�!<���_�(��'�Y>��N�N&*g��1�5-T�+,j�@�.i}s�����;9=K�Lg�it`�[��v���-V5����曯�?�G��)�HlڗMX�Ţg%�����6��r�ߧ���x�R-:X�,��^h,��;��!~*m�H���.%�O�����M����򺜻c�ҭ%��D�,�	�dZ�3��J˕0��I {��N��
KC��g�6�t6�O����*[b��.��#H��j�x��)q��pss����h���ՠ�A㈧Lr����V6ܢ��z9}��Xy�$��A�HB�t���fJ�`-}��&��M���O�v�x4��`�O�3��(���۶�d�T�ً,[���}��;���p��sM�蔽Qp�{l�CdEъ�c>��d#o� 4O݂S�?�E�*˻��
��6���6��ancD̴.כ˲��ӌ�]��"�fe���𐖰�w�5D�G����l>�Nf�Eh�%k��1���M[Tp��NOSf4�� 
��|Hk�YO�>UWM�{+$���Z*>�a�H�v������!`��h������6Ē8���-ا�M?_��	�T	I99c�4t�!-F�����G�Wϟ���՞�����x���]>���i���)�Q�a�3��^<�j�hO`2�a��X�\����oY���Kc��˄����?��+j!�&�A��Z�~�gOW�t�ĎNΒ���#b)��"�9: ��Y2��
��`r܏���BFи����Ɓ2O&Q�g��w��%�777{)P����e!<�z���
|��Qġ珒Qc���,��B�bǖ�5���h"��O�,��
����-�>:c�a(y�����2�^��,R~o���]�-��(��i�����9�`�7|������m4^[��${u�Ng�>�x:_4�����hB�/��p�DA�O����e�٦P���ѓ?�K=v|���Oj�~s���j��^5���A�(�ܤ��-���:���6�˻�RiN�N�O�"[��j��iqPS���$�j�f^x����1N7����Q�+�C�І�\~�26�qS��B{>/FIhx4�E-��g�T�-��i�1Guḍ�i2b� q���%�{	��H�4�
u�٬���|ux�b�h�ISu�r(�d���J���z���O>�<p�H��O�+c�Qcskiu���	Gz@*%�s��r�{ǩZ���H��%�����fyg�a-�8vg�n�P�cU��1�oEv����O�R2NiS/�T��ʲ���L�R�g6���'�`e�Y�����`�>|�3E���g���(uMF]�Q�X��:���.�PǍ�C��8$�&kr�:yq�<��uZ�oYK��塵�'B�ۻ�������%���aBN.ia���.��VK,HՑ/Rne<����Y�Z�ϸ;�����B�Ge���fO:�XE��^e�Ɵ`o������a�,�'DN�����Jغ���`6�p<!�)@d'?�Q��ć�6w"hv�˪��}a�gʿlk7d*G�ZA�'k�L�"l��M�w�Z�\��^~G-�̈u�ɞ�.3�x9;�.�\�P��	���%d;���85?�Qa@�K�l^��ڹUv����X^�敲�tr��{��9�K�7��g���Ō�`��������/�_�d��w/G!/Z�4�?:���?A��H�HKe��Y�=���fhR�G$ �o��
U�A
����15���.D��8o����$}�KU������yU8�a0���j���>�Όa�P����\/5˟���9հ����WR��g�^�� ّ
:�{��)g����p4�U�� ��eV�aQ������rHꛛ+���hq~~�����hll,^�g�-�h��+cݕz��2��>:�C�/�~��G�a�%=iF�r[Ǜ�s�C���{oBȿ�����n����^]z�!�X��s�_�fB����򗿄��l��j�8#vB��|\Zǩa]���9��j1}J���(�'e�=�{�?���1L�a7������Iu;�ܸ�g-�L(��@ա󥲉�������*�-�*��L���ֱF��=]ڐ���P�c��+�G.�':0C�\e����z&өZf���J�m?W�J���Jez�������^�b1��p
Y�v�+�+�$��_�����u�����jX���#;ᴼ����zｇ����\�]�Y���)��B�^��ԲӒ���p|��b������]b�=>}&�a7�I1ܴ8��fc��tlƟkX�HUz���$f,��!3���,���"�:�.��4�i���"0�(0n�+PwY].�#cf�#�#j�d졔��}�e�lDt�ο�կ�b�'�xvW:�l�ħ���P��h7�� �~Ȃy��5V��L���'J.ݼx�b��e���[�~��A�Չ��j�C)6��Xq�pͿ���|�5;JΔ�c�޸�f�g�;�m��S���∱�ﲊ�7����YƷ3������8�{�\OT\ʤ�6�W�/�I�xԍ�
zR�go�w��X'HeO��;�ƪHǰ7?u��fˈ���8;��@��mDۏ���J9*�2�H����0���Ty-����+%_��G����b?�a�P���QV�r���W�����ɺy�G[�h�����Z7q�hM�x"$���j;Z�P�����U�BZy�����c�aN��:kR�ҍ��j�RL+R�s�U����.p�DYI����b<)}�ӧ�+�Jm_W:j]c��+�_sÅa�p��p||w�Jʊ;R*3ID�3����R�Tn�hm�`k�-V�H9*Ϟ��X/�:m�j;4i%)u�%�r�3K)�:1>��=)���c�(�@޶j�||Ï,ly�Ňq�66@�/3�܎O��'��lEǃ��B6��h������Ɨ�>��Nx庴��68�.���wԂ ����//O����#6�P�_��Ǖ�t�������(=��XT�2�U�ꖈ�=���_����S� 0�p'�I/�J���������1��S+�u�
����-��~��e��-Q},����fJ��j�s��q����fS�����K�!����>�o$�~���Wu��^7S��gV,WM:�R{	�t�'�o���'��=T�;$��{,�ڗ֘�X>(����$)RdHբot0�)T�0V���p��r��wL���A��A�*�xW��	Å�*��}�M�ܦKS��(t<��%`�7'�&tVä��{^<%9T�� �S�5n��r<	�j��̇����F��%��H�V�;�(����+<���ί7�o����J8My9�%�?ዞ?�s�߸��|r���{���-��+	���cz��6��
]8��<��̨AeI�q��ec�QG�Y�8G�U�l�G[�.�����_����8�	��KVU��L$����+�z`3�y6�X��x[	ĦG�ɐ	�T��'��a?Z]��Dd�'�%6}���_��F��nn�/
q�9u�8�~撔��`�>/֡��m�|��/~��t,b�	�� �;���m�h+5nd(fYzeSy�>1��T�ψ���g�I�8�7���5<b�������>�Q�][��x�K�_����"�����-a�t}9���l�j�4�)�8�LZ���0�8����˾}���P�}U���iJ���y�Z*7�2j�{|�{j�oS�cȌ<�MJ9������?����lVl������dUP��\��m:���x{����T��F�vc@�#�/a��SYd<�#�,*��ڼY����c%S�F�D_!E�v\��溧�s
n���0+�S{�z�tД?R����@�'YUD���@H �r�Ŧ��m2��jw[��l����i�O.��W�wvR�������mk��~���q�蹳�\�^xУ��[ٳ����w��;o�링�wH�����!���N�3R���$�zg����r�}��\���\�޸T���u��B��Kq*�s���2pR8�=7�i�,ޠ�ޯ^�z�왝z|56(��
V��k��};����z,tdڞ^)�A񪀡��M=t�����=@��L�q�}��W:�X��>����Q��}�ѭ��/_�7+�B�",�$N߰%�.@�L��$R��=e�=�8�� �u0j��*��{Ė�~4��ifAw��i������l����O?���hfՑƼSF�����������A�C�8���g/;z@#
۫�z��~�D0�4rE�����g9M���?=9���m�$ƙ���Y�h�����&����2��}����(r�iN�{��>������$��3��'*�4W�Z����iB���31eQs�!��0;�ςF뭠�H���\Na�To���G	�Q�3�˽�8�T�����pu��ZCk�E<����p��jS��ν!/uO�*i�u��tU��,�4 e�Hx�N�\v2�=#�9 ����v��~4Mď���1�����KY���?�� ��p���9UUm4XaG�|G�X���R
}�"y!.��Zs�h+o6���L�������ǟ$�_���}U������7��<G-�!x�)���0�Yӌ�U8
�2��&	�E����뗯�˕�>X�;��ڋB���%�p��c���-�c��
'�r�ڰ:Z�ۛ[���S�X����d]F�|��&>8����|�ʦU(�)"���I��)�|E	GV����b�(e�z�h%�0#�:'�3J�3C6�W	7���nCO=I�������o��:��/^�x��Ybz����9�ё���h(�P�_�*�Z.oI�0e��Ś���ȿ���<|@�H�����3���gQV��}P�ļ��$
9�u�/Nԏ����P�����t��=:��=}�ٳg/�8q����F��x<e�^<�鴁����j�N����,#\H�tm�V���@(��)�q�2���:}�w�U[��	�l{Q�=�ah����^\_���PJ���T<ܣ��mi��{��;R&)�nW١�E�#7��'z.���FE
'�w�ݘLfP!�?�c�N��㓓�(+��f��ً��%�AiJ�zn|�m�X�����s�����F�I��8�^�~�HdYq(T��Eb��F�۱�wB������J�LϬ!�P���]�KS���q&�
�O�Y˼� �T�5�2��v��#^�rK?���p�s�5րD�(N,�m9�p	<7P���7�}�T۾�ah8,��W�-G��ZUv�\�������puO~�|���͚p��߲�#��/ut�+��v�v�\c%�����r�/\պ	��P���:'�bz���#.�әF��Y�MF�d<��6�]����Sb�ʎ����3Z�q���j	��].�>�T�$�^��֫�zI���y�\�19�yѓz=�IN�����]��;4Y�snI�8�X���n¦�4�f+�S�O4
]�aǑ��{svG��,��5w�#6�#qt��f1$0g>����1�H�xaْ��(ʘp� ;��֙�#�j"ϟ�'5��������@���߬ne��B��t�a��Á���}��=���c�\��%�����)D���`�.B��l�0=[j�z�������֬~� �,�͟��ǋ���
q���f;�+�l��\�$�:��7�\��ȶ�ev��Y�'X��a�����m8�ωK���v�p�	�=֣�>�.��r�Y�Ąl�-���뛣��օ>Y2۞p�D�ZU�� �n5��"�Fؓ$8�d�&��u����Zl�%/g�fi��'��d:������_l] p�pe�uϠ��e�p�8v��^�^�v�8��M���~�}
�<�0rbnaյ�<��Pg��r�R�|��[����-#Xc�m5�8�H$IoA:ӲignIkUX�;��g�+��l���x'���3�KMk���0H�W�[C��K&G�ى�i���l�}�����9����~�9�@I��G�b�d�ggW/ސ'�]����|��F�z}���ǜ6yS��uߥfdO%0��l�5�%j����b��X��(����~�C@�K��Ao�z��h��Q�xB Ć}��'�R���["���������.e����p�Մ~����IV���`�c��T̓1aY�F!��{��^o|�N��+�J6�A��i�ݺ�n�<��w��Ԉn�P�-����맧/\��6C�Ѧo����������{$��I	=\���aM+����|L�<K(��N.=���O...���X(0vp��3F�H�o�/��c�eW<��
k�9����\�q�1/w���W�<!��"��i����|ͬSUR�n���8�8�Gg4��0Na�g"��	p*�P��ѵ��ίm�Jn}�����͐��ĝe�
�y1'�	��Cm�j��I�L�x��:r��j�p`'���0�{.l����~�V��F+`!�}W;�mY9V����T�3cgpq0�ka�q^����k)l���m!w�<�3~��cx�_�1��TZQ�H<�5�=UEH�����.E=3����~��ߔ�>��#��D��os��R�AҺ�(�C�0��<w�p2	[�t����4��Ʋ�!���.7YÚt`&��8$�3c��f��V�l(���Hg�U��֓'�A���v��b�q욼"9�}?f/��	�H��֜B$���Ӎ��ژ��I.,��͏����HYQR3��|��^���a�JK�[���g�8�A�m����!�3���~�-�6F��OOO��T�z^ܞz�]=(!�c+r�6����pR�f���zY*�D%P�j�r�������H�Ny�!R�P]�m?�;�g�q5|(�Lqk^֣	Q�e��CT�Y/���´�<'GT*kq>U��.����^�Ml�4��4"�8�7��KX��cɌ��z�����V<�}��b��??X%�q|���[l�c�DI��ܚ6niG����ڀ�0���,|����Opvv<��|	����؉2�C�@�@���N���o�#x�r���mu�RW��Zj�K�i����on�o߾�x��c<B�������n_`UK]�C�Nߕ�4|�y�����5w|$���t2���@y�kh��RT� �n���U=��l��Ĵ+J[�`Rw�CyrQ\&ylt����`�9qA�l�t%�w�
y<]�շ"���'���Oz9�r��*EJ��m�J�� 2d+#���f͂��c����<x��ϟ�����'�bavbH>�n�����#��m�f[��~�R��`[`"�g�d<l@\�ȧ�%S;�쎁��B��H�Pt�T�����Y����<D������l�={C��­!�"Š��}�um�F��)ͪ��!Q莳Nw������1//Ns������!݌��Rb�u�#)�/_B��:��w�_��W�j���m��HB�\��O�����ggg�{�%q�iƊem(w�v�zC��l7+IK��`�̽7�pN?ql�þ��� \��NC�����S��}�ᇝa���HVg(���L'� �LA*�d�A�pL��0Qg�Ÿ{�Ӑ����X�ˤ�ߵ�:f�uZ	�/X������������+b~	�3��d��y7�$�����~j�|�!�O#c�F)g��1�^a�NOYī��U�As~�i�XaW��Zzn;Uut�F���<�a��߼����ۍ���Z��#�!D����,0���F�XX_��J�Ҕ�7_�tE0�D,bB�HkI)a��fD��F��g<?���*�Ъ�.�!�ƨ���Wt/�ӱ!����/�{x��w�$Cz(�~��6�i40RG~_h:R���@�~G�bG:���5����w�S��n�Vc��t{x:��W���t�G��Eh\��"i#�8��cċ�뽶&vKndx��J����G��A�e���aٰ�B�!��gC��<㎨A=k�cV�z��"��˧Lm��˧߽~���Jl��BP<����	�{\]n����ٝ>y:���P�F���v�ꨧ�S�Q���?��Y������*L���}rh4��������ٓӍ����[�C�j<C�* (���~aOB������+��C[��_�5=�����t�Fl�*M^��}���cq�1�U*�*H	P�Hy�7J��J��1��nn�&�ow�.��8b�N��Vtu�ym-ɮS)5I\�+~G�LCV߄����ni��M����z�A}!�u�E��qg�MI��"�$A���|����6�#���>w!d�G����\��P!�����\6�1�>AW�NO[�~u���5vhU���U�����+�����B)I��3mNg�KO\E�m����kS�k
;���˻7�Z�u�q��Mݣ/�1�i��R$�|����Źl��<�ti�T0�&W��Bj:V���5>����)Y_3�����I�~�s��~���`]�t�7�<HՔMi��H*�jz���<)O��q�U;}�f5� ���t�V0(ͯ�����x�"y��:��l�h���������h=u���m+E(�%��)ɛ>ee	O
�I��j�5�c��m����t���8�!`LҀ�jzb�!O�uE�5����./���û7������ԸM9�$~�����J��J�Ժ�=-����a���v| ��B�6����f42o�2Z�e�'��9����;0~�����$���mj����m�+Vn�y�]RL6���\ڶC��Y*:8�����A���6�Bf��V[�j~���8h�� ϡ/��(��?�E�U�#+�;C�x=gT�sI�OGFU�Zm��$W3���߾��dEd���rm����_�aύ�T�Cu�ȂX�HCI���Һ�K�s��5�+�� R繍uŎܞ�0�$5�;ϟн	�r�(u�+��6��W�NK�a��{����LV��ΦrX����=��h�<�Nn��Tu o�l���r�Ū�Օ�����vDSu{��%��l��)=7~��ԚL� l9	��1�='�?6}�`<��m�JXQE���՗��|����b����S��Z<z�H����D��$�T@BE��!�ɲ�]�Պu���َB%m�4���ɻ=�I�C*e��k������:���!�1�e0��S���	�U���ꫯD�eQ���kxb��%ڗ�H�����mT�԰2
7���"��������?/�VR�0�)�~�&E�iM�)U8��^�A�H�ˈC�//�?~|d�:6�8(�.x��<����3�CS{���1�?.h6�f���y��;qD��z6A�9Q�U�����E[g�}��,6Y�G�S�$n�9��甓:�H3��{&�N��0s�	]�����भ2����W&7��<aR�h��8�O��rz��j��LH����IM�<�Z��8���I����C�-\KVUZz�ț��h�s�J���9A��e�È�{��1 �R��Р��%
˕߬z���x�\���*�ǵ�5��w��[�ֳ&_Mk��ȹ�ۿ��_��7,G"�"f����6E���KW��l~�_ׄC��uf�m�&ˇ,��h=Ӄ����(.kw�ǋ�c��s�v_W��f��0��$�F	��8ֽ�kѬ�{[3s�:���)rh�W/��Vwu�G���^�µ��%G�t$,v��T��r��{ݍ�к��*��g��s�0/��~yqb���;�Mc�ke���U
��Nyո�I2i��F@P1�@�F���q�⠬�g�׷���'��T���I��[�z��͛��n}H��q}}%gn�6׆��A.�2���e�������xY�-+��gG���MzȪ8䑑ul��v�3l?ei�Z?&�bh���iq�QK�XZ�q8^>;^�A\�\�8!��fްh�~<������e�,/� ��gU�� fU3G�Y:šJ��o�`�^?fM1���w�KSWݠ��ݞ����
�g���r��b�D���|6:??/
�"�V	�����М��H�Re�0!a�AR����2��ev�B�TqV�i���֠��Ԥ�����-�eÃPp�k������pע��+8N��fu�fH��zɥ@�X��'e���些 ЏI�ղ9]�2�{��Ab+?����'"ҥ�q/t$�j���in'�̳-�%�G��]C��E�M���yq�?���e�fTW�ԸdA�1R���I��h�����&]��ݼ��4�zH5̡o6�C̪αn��c܆%��\��������5g��$���|��Mg�ǰ�o��%N�&��\U�M	5�)��^eRfe�gL�G����n��ۧ1v\a$���<T�����X|��Bl�P��#������x���)����7�|���s����[�3��Fq8�����"�H���ԉlke����DZ����#�w���MǤx����.�`!��;���`���jβqI<n�+��	qҕ���9�oR�������NVP��j�͊���Cy:#U�=ԭ��M���۷P�_�V޾�B��Y8|����r,]��R����`��,t�YĈONO�d͙�����˗��W7ףIb�V%l�z"�!ؑ��(Ϙ�*��<X�Ik�VDLk9O�0�*r���Y���r6�UX|䇯�ޝ_pH��֓�r�[o9'��N��e�#�ȗ�[�]��MY�B" D��}��ib{c����8}�Xn�P$6?-��⢑I��zh��;�]&�v��ɵ�8>
9M{�߃�*A �%mܕ���m����7���u���+x�#FS4e񌢎�ǇC���;��GGq0>��Mni�4f#� �M;�Zµ����V�BY���/�2�^aZ-��3��|�3�a}q� ���S��#�`� M��#�V�<4U�wO��5��B��@{��E>Ga�ƉF�'G'��#Ϗv����F��f���l���R*߻��y��ɇ�4���[�s���xZ5c��}��o�5N�ģ��� *e=\.c�ׇ����&�l���n�ʾqı�6��dj��V�b�1��*sg=�a|x|��mj8�7׫�rG��x�d����[�9ybW�1X-� �ҸT�D >��p�ɵ�δꁟxn�ڨ����A���?)�:��4�������w�/�����H�1�m�
��������ve	��Xse��9cN�8/E:hYa)[�-פ~{��%�I4�S�PP�r��f����!�
(�sZ�;h�3�$f]���L��](�0��<�ӡ��A�F	�ied��	"n+xIh<�J2�ӏ�`o7���������͒��������3d�];�m���><�P�QKgODI��
#����P*�����6��OiE)j̲��!2ڕ���
�v*��ǐ-�TM-�v�͝6��ґk�N��O�`�Q��A�����E���t3��N8� �v{ˬ�z����Ʉ��f��C+ݎ�V��d�}A$�V&�5��yr\�j��
�޻iZ�j� ���t{q�\��6�(���e��L����k{f*�Fި�Lb��N��xm4b�N��o�-��<y�P�c5�l֫��tAl�g6(,y�������v�����S	qt�წ�A�Y�N_\�Y;�e��M�B,Wp>[8�..��+.������� ��}��z:=��("[��EY`}��veN>[R��^�����%�sqV*�pe?����A0ݶhk�]V�v�(�d%#��䔭ja����'������3���*��*)��1�b%��c���qH�o~��J���,�Y�Pa���X,� ��y���??�� ��`��{/=S��J*�;��k�׵쉡��S�e(r��0(�#��F^:��dO�,��$tN�9p�d�"���E��h��ې��2�dh'ҍ�#�\	�����SH��F�:?zOX%=���������C1R���0��&�{����oY����!%�a�
j�)�iP�"Z\*�6������R�|¦k��B�N狣�S�o% �׍`���kH.ى��zg���u�t�OȒ�����i� ��A�[,�~����_����jf�3�ժm\z�t��!	(��C5$˕�v��������vS�4���p�sCU����U���񱔗r.�����4�m�κ��R�>)X�xU��~�7����t�ӏy��P�����
��p2�xiz�x�b�O�J����A�얊r�E;=e��Aa�yYeU�-m�Q.��6"�9f���#| ��ֈ��0Un��ad�#j�/������֐����P����qLj3,s��&[�	�5�?樲��c��_0��*�ju݀�/*��f�cem�U[ŕk�@߱ea�������$,˫���޳���N4/�i�N�Ny��0�5�G.��ƿ
� +��W�&#�]w�j+w8P�M�P6pꓟh(8�n|��W�Y8P<�,ƶ=�� �9�Tv�H2��w-���w�7�o4-#��/^�}�V�8�xëW���o�WۺRX5Xڏ���@n�.��X�p%J��n��y�������f�N�o���I�q3�ٷ��1���F��:p%%?b�%6�P9��C�k(�M�xV�Z���2Ќ�]HXq]/-_�g�im���`X����j�`2x�Q�����\�N�2pyv�oِe6ݳ�1���[>7i�憼��CA?�j�Y��8reٔl�CfWur�$\�G�:�
�F��w�E��AX��bA ]��%PX�2C
������L�sl�!��M'���j�vj��ӳ�3�J�J˩�L\B��7���?z|i���KkC���C�Φ���3�JM��ґ�Kf���oD'#�C-oFw.g΋����3�τ2�(.����ҫ�=����i�������#@1T��%ɩ�����zR���Ny�Z\0�"0������w�b�˦�6�۴h�f�Pf��5��`�p/^�P8�'����@ێv����!�Ukm�k5��˗0���5��0hE��giu֍SM�h;����Cp0|mO� �#K-���`K��15�h�)z���B!%���"��@U�����@!�Tu8w�7B#��!~��Z�Z)І��Ɣd�%��W�����V面5�K�X�]z�=5�#n������-�l-Q6����.M�K=oa��6�Y�B��_u-��NE�ӆ�����{\��Eo��9��4�V�y�W��e�_�.oV���k�Ŀ�V��R-9�3����[w��w�6�:H�s�b'����X��Vk�{]��{�(l�����8k�|11��w]����As��l��
PP[C���*k�����6q�	�[È�滸��d@E1=m�� �
����h͒��V���]�.�	S{�Ms�xjX|h��ˇpx./ϱ�B�;om�xS��QMy��S� �#L�C�zQ��[�`�*ɴ=3�K�ޟ��q�
�T �J���d��1´<5�P��q��+Lߪ���`�1��ӟ��'�����c���V��d�a�]��A0�&�_�@L���Sn$>���Y��eU|Neql�NVu����`������~r�NB��>�/���$
+��ؔ�\���+<n��$��O(�+	o{���ׯ9g�>�� �s٘ǳ����RҮ2�^�Q��nt0��g
��&����������Ң�L(W:��.3!�/��\�f���H�l7ި=��	��Ո�XS��M�r�1t<H�Cq�"ݤ���~��lq����\��)�'OR�C��e	���a��]e-�V�m� Ǉs��=���Nbٽw���	3��lߑ�w�֎��{�M���f�i�15����I��7��i�W[1V	oK}���Q��c˾�DTjV���|��9�X˛�O�B��F6k"G[��P	-��i8.�¦�����C�^�pf\���ӁVOg\Y�|0����u���)؍O���!J��k<�zuC�Vk�%G�rE��wϘ�@�<7��$%�^Ҙ�xЩ赞�����<.��4�bá���'1�b�3��N���QO؆�u�E�]����MN�i^�_{_�Y6Z͎��D)���L�ѐ
C8�j�����Ռq"U,c^k�xGg@a�gH�PϾ�^��a��J<���־<y�O��ĝH�=*S���zN6Zar�Z:���T_Eףc�a�4)Q�˝\����4C`=���3`�~�l.J�>D�E�r�~����7����4ن�~I�l/V{!ZCh{EĽ�Tk(���K��I�G%�ޘ۾�7: �ñ�(��9P|*ph-y���/zn7���)���Ç�8�A��WS?~��D���֝o�*����/; ���DL���u?	����9n��nӍjZHT�eQ��ROn�q�����?��������)�6�nBD�����r_�z}k#2�Y���� cV��Y��n^8B�=QQ��W��[5=����C�5<���>�\�Ê9�m�a�c����FB$�3���P_��o��j�!Y0�fn�g��i�ỏH����Z��n�q��"���B^K�M���h�G�YO��5|�N�zĢ~����t��I%�Y�3���f�4eٜ��Sj�C��8�9������9��Vۚ������֤��������0I�`���˳v��_>��`q|LB4��^�o�o^�ۛL��-Ħ��o�(�s�C�����q�2/��&��V�Dg�m����7/_$a0����^��沤�qΩ�b���~�zhw�á�v�eG�1�!0��f�vYJ:K���(t��	���\[Ǌ��T�Þ�)�����*)������f��R��6AOM]����@�pS� �b��v��ޜT-;�UNZXʷ/�ym���4.@��~�4��?
�����:�}��I��$��}�9�A�&���C����#��l�Y��Na�����$���8Fϻݮ��gux�ut��\I��,(�0N�����9���9�1��
�)�B���qc�nkI���3*3� ^����-m���rŉo��<���&D��?!'+��m���
�ݚw�'it�������s���=߼���KF!Iyb>]�7��o���Q00
��[����ХeQ7V6�ˊ�%���g������]���,�Zu8�v����*Z��(�� ��Kʞ-o���U���G吢g�Ö�D�@d�q���X�B��ZTY}����Y){b� �����@��t��q<�
��@*�E��Ӡ��+�BV\8,�����  m�Xd�~'��F���1;���p��mm�[�����@�,Wp�ے@�Ͼ��ȬO)����t�SMìa�G�j������r}��������6�{s���/��O�7� �E�Bn"�ɆԴ��1j'�L��VuId���飙c���ƍ�%��I��t���1�v���WR�,!��N�d����3»����/��6۱�esw�/�5�`ks���x�R@(� ���&���(#�P����؃t�����ʆ�m�!a��R���|;e�.��]�~�N��.Z�#%smt4�:#(4|�D��Ɗ�K�1�γ�R�tNX�zu]�k���W/_�y�y��;B�Kg�P��^CE����5��5�/� NO'����ͩ>땉5~�u:V~��R,��|��N���9�B-ur0�[�����Iy`�h4ƟQd�ܺ���|��E�ƍ[fe�ck���l�0�x�Q5���Q������]]��Y�ns��n˼����^�U���]D!w��Yς{mJJ�vY s��D�y]�A�W�	����7.�K�}��!�1d�`h��K3�;��@�z|L_(�t������]K�Dg�k���j/�W�7?;�M���w����0�w��Y���j�TC��.��>�����'��c7'��'�~�����8��gf�М0Al���x������ꫯLǳ��LKr�Ŗ�����m��p�h;���ұV^��".:u.�\�ұ��#~g�k����F3��~�w5��f�Z�j\;��]��:��4vl�"���F�M:{xA46�$�T�O�t��>��?�&�"�����Y&�rWTӊ�}+����aT��ʺ,�F�h�ү�u}{{�X$;f�̣��-$q�T���ɡ[����@P2�8��������{.��$���5�������d��/<Q�x&v;ݩC����.�������W�Ȓh����MO��¦u�,�����P~�߷�Т��񗹚�����$k�˂��hu⴬�R������'�vi���A�� �ȵ����3Ab�1���l��	^��$��lQb���NK�1��i�4���Z���^_�f���<��+pK����q���B�:_LTaِ	ăb��	��~��t�t(Yl�����������XlZ26���αVN�~���&�4�Y���V�i�:����ͪ.[��N��#B[Ⱥ�u[D�E���b�=y�+���������+\'É�o��R���8���Q�WYT��#�x��p�l�-+W����z���_�n	�U����x�=XL'� �������������Ƽ#r�(�\uYMdV/-�s2N���*��*1�:00��3�0r��g�4�0��]��1&�5,Rk����t2+�pr�T-��hﲪ�c�0ԃ�WxB	9e��r,ְ��~���%�_�ެI��<�k�Y��WW�V�  @|�o��E&�I��o�̘I��@J���tw�{fD�v�����9� 5Ќ�`���Ȉ{�=�[�s/٥*+�6�U��r�>���/��A>����1�E��p�!�jW���r&�T���x�#�	s��n�MY�����IQ7�$���^o�����ۅZG��1��g�j(_/�]v~yvz~��u�ׯ�J$�XM�6��� �Xn������W�K$`�O({U�H�����u���?~lnH�.˃��_|��/H�&L#|T$�ݨ�B�AD��^Y�P#S�U�4��J��u�)��"ㅡ�L�b;ޘ��K;68l��:���[��՚�����׀t +ƴ�N�e�hdeIE������Iٴ����ڞ�����;�+�YI�9L�,*�֌�0�`�
�=%{0����>}j��>
-q��$zn�={��C�l�(�gQ֊���N]n��[ċ�6��>ʱ5��n�;��Sq�w0m!��-)z%�("P�&�������X���l�l�ihsH�C���Z'��u���t�4E����s1Lš�m�\fQh���	{b	�jB$i#&�N�ʋ^�2ɾ�Ne\K�݂�H�H߅RH�!�}$pVH}}e�CFD� ����v��[/��x�Z�'�%\n�f�oP�������89Q�)��CT�2�|s��Z���Q����_�"V�K%'j��Y%���o�B��w��ю^�B��G�ث���l����5s1�j$6�=T}*��?o�֊�Y�O��rb��M�_��ovpqy������@�W���xUx���*[��N�+�(W�JK���J�� �ݔ/^���ѣGC���u��(u�8/��h�ZB:�H���$�`ZH�-[Ԏ�y���,��6 }�1e��Յ+�_j�%׹��D����gg�0U�.�/z�ؒ�O`��`���	����g��@[n����n�Wv��i}'������������)�s����0;/w(HyJ�Ţpg��n+�`H�K����K�`�?@��R}'����|u��5Lǳ�5���g��D���a�t�i�"/G�s*Rs4�&�&'����{��H�%��;�W�m}�"��FS�kG�_O~��gY�[0>�(M������젅�qR����D���ek>��|����陶���ڡ�3�W!��ZZIp�� zj�4��L�&�~F�AD���~���x�o�USvr�-�����f�,IÔ�M,�\�N�>�<�o���[׻jn��(��`�e����fF�������fʰ���{�[�W������ف��q[���D�����z���e���R�m����]p�i��T|L���Y��9!sN�\�L4M=�J����K�3��!,g�;���E��\6�P5p���LXÒ&fA���R�ϫU�j��Nt�0Wֵ��Γ��k%��h��b8��k=��eb��Q��T��5 ל���y&�6��;4wi{I^�%�0��`�Zv⇏8���<>�'e���ESl���΋�+��RG����[�ݦUUQ�P�ic��;D0=2s,(7�ݫ#(�RMP�f���}�}��`]V��A�/o�7,�dF��Cy�Q�\�}�-� J�"��Q��p�[���X��:�p��%l&��R۠�3�nK�����|�@O�d7�M�Vb�[�gԯ�m�4E���9�j'����[�$כ�-Q��l�h����P�<��Q���<��p)��Iql-�z�,�s�i��U%���;������7f�~���������+�){v�3D���G<�E_��۷\]�Y�wmŮ��j"瘨RxY�*׬d!��*tW�;%N˻j=Uw�[ڊ���gh�r�bچ�Df�<��'UK��I�9!Xo�ߣAo��ٳg�YеX��e�k�F�-H/��m�Li�#�Y����-��S-��Ǉ����hw��%�%���E�H��:8������kD r�����_K�`�w=�e�4�D��rK�������h2
ޡ%�BQ 4d���˗���<�˗��X�Κl����B�!B���?����(7Ot����ȶ���Y�)�ОWL^/�3��X�l�v�"�?!ԃ4q3���z|��XM&&D���ܿ����
�U	=��f-�WT�޾Cy�Q�n�9�2�R$^���VB1Lȕ��&�Һ	�{���������vU��������جA^1�U����0��$%���G긋�Vo#f��h�HJ��a�������a��O�+�7.O�kʰ���	�H�6[��#X�������X����+�ko���%��#�/m���Z��E] /���>�@�8n�;�ϲ��NՆL����3�81 ?U�,.ֶǲİ�׋�;U�ɻפ��m�u�ޒ����! �qB���)�ao"Mk* �g�'����yE���2ڒ�Iv�39݊>U�@�j�1u9\0����~�G{^_d�Q�"��F�4���{�{{�YA��;5��sƹ���L�G����ba��AL�481F_K�8�@�v�t��dՑ>y�u]��%X�d�<xPRE�>A\�!T��nr��^�5������� "�/��_�_�)%2�
Du^v�ŝ`Ϗ�3�뉋�*�D�.,E at҂�[��O�<��칙��>����<����\�A��$)��	��g����`���Ѕ����ݝ�&l��%��Q�h���^�זPN��q2���DCݻw�.)�*��*�+k{���y�V�z��S���������J�?%?x�C�O�{[3�[bn��?X!�I����?�5���]=/jDl�ٲ�ݬ��I���s�$,v!��a�� �B
܌��	XA��V
����h[�S�����mJeJa3Ǎh�,K'�Gy\��P���Pd��c�=���N�>?dB�����K�מ'&<���~�~72���a�E�b�w�Ī��Q���KD;�k�S���?�X�������y�/a�����_��w~��m�3'-�~Y� �����|7�!^�<�!!�1D^!�l0I(��ؼr:D�,J���ɱ}i  ��IDAT�c�z��{(�M!�J���^U�翨~љ�؛�oߚM�ó���雫�#�鳨��<S�������Q��~�ʅ5j�6��KODNQQ�ֳW٢�Q$q4�̊m}~vU�\y�:���XTnNe�68���JU����,�*���R�X=<2'�����'��X��oj��q���oc��K&o����X��5��恲<��w/�r̚�b�c/�zEH��2$��#a�X�F�4��E���v���o�}��@�q6���X�_4e2���M�Ol/.On�IRp��l�y��ַ��j-\]/;��MyzVW�@��Qf��;uѴ���n�v�G6g�%oU���j#��ʎ��Ͽ�Sc�)mWԾH��2F<��yE���PNtrXw��a �g�`��t���읝���_[�8�D����i'�`��zkw:�r{t�֌���,RG��tf��v��=�Ӯ`{ʜ @��+ �R@w��p�#�0���%���˯������{�`�W(7&H!�H����k��f����Y�^\%D�2 ����H�ff����/ߠڙ��,�t��~�tED$�^c>�_�f�4�V��x�� Ҙ��4"n��^���B갯�����?)#B��� �ݮ��6�i�^_\�~�jqq�tB�X�%���g`ۻevr8����|.S�>�_�o��3�b[����i�F�TeMQ�*��y<��]`L5"�7e���ZFЇ�F��){1��r�B�1)��%vf��sUM;�ܓ�7��ٔ����{�`�*���3�/�G�|����������Ԟ��2�����b~��	���F��) ڄF�1�S�3�zwy���7��lS���x[V'g�r��X������z<ٟ�gy������x����ɽ\UF>�!�?��=��[D�\l�l���qơ�����۠��ͼ��\�0�xuv��=�z~Z���@��U�tlF�~ZM7]C��rJ�sx����te�yn�.r�xR�T��jc��v.�6�*��5�B���\��t6��`��钛�#��y�����Muyzy}5�L̴^]��)�۷E�v��*Ywu>L���bJ媠������;P�^_��%g{{��Q�1"T(����B�<]�6F�m.i��乃3b]7��kϥjLuP�u�|~mg�'���Q�@��$�F�z��!B�s4M=�G�v�ܰ.��]��P[ã�rlb~v[n;[���+�fc��P�l}�-��S��ZT�D6Z���C��?�����a�{j���3�0�u	hf���x2�����w���~��_U��!T��'۳����"ȴGZTzƮo�������T]6�BE��m�������1��f)j`��z(xF9ػQK�z�vZ�\�זRR���q+���%��Z�v��!�=��A�ow7��źz�����wF}t���r�L<s����|�欶~h&�)�b��7k�!��[e�������/.�Gǧw ϸ�����9�������]�><e��r���d�k@�;�&�K��D���E���*{n����ݻQ>���p�h�lYY����-vk{���ǘo|��]Iʲ��Q�A�؃Ju�ĳ��;�:J�N��'��2�j^q�2��VU��������҆��3�������d�J�y̪-6�`?9���U�Jo�P�5?:N��C |vzj�����T�j)�N_��N�P��֨���-´*7�y��Z���S�j�8N���t�g�I�f��� *���|�z4nh �؈�&�8���|��a���r��G�ܬ� ��۸�r^Ƕ�6�~�X8� $��,4 �c�tIl_�G���vC�(׋��t,R�
��f~uad�^��&:��$��ZN]�tL�fv��MGs`��ѣG�9ϟ?WO���ȏy�eR�7�l�\�(U���5b���fCo�j����mF#em�>xpǾ������1����j����i^m�T'�>ce,�U����v˨4�ܺ9��S�_�f�FD�ُ�)Ԑ/��Zgt�����gϞY�=����0Ɏ���'�nkh�ͬT�1t����'|EONU�!�������P�#��zRv�WX�M�v�	�.vB:��kh1j��1�����|C�s��64�fE=�T*"/aK���MY\^��7K��%��{�j$���l-�'���������Ez�P�7�6�K��;��(Q}��˷��JH�ʯFV�Q>~��~���0>�� �멨I��ئ�K����{�Η�L<�t�,;����:����~?���}������Ӷ��)��ӓs�}m����}������PU�؅%�B"��R۫W��3�T�.�k9S��F��vk�m��L��@���|���������3�2�j����X��o��'�޽��Np7��U�`�}���S��w|}������W��ߪS�����)5�ԝ+��D�� �_�Zϗ���-!��]e��8���b�Ɛ�X�� }$�b�x*^�ŕô���
xZ�Z{PڵɎzo�ţ*�tN]ѱ~D<��D'�:�9�l��1�dwYB��&#�%?�uw&<r$ѷ�/��o�)ޑK�|�j����{�3�u��Yl�x�����:xv~�J����n��������yc ��kd�~�jd�3���/�>�~P��wSϢh�?��(Ĭ�p�#�-nyN�̲Ȁ��}��Q�O��Oh*������v�R'��'�ȩ&�[D�j�%(��yU�����߼}e�u��f��Z};p�^yP��C�P�<�"t!y�U�9�U3"�Z�28�C`�6��r7��F�Z�nxv-�U�ؚ�w�즚�B��K�y�&�#>2.<Kz8�u�7[K���
�7��������33we:C%4�!�<�殡HY��9I��fc�ұ�V�^���a����䒁4Y�kD�)���sJ%q�}��O8�n(���M�0)�����ۛ��V�Ws�U`j��E*�ђA-� ��N�Ǯ�^}r
hl���T�PZ�|��6�[`yn�/��D�	�?����ԧl�ŉ�Z��G�L=����z�tj�g�;���*/#xcK=�p���l�f�B�l
��4h�]�_����:>:��M�ed���Ы���&��w���v��<�#4����,"�H(��h�Y8���������,.ڐ^��w��r��H%ʜJ;��
�������,6r��y#/si+`�9���ٷKذkf>��>�²a��A�� ��l�b]B�����N������Q�LQn-���I�sn��(vغb+y�'�cI�L-M��Pɭ�UA�5}�X�ʵ҂!��0f^�y�yY��zsttt=vxs~-�$��إ�ȉd̓s �ִ�Cmt;*��ǃk�IU�V��zVa6<���[v�@Ԫ|_�2Ua��D�d�vKagi�_h<���6hz*r�#�{XT��HIǳY�[���WvI�6	BI�
9��篯�詤�	������!o�i�˛�SeO1�Y{�g�Ì���VԍW����PP�u�i],�����	���lb�7)�"%i��Ij��Ǚ��۷G��h�ʇ0�=I����
����C�B���=�_���0g%-�����);��n��k��-����h��Ǯ�"�f��s<�T>n5�eK�p8/z�@9*ze��O"7�����7�|-����i�&�gF,4��"���͛�����8qܦQ��<���˺�ފ\b:���B8����'O�y�4����!Ce�9+�р~��S<w#%u���0Ϙ�]t�f�8��s��m�Iij�W�M�}o�,$�ў&:I��!��g˟���O?~bN�~t}���o~��l�����+-T���JwƩ��Ȓ+8��~`�׼�o���1k�#�HP_(��
ONN֫���S��q��:F���nD����������^i�`��b{���h9ip��	�^�`��0�G�;��Z7
��A��_~iUA�ڨ�;!�8���rBR��P7Wfy�:�&�-��pn~��W��'�i�����ɍ���<�ZJ�%Q����iLt��Q����d�>u��{3�eM	���&��Ƚ�3��^���\I�*4��Di��1�͉d��y"?�SH~�ד�O��9T�Gqڥ�z�jvxx�xW�kʪjP�XƆ�#m� ,U;�4��s����/�t�)�I�D��dj�y�T߅ٓ�r��W�ln�Dt�7T�@lI�i���d��3jdk�E_��=��l5q������ ���^�|����H�4���=�Yo��$�>-<�8��L�]���)5��XI��[��*A�w��A	�}��i2F��-Uq��J3S�����%6XBІ�O2ڲ�	9�V�%'�D��a!Oac�9��r)�w���1y=�"]�OVt��>�e��G},o�����o����E[�i���j,9�;1,��u`��K۱q`]ǈWl�f�P�#zт��O���m�َ��vA���"��
T4�yΓ֫��]�����?��_��`�+F���c!�j=�P�P�	o�<���qگԎ��1�U�,%�|��f�_�~mf��#���Ϧ����_�򗧧����
�n��!��:����=#�����WPGU��V� d����4�J�����+8u�O�X�b^/#;���s���3% �o��{dP�Kl���jq������~e�����o���C�\��K
�����M����f8����f����G�>���ջ�{a��\��W�Edv��s�<��:�3��ը��b$LH3�5% cd)W[՘��V��s�*^�'��u4�#����ٔ������z$
tB9�@N+�s���_ �����������~�R.�w�L���P���a�B��+��H���ʝ�E�d&��@D���؋|{JQ*5J�^pBu)�j<���&JDU{�X�g�VE��^�^���yryr|���%ȁ�VC[*P�S��^��8ߪ�������������>SHz}u���$�����4 ��P�f7��A�2O��)�2��e5?��u�o����~eq	��>�i�0+\����\�-��-�C��$���]����{��2�i �G�'��4�!�eђe�}�q�r-e�w�f��k(��>�-��* �bU`& �@�gM$s���<طf��IԦM�l�ԫk�_����������իL�ZS Kj܎S����n��r�,0nSvчm��F��ʂ��4f���S��E�W�һt��5�J���p0#O~��!v� !��l��6����6Ǎ'' ����R��<�`���3�i�(;�]�}nf�|r"���@�'té�b����zy]�����\#6��^��A֥70��jp2�n���x�P)��������aX�lO�x�(��ߘ�ۇ��1��%',���p��5����z:�c���%�骓NWH�<0���XjgKnNle�tuYW5sl�,�;yw����������0SL�;�p�,���++� �^~��Ei���a�uj��Z��>�/0tVl7 ]]Y�\@yc��!�#��Y��nga17k�IY��5̫ښ�b$�Il'W[��B]=]a���x��Z�K��"7 �Uܷ9fp�[�3e)���>��û��*���tV�^�E�y*����p���^72O-7�j(�cج�lm�o��>Gl��"<�P1H ���/W��N�#d��Q���y�����,կ�U�XB�#EޛY�"�=��l�8]^/N�Y@�ݬ���QJ`�۱�QK�B����f��OEj_&7�w�}Y� l�QR�ʓ��.4�����"��U�m����bm�~2�O�s�w.W������pv�(\�Vr���:T2�A��:�%D%�Ӓ#��r~i� a�(�8;����־ř��{���&��dh��]5m���j� Ԋt#��@6M`����s$�1�#�)z:e
(c�J�����뒜l��Z�X<. ���U���SZlZ]-�f{SpQ��1g��{jW߾���WϿ�GHtm{�@����pPS�6U=�mߟ�0�e�*t�KP9��i�ac�͜vl��Q��t�̡�-X��L������lvR0��q�A��i�;���ݔ��~C~n���!��)$2Srͣtcp4������W���<���W5XOd#�hU�7��E�r���*kT@7*�c�"�� _�_�899��j���*3v3�c�*�Y��4+Zبgg��������m�����/P�ae����s���hGUf~�M�S�t��ܒ�4��.�ڪ+���/.��zVc�>��0�Z�;3	���۪ͯ��@�Ԫ���El{4�￝/�8}m9��G�QS�� �˳��&�]s�S ��Ѯ\�v��Ct�w3n�xl�+�L����?��K�����^��Uw��E�R�����v�f��{�5q+�:�,���8��;��2�]���w��VT-)�4Q�Hy��� �Yb!#�7㍅���r�i�q4U	�����Dy2�CD���S-ё���W�
k@-Y2*�p�?�Q��^�$�p�Y�#~=F���5UDE��ޖ�촪��''��Oߧ�T �s�.O���.֫b9_XƁ�q�pFr`�xH�������f�J�^նW:K"�����&R�1�|�Umv��O�-�+t�Y�����M�fRf�'�+r�j� Tc}(�Z*���N���'�Sd2fgо76�n������~����ǿǥ�<5�~ k;��^���ga��C��I��M�JydAK�=��i���`�M@�%�Jw���1Z�_����\/,b.��/.��
���/�C��E@δ�@�'f��ݻ����>����5�9�^�b��ZC��ۓߏ[Gj/,��bň5Au�4�i~�N���	*����/�I�]/�`2Ɇ��z2��ث��5�<I��9wcm�DAa��'�4�ʒp��B�!���$�����݈>���#4�FJu/(�l�`���zu�=!��XZ df$��6A u���4�9;�5T����K�;��U3A�En��f����2R֪�1�}l�Yhm��yd�
ٙ2�����r�Avpԃ�c�t��T��p�j�v�����VYm%��p�v@h������,.���9}��!W�R{��b/®z�V@�I1��)vk_~�������N�v^�x�&�Ẍ �W3[ǳ�����Z{x�~�@�v�ph�h���3�3���������O~�;�o�?��c;�i����lA)��2��p?}z��_�z0�o]����D�8�_�m�νb���0R7���o�/�%��J䚒��~s�7��~0��&n�A"����w>��ӧO> 0�"tv����D�8�W�w7���A����.���b�P?�������òX�@� TW#�l�\P3t<��99;��]S��1?iI,|�[T�E'�F�o�~�s�^�L�h�P�K�6q��!E� ��+���r�n��+O��z;%���A>̡�#�Lj�t[��/����y�	v�g(��5{�@�1�g�	ٵz>d��X������)J(Ypw�
w�i���!��K˥j��7���'�*��H}TݻD\��PF�uiA�y߇�hAs;�Fh-�T�
lP��p��γ]'�+�[�$� ;iFe�vɅ�C&	P�t�a z0�n�`�/��۷o͂��4������cbg?�s���^E�A���K��a�:�1i�%��`���x����>��jq���VA�]��a�S	l�
��v�~�(^XN$������J��sp���������\1��eF��5�-�|8��WZ� �Pm�g�X-��<�Ek�"J�~��+0T��FD��HNFcj.�EN[|2[�`ä�0��ih� �hZ�Ôh�ܤ��G/J��i�XD�����]	� \�"��p�� �0j#u���rx�4C~+�"�6���(�EI�!9�b�{���h`a�XÐ%f�4%��m��~�x��c ?�1ף���Ʒ�R�`�%@��������@Q��]f��X�qmv�U[���hc?W�]�F�Ȟ�o�<�c�)�2��^/�!��\W�͖e-�Ƨ�=�FS.�f�֓U<�B@�L:d:�A0����7���7�Γ�C-�%��*J�������H�Uc�~?~�G��W�B�i�-����AQ��X`Uf{���b��ȶC(�UU���ڟ@a|o���<�^pC;�ڢdx�<]�p�xr�.����
Ȕ��~�.��J�-�4�U� ('t��ef�~~~zj˻8�M����Ȧ�9֖��uۄ��AO�z"�S�Kʘ�Q��ȸ�<��G���X"׈�C'���z�T<Z+UCCN���H�|���&�G�;�8�h�����=>~g�7���b��RS-�ܩ�{�p���5H\ܜx�l�8UD��F!���V�H�m6-�U�pC��Q��K��O۬�isA�d�H-��6�4��'�K�KQ��ĿS�Y*�Xn��4K�lHz����v<��|�S�e�8e�������B��k�N�^/+!Dd>��OJ[!����A�TS-(Na?|��٣G��cm߾y�������-KJ]`��e��o�xD��-��]�!��^���9�kG�מ(��� ��R� ?B��g�y\]A�x�j��Ηo^�UJ�PPhV��
�O~�SuS`_�^C�8�9M�:2����ξc6$�$�ў5!���' _���L��5���a��	r�� ?�H|y��&ԤT�Q7Wx���;�Ml�ڟ/��W���M�~K���ت�Ɂ�+��S6��}�QLF�u�~�Cj��~1 z��0?S�oI�s<�L���$�����=m?�Y��(��o������~�'�8�Z��qf9��&�'�i<�s�e�.���,�����~
�Reys��T��<א�kv�v�I������L��s얷ok[Fe:jD����2ը�]��Rt��	<�+t/tZ����ۗ�!C�寤5_#�(�{]�l����<t.0�����*p��!�n]}h�ZO�q�K��.��&e��y�!VUY��b�~|��{}
���
Y	gS���I��ޟ�F�P�tR|�d���ۃ�s�9!Y6�T.\W+�N�j[k�*䚝}� �J�A[Lbku�Ν�>��(:���	��2j�)fZ։���t�c8��ݻ�-��
��Ƴ�9R)�������w���/���?(F�y��t#�&��+��Wnk�r�q ~�5�=��R_��Y�h �\�U���m�o�^XN���O�Ϥ�PƧyU3X�]�.݌%�oƪ�[N5gJ���a?��܀��5���Ņ���ff�!V<���v�᱀�2B�͏�(�L�0;*�W�"��Q>��|��'t.�6�f������H��T�������>�$K�G_>UU.XZ�k��@��v
m��>�L����i�	!T{5x�{MaR�_)CT5&q�>���B���옗P'�������#pŎ���PA���ڟ���_��Gݔ=֧O����S�GD�zv��y���:t�����
����\c�%�t��b������>hI�������r���/��ݻ`v�ާ��U��xk7Ю����.��@���x��5�����+���:�o�"���W����#�\U���
U��zɦ�E���C b��ٻ}�O��m����g�}^�>��_����?q�e�t.�,��tL�����[��!h�]�Nq�n�.�Y}8�ڋ�I�~�N��e�u6�~
�	y�� G����G1���!�È|�����O�����w��X�	��L؅��޺�gA�^㧮����_�`�I�ݽH����˄v1�_��۾`���<(�9c���b3��ؙL�\�27#5%b7d7{�0'GM	k�E�0n�˻}�� ��9��b)�(8KU���5��%{��-}������ݛ׶5m�Y��3�Ō���S�Ѳ����ز�q�F82�/�4� s����I��]�?�L�Q͖�ĚǑ��)M�^q^���ױ����H�XT����D�G�$�!��� ��#�GK�4������ �JC�Y[@6�����<&�I5.p+��'���]�����\9VA!�4�Ң��W��؟�cb� �	e�A�,�k��Ǐ-sɳ^��<��""&��e4	狋$�p����Uѳ�Lr(]��q/3�{]��,�h`�c����S����X/Ps[_�T5p�+���Iv� ��I��_��GU=7?E�㐸y�Q05KFQ̱�q� ��;
�ff��jr��6�hπ� #�]��a0K��߱'_W=�)��W��>��5�U<��9O�-��l����x�B bK��$ ��l�(�/��1L�CO�
�t��	��_E�)t$l���R�~̢:�&Ts[̛YbRV�rj�~�����j��1 � T��c ��}��2B��gO�\��zr�����_�MYT-3�s��r�@������g�%}��犌���y��2^�m9�;�Gyqf�stt"*RZE5\��`�q�b�3���PScM�3/�H��,=�$�Ա!��\�/`v���5��%@��&��P��pB�l��d�IFW��~!t�VH54��<i�S����ڛmc�b��R+�O[P�`�t4&w�2���*�Z�UF�8��F�YKt^�7�WeGo�F��E�4Fj�K�!-Y�����7�����}�^m��1׃<����C���5���4�$��g�Uo~d5��l0)��r�Y����"�0���3S�ڜ���洏j�u�Jq�g�6S�Ŷ��;#�J�]$TaRF�qȇ�����>�S�#|^���7Sɳ9
38dݴ�"Մ!�Դo糶�z�q�Z�]�9�Hc��jq�d��P����$�f=�N������GVf�`7Ww�p�8��� ����'��)�QT�\+�%�L�"�Z��$dۨY�<��	�W#�TO���O�޽k�17�W�W��s3��р9p��?ӄ����C��X�@����<�a�����<@:}'� �3�����58�׌�h��c�Kb�K�>��e��<إN���Z+�l�Rh����p$�t�wk��w��E�������d:'���jC�P�c���t5��ȸc��J�O&�Q�ާz��vNE6
i�9Ź(jq� vJ$J��,��,�i5ۣ7ϟ={�V��/����6E��^_��)5}-D���w}��5�����vd�͐����!MWk������a�>�C�B���UQ	[�^��'��Y;i&���{ih���ͦ��<��f���yW�em^U� ��c[�ck�'ɶ(kȘ�a[����:�Q�n��vENj�h��/���C��n=��� C9�^�p�r�4J�{w�=���dʎ��CA��Qz�f�4�������_޻s =��wP���k�Ļ��.;R�i/�$�E��Am�YΡC,NF���,�����R�,[�z{~v�~a��;�K{
%��q�L-�H�1�ͥ�|A����brL�c�'m�!?����(�ꫯ�.����3��%���a���Q7(��P�5o;�S�PDd�*��G9;���L���`���j���*���Vi�hT�M�ꃵ��
�>��. g�^_,�*�7cr�$NҤ���ѣ����Ν; b�F2r~	����j9\{vp6�A
uU�j\ �f�E�Nd,�2�P����??x���Y��ϯ����7_�����V�O���^��q�械��ݢ1��ʦ���9��adRL3ؐl���eU�&��n�6����k���c%�W�bs���}�e�mkaxo,��LH�\6�.�wI`j����=�>.��-^����!�}n���'�Dh��	1��Db��ss+>d�0؍3��*އ��9����E��6�C�v�tfU[���n���q�t�X�����O���7��k7��'��>�(u'�������`���+�ZC��p��<J4T��#�=h@=��S���δh�TX�Gu�T�W�[�]�at�'iQiRw�-��̲�X�$'n�s$����=�Z]\��`�Z��O?�����h�G�޳����[�[o���a6�&|o0T1]�P]QQBeJ�M�V1eA��綍�������ji?[�� %p���rK6�`��y�m�g�����.Z�49��`Sd�DDƾ��̮C���~�k,���;>�[u�o��_� ��/V�@;�c�<��,}�UȇEv���{zr	�=�S-��RO3׊ەS�܈vx��d�},E����'Q�} S��Y��=���mjk2iwm��\e^�|˼��:�fIF�ow|���+�������ԯ(o׬D�p��s�I.X�N鮊ӝ��5z,n��(5�%�?x�������*Y�����@S�@w=bV}3������ᶠ@�V��a�p�t$0�vD���y��=G����-*V��r���!-�%���X�ӅhST$U��]Y�0���ݻ�>�̌;�13�t�	�+��z����
����sb��,�����P�J��@�G���Vl�l[`5�`q�Bi`ũN��F�g�w�f�e��g����1�5�����Vsz������L��vR��z������Tٵ&=���
�H�xq�*K��syN�����E�9-�1ݪ�%�pi�Y���z���}@9�ql�R�o6D�;�@vi�܌$�v�5��5�s�,�s�V)�:]'D��JHac�$�'i�DؒZ���T��gd��H+�5����x44��O��<��;� �th���	@�ZԬG�B�h1S������t4�?��9��e��K��Ϭ��4��W�c�*��M-C��}5P�	���uR7Wk�����z����l'V�VĬ��u.���ɑ#[���f��a'���R��Ɋ
 ��.�����cG���?Z6bA�|"a+�D3K ��$m�CZ���������P��Ԟ�K�g�"�T��Ů���
; j���'t��Fm�d�3�˽c�:I1�c)D�a7�ڎ��������M
���V	�8�d'��$�K�5Xn��7�?���wXT�1�sL�g5�{��hQ����(��װ�`S.I3T�rG�:�-u��Ϯ��)�ųk��'PWT��(ɜ���$�Y���:{d��:z
����KT�R���<J5���7K;��� ��v�l�rc��*�˚�4��M�:�6Tg���_��v͢�/ F(0�s~y��Z;9��I���YoUEj�0����G@�O�c[ϮQi�5�	�Ҙ�0�}�R���8)d
8O$� �d��x�y���5�?����%��n��s<��/��_ɷj�Z*��vl��\ޝ<�J�*�.���� \h2E}���c�	R(6k5Gxp��T�� 
�Լ�b��<��ƻ���˘���K|^]��I*wj�k\^'�x�:5�݋��ӧO��/���w_}��
pJD|A��&��G�>�?�Y�)Y~�§���Y��5�k;;�Ҏy7~�D= E���!�:B/{AY�<E&3�D[�������G����Z$�U�?���٘���U )��#&f�6�Q�+�P�: Ϸ[���
�=�?�JP���O&�>"0���Β���Ft��+	��*;dPY2�k�M�j&^q�g�����r�"���z�(h7R�V+�Bua>�������1�ל�/��=z{e�5�y���?N"{&y��}&��{��f�Iʙ��~N�����N69��Օ;�#�UO����X��:=hL�Ζ )����`���v�c��W<�HXE=��XD�FZT���p(j���˖h<jt��~�ճ�u���a�����d����g��ݹ�(�C�پ6$#"���x�ⵊӡ�LjAxv��Obq���2m��v#�}^�bGĔi�JN���-1z�0�����6���W�':�Ija\ҏ>��������o���W��y�>�n�y^�|i����]�_+`�nL�E)�3�fy�q$�9l��MJc&5.�aq�:s�<Jrkf,�D�Ă��m��dI�P� �E�	dm��'����#�������MH&��G:�w܀m�ѣ)׳p�Q�T7K�f�!tiWk�6���x:���O�ӟ�����������K��۠q�(��Yˈ2fq�uY�H�\�M�[�l�(�T��;���
�?�yD_o�i?��io[^��^0sŞJ�XӉt4xk�a�=aHq��=5��8;�y�}�����P�Q䤍��ݻ'�ֺ6b����ms��O?�Ԟ�<S{��1��mY��h��CJ��~ �����9�m� ����^�R�3�<#A-�e�.ZS�aٛ�_�TEJ �r쫡����s��̠E���ždq�i�}7�TJ���n���'�e*cj	�y&0cﱺ1Z����j����;Q��	��o�={�VJz��g,�."&Q1y����_�o�}s��������n߶���������/^�>���R)�6���x�J�����S#��]�l�v��m7�
`Lfy����}��[�9���(�lI�j����>z�h�d��оu���n�͛�,��WX��΂`��d����%��>������.\��{�Y����}3���	�K�ŲS�oĢ��[�00E_������{�����������ۈNA�p9�%�J�jŜO +
D0�������B�� YH�L 0�)��L���i�d� u�P�ؖ�yK�kX>� Q��N�C2�k]T�kƦ	�lK��{wF�C���y���ԍ�F�g�#d=�6���}:6j�^n8�g�=W�u�e����OXWK�Ga΅JHĢ*[������R��(��rC)fgG�[hEC�����F��y�hӗE�٣oN����������B��R�*����0��/I1kj�3��Bo�$I- �G`Y+����̯�׶��E�I����u���E`q}�ȣl�\_���\�}����8��ho�U /�
�S�����͖�pȿW!,�F�E���c�!#:R�0%�F�5��瑤9lQV������M�<y�?��9����P�)=��eʾU[�F�t�Nfe���q�(��f4�Vu��H����Ջ�������|yZ���xt�7[�wm��S����U�=�Qj'������It��U�In��;[ۡ�[X�N/ȸ-H6I<R)P�Ģ���pP��k@�Xl����\�'�̦�Y,ԉ��d���d|i�h�W��@-5������o�ǒd�t(��q�-6"��hǘ/ 3�]yYY�Y�����v�6�ᤌ��(,܅o`�z�¤�}ʀ�⎬�yj솆�#�ج��l�#b@ ��o���P����d:��ɓ<�x���6[�=E�=/��^���$#��0�x��#F�7ʇ#p�$ �9�����C˒..��k�Lx\�k�!䅭!*�s��ȶ+�W���������v�̂=�!�X�\�[�ζB�i��)�߿e�LM������Z� fc  �=DC��U����*����ݻ�����/8z|�/R�6�v�ݻc����1E]��ئf��B �.'���
٩�$;��͂i3�<*K_���\���Sps{3U��7!�2��Q���&�-!��cϯ�S��X7��Ae0q�^Q�Ŗ��HA�N�*6�Z׿�/���������r�U:N�%��4W�x��Ll#���oa2�ǳI
1�~B��t:��*����HNv� �-U���b��[��z��uB��e��,M]�p[j�'��-L�$kcKˋ%cJ���J�����X�oT�ox��d�4��8�G,i�qD��Sę���ja'h����1�U�DD�����!�1:%��mq���M���	��˗��hq�iZ0m׎1��s���l�8�����%�]��Ԡ��$�fzVg\��h�y��L�Y>b��T����!��7�sۣ=,���K6���aE[���>��4�k��*���堵dR	
�4ͪ:M��`�1��u�8�����������}������r��6޼$�b��6��_�P���hoq��r����ٜ(zp&����;O3r��[�6ROA��9��(b�l/yE�s&�ڕf6P���,���ů�˿,��?��?�������;�����_����ϭp��/�eNA�pJ`�Y����L�;��f�
�c]l̸���������܈�-33tyV�D�Ro߾��/��R0Y�ee�([O�rѲ?W�Hބ��h&���zS�~���~������TQ7a0܂��3i��9���G�n1�L`��ك����ެ�����k�n�޸���k���m_Nv	2�jip�D�X�9���2.�W]�k�-	n"� �[��V�fm1]$�/���dͦcjYT	�2s����8�����D-9==�~��`4Xm�W�K�a�}:��I���Gid{��|U���㪪>|8� �_����1���>�6g��ە�.��0��B��	�ͦicIF�縘�ޞ�^�GK����{�
�ぅ�-��uQAq¡,S��<%-tg� �X�N'H1P��k�)l��	]���ri�`�ŽyCys2e�t��yA��ڞ�;y}T�Z��^�������G�>��%�� �usD1f�-JH1lj��B1�';?��{��:�MTzXm��wv|�xp�[u�h��ir��J���Ǟ�)v��r[�t�"��� r���Ø^��T`�k�)��ނ�lҏ������۷oa{������޾91�̂��d<�D|V�uz�z��
Q���f��Ϸ�f���!�1�/1�gK�����o�m�TZm!�f�y���f<%��ݻ�E��\��5O�t����@߬ٗ_e�͞
����Қ.�4K�h�Q��8L��0�+l��5�~c�3P��5�]-U��"mWk0qtq4	NbN���'��_��������b�/�@��)y��d
,N�+���ic ^A��lJ��������R��庹N��9���ޞE��m�^��jqr��T��V�o�z�U��==;�[�ڧ�zkF��+3����|�[=���lz�f" �5n����=�o�r�1�N"`H���s���F*��u���DB�w�6�>v��/<�3�C�
X0!6�i����f"�!�8�ړ��+j1yav��-�Z�,B�E�iכ�^n�n���G%�f��;�IOa��*;Ƶ%my�Z�m2�C]�7o�h{D��I�[�U �ć`��׋hڶ�7��#蟂+�r�KL�����F�y���z��kjy��oo�'���K�GKGF��Pz@d�$oGZ'�hI���h�~trz~y5 �d��~n��%�����p4_Ν9�K�EH�S��1����qi2��זZVe�o�m�؍`���fa��U�G�A>$�Y߿��Gپ�����feQͽ;w?��c{ݹs��3��dq,Y�jkahX��ә�&�57���f7<3^ W�:	Y����{��nI�Z�q,|�+�)4��>�������5��أ</���\�h��p��rK/�2m��Tj�Y��%��NNO��ucV(
�nD��V�L}e�c=���0�{���=oQ��{�'��G^^0�F;�o��y�P�v��}{��P�<x����P�ɼ�N����j3 E���o@�R�.
��e$�X��C�y���-Z��ᡫ���g����������RHD��V�ƁW\m���A�-FK�o��]�����뭡Q�������Z�ċ�@��O
�
Q�bW#�����Eڣ�W(W�G<��Ώ����Hz!��,�>��fBQ���V��<O=~
�ڪ�qa�`8m�Xk{5�$��G�W���"G7��	gpehp�R�Y#ߘ�0^������,�(6�B��.ٳ��ۗ�"`r��=oK���?��1+D��v]a��G�h��Ж,n4z���d�Г�����@��!S��b��-��(�:@����;U���Y����Ҷvd�P{�a��;�� ��ޡ4��IX��Ӏv�Ї=!�U�`R�^�xa[����<���Ç�դ�7<7�X�E����������INǐZ@}=�Ǐ[�2�H�\�	T-��(q��IȚ�&�<q�T�W �H�i�uc+1Юp��-{+����;
E���
��� +(Y;�eT	z��Z��PC,����$+d�u{��:�2�8Pg
d��E[�j���j�K���`I�E+ *�-�0�)7�G<�7?N!4l������[۰�������^�f�'%�e��dr���+5�D>0Ftk��B=����h�'P*�?��?���϶��H��u��^L��x���s��0r�#��ڸ:������o�\���Ŭ}+ I==�s������e��92=Q)8�O�/�w��2���k���b��V�N�֪Tk��Ö�V{�#�K�Pޢ��|%�L��|	�4�#�}$��H�#<_����W�y�G��J�����$GL��{�#�s-��Z%��Mcb7�\b2��~���/���/_}����Vc4�p�}�rNg�*�0zq�6F�zS�f&��C��k����xfn5q5� �����wb�`i��(..�߼9�ɺ����o��Zh`4�����<P�Ja�ɞ�D�>����<��,���D$����4�uu�
���� 
$��FP�1N���"2��d��Nf���}������m�)�M��i�ܟe�%��Vh��
��[�r���C��]�F��o#�k��u��'�ڢ)����v�D̍e��9I�`+J�j]�P���>\�6�6�	C ��~��~HE��횰>Z�۷�}W&��e�q�Y��s�N<�IgY���3��ā0� 9�B���cq�ɪ��iBMc۱Ble>_@���f1��C�Jx��b%@k�K���j���:�@6W���DѪa٬������һ��?���*fh���?�\N��K��:X�]3N*�М��Ο���K!��(ɑ0��>J�	Qh�ۂa�����-�:�k� �����m�FT��~�D�Vc��amG=|�(�����d7LΒ���&eh��܊VX��U����쇯_�V>�p ��c��׫R�T�hW~�xU���x:{��&n���#�������P�2j���ju6�p,����������� �/�����O�H�J��g8��/��hC�9��y���,��!���0S�#��6w�c���;����3u��m
�J@�d�(�a�V�ZM�����~FGϢ���5�,��=+TU�-��3���}��0�]���_�9q��=����8Pa�>Y�@�c%,�)�0�&ct�k��WV߮����Yܗ�c�����r�v��4g��H�����^GT�3�|���w����מ;/�]Ϳ뇜Iw��v�ݻ%��3��G���U��:��1�I�r��$�O��?���V)�ZJO�{�[�q� j\iw��;���c��0�)��]�5!��X�
���޳����p0��|���3T�F����0�K�5b�(�<��"���ѣ�J�f'����vMֿ�
��n���ߚ����+�PbK���F��&B~eo\�):Òg�hF�h88(���M�}��+����& c}b�8�y�o���}�;��NN����g&J<_u(��^�� >iwYS��{SaL�9�!{/2�(P�]$H�	/��i�dѷ}^x��������0��d�߿�0W6N�SEKvHtVEx�s��W��"z����|\r��\T�dǎ���9�6��������u�}{|�����ϟ��,�(slѥUm�#��m ���6�A�Ж����*�/�-��;h-Ĝ���=d,�/Z-0:��ZA֚ �:|g��L��j�f��fd����3���T)�0����.���!Y�ev��Ѷ�t�"�E��Iͬ�'գ�ukzG�?��kI��§وְ��~E1%�vۚ��|i�P[�96dt6
�"�R^0�������	[���"T��R`x�`��#��um���b	dx8쯽��lӢ,����j}m�[N�oCΩ� u�G��D�ɸ��i��#��Q����$�?7hk��*^o1GoIV������[���A5Ֆ���|��N�2��z���ytUH$�c�B��z�];�+#�1E������xV(IX�Ge�D����ei&֛e�b��A�D�����e cG�'gv�����Yc���<�
�H���ЖS�)��5�'��9�`C�����E��պ �\\���c������S׷�+'TG��z�^_��ñ1�o���+��0P\�ј�	��:G2+�����M-B ��)�O6{(3�RԤo���n�f��_RŲ�B��:*���=�@k2���ԅ����Qz���mu2#�:���{߇&7�V��޾9*�9CaZg����Y��=x��F'㞴��TmD���q��Y��Ѿb:�Yhke�h����o��@?��r��G��.9[:D;�nx%���,^�D��a�:���!E	y�.<P!5�����@��������+�E�W��~Ë�����)ʺ��ѕ"�H�/_�Q�.Xk�^z(&�b�HN�s�|�U��Ed�
.�hqT��/2/̹]5o�̋��)�G  H���TN�X�wLk��0Pʗya�֑�$a�ȶ 1Ðu;�Mv���ͽ=�2�wE�JZ
R7�\H	g��qr�^)�U6������������v�9�z;���mg��q}m�
�t���l=b0�!��5�Z�ժ ��x���{�u
�\ܫo�c����f<��U�hH�"Ɠ��,�՞L���i|�)��~�x�$]q�9&��b�dFuLF�
OX�j+b`�R�B+߃��h7n�����&s�+��R���lw�1�y}���a>z��˃���x
����K�/�"P��0�9� ��XP8�Ň��Gz�H+F a�2�}���]�OѶ$n��I�D�v�}2�C�����+K���K���J:4%��[�F�^����ذ�f��2vDޝmB��X��k�(�sqeḩ��ä��������8;���W��mץm�<��*��p%�LFz.d�'e��А)?�]a/�����u�h�-Xa|&n3���Ur�G}g{ecƽR�����(K��kq����������/^��"g�����Oj~�Y�2:,��b3S��ҧ �MGx��ե���}��d�W��>}��9K?�����y��������Ŷ��D�<2m{�b�1��22�3U�f���W��Ew�o���Q].������gy�M�o̸��S.[��\���~o�������}�'�|"��X�,rʇ4Y�=��deO��щ]���o"Dn9c+i���/��;S&i��>�o-\�F��IY%�lx�6�^S汥�E�l>EմJ�T�ZF�3d$;�ɍcʢ��<B��7�;a�&`ޝ\?~ڲ�0�;�r� �!����̿�6�?����؜.�3q������N{���;8���,NKr�x�����lNc%Ž���IT�m&����v6�H�(@���nJ��G3��v^m�M�'����W�G��4f����S�qTD�_��m9�=l��4�0ʈ5U�]U��� ړ���&�9� ��F��޽;��ٶ�͗_�q�pyfG�.i]Ւ�)n�'��Yڝ�n_���S��CyWGf>�V�
ǿܼz��
�r3/���20�) L�&N�(M�0�mJcR�g�̳���g��13��T�2�Ô�*�Pv�ji�3��<�aB-�EEhJ����/���^AUHcп���D��p( ��Hq�.UYFGx�:�?���o��������̨��	��2���I�U`+W��O�pOb3A�-�m{=`Q�lV�_Rs�I��v�-����� O�;�@\���ߝ�v6��ma�1�P���O�~���?�m�A�ތ;��B\��t��k��4_��fV�>\l�E(�-T�p�ӝ4�:�>�P�Þ]r�X���%~���+Ԍb�C��E��Ɯ]_;?��l���"�Ps��[3�]���<qMo�d�}ρ���ٽ�~�ō�,"�|ѷю!�ލ)��p�w��;���`CAW���'{�A���\`��!�Ձv��4���(�w�nOLצ@94�N���Un����D��I�����%�n3�
���W�U	�c1���TD�R�i�$j�����m7@���~h-��2� ����=q�1��W��Ǐ��Q���g@��$��lcڷ|�5�l�)x�=��,�)#�Kث�T�C�o���y������4
�{�.p��"���{_��}!)��D���"���=j+��Rj/���z�V0n��@7t����$��U>��ҕz���F�Y�Er��1����C�,տ"�|&�
Z8��o�_Cy=�
��fI�뺬�zyۼ7� H�E�h��B�`[�݊��lS�	�����Ԟ�{��̮�$�=μ��ʼy�s��Ts�V ]`WdBM�LL�r�ծ �����x��ѳg�\ �J�1�c��:�a�y��9�,��7��_��nZޛ8�Em�P����e1�BNg��/>W��Q�����҈ �<��ǊBtGtǁ�5jM�]r����9G'g��8l�Cd�
3��./W�#9SO�.��%�NCf���޾}����7�W�C���Jb���,d���g�@>+�K�̨ؗ=��K�ò�4	�4E܂��.X�0�v���p(��c��&M0�@��� (?��@����l&���~�%e�`L���lh0lj���ߐ��	����2ڝ,d�) rN��H�Ui�Z�8 ���#�3)��h.��̌[6�,�O� �l�EU� ���n� �\S���׹Κ��<9��h����4h�G'E!D�Xᬪ��o�%:CB 	��AIҘ��8|�06�� /�,�Z�9�p�aY�q6���֌����]�*d���h���e=��`�Ù/+�S&G�Ǝ��n�Z�7t���L�6��\�TbY �J@8\3����Qxl����cbs�YZpŲ�����ť��0ꄹ�T�"�oJ�ޢ�f��.���r�^�		?eA���̀i�'4p�X"���Ům4�p`�+GLE��˛k�n.��`a��U��IA?�37�l��K��,�9:f6�����鄘�*�H�)�k�M?��-�����իWi�<ȴ�y�D�L��`��y���yA� fA�B�V"�R.^}��PҘA�۴>?�\��r��f����U�hy�]7F= v���AW@����ܗ/_������W��$�����S�ShH�B�F#ńMd&�g���I?�,�A�n���ؼ��N��du����s��ز2b�1�r����ƪ��b��H�l��*�� 9�]0��|3#���4|���'���Y^ί�����nЈ�������uB��,@q��>�I���0P&��D�75��c�P�@�Ӏ6xecB���ϒ��I�&&����_��w��8}��t��� Y�^f�j�E�0�Ȅjܾ�>|��ꫯ����N�SV��?�\AipX
��KDٷ!ZyɌC\"��(c�O��n�=+��c��D�s;9`,:�nҐ��=nY��2J��ĩ�~f���t���^�xA5�X�7s'��e��_����ۿ%�|p�|��N]-_K���p'�[���ֆNL���))r8j�L<z�s kP}�Z�2���:!��*:�>>�����Hp!!��'�h!���M։,�@xy����߿����O��?����Π3|�?.�(WǒUtފ0is�Dl�7RI@.��K
��[�s��=�X@/�2��mP��wl��✼��d¶é�0wB:��\J^Q��(��!8``��z���O��-g������g���<����,A��<���v�f�H�N��/��_�&��,��|��M.�2�|�|�k%��"B�灖Dr�����>�ͩv��:��BːV) y�$%��1V����xp�k5MC3h��<G�N�P��������Q�5�k~���1��gs�@M����A�����ed�ĳ4-3���J��32�DM|z��g�>	�GwQ�r��O�<����kt��<� ����|���_��T�*�=l����2��y����}Y�T�y�m+�|n'��<ƥ�ǟ���Qy���6t��D��e�ܿ�
�z<~��6� �T��4Eo��(�O?��,�-��q�޾�д K��!�����/�������^����t혧F�#�	"�Τ��CǑ��0קxfx�(�q��KՁ�q�G�5�&j��aL�G�9 ��H���U,�!��O�0�)���� ���&��G/*zrKM����0;љkr0�`���7��4�̳	B��O��s(�؎(�4�1J��ԉ{�ώ��π���e��$����|�B�����|�����2+��~������Ѭ���g����/�D(���$�O����?�[��~��7�THm���Ԭ�|FZ��H�n(��QT���l��Wz{T��&Г,�R̢Rf�L��EVHG7�x���cu�0����!/�!�ğe��D�R�!R���T���ێV��/��Sו�R�!�v�a+��vs��zז~���~�ro`bܡ�����,���Q\��3���8ĳ�K�pJ��W��%�A�M���d�Ͷ�r��'�q}t�9:>��1E�D5;�+/D�t�U�{B�S��fۀ[7��,��� &aMD�NU��M�:����+N�O�A�&��1��2_=����|n��Jl�1�����k�&����q����N$�NXlKY����d�����G��N�J�>)�s�Z+�����������.�EU�D�i�yPtF�,�g�}��ɱǅT�Q�E�df���F�|�"�7�җ��}��VKS�I�tK�$h��j�hFeOD�F�3��q�*y�I�sqY<�k�l"�{T���o/�E��j���A-��ʥ��#LjW�9�� F�����w:C��r��3��ɁȗH��Q��>I�t�������� �F�0N5	Xs;@����&i�~�v��[�\����zQ����-6T�Td��
f���L�;0$��_t�h�4,�����Uك��I���|��hF�&�
�0&D^Y�,_�p�)̓�����zR��N��]3��p!�Z�%���QÄ�����)ֆk~`��J�}��DӎڣptvF;�� ��>`��f."����Q��!�Q/j��pU��%�]c
�gn��L�ugA	�B~S?�M ��t�Ad< %��%F$�L�X�&)�<؋�_B5�V�'����	ܒ2+��hDe�Bޖ=J ��N����,�l���D��d������*��x�N�	vL�Xټ����9�q��c��:*���JgltE���N��P���Dw��ȏ<R��z��"�;tp�w��S.�����o�u�����ӧOq�u2ёb^�l��L�(jl��:}d�-������h�q��+���S�v�����gj�"Ix� :��,�<fЬ:��S��L���:�O�ʺX���
�.�O�nw��l�~�C/�lh��6"�2�n�!7�wV#ɍ��Ա쓙���=��`1&��Ŏ)i�de�C0ߍ���Ňb�N�����Eq��%{�+�K��\�e������r����ঊ+T�V�8!�_V��J�=��O���T��L��bZ� 6�:㌼�*�6]�Wl��f��r�t�׫Wo�qz��]���|�駫#wus��ggg��eC�Qo���v��!���]��v�����ե�?�27��LF3�Z<��ֲ�̧f�)Eb��ӲJ�E&ў���'&�C�@�T%��~�.p��&O�X:'��:�3y*�
ڍn����o��N��jU���+	tѦ7`v��O��2aR�J2D��(�a�]^-������	Sw�Jo����!����u���rW���zyt~���;]a���85�*);��P�L����"�CO�Ӈ�B�"���Pn�r��JYQ�8��ɚO��7
����-��ϟ�p||��~͸�o�S;b;���L���0�-��ʊ	��ɠ�#�����eh~�<ꈸ���ϯ%�#�>�4i{�`"����2G�i��r���NA�c+�,�%�}����o@��.��x0��i%P+�NZ�d�X�����������>??g�]n���݇��Em��.�b�j�K̫��K]9P�zʑ�������+"��d�Ԯ,LIăo3�B/��k�\u=�̼ηۻ�	������\UO?{lr0m�[M��$�!�9�gj��N(�h6�g�nb�%1Z���F����Ѯa�3nC���Wo�.oĶ�߂�2Y����%d1��i��0���L�K��vSߥ�l�|.g�T������ϻ�5y"�n���Y�srrp������ak{���T�$�XYmW��B������<����'���m��I8� �H�e
S�l��� (	�s4�VS�L�K��m7�ĵ�W��c/�	I�i��TM��$�G������S�Z%3���>T9l��z�b�|��G�`N�k�X%���m���X����O~�ӟ�~�X��oW�
�L�ǳdQ�K�z��ٳ��������d�1/c`Hn%�Ov��V��c-�'�`V�U��(�#zR�-�%%���䖆ID�9��G�y�P�Y7hL��8���^1A�@�#'�9N�:>Z��Ӡ�=��֗���͍<�b��哃�����.b�%�ȵ?lc6-l�&挋%�x�F��1gf�
���Ǐ�"a
�B�Zm�}�o�!GH��ۅ�g��1K�V2��o
 rHa�}�e�\�p���I��\����Sw1�,IS��'ad����M2ɤ���Y������˹��rQ�{��%}�4�����:y��W�|��N����fƫ�-�3�"��g
�q��Dw[l�hi�J.����9f����F��ú��0�
t��KS����d֨��!3���7�~�H����Y��ߌjɮ�a� #̛7o� ��^�Z�}��N����JM��[�ţZe�y������\n���b��e�x�y��$�y�@�n��j�UD���m3K��<���i��8vu��^��e�=��WW7p3��h�/^<|�HT�f���:�A���US���-�phrDr D?B3�q��E���ݏ��	�6)xd��㎛,�U�y@��2�QQ�К�E��^2���躏+�{��Q"p�2�R�"�/�R�s{��F)i�T�j��M��Ƀ�=|�i�uW�l����^m�Cz�Y�a��WLgě��������W׉���Z�I�c�Z��!�^<�&�"�*V#���ň�1�q$3Z��m)O����˗1�@�1�;�@GdG�����������59$�5�[���E�B:�5v�PÃ)�?M��G ���m� O�F�R$܏z�E����v���g ��<����L ���ai#ʲ�24Z�B�ʲ�E�����a����JXI���gg�h,�$��KL�r/��2�~*��+ϊq�G��iw���	���0%�S�:�������̲�IHR'��կ��ubf��G�w\�g#qL����D�)Ӷ��=�f�l�h8)c��)��o�vO�N+3d�lx����U�e�����#C� %J��G���SVU�yD�?;;S�[�*Z(���rQ�F��CLp�EraѪ�U��z���D+j�"'�~s��S��,W�����>�M�66�c��w�?�o(*�e6�Tƽ�F*��<}O�����!�d��d+�_��r1�Tb�=���FŌ,�5�;�Z�m��Nty{��A��(uM��:��#�!�R R���z���[ˡ�*[dah&|!u�&�t���>����X����<�@�i�\�!05�ʚ�@x����(i���ԙ�$�Х����i��A���ٚ��Hs�@iFrJD�l���*����\T&��9�IزZ����E��I���� ��'���H�hU���`�i����3W�ҕ��F��'�͛��b�#���ߋYd/�rU��D���N��e�[�_��n��}�ͦ[.`������X������Մy�|m9��r�g&�J�{�@�����C/7/�|��*����[+J��C~�6�z/����7Z~H�и��z�>Iur+]�Mh��t�ܻ�!WTϿ�~/K�^�`���A���'�($D:�t�S����`��799}pNjNBk!{㿀̈Z"��]�,%����,_�NON�b�"�\Sx����������ʍ+��v���k��Q]Ә�$�U.c+*�)���^��S���=�����N�pE�*2〇�8EJ_��`q<o;����޾}k����Ӛ���~D��(Z�œ���k�%�n{E{���C��}�Kn���t�dg)���d.�S#�Qi��2�5��[�3��r<���'\
X��(~��W<e*!FC�,X��"�IO�o�f�OM F�s��%n��~����,���N�l�|򉬉,�H��>V���LgʑD|x���Z���r�-@�$r��A�R���0'M�L����O�x�<�=m<��Nw���0ѽ�;Nq�Ɵg��t�	�)�h%i($t8k?������E�]�3�&ҝӪF��[J��W��8���gH��gM@CG�p3��-t�^iO���+�
�~��Y"B>-���Aksm>p��/���%��g�?�߈-��<�ϛV���p��I0�Ss�'���qD��]����opf��ԓ�~�*��t�C�}��������A�;�5�մ�y�=�*��PDz�X�j\=X]\<ܼ~�Z��ի���rV{YeLJҌ�q�C�����(W"~��<H�ܕ43N�1�	���kFyREP��n�����!W��7
ٻw6&휧�uwƽ�?����q��~t�L�������B_�l�����Z`�x�8��)J^�?�!���<8�W��ר�Z�����6����I�H��u i^YI8T�Jk�A����(�'�5�vQbҼ�4�5�.�V���"D��B�t�u�����]���9� 
�rDb1��㩠�d���ې�:c�v��3:��q�[(ߊ�� �Ic�&�����?2���[L��&��6�ôk�u������V���O���)���O���Y3�@�G���y}S	-onnd1�[L0�u&ޔ�jW�L>�Q�
��r�8�<����/��8�?
�x�htm���sٵBޙ�Mͩ�,���^L��A�{�&b�S��m7^^"�{�i~���GQ���ܗ�^�W
��L¦,p�.V�b*NO.�D������Z������;hg�s����|�ƃe�Ho<�?�BQK�/Tu�`��qp/3u��ͮU#�n6;%��bf1� B/�H��js�MR���(��v�զ?H�`�,Τ�m� uT�,A޵���ݑ%1��)0f�ِV�jU΍�9��X��ڶ#!�������kM_����v��[��\�\K9���J�Or4FE=�MBV��v�`/���i!պȼȿ���pX��RZU���wjP�%��iwg��U�<�g�p�t��u�x����h�)�K��$���ZM	�Q0�;��3O1� �#���,�Gė1"_,n�8�����h����3�{������ypP�@Q�SB���lw�P˙�I�������e��Ћ.(�PTf�8�C:�jP9NC,�0��\]\���t����_�!24��3����ֺ�"�����<G��z' �v+;8	�(T������qP�A$�^�·����`L2;jG�B>?����G�0��$3p�c��h����l�`�AL����B�op}����;1���g��)*��/��C*�|��U�>l��Դ)�Ev�i��|�Y��3#S)�Q⍬ ���Ai,�*����!�nAZgM6�1r����侸 �����ޏ]&�5z��d�(�s�j�l�M�v��GWm3������^��c@�5�h�	��8�	4����4�A�P�_�G\'8�����K�]�֩���#p�T�l�4UKZ�Q=o�wi����f���Kt'%��S�wa����٨��Y��nv����s��ƀ���n.W�$��Ϡ� P�s���MW�!_2�i�cE'��c�ZeΔ{�݋�a�#�QA.F_���3�p:�!/�Q�<GV��N٭-�����dZG�����]�O#h���	�.�E�t#�ɡ�E5�b1G��f�������rËcxq7�;��8��>�EB�����V;QT�Ř�+��O�d���L4b��OV,����9_Pg.�:��$�����ڬ tf� _8���Vy��y����V������U������+m9@��f.�=�O<_��]��e��!� �8��4�*O�Ԗٝ2B��{y��[LEj{��!���ӌa,!�|�w$JR��|Z$��"�ނ�`���=�	:�1�Nu+Xi̥�L�R���4�����0@I��������9�O�֑���8)d���:� M������n�P�$�%5����!^�a�����y���*o;���*W]޵o&���M��)'a��RTJ�� ܡ[�8��j�t;�r�E�w��5`�Ty�F���+Mk֕����n�4�_~>t}�L���՛7� t�?~�x{ww�^��tu)������_�J���J�ľI�x�{`�e���xv�����n��c����᳴#�Zrey#?��`#W+�Ð�v��A=R�@f\����6ɫ�[�].%����$`݊��v��Q�wD�\�FT��'� ӹ����9����H9@AS���~ �

<��WoW��7���������/��2ּ�f�6U=۝'�w�
��g��(���۶[L��x�]g��d�r5��D��Pa(0���)�/yOUԽ��;1{���T��,��8e e�D^� OaZ�		G��X�qa�[�3�E=���犆R�1q�L��h(2Z0���+�Ǚ�?���"����$��S �LtS�={6)#'�{�և�a�iq	�TK��Ww�!w!a��4�z���'^�F������郳��$�Ro7��Tֱ3Z2�����O~��_<~���͋X�S��@����d�H����re2���0�O�~Í�Yzv|��L�PrtK%$���k��
 s�L~O��l�PI�!���8?ef�YZ�_�M����Nw��'寕���AK@19z���x��:��kSۊNI�c���T�a��FO�n�"g����2��n�v��ɾ)�3������٤ZӖ��ken�� ��ζ��H�D`�d.pHѪ�4����0����n}�S^t��H"�QN /ͤ�K#
�p�(u �BC���uLs��ub�����Υ
d%aP)��r����y�$	�O�y�`�k�@��iU�#칿&P6S��4}��+Q}$����E�څ�.� �Q�ٝ�R��wۥ�.՘��2�u(є_D����cDD'x����Ҳpog��3x.��c2˩�Ы8�$������ӟ�Զ`{��J�(�&�`��m�v/G\q� =�=���R��x����8M�h ���B��T����j>��'e�I�'1�&�ޏ�j�rNQ�� ����_�Y�ba���O �`0�h�Hh��D4�\r]�;L�>q���I("֊-$C6^__���sSDf��^,jDb��C�}�F�J�.�n7�ͷx
�z&t�Eu/��`��8_��I�:�r9b,3,�-j��<Ͱ�z�ڝ�@���)פ��;MC�nc�����p:�p�s�/��o�@���0�4$>d�]���������hb0"�Jwz�(?�[�' �n�h`ғ�GB ���nѲ�%C!L`q5�F��H�F�s�RA�b�����*W��0�l
�-�G��z s.�����p
����B���A>���JY&�<j���LA�z�jq�K�qGE��ԷW��E���q�жS�<����I=� ?�"q�S�@�Z��wG'+�--N������D���S�x�����0�4r�d�Ȋ��3JW�e�af���@�ӣc�S���l���~��%G`����y���;���M	-������\9��Z�&�V�&�D��Ws�ѝH���3��X���)���(�'*�� "=\��eڻD)�����zդ�dK�$=��A�R���tR���!��0
�Y�p)���g�Ui��"�l�\n#Tp2�Cx�D�Z�����g����w�r=T%�(�9�36�i�"}�˴9����%g���b�|��so���w_���������
�CI��O�I���b���n >�BU��%��F_��a0O��F��C��A��y�	�/��߷]ӳ�W�2�t�}5��A���e[��K���"؝�}6S�L�^\`�z���7*��qM����{	�Q�"�Y.$�����!�1��0��q�t�=2�)J��پC6���1Ƞg�Sφ��\9�&z�����*�/���h��˗W�%T�f#�;?_)�£�;7���S?K7CG�;��C���n��`j,23P��
*"���"�z��B�P�*�Z*lv�0j�}�AV2���D�ra�E���΃#��U����Uv��{�
�J֒eXE��{B�HuJJM4�na%�~�G�l�OQϛ�h&Z��wD�D����1z��%%ꟈ�D��5L�ڀ&��b���A��:!:�./�w���0_X6��*Hg��у��
pKU�[�
©��h�#2e������ecv�'b�lx�����X�2��i�� Bm�*�0�ZD�a�VO9u]�`ޝ��^��nw}~q~����g���e�.�����h��Кt�y�F>.�z���w�F�aoZ�ltW�k��Ԭ�fy���ģ`��*�,�ʠ��u`������h6P�Ҙ�=��������	@��H�"�I�I�1�c��NZ�^� 
���˔܌��L�ŗ����ʓ�Y��������dA���~��ײz�LqWUcx�JqŊof�$	0F*+?��óF����u�e�VKgM&@b��p���0	��qIQ5=�3f���I,ytA�)?�1��!y������Ѹ��I�<�I��чa
��<�:K���_�-q���1�F�Ǆ�T��V���<y"�*o%��g3��ʤ(vʿ���	8����S���b�hK.�Z/4�g<;{�(1�Md���̞�/��B�#�u���h:#[��Z�5���Ng��31T�oBFOw��b�ԙ�ڜg��Gz"M��@��Ʊ�-X��I�+����Ss
��஁�Hym�?_>�@�(c�K�
�7��H�]�5�K���O�O�.N��"��_��x��9�����i��ɳ*{|�@�A��w��e�c���9f4xtq�v��7��[�1tt����)�|�ښ��:b
8Rc�F��w��ݶk���&�[��Uc�sk��~��1�jL��lӰ�Z،a8����S�%��R�1���c��u����X6Դ�X���@�4��:�,����hC�=l}l�J� �b�#MӪ����L�j���;$��WK�h���S)O)�r�ײ.�}?��E�O`���o�/>99a$'�m8��G��4�f�C�愥Y1���'bl0>�}R��.�����V�v�0?��$S���bzW�x��#``{j�XC(�}$��/�� �m�`�6���!neJ@fѵcV��7���Ŧy5�|{���������m���b����u"�� �v.5�),+\W)�%V�
&S��Hg	�/�b>+���P�G�'���o��n��)���)9Gֳ��M�5�MH�[=>Ô�߀����V׼�ӗ�P��� JQO��K���[��'℈i�ۨ��Շ��������`O�u��?��޾��wH!9��ZVh)�c<O�R!����k�0Hg"LRB�2̓�ǣI��Dߝn������&?�vD�h��m<��r�����N3D�c�YTN��7���YB�z@-7�؛��n�D�o�tǳ6�O�����Qi�8M�]f�S%��8msˣ)�#�6<cϥ�걉�� �?�ɞV��7����˔�p���4��7�F��t�%].s���F��G$�Z�T6%y�qd1���M�
x�	�:��i{�3���O��f����3��x��v6��;�Yt�@5�j����!
�ҹ�0̈|���(W�
���53�hH}�f��&Q�~��E�[+;�(��J ��I����/Jd`;'X��������!�^4���LEqZ�0�b�E��syy9޽ә�~Y_�%�H�vºC^/M^U��i+4�{�4r+M��J[:+��K��'��m\���J�Kw~�Π�<:/?�����ֵ�l{s��	2��
?��	VҟtZs�X��PN��#�b����C�@��q�D��j�Bq�>�_�α�W�y��)NN,�؈^��<�,!�6U�GS`����r�(	�v��ڼ�\g�����eM�15�Yr�**�I������@��h_�<]U/k��2A����`n�j�<{IUT���G��`Є�k����谮32�&Kw�8'�"L����i��'� b���ĩ��2tr�� �
�g4�(�$�]�5C�Aξ�󳓋����Et���ժ��&�m;��m ���L;zy�:Z��
������ `s�'1gj���˴��̌v�� ��&���Ny�h�=�$勓���e���L�G�O:y�X�Aul1e>-��JQyT�D��A�&{825[�nw�N�Vt�����Me�DO�1�&h3��D�Q��#��2sM�"U$x�.x<i�V9�8�ݽ�d �F�Ø�T�ej��3�����q2�����5.�l���Q�l�(!���C$J^���ڵ0��N�n�w��忬k��ވ$��Sq�;�KE���2'Wu���˝�c}w�Y��U��r���&������#l��+�<$Dw[U^�t�*3ggGb��՗���ve�0t!Ʃ��Ē��7r�z�"�����s:N�7�Ȭ�+�
E��P8�������Ӈ�d
 h:�)��)�A8��wU�
������e^����ux�F�e�� ��:��iiv����d��ۤ������Y�L����>���r�P�R�tv��켺�"�C��G�c�Y�M�բ��cI�ŵ�p7�'m�Q����gh[t�+���S_c>N�[��	�wp]�i�O���V\�I�K:!p�1ˑQ�]��\����{Ι��u &s�du+\B�a���!z����A�ީ��s�M���:v�t��(���@�U���m�A��������K�aY�b���~���>�F��YU�L�8[���=�vc��G��,Ǫ�(ϛ��7o�[GH����O~��m��,挢��h1�C���{��gg�`F�����Q�c�ii�o�X�$9}����T���?%I��l�  �J�"���	V8�0�m4uH���~���!��j��~�(RO�3��C㉜��	�8��{M�N9����vo�o��Z/kf�0i+��� M�mV���}��.m����	c�}����,�P��A�A\Þ2����9����K��`��4a�wG�'O��LCw������/T@��BrkH���x]�����Ǳ�J�1�}]�@�D�t�Uzf�6�-ł����Qw��o�O�T&��K��6���
f	�U���9����W���	���͎iXC1�ݐ�:_��w�[Q*�ގ�Rs8�+�b�yt±`9� 򪐪�A�-�&�1Wxi�����C~|���?9yx�<=N�SS/'�t��O�\f&u7�i{�Y��aۉ���f��k`���9�}����r�H��H[�g�TL�2#�~uӬgd<�L��BSxy'�[7�����a��	IĘ�&w��Az�sd�������0���0!Iόҧ�~*���\dT�LR�s!��r�b�K.J!΋Ӈa'�x'��_���dB�'�c�,�f��q](�{t:�k1��]�Yo��p���_�3_k�c5y�bȒVQx읢���'o5�sZ;0�1���r�y���wĚȬ{�c\@��=)�����gW�O"-��(�T�i��Ɠd��4���ɉl��`�)���EN�_|!���믿��oXJB<����"��e�u�/�,�m[�f�H\��+��p6?~<*qFL��L�9P��H��<�*F�&�8��D+l1�0Nm֐�K�#K�/���I/V�P���祔�X��HdT��q`�	N�fa�y��	������x"~t�] v%�z�0�� �	zF��#9*&�]-h�&!�=~UU�=�3/�P�|8��SF(j���B��X"&FP�T�Z�(��09zPn�tƂ���봃Bc�i��#ά�%�� <�+��&���
�3��3:ă�'-y'�V�}¨��C���4bpо2���gi���#v
�+ ~��G�ŠN�Lvd����f���0�2��TnS����%0��>�g�<���i]���d:}8vs���d$=7MXYԁ"����cݘ2��+������[5ŞD�m�fL]�4�(�����3̻�L�l�z�������$֨y��:�G'+,�S�>��HKT)��fu� ����%��J7&�%�>��6�������IY��15y��@o����\YH�i\�h�HH^�DK�҈{�s���!�3	�Q����`"U��P/�$�����B���P�ᩏ�1��Xک�"Z�xp�ff��d�Jw�HTQTtOa�sJ����U7.	m�\��� ;V�YO����Wǚ0O�xy4x~�0�ą2C�Tw~Lx@(U4��Tw��N�H�@���W��	�����5����'7�e��P���Lq����R:N�VO҃��D�J�&u��%p��}�� ZE����� ���O������+�T�&©���+�`\m"y���Ҕё�Sr��;����O�>QKp�N�@=#:�j�ic�����Sj�)���F�Ϲ�1�0��#�q;!��Uh��u�.�'*ɝv����"�}|+߼�}����c�)�)��&\,��/���Q	��(F��6�p㓹�ˈ�1�P��{��z�릫��js���t��,*�hh*���Bg8�"�L�@�B᧗N��M��*�?�t��׫�k	V�S`���@H�zm��7�E+#���s��3���%�OyE���3�q�ˉ�V�K�`�\I�B����W���$`0)<��6�Rt=p�U�ǌO���Pdyrf���#�%��[� �)J�:S��.����կF�p�R{�>���A��3(�V��7�\�.�|MH����0�T�yQ����ܽ{��l� e� }�a(m"Ց���cp*�<ї������w��Gpt(�c`��V�U���*�H�0=dJ*���X��e�NN� v��c�+\��ŉ��*�g�Xi��9�'&�$� �yFA�F��	�FY[�1�.�p"ۡ��[���Y+�Z?�X=�N��r�:�Lvp0�a��v}��k쯢x�ԓ�!È*�<T�-+r��K�sy�m�׳@7(�~���Е�������?�r8�� �΅�U^�16LÐOx(�:��sѵ����8��5r�:������#L��r[�UF̲d��Y4�����ѧx�D�N���<m�s\#h�Й>�����3�/���@�A/b%&�a����Zk>�s�V`�(����H�K��0�I5����(if��#( %��G�L��8Q�LEuP�X1��ox�)��`|�D>����ahIX�y�H�h��c�h�LH��(`E��0�Xbć�L鰶�C�O���Vw��+�H5�n���d<���>��Ǐ�K >#n&��~x����$��Rg�;���,�h˦i��AUI5pP���.4ǣ7?�&DOt���cA���&)���s~gpD2𤄜�,��i^�I��1�51���X	��� ��T[`F���S�&���������č�o���5[fs�B�V����������O��5|;�#�1�߅\�rsLU����Gq������27X߼�b�+�4+]��"T.�W��ԞQ���f(��δ,�S��0D�P+#�q3&�Y�`,�S�$-u��rR?������s�q��
./S����]GY&�k�$�F�����R�����D�M���J�7��̱Nҡz���wK�+�y=�gʯ�^$�}0i�$μ�������4�=�<Y��7��S�ͨ.Zm�f�mDS���_��F�����l�Z*�$L�{���qQ��땘��bv�1�� �,�xf$c'��3���ޱִ�=pS��	}LtS��Y3�c�\g�|���g5i�ّ-%�u*>�Ċ��=�҉g�w�Y&��S��P�Q���R���Wz��������#�Tg�:g���?��<���Crp��~��̤��Ǉu��j(*�E��Ĩ)@�G��$�X�Oa0���6t���#���ey3�1q"0� ]t=������_y��=Ԛ��Bs����&���H����! =;�؞���������,�|Q���_��O�28�۪Q�$_m!���! p��b,Chq�p(���a����zV�4��,�8���A`�xR}tٟm�,�fYl��ƒ0*Ԡ��V�Lǽ��?��+
�hn�=�K��
`Ғ�΄���������2}��,�E��ĺ�dٓ�4�r۽�⼮���	<�r�"�;]&,�,�HG-���'�&l,Ĺ����>�� 2��kZ'���
����	�Q4��t�bR5>B��&�W�0L��P�f�6j~���3���+`DU�3 C����Dr���@��0���Z(���~�y����w�Dph���I^�9�������]�י^��G6�q!��~�UmB�/Eʸt��=��V���R�7��bEJn�L=NFa�S��XN�FJ0g|e%#��CHد�2��&��r"���7�U2�!��Sb8Q�P�,1�Hf\lQ���M�'�vPΑ�a~��17'���^߰? m'y?����G��n��~ ֤̃'�t	�x҅6�1�7�ٹ�<�lؑ�E�i��_�G������G�m>5�	'?\<z(7p~�п��/�qE7t\�4�f7J��G�KL0�%N3��G,������i�N_13�57��и�(SrtWx!�(�se(�~��E^�.2�=S-�v��=Yp9tH����N���<����R�m0�!��M�6�/�����}M:� 撨���4:���,F}iJI9�e ���UЍ�Y(n��QK�m�5����Xb~u��]�ª^��҄�����m��o�z�^⽢@2��X��h����Ŏ9�x�荽'�d��E7z���bM�F����^��v��y�zz�1+4LFS�M�-��ē=�1	�CD{������%r�%���X��ď����x�;9AȲɊ�㨻__�L׫��9�(S��q�n�X�}ʅ...�(ȭ^]]��ttl	�|���͛7�Q����͓D1�b�\�>/ʇ���ʧ$��d�@n�j��WZ	9����Kky.���͕9��
joZ&bH(�˛�oDb��'<�h�p�4�C��ܷww����_�{��۫;�B��~�)A�[�z����~?2gQy�J�%F]��cB���d�v'
������QѸ�di�n��Q�	�,�*���U���������ŋo���Yh<,CV�P��w��v�����M���H	۴L1N$�B���~,��j��������~	��XX��E�����<T*C��󐇏��������^7ɮGu�^��E=��:�����K���d�aF���E��E�v��.��J�xGG'�����˃9�U��4�)��	z��i�7l9��[��2�X��S��$�hvӇkhYV��/M�l.��v Q'�S�]sr��fefc?Qo;=^?x�__�;����{�&�>S;zU0`g�������u�X�"p)���^'��mz����"�**�	�G��z��7��$az�E�D6>��S&^�Pg��j��/��o~�_��'��o���o�������w$��abi��o�q����a �&�4�%�_�����S��l��b�� *R|0��"g�t,L��B��m�(����V������;�%���%�vj�i�G�NN^/�n(����BCm��b 9�s��=�7D�'[T�XN�bH�>ٷ�M�jH��o;�Ne��j��|���x�"+�����F;zI���C�������U������uV�    IEND�B`�PK
     ��Z����=  �=  /   images/28e7f2ff-99bf-41f5-8f78-c92be5544a69.png�PNG

   IHDR   d   3   �:L  iiCCPICC Profile  x�}��Ka��ʆ����h�J� �5�"谂��<O�����-ZC�?Ƞ9hH"Z��!��&�������3��ޏ����󾼼�?�1V�P2+��K+�U)�
=�4�f1U������/{7&f5����^�tz������՛5l��/RXg��dbu�a�w��,Z��"8�����gnf)� �!��%n˙?������Al4��E1�4���Cʐ�"�G~��'�A�2,�ˣ �zb�	�,L��L� LRĝ[��o�On{�/�t�s~����������F��@p]c���Vɟ�o�@���5;Q��q���� p 4+�rެR�pi~)j�^� �   	pHYs     ��  eXIfII*            (                  �    
   �       �       �   1    �   2    �   < 
   �       �         i�      %�    
      Apple iPhone XR H      H      18.3.1 2025:03:10 13:59:46 iPhone XR H      H      # "�       '�    }    �    0232�     �       	�       ��    359 ��    359  �    0100�    ��  �    �  �    k  �       �       �        �        �       �        ��    �  ��    �  �    �  �    �  �    �  �    �  �    �  �
      �    
  �
      �
      
�    "  �    *  |� �  2  2�    �	  3�    �	  4� #   �	         1   	      2025:03:10 13:59:46 2025:03:10 13:59:46 +01:00 +01:00 +01:00 "�  3  '�  E~  �  %O               ���2Apple iOS  MM )  	                   h     	        	      �  	      �  	        
     h  
     �  	        	         	        	      
     H  �       �  	             �  	             %  � ! 
      # 	      %       & 	       ' 
     # ( 	       +    %  + - 	     a . 	       / 	      � 6 	     e 7 	       ; 	        < 	       A 	        J 	       M    .  P N    y  ~ O    +  � S    +  " U    +  M X    ,  x    " # # " #           �  "   " # # !         � ! " ! # # !          � �! # ! " ! %�*"�"� � �" ! ! " " Z�|� � � ��� � �" # ! !  � -� Y h � U%� � �" ! ! !  � �C� � � 9� | �! # !   �� � i � IG� � �  ! ! !   � 	� w _ g 8� � �" ! !    � � � � Q Q � � �" " "    � � | i _ E.� q �$ " !  ! � � x 3 ` (	� i �$ # "   " � =� I ) : ?� c �# # $ " # � ByA8�!� W �# % $ $ % � >��/��o : /% % & $ & � '��2 ��;J  | bplist00�UflagsUvalueYtimescaleUepoch  �e<���;��  '-/8=             	               ?  � �e���G )E���=  n`  �        bplist00_Ab0ADS86MCAjpKaa8LFhJJlP1mqK                            '     �  q900n C4B2F7DA-8462-48A4-BA2A-55C71892FB82             6    @� +E  �CB48AC14-E04A-4371-B2C5-73D7213C0CAE bplist00"A�                              bplist00�Q1Q2 �
�	S2.1S2.2#        #@=      �S2.1S2.2#@3      #,5:>B                            Kbplist00                             
bplist00                            
bplist00                             
bplist00                                        	      	      Apple iPhone XR back camera 4.25mm f/1.8       N        E                 K        T        T        �
       �
       �
       �
       �
       �
      /      +        d               i  d   � �         OO H  OO H  zQ��  0�IDATx�=�gti�%D x� 轷���R&]eUfe٬�����gf����sv�̞���tj�m�dmuU:ue��KyC��H�;� Ax~�u�#�����w߽��1O�~�k:e2}�񕭵����T�x���(k6�Z�$�f��[�>�ol�X_��[�M�W_���<�\�ڍۆ�^8�!حiڃʢ4:���6h2�+�+�C����q�������;Z�c�fΥH����{[�[zu����|���px���^3�`��K�dz|�Cp�8jiq9��|�~�N(��������b�T|?�����B�Jek{O��}���k��������3��e�o��f���N���M��N��	�]�tEV+Ŝ�5��JY�^~}hhAb�g��v�X)�l�*e(m=L������_��=�-2&���ކ`(�^�*sM��JI7٪��k���N�kiuS�入վ�`S�o+A��Vև��˖$�(����Z̝���Mݻ;���Mά󼻫�oe=23�\*�z��SG'V7ck��x����������d&�55�Yk���5�����M����٣�O�}�����ֶ�����7�>98�c6��#��x������������(�뻳�T���er���&��z�����6[9�.��&��N���wo�����^{��׾�M�X�}u�k���C��W���P�����'���_�y��Tf}+J]���ӓL���҆�7�:{���t�`���s��bs�⩬(���K�Κ9�~<Y��ՍE3��'�n�5�.�v��œ+���j6_h�l�C�}�a�"�%���j�sP�UE7�w���Q��I�X��As��R�����XQ���v\V��酲47�HY=�,Ee+�
v��@o6w�PQ"��^F=P�(��7w���fuD�VdE�r�����(U+7o]�������������.^dN��p��3Y׃M�d2708^��R�L{k�O{ Р�&�Zm�-��,<K��(��=[b9.�.�c���I��m6Wd#ۧ.�-z���~���w���~�j��*�$�s�[!� �:�Hd>x�՛T5-�-�,�5�D��N.W�V���77�ZV7�v���G��������U�ݝ��D-Q�}/���r{C{�C*�{P)���ay��Y^�s)3k)+�Q䝖�,�y^3�j��<�y�Szk[[�T�lvH⫯}SU�������陧�T�I�s;�XwG���,�UVdNUdI���RE�U]����7O�<������ܜ?�����m6����*�x�ġ�gNeS������ԁ�?�����x�$^���������5M13����������	8"K~�;�������/:�.��;��7^{��v��o,<W�����e�\��X�y]GdMo5U����w�xC�Z����k*�LUʍ�Ʀ����p8��v�c'�&���>^|�m��'�4-˓���$�|N��fw��A��b��a��1�|v?�ffa���G3ͲL&�{4��eY�ɤ��$��BŠ(0��k�لO��N�߷��E��nw
�h<���ә��H�V�^:s�f���w߸q'�/L�uu��^+/��R����>1�O�f��gf�M4���0���k�I��ՐDpl|t'�}����#��>�k;�MR����ӧ����_�c$r����,Q���_��{�(.��MOfr��3����V,Z����bahx��r�ff�D"Y��>��l3 |��l�����ҙ��eUU�7wk�/s���aC�>[����i��_���c��P�*�/󞮩��������vG6�s:��x����#&&�{G�j�	�"ЩT�����}p�~C�/�����_uM�4�õ�ˤ��b����^�e�c�L.�O��>rc�r�� Xw�M���]�2p��ťD"n��]YY�i���U�J�@�ʥ�{�eU-J���T����ش����{X�6�t._��@jyy�l��Z6�ݼq�Xm�3��2�\v|l��Z���m���Uk��612D��	�4�&�L�(ʴ�����eE1��7�I���L"��9�T�u��"��0�̈՚33�	�Ԗ�WeE5�fڄ7�2�����¡(R�b�P�8�E��rx��4���Y9.8�l���C�k>�{d�����׺{��Gvr_�)�L�T.O��
����d��{{���aԇ��JePU	��	$j�.6`�\.O?z2��e�/?�M�[ZS��(���`�A�O�;�-�v�"�!`��9��ΑE�1C}�_��us�����z_W����{��(���O�<�k�^k{K�)X�I�mc�y|����y}}gqi����k�	�KEڨNM�(�,�=�[�aX�f���_Z��mkn��S�}ݟ~vut���)p���J�r�ֽ#G��ld3���}hp`vv���2�����rLS�9��T��,8d{KSKK0��/�̕,+H2O$~��@��fQ�'ӊ$C�����W��Z�B�(
��	�!�1�bYz��o�Mc2�T._x� ޠ���P��D[ �2K�}���nhvY��Lg��������>�>4��꥓C�ܯ��פ�@�����\`�VK��*���$��_��5���'����4?_�5��o�h�D��T*3:4X��(4��Z�I���g@P�R�����5h���R8E���t��M�b����@��SG?�0z�Pl�[o��߼��������2�R�:+�Z5]�(\�^��I�7����qx�;����5���NBgf؏�|��8�ȩcW>�Q(����s�l.��j*�0l&��&���L�j�,��y��t�������Pk�B~'w���)���ǉd�r5�+�n?�����ޫ�E�h H�L&�LU���!U�l���;�ܮ�� t����xS��=2EEc�x2L%��JMe-��"�<��8>ѨV�MM����Ύ���eI���k�η�:A7HI�5���ұ��Ͼ���0�T��˽����"cf�9�t=�� �-���_NL��ⱕ�u����JV�#��OY�Ɍ��<ǡlS�|M��>��1c�PQ嚌�C4��)�n˦�86���ҩ|E��
K�*�qCWh��da��	�3��P8�/����~��q������'?�$�`��@���C S��+��u��>|2�&&��ݸu]���Qv\I��G����K��Yv�<>���n"�u:��M��ׅ�=0�MF�Z��0�\���!���L^���Kٸ�������^�h�>x���9QP
5�@<6B�z4Yem/_>�rز9����/������_�8�p8�-j������C`ϟMd��j/��V8��ӹo�b8$�l`2�D�jp�Ț'�����V*��]�:wwv�-Q)3�/U-ֲ��A���L6�p�x��󶱁����R�����p8jU�Z�U��E�Zm:hԔ�o=?0Y����8���Kg�&���t!��N�$�P��2��;\���O�iGhgG ���@�P��'R��X�I*�T|2ͪD��m�w3b����(e�!�Z5Je*aI�fxx���	��YI��#��r�õ�X(F\���tw/�l��v�oP��o޾p����N ������z��L(K�r��j[ks�T��$����fm�������v��3g��x���~�Ȱ�	��B�_|qVCJE7������M�qݝ��E�4OW������{����a�I0fh���[,Ld?Yk�`�)������
<���.0DZMb�V,�-�EU��f�`�pH�G'2�I)�{��Ý-��gj�p���MU;<9�_��?-K*LE�he~��W�+�A���~_}�I��� ���C�kk뛹|^7Q�Mp3��D2&�Y��?E���jokz��ikk��V,���.=4�0�lpx���٪T�h,�7~ t�o�f�v���M\M!����˛�L�VC������?�j�[�V�4���ݷ.�U���,,n±���߽�s�#�Կ|qTz�����n<���Y6�8<�t;J�Vk/,�	 ���k�TC���w��9�IZy�*��V�����m�����=���ʕ`s�Y$p6�
�%l�io/j�/�@hae8�7խIUU�p������`0�t�w4K�,m�"�Ͷ�0�R��/f���; ����_��%h����E�_��]87�١`$=2�s��t_OkK�?�[q6p�����/}���榆bQĂ@��CC�����7����P(h��\��������x�>��z�X��d�W����(7$/*��&]m	:dY���%��Ny�^�޹{ll�g5t���o��M��>��zOW�����`3�P:_)�/E�b���}��(A8J�׍�}�t�v����o_��Z{{W&+޽?�M%P����F�"�A���A<U��0��FǃΠ��5��6�=a�2���  �I�"��h4u��0lAK���6k������;\v�X.�v7G��Ϟ�v�B�넍BK\(��X��V�� 6'f��R)O����T@��- `&�v�ƍ���<kB�P�(V�����7^}���C���Oy�^K�X�s](�v������R�X�<9>�'�m�r'54����l��D�����/�'P�!Հ��"�5���tb��s�)h�)��:��$�J6[|�h~h�kt��΃���-������.�m/*��-�OW���C���/�@t��t�3�kh��w&F�{��HW)���;Mη_=y��jify|d� ��#q��98Щ�:m��	�zܮΎV�J���s���T"��E�����,.���������Od����BaT ���=���j��UT�&ݾq���9�%�!ׁ2�<�<�Ѓp,35�a��w�8z��Nl<��@˨kz�-(iPU�<���o���opݼ?9�d��pbl����5�QX鵍�rM�l�DJR���_�۹�oii@�ڍ�t6���r�!-N�������S+)c���k��McW�wݮ�n�47@doۋF�WVF��.�
���4G�7�6��d�� 12�^��@S2�����H��ߺ��K����_��#�
��~��@���r
��1�}i�ac��b"��ҩ\g���*^��Tu����yVQ�T&!�kE���k��"�	�:@W(����_|i
���d<&��O�a�#���q�����O�9;{	��jW�r*#~����a��^�~��������+��#�h'�4�,Tl��Ua��x{�b�(��8֤Y8�	�	N��X��N7&
dj0((2e�9��$*���Ͼ���ь�^�5���kQ��F������u5$Ro�TM��d4@�v��n�MdV�D�+\ؕO�]�z���q��0m-��'���馍0���Af V�A�m6\�F��w��w�j�����6�e�R�,�H�!C�����#�0P�ZU5^81UG»��}�<��ne��sss���2P0&M�b�p�j��	L�\�N*d����x:g���B�z�ִvb�1@��_�_>-i�"�QGMVaXъ�q���a9���D�zD���$
'����D<aY�nd���*\�n$l"�X� ���K���^�c�*c��&8�5Q�:0�����������Ͽ��~�a��~��Ԓ�hUVk�AhT�KP*��mGK:ɥ�n�<��U��jD����_
�F�Ū���)���kE����������j��=45N��Ӥ�!����;�b�M����P��|�A�J�����?~Z�ˡw�_-L8��z���>�d���QF�Xi�{���X��,�G����p_+���W�>'��g�UEQ\N7��,m�|���Ge]�AHAw8l��5@	�G�7��W�P�<�vt��X(�l�K�U�<v!� �F#¦1��WK�b��E`��`�φ�`�8o#ISL=oƁ�6��N�BtׄN���f����/�K����T#%P3�/������%�9gY�1��܍A����p{G+. V$D� �7h��D"�-,���?(jog����{W��-���	���H��f��:˒�Ѧe�8�aÑ�3G�A�R���T��X�&'|O*�y�������$7M�/<��Hf��^4Q�	 �C(��P��7:Iyk��amm�N?�)�kD_̷���_tפ��\�,,>�������f�~0��L�t�U���AO$�z���r�$�,�\\�&�+*��s�w�Cg�2Z�R����R��V�B�DH���t�R�"��T29a̪�j�af�#I�fm��t��:#���,2� ��9�2I����pY!��Zd8[ox�n2���ƓD2Z��}:����=���cX�2�0�:��:�!p<Nnb1��7_=���)��Kf����W�R�!nn���Ʃɑ�cֶKka�~i��A1!��!�/:a(vl����xV��w~��g�f�||�X"�y������(�W_x�t{g�+�UD������L*}��#D��'M���ݪɌ>)Oe�T아	�<��N^#{�ʢ>.����a�()K"����:�g�!���Y�o� A+4�@���B��B���Ƕ�=0e1�?��+�\:�������D^����Y����z{ZVV#+�;�B��5���*�S<��uw�����G��(��&�ˍ�_8����a��ɱ��^�������CG|��u�φn>q�����_^e��_kij$�h�"�X:���x��Įd	��R)�t�S���0�r�`jU_Ba�t⭈��ê�'�41�0#�d�B�	����AX�|��2�
<�'.��Ti�ﵓ���Lܹ?��~�!�H�[���NO�v6ݺ=��ǷeM�p���Z98	�L�ICA�� s�ՊBs8�bY���������B	�~�r��X��qIb>��)+o�R�����ȳ���gJ�T(����u���������b�Z�1u`R�T�sWN��%#{ѕ�E�nC;�hu+aP�Z��y�e����������	�x��%���I�NT�x����}�/DJ�)6�rh���ʧ����eA ����T���3S�$/���J�ot�U�f=���V�s��L���=��"�%�
����������?����H�+k`a�3�ռ�c˕���8��f�7+���5�}v�F *��e��^�K��D2v�F�Cˉm��d8��v�B��"�xl1Y�W��������c�ƍ�(�U4󰆌�g�yn�e�*����'��ȍ��(��4B�p5b���vx�v�IRI�4�L��Ѱ%��0p�;߿O��}�����`AʡRF
���Z�2r��p6pWK��{ߺ��Wg>�U���'Yr� F�H�s�T���xܛ[��B�E}P����cG:���ɷ�����O~�r8o�}����V  ���/V� ��VG�R�Z�!�>���/E�������m�6��O��X�[�73Eny���&S]r�'4�^���i����^�)�^�d ��)p�
��՚�ŗs�r�*v;�1D\p6 ��X�z%�$ebaY����d4n4t�m$Ylmi�dK��}+��rE4����^�|�+�b!�v�GG��/��?w��8��T�^8�X)m.-�;{B�jXg|b�Z��� ���|&�Ƨ(�?H��O���s7���8�2[ ,�|��h��ɲ6�E�U��*L�	�i	�0���T}tEr^��L6�#�̤2�����c�����T3����R����B�z��B:�'l�06�U�jhY*�
J�B�C�=�Á�Â��v	�RE�ufe}����X���#s�����s��)R5����Ew7ۺG���T5�|	�7� �ǌ���7�J�4�z���ܚ0��d�,��w95I.�K��bài�tAT��NZ7�+Ѫ��ɐ�>���[��ALi��BM�h��2A^�ϗ�"����Z�$�~�̅oݝ�38s|�_�A��H�8+���}�|������l�̮�Jb&�.#�.����[Jns��84��(�4:�JKGWYT�l�Rt�������{Dg��$=��<61%'k�.�"	T(T�굛'��֪6��x����2txꀻ�9�~���

��}3�i�<���S�{��i�~M�B��j,���_���s''ŚR�j�h"O���?�`��}'��Y^^_�P2�01�*�D�O��B��,id��n4���}���.�?s����x"��A��cg/�����7���?yhxms����sD�T�@�.cc�$�B�iT!P�L��c}���O��<�y�����~�[p�tS��D:P$3�0�2�@�ʀ�677��v�˃���1�h6<t��w�5��v#�����Q��L��aw&�)�JWGG8imilkmE�ry+-3�B:����O��n�����+�A*S�䫄��j��Ơ�%r�99P�H)u�
�J���6z��"�1���.�G��~29�����i80%Lh�Z�	�*⮠�R����(+g,c�<n�#��v��+t�������D���>�V�C�<}�����vC��b/ԣ����u�B���Ǖ���x����F���F�"����lll���ujkk{rb�).����;<5��☼����ǟ]-��
�z���|3�?�KVo��ĉҔ��E��u�EX����ӹ/o>��� �4�$�P� �+ߟ^F[C���8�uM5�2�&��Xhr�W(�+8�;Y5�V�6� 0��o����{�@�+/�E���/�ʺZ|��t����^0����<59��eB�g�ٵ����Q�jey���Y�;�������Z�s3�^��ܙӷo����v?�[��w_�� @�|�k��<�_:l��`eO}�N�!��T�F�VĒ�Ѻ�xo�K�Ă4T;��
"kg"�G3"����5Y��F�W�ߪ#-���E�4
�qn���aA(�Ųab6vR�X^�6��<��^^\�Tufz�!�-���ѐ@Xa�NN���������5�|?�Ֆ1���89x4����nmnn���\���o�y�%v��T�[:�'L�ӵ7��!k�R����'��wb����́�n���%#=���:lit�I��=$��H��|�><3Uj�)	\�O�<(���*j���f�����B��
�J5�`q��<�=[� � K�S`]v	%��^��t�8��~�����䃆 ���m�z��l������Z����p$]��z��Ȫ��{�)�>�0_�����Ċ���#G��������v��߷��`"X��X�9�N��Bntj��������-{C0�ɧT=�st��)$	��C�.�쮫���Qj�N�	�=��YXO��Ȋ������6�BW�,YY�?����F"|zW���y�4���>��I����ۛ����s�W/>89z�ƝO�͟;9��W�>�����w����W?~��O=N۫/���\�]��yb���6�0���0Xy��ai���*J�a7z�w�5��J����%E~�`���$�|I�}���^iz$M��`��p,]��]#uc��#��md�c�
�lAl��e��>���\����2�����R�"�
ź��RY�{�f�ʣ�t��s��[����]�R*9m �ɛ�ŜK��GW
9@Sv�)rP` �yT
ēK�u�~�PEL(gl�+#<�!��N�]�I
��1�E&n�F���];q������=���X9+�@I�����O���[l�x���9}�/oT����I�
��J�F
2}�ҙ��f<.��`2�����F��/�%Oj�-��>�%�F&ɸ�"�����^��V��ڮ���t�*+3+��ЮF&���N~7��/��6>������d��q��zlq/��x�}gfo?������������Y�o�o��(֑ɑGk |��W%Uk�b�mR�5����x���	&�:x�@ww�]@FK�(פ�X�d�O��7wق]���A+L������֍��ЇG�7v�?��]nr;6[��ġc���+��Oc�w�&UO�s��Ѓ��O�q������u-���ށsik�;�o�?z2o������D[���~��p�(J��?~KI�
�x2�A���MsK!u~�F>��Hz3�5Pl�m��z�<*���ѽ�~&��n�V�L�]���Lb��O"�d�����E�`%�����G����F�g������V�F��?��8��e�y��ҩ8�F���T���ݖ���6MsK����8��P_gW> �XZY�;-�_�t��9���y��z4=������`X�h�����JU��}�}}�u��k7A@Dl�����L�"��Ҋce��h
g�~0ȶLMF�:�t��7QKE�X���Y �<l�p���0"[����^<�)k��;w^���2��vh~aA�jddf��P
y���IE!��r����U�՚���ԟ�5�gr�!������� �����⚉�8���3e�=}�"�\�ֺ��P�w�=�i��c[;z-����TMi4�Z�v"V�p��q�g�j劥�Nx����1s�9��1��˗.����r���<x8}���?z�<g�����w�=��?�����Z������<�	�~���|~Eӓ�ܳ�y��599A������b��nin��"j�T*��7�6ފ�@��G�ϝ9u`b	(UJW>����SN�;�����r��#���v�zz���ڣ�Ӱ&+%��'O}��oy.����������s���G56x:�z�۳�4ZDo�𱥕�4P����w���8c����Z_��.9z�[�>=�tnvvxp�����Qh�>�������N�`X�g?�[T��>��-45 �}�ݨ���Fx���O5E����e0��])�p�J��B����1�߷��]�UǇ��T �x��D�T�߬�O?<40��������[�������[�l����OMXXKKG�X)������(�Y�N��y����_��������60�j
�t�"mfE�X`�3���ַ���O�c���]-��=�30<��ޅme2�ƀ?����t`h����W��5�m||�x��D(���r��:�y�~[{���<~���9��/����mi�j�x"�l������=(FV��������;f�eXӅ���knjڍ����ݼ.om
�./��Y3����X8��Ph��m�U�B�XȥR�����C���}��?eK�{�Y��6��������7n�<�6t������j�\�z�Z<��]�J�[Mjll����N*�v���P�w��Ќ�]����rs��ر#&>�B;�h�岙��g�l���AP��߿��|~dd���=���r��$��wB�ۻ���o���%2���e(qOWS0�������9=n��au{[�b���C`G�{��m��<�{�l�Y._<}��K_ݸy���9�����c��v�P�$qbb���s�Ϝ��?�˿�Շ�\�~��#�����+t�[[kn�^	�S$��G��lm�,/�(�?�m�,�˒l�+[Ã�o���l�x�ν�施�=�
���|�}��t�eq~~�n�;Q���~�a<�����|�ɉ�L����4( 2ݏ��7i��t;D�v{|��a��.�����/�wѲ�wʵȢ׋bw�xKSs���2����^|���;��.-�����p�ȑ���ɣ�]յ�ǎ��l�v�u�6Szmld���i���ͧƆ���nd�j������9�j�y���QCS@�(�Ս��G'|^h542��:81���a�p�ΝIgr����K���������o�~!
1��Q(��Z�P���t���^.�~��߯���{o6��2MM�\>u���5Y	�E �\>����C�Y������'K'�d��6�.853�pv�<�^3T���J�lݯ��-��f��-f������|*�ZX�v(26:�7~�ڍ����~kK�٣/m��p�h��-,�M�x�*ep�׎�:��bUk�z�"Q��w�I����tjmu��>��%$ɸ�ʑH4e���Ϟ��;�����Gz��{����:��Άf�7._"�V�EQ��}��p!�`��ŖW�'&Ǿ���1h�/^zYV�Ͽ����ֶ�U�<pAWk�QP�x*Ǯm۾�s���㪤,���]3��{��׈���6�,�,LO��j,.o��h��&�}3M��jM2��3(�R��jՒ�<]�\]^M�l�b���g�����2���}���:�ˢ�j{�dN�U�����A�L���[��-T�^"-��q}��E�WwG�����P5Iv��++��=�cap�%�^X ψd2���ˇ��v�փ�8�@����ۙgK�*Q�v���'?���j��J/�Xͭ�    IEND�B`�PK
     ��Z��:�  �  /   images/8d902f4e-ab09-4493-932a-1f1db25b6d7d.png�PNG

   IHDR  �  �   �Xa  �PLTE0/0%$&\z   ���>=@)))�Ɋ!#fffJbm,+-@S=>B<aq" "̀
�}�}&%(]{�Ȋ Tl:@G112_{���6r�.-/���ׄpF+���ւԀ�~	�~�|
s���y'h�<o}����w���Bs}&d{�٬����Ǌ5l|�����]{���������\a~�iaR;�ʌԽ�^M4����ϖл�x��U|`O8\K0���������*f|!a{K��|��#e�h��`{���a���Ɗ���������������������d���ĉ0n�������d����Ѐ���ћO��C|�������-g|eWDcT?���{���͓�̐õ����������s��k��0i|�����ꍯ��֧�É͹�������H]dVB��ޫ�����բǶ�����޷V��,k�p��`�[I-����ӟؿ�������Hu~#c{�����ښ��m��>x�����������ܳ���Jw~�����ִ�Ր��3D��ᢾʣ��Ac_�۰˸����Py~\��G~��k�k2'1Lx~5af���RmIafYF���My~�qfiHfYG�z4q� ^tvg=�{B'�sЀ�Υ���PckWdiW8BH.8-9.�D �  �IDATx���]k�Ppy8��~��"��+�ť�j_.V�:XY�X��������ε��n��6���D���x�7sl=I�IN!�b��Ȓ����](~`���v���]0g�����zsvy|-S�'���V�V��5�s�9�P�� U�iN�O"5�*�����؟?���|9��_�I2wF�����˂����Nq |h�Q�qw7�.�X�n|^ˇQ �rXjŎC��T�:�}�U�Ie|[AG�����G4>��-b�1���>�h��W#�X]��s�#j]�	�E��~�>Z/G^"� >/��Ӯ����7�5.
Le�~��G��l|��0ձ� =��4�D����|���B�⟠=�.�a�<AL�m4y�l���r����
�b�!�
���cw�@_��lsy%	g�\dy����P'�}4��dZ���s��\͇�[xJ�6w�A�Y����op2�M�)���@�Bu������-޶	lguYb#h��*H���n�$"�%ԅ���E��n)"��UfU�ju�4/Fɴ��+}�؊�2��DZ��ו��.	�,w�fѼh	�Yqdj���U7=�M`E�^&��;��y�Ed)�`�� k%6
���Eְ��b�{O"H)S��4E��v� i�*����vy36]1p�<ŮdC�U�f�XD����%��Q`qB�����,�:�&���*��*]���@�q��j.��%vd	� �}"��'��Ut��:��$��$�m��$qQ [����%b諒|O�ù&��[�0�Y�:�I���d����3VD"61���f<���"�
<���=8c�9�Id�;�VH�q�ԇ�G�|N2��2?�z�l��"���/�xiļ��u����#�8H�M/����X���|�yC���dv�	�da��I�9ANmBP�ufx(*�yxﭷ���*W-��"��8H U/�������~�]Z8l�WTnV(4Wv��+�>}�-���뷼���*qPF����&qGj�E�[]oW����V��X�-��˿�1�-h��l��`[���ǁ��Q�V�Z���o�=�؜�3%QV���\I�Q0
��Rp,�p�����{���2��"��(����(�$)0��H���-�+:x�>]āf+�A���l����罽�7_șaY�-�aF��9I
V��$$9$Z�F�P"$X~�^2������2��#�w����ڵk7n���co���!X�WC�&+�RC����. ՉL#��6]�R ΰ�rCH-�qK�A��HM�B�M�6��EV`����Oq����秶����?��yҗ�j��jjWade�~٠�, �������´��_��~��� ���<�:'�?�wcފ'���Bꯏ1�@�8��H�P"�8�
vM�[��ϻ���2���m��¨�e������>���%��B��M��N������`���>�ǝ�n��Un%j�L����%fTn%j�L��n>ʧꛪo�2be0��gU��;w �r���h�=Q�v���6��S}
Y'�����#����EjyFj�@G���<h�<�X.4�:O�7�Ϭ�4�:��瑇�4��K(�)6�����=u�`��a��c�N�CE�����{����xq��	�>��� �����1 s�Y����K�qԵ�VW�ɽ� �s�z���P��1�����O��6����lz�Q0WS��m-��k?;5tq�-��+Cs]K���57te��A�c�����v�o�0�N�N�P\�*�)7�s�-�?��0�a�k��Dv��I����=���#0�_�ȹ.?$����+��m��	�F�`�N����ӧN��w�aM?���I�ww��:u���;�I���$ه�70��md.��3?'�CO����'���L'�_�ȃ���(�D�>�
 �Li��R��e�`��� �����H@�ŷɡ�[\w��iԃai�h��AG��V�uZ�����S��7��LUo���M1!�ā�䏃��zm�~g�'��1b
 �@'FoFH&�+@�W��1+�P��A_]}���W0�h���t��<���N���Gs��P���n�-g�/�2Љ��Ib,d; �m��$��������t����9�x�h
:�����\�;�cd}O�+w�j$��Y��L0,�%��MV �d5�õI ����>�iTh���$aMBg+ �J5�� eB�Лc���Qԃi��,��
����G2V&X��L�R!��i�"�d�32�x9l���SB�����@�����^ z[�JԴ�]�f0��ka�_��Y4��v�4�Hpr0Ѵ���Ǹ�`!S�:�Lv0��ɻnG<�Z0�`ـ��X��}�`�X��8��5��<�`U���ɦgۡ������zi0���r��i2���� v�������P��f����b����*ZB�Dޔt��~3��� ٣�4���/����&��� t
��`�d��`	�d��Oׂ����(-o紈�&+�^�N�0����|V%����N7��� p���qA���V0�����GGoL�M}1�`�+�R�`\»,�T\���l3�3#+�F�	E3`N��#�V0�  q+R	&�b�9���8��~\��@#�a1���%)m�'�r��͖�(.�8�7�,a+��;=�İǢ��ba ���WV�Qk%V,!0x"���%t��l��h>��rc�!q8�!L��y �MPq:�SS$�AVy��F���"#�TO��m��v�H2������5�Hɖ�E�G��2Px����C�`�O���2ر����x�`G����������������������gǸ	QD�đ�I,N��9"�~��T�f������������{��_��#���~+��5r�����8���8l�Md�V�Dl$1�yM�62; ��7ۘ�ě(�M�	l�M��f���60;,���a�$���g֟X�M���C�'Ɓ�gV�X<1��N�����&�`��!���҉�`��A��?(�`��L���0�³�&��uS���C�~�W����`����Ug�M��&�5�����`��d�db4X��3V��+&f������`�e������KL�%ƃ���j��ز?`��,�؋�;:� `(�����O̶0$f����XĀ�",1`���EX,b�b�,�	X,b�b��XĀ�",1`���EX,b�b��XĀ�",1`���EX,b�b�;��",1`�;��b��XĀ�",1`�?f���),��
X�g`���EX,b�b�X,b�b{{���7``����=�M{`���EXlw ��=�EX,b�b�Xl��EXlw ��`����0,�;�Ŧ=�XĀ�v�ش���� ��b��b�X���v�XĀ�",�;�Ŧ=�X)��`�R��b�,�;��JX�^)�X)��`����`�R+E`�R{+E`�R+E`�R{�. ,�;��JXlw ��"�X)��"�X)��"�X)��"�X)��"�X)��"��-�b�,V��bWr�Ŷ=��1,V��b�,V��b�X�;ƀŎ1`�R�V)�R�l[i��R���t��'0Ͽ��,���5�(
�hR�i�½�m[A��1�3g�4l��Ӱa6LÆi�0�a�4l��Ӱa6̇a�y�Ӷ�u�þ��l�}8�Ӱ�5�UÌ �aF��0#Hl�$6�f�3�ĆAbÌ �aF��0#H\0�����>\��v=,s�ه�:�kX�^5L�&D��Ɔ	QcÄ��aB��0!jl�56L�&D��Ɔ	QcÄ��aB��0!jl�56L�&D��Ɔ	QcÄ��aB��0!jl�56L�&D��Ɔ	QcÄ��aB��0!jl�56L�&D��Ɔ	QcÄ��aB��0!jlؓ�;{m"�8.�L���(>x�}H��@IB��-ڈ��X�Z+AKQK!P�h�Pkj*��>)�/O�h�≷������dwg��*�8��R:��䷻t[�jD�
T� �U���0�`��A�@5"X������f���0������
��8܂B��C���MM<r9���0W]��&��RS`E���W.�=���` �]�3��iX���q{l��^Ul�i�c`YU�	����38k��Ui0Gm�im�*6�r�	��*�3qZ'b�sҵ���`͗�K���S��Y�{
.ǘϮ���R�X�����>���ݝC��C��_��G��j9F����
�%a9)��D0�:P#��,��PW�(�$��ʳ�u��k��-P$��ɗC#Ҙ�<X�	2{�f��]�������6dHe͂y�ȶo�������cŲ��&�Nې튏�sͤl,6�z�Bg[�����I4�����G��A�}�9/��u��Es�,#�r�Q�z�#�����/�=�`��u��'Ir��V,� �x�ء�>�-�WP��N���'F�ĘQ�=1T�{��/Y�;|pj��`�<��HD��>�*Ҹ6��@lO5o���C��b�{6x�*�:R���\�n��m���J�ի��|�oҹ��?w�z{�ru#H��P�&ZN�"�n;7�C�ׄT�hET�b�:���FE��FE�Y�t牞�nT4��d� Վ�m"��Dǻ$�Պ�{:��t��}I:ާD0��IwPj�y�OT�eR��� ������h��G�I��+�`����
��&ݢ!b�<�n�`<(��Cq��h�eP�I����?ra��s�}Y����xw��:�u�˃�3����]�#K�b�s�m"����U��Ny���r(�c^��_�	6ƺ��P�+C��0(sm"O��v�g���`QeH$���$��e}Q7Q6^�eI ���E0�`G����A�~b,�����k(�Ρlcy�{�9�e�D0�`�P6Ț�M�Sl��l�B٨��	e�,�(�kAY��1s��,��:b�eiM0�
�V�F^�x�A��w+�vk��VY�������eP�5i~#�`7��@�(�`\��P�n��1�� m�ߡ#�h���y�(k�7;�p �� ����d�X��P�U�~Z��F�`H��)6��E�8��bD�X�y�V�C*!�"w����x��u���2	�$�n0G��q��څ* �q��jL$���>T���`����]����ZD0�`Ђj[��sq�&�E�F�vŰDc��P��`_#���,�q��Xj�|�s�=ԍ%��`h.�D0[�]���f��lS�H- �q��W�TX�̋I�@�Fm���Q;4u K�����o�.�ءc��v��:��8�v��Ӣ�EO~Q���_+l/��K��x��hӦM�8�Q�~ds�I0��:Xc�Ve8���{h��7��2|���	�fo0p����>��Q�3�?@���|$�:b-n`S��/_#�� �1�qȎivY��3�\{o�E���� "؏Q;�@ѩ��9�Ì�:B6xW�$�I��A���M�!�l�ɵ>5��v������Ι�"t\�\���a,{�F���6��h�1 ��Q0��h�10aC�F��6�  �]�l�~X    IEND�B`�PK
     ��Z����(  (  /   images/4c416a15-58ad-47dc-949c-f0bec13a5bfd.png�PNG

   IHDR  �  �   �Xa  �PLTE   ���@S��Ԃk20/08BH>=@WBs}'1���Rm�Υfffm��pF3D`����a}���'���[I-�wb�����>x�������<aq'h�+���x���Γ�༷z)))���\z���bS=�Ǌ���T{0n�M��%$&-9.+f|���̹�<o}����y���&%(��ڲ���ݴJbmւ3k|r�����:@G���Ia�{B���vg=V���}fiH5af�ћ{��$c{^{�i������eWC���`O8���Ҽ���ܷ���sAc_Iv~�ĉ!#�٬\i������~	�}������#e���抗���ɫ���Ɋ6r� Tl���112���H]]L2D}�ؿ�s��������Ƕ��q,k� ^t���\��.8�֥Tdj|��fYFLx~d���k�ӟ���̀
������b0�   	pHYs  �  ��+  IDATx�흍[�Hz����ݒ���]�8�� �QA�j>ʓe�f��&��ڇ\
�/�,ߦ=�R���%��/�d[��f${4�q�$1AK���;�ч��T�0� a��$�IFE�B#�љ��z�[�
>��Ł����R��믃�M��6�B9�Q�1V��@�_V��F�����|�Ŕ�<�J3�
��]�x�����ן~�'���ldm�CB ����6�뺻4�
˖K��j��ѫ+�
�.�oua_�O�J�䇪�O( S�St]�Yú2a3�Ϸ�(�( C2�íFv=З�Ċ0#;r�Ta3u�o�cF~�~�Sv�ф�>ߪ�Џ1��k$��Z?F6�oNo���o/{Z�+ �{|�Y�����MuiR��N��ag����L�R ���϶v�ۃ�xW�Ia����]3���d@K���(�Ý�EBX/���$�2�B�ĳK��g&��i��F&D�5�:x~<��{��h-O����I��B)��jӠ�ټ�vh-�>����ʕi쮩���:�*���>��B�'�=���+,_@���ɱ�ᦘ�P��֬s�w���Z�FSK]9�u������d{U�e3!W�
��<-ܘ1�S!�aC�e�/=1�,��z�,����]�g�Lse�����z�j��0҅�����z�Ez������+l	O����̄�)�����#!�ǩ��)��\���J���B�Ʋ�Ŧ}��,!,_� Z�;˄8�0�%/�a�1���c�X%]�Rv�@4�b����C�G�hx����7�/���H_�8:c�r̎R��Qf(k��4bA��!�pc)�Jdؚ�����ϜB��w��������yu&0h^�BhoK�ܰ�Q��~��i�u�q�8ج=��DPJ0MD���:��-ͥ�͡����tsQ6n�I�+m"��~���S�g��G�;gy^Ol;���O8뻝Ї����m���·�Z}o�����w�۳G�t{G�5Y�~���sz�@��Ne�֭�jZq�z�51g�HuL\�0U��-�#΋����y{''���6���<^��Vt���tl��,na��^5�pK1]��ݞ�0�^+������=�]��T{��>r����S�k���΅�YK쓣�l���(셳�;���c�Aa�
[laN����J��]�jC�y{�<���_�L����i��o(�i�ҹ�Ha,��!�����WX���e=�	#����vR�3����[KX{���g�	��U�\�2�ނ�9�.����>�ʕ�maq���/X����X��<�]�L��pD��)U�/\����ד�Y���`6��{�;�p�~ԠQ"�1XU�bS�D��%Ã�ڄp�Y��n'�Ĭ�3�|a�{Ēw�éă���Z���vb��;,7�m��:��TZ2<���;rX'����6�s�-�;c�C���=�����hV��&tzwukN��r���͡�d\�^I`�v���r~7Ѐ�5G-lq�a��؜=��@+���Tb�6�$a�{���_N�p�'���ы����E�������@]X)�S�܄M9G����O����Jb�ΈM�6�k��u	��PV&&�h5��-���C2rEJ�(���I��8�9�H�L<�?t�2�)�Qv r��0��.շ�b	�SD�Q�#���Ϙ��MVi�cxO:+�����H���\�{ ��MR4�U
s[�����+S|ʽ�a}���U�b^c�^F`8uD��Ű��F�^axgO?f�����n�d��o3p����������������({!�C윧sj�h�WPHaƪ�k��~l�SB�PVʵ[�	:�,s��=j9 �����|�{-?c��w�}&:>PR�3�X=��#Ns���^�d�mc=�a�[c9���(N�{%���f+��^�P��:��Dq`+���nl4l#f+����473Ű�=ab/�w��[$A������g�bq��ae�K���jA��F����K{bm����%�:�uC�ˮ�r�X ����tup�>�H���^*��(�]�V/^,�������E�]�'WoA\�vB��!��}�����=@F9%�$�s��=��=���g��q���������B�G}�G�ď�_>yh=�����ޓ���8s���ks���6�6�F]����Z/1j��sP��;�e��A� ��n)��.��|�T��P}���ډ��*ʭ9KCϙ�ܺLn^�1lx����uԧO&7��nS���x4۹<65n����6���lw#��R;:��9����\2yK�ܭ��>���H�K�M_��g#_/��D�x8��|?�O)ʱn���̙���=ǖ{���~2v��[YУ�1�ُ0^��^��S%-k�����d��������*�cFE�����Ϟ(!�Tw���1���BF�OV�����q��&L��o����V��(�M��͚0�~o�����'=�����uK��kCqq�n�e�[¬wu������X�ݵ11�R
���	�X�U6��l��5��f�v1a555�ݕ�*�3�#��<�;=;���cv�^��n���K��cw*5�}U�%���Չ>�9�U�p�S��7V1��4�%S�rf�M�&Ma��	&,���<:6���X�hF�&��*v�'���}J����IWSzbc�f�#,�_}OLv+��d������������/J�h'3�o
�;�3� [pc��H�(��x�������#e����@^и�?�^�ΰf����O^�؅1����_�x^:@�Iv�u��Z.�y���j�Q�̎=p���7���]�^�4=��a�ߩ>5~�W~�>k��<qm��G��|^�������L's1��\�miW
S%�2�ZN�R��[�Ӿ�ݱu�'5a�ɜ-�t�k�ѳuk|P�t`�O�#�瓖�g���L'���@_���^"~k�*,�T�JuV=R�`(ŭ�ǩ��ޭ"�@la�f�jc��K�w��;Ua�c�~��f,v2���s֘�O?�Œ�}{��7yv�;6fvNw/7��7/w�u�F9�O��Onn(�/c�G�gwͬ��^O53y`��6��솄����N�ۚsxP�^����4�{D���M����=p=ݏ�W��ovgg֔p�_1��>/��;�sd'{�V*3-=�L��=��0�
�'A?DaR�$�+��5@\>ar�$�I�& L2@�d�0� a��$�I�& L2����!�W�p�����XF�6��Յ}���ʴ6�)a2����&a�i�A�&�1�=h�$��hH7+L>c?i�@�ٌ�ǰ��Q�lƴv ݂0ٌi�@k�ark���⎳\ƴ6 ݚ0��im@�SS`�/��%�dL��t��d2����Ӥ���y�ɟbi�$2������d��gY�I_ӌ�IcL�v�tHbL�cx�$�4�I�&�1Mn�����y�RӤ&�T���v�>�Wc��0?U[c�̤Yc�����$&��W�7&�#�0�i���a��8�B��Otc����&�1MZB�d��Cx�8�mL��th��6&�#̻mL��Po� �1YS,�0��ir�U6��I�w�c�I�,L`c����)0�7֘&#����1�p�����4	�s�DA�ɸ��"LTc�|�#���$L1n��Ә&i^��4&_�q�I���4��yWm�i���(�1��}�4�I� c���+L@c�\p�(�I6����+�Ӥ"�]�p��J�(>�H4c�LD�qT��*��Q͘&}��X�dJ��>�O,c�<�#&�1�R,���ʘ&~h�H��I�tt2��B�,�1M��g0veґ
Ș&	QR:�"Qǘ&騅���y��cL������@�(�4!���C� �4	H�!�5� &�1M|��#-�0!�i�#N����I��4�I�$��G���� a^4�I�0��d�&4 �@���H��d��)�(h%���)FCFC���HE�0:���0:��@I�A�04Aa~hb%�A���a�hB�|3Š$���d�?B�@(���b�aAh��фJb �p@���F�q��:h�V�R��C(��,� ��	��&P�#TQ�k M @X��bPAȰ�Є�5�&PCȰ�f��D(�"J�A�5�& �a4!���0�@�5�& �q�w@I�� @�]-z@�UТJ��"2�JD?� aW#j_P�H�)vE@�lD,J�U��(B�]&�
��xu"-��aM �d#BaP�!Ba�aM�$#�q���LdX��0Ɉ�(BIl���A�5��h�"���DdX�0ɈB��V�@dX+D0� a-�_����.2�5�E�"��AIl�� �Z�sQa-�W����*2�u�E� � $���0�0p,� �	��AId7a�al�VA#x	���
N� Ø�$�O7%�\�A�1�I��%�%�A�1��F� $�%�n2�1 L6B%�5!E�0�0�U��S��3
& L2@�d�0� a��$�I�& L2@�d�0� a��$�"�ƍi^�m���7)L��'^�7�~��.�7��!�VX��1�0��d8F2��"���c��A�1�c� �X�/b�aL�1�0��d8F2��"FV����p��?�KӴ���+�p}Y�Eط��|�w�����_����O��
�$,t�K�q��/�Nᲈ6��I'@�E�1�_�@�E�1�_�@�E�*��1ve �X�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b �	�"�/b4a�������~���mt�D��2�ۓ>�R�q䣛7o�KK�͛��7j
����o���������򙬟�z�����k2�Q4�@����5�A5� �0E��ʗ �n�֏}Y���|vM*�]���5��� �#L��0��v��DD׃�#L��aEG�L�bQƩ��L�Lo��«T�Vg6��yM���������Ty-7A[ XX�MJ-�%�«�МI4��MX1��f��x[W�éûL���՚)ۗ���#��a���h'��+�����0SX��L���3T�nUM�3�W�ʡJ�UQV(������q�m+�kx]�fl�=��l�(�����^��􏿰��w�x�I���� _V��,W������Iÿ|��o�g��ʀo��r��~a�d���WɄ}���v̨u��v9ƨ�V�5`򘙰�x*�����[]��"M؛|�JS�V��⩄�~���~d���;UK��%w�C�󺞘_tK_Q�𻧒
������L��*����_�.N
�/��.�uD���C6�c�U�?�x�����
��2��ReqR��ğo��;gRy*����0&���eO��6^)����G��{FM���:�?�6þc��F
O"܉,�E�!�c�Ipc,R�Gy����Q�|����4aq,��u�h�A/����x���N`	b��:��!��ӏ������Gy�0²(�>���W!���_&|Z��e�T����a�Ƣ_��Q��	aF!��V�G��Z���0T�}�=���°�n����k���u�;�FC)��� JR���*�Mց:��p��.��
�rZ�o��R��)�Ә�>�6��mEOs��o: �	g��a���0�,5�܊>Dm��W�h+֛��U�1�<��naƸ�B"�g���2l�U��PA����7���oP��3�6���{�Dꁂ
�>�,�ax���t��a�[���%o���WVhnEAX������������аe2�a[N������T���>�,��CƦ�9c�� ahf)�v��q涳�js+*�06����L��qH�8�x.Z@)��t=��M��F�@�Ď3ւ7��F.��V��Q�Pќ!^i�<�b��L&���&ON�_�>��L��t��֜=,����.����3�F�P��� ޅ�����s�\�֚0�ˉ�_����ҖB9	���+�X͞��la�'����
b�r�!l[�6�:�R)��j��0F}����}A)b�*�t�°	{��F=�嗙`�a�
3�pcDU|���z(y�/~j���=e��?-���X@�C;�P�LW�/��^����9�[=G���]ם�����!\�����Ӯp�ay���·�����=W	�r-�W�ӗjf�늫�^L���~�<获Z�Ӯ�(��X�� �pW�ҷ�0v���K����/�u·jKw a8�ú�F��_�\ט��I� �E��^�W���]F
��W;[����U~���?}�'ʷ��h�߻���{_�bS���������?&?���߳�d��m_}i�wc��&:Z�"���%���%��y�[����V�  ¼E�[���]��)��~��T���p@If�jl��Ύ����R/1�/�2�w a4�k�p1��N�չ�e���R���˰��
�ctN����xf�w�;���Ȍ���#��|1��V�W����h���0�����.a�̍Oی?s�ܟqa�W���$�I&�& L2@�d�0��:|��=#    IEND�B`�PK
     ��Z�/��� �� /   images/b5c34fc0-5882-471e-a80e-5adb517f5654.png�PNG

   IHDR  /  �   �Z7�   	pHYs  �  ��+  ��IDATx��Y�$Yv&vl7s�=��\++��WvSl�B���]?No��yh(�5.��fUמ{��۾���5���.��0 �j²�"�����g��z]�=n�����=n����������=n�����=n�o�q^n�����=n�����V�����=n�����=n�o�q^n�����=n�����V�)�Ҷ��^����^��yn�s�VU�<}��8����n~��'~��c�����mϵn|�������o��7}�����G�W���7]�o~����s?��{Q���s����G�k߼�G7��������/��~��9?o�z�W��ρ��eY��z|돎��~X���)���@����$"�_Y���+�?Eso�w�K�	��u|9��he���W��|'���V����;��&�sN���:��E{�:��z�v����۪��>���푦׿����?����H�=�������o�a����4�� /�g�r�����Ӣ����������깶�eS�nk{~���6Vm�m	�)�~����K;p6��e�Ȯ�
B�v�j�n\i�����u��s�P'�[�ں�@m��l��Jܢv�]|�k|/�߫IZyQ8��xR�����Z��ǫ��/�><	���,I͍X�mU�[�W7|B�u-�vG˵�&��q���3c=��>?ۮ�0,��)+7IS;Y-�t9��͑�g��o��mܿsm��8��g��c����������eY�\^�;���zM��2+�PJ��Kڢ���}�"h	y�����lm�*�p~��9�i���0R�v]��m�)��*�Ҫq�j�����g�m܏���s'�Y(N��(ċ�d[N萚�V��-�{č�I��69J�-%��4�8�V�$m8�m[7q5�����Xx���wm�ˣ�W͘�+э�}��?��3����T�[�
P� +w�ڙ}�~A����[�Jݱ�q�u�)��n.1h{��/t,ǵ�����S�����e��e��@P����-�]�s�������oʡ{oؒ���9]�.�|�����~�I��r�0��l�m�F�4�ʼ����v���M�v7빏�X�l��e��k�e�zh���ث��)�T�&Ib�uc�*�u.��ܮ��O� +�M��M�������u�YPF�*���MՅ�ͳ^T���U������i�{�k��`��[>�jIrm,����2�l�l6eӆC��[�\��j��ݰpۦn�"��q\I�7_@�����gx�/n���7A�%��f���iI���s���󟟷z�?�s����벰�)�mY�T��������_��ޞ���d4�\��9D�k��Ձٶ��N��SHڬ�-������<����ןC�y���}дk��7�����7�k�˷�h�{c\���8����;x]���|�X�alP4B�q��}�Z:�ac��O�j/�+|��ն6�g��;�m�s�J�՛�!�Ͷ��tP �-P��y�柵m9�����מ�f����?G#ߕ��(A�b�9/�����3 � (����ϱHϹ��x���'���\��Ӫn ���AP�mU�?{4�qoP;��4%�T�_Y�g���V�P��]5 $mi��ߺ��s
�20\b�Wl`K6um%��S��SQ���q��y�A��a��%�+�2(�¯���D!HKO��(x׆>�Ɋ5DxeYu�Zu��}����Gnvo-P?�,9�P�ڍS��4��Be�Q>p=�)�M�I��2k��Y{qz�_��z���-���db|^���sA?Q��1Z)�����.��!��b���3Y�m7��Ֆ
u�ST�B�ð�q]̩�En�Q�PP^�b�d�jT0u�U@"�'�K�Laט[��f��q��{�W��Uk�( ˁ� _8�ES�yY���޻s��w�^���̃j':��Z�,*;(L�p7��I	�ZE�U�6��BX�+>6�W�&R�V�4la^m� 1�.�n7����h����)	L� %�g�N6�0M�^U�.%P�e\@��^�h��=3Oi�Y�E�@�Y�+�.�Ұ�t� ���LeN��A���)!ٻ �B����X� ��� �U�3y~��l��Yo6��ɩ~~��x H�a_x��6Y��<K8��:7US��奓�3��0��  �Vj���*;��)��,M��z��(e���*���!�]P��:µI%05l R�L{�f�UPNdPJ|���G�?5�tڴ���U����,[I�1V ��"��s�7N�Y��V> 28�v2Y��e��I�����:{V��"/�����cnK	�B>�u.�#�u�Vo��@a6�s�H��p;���B��i3��q幐M.�E��,�]���צ���N�@b]����ȇe]��������
a�%�82�8��� ����?�G��o�{:�C�� �Pjù�ah�+�6�%�" \���� ��3	��w�Ź���/"\"R��U||P�@ f����
��O~�+�z�{@0A̽���؂�'q���x�I�cc�igY��l���pg�����ݤu۲�L��� [R ��a�~�i0]��^��16�Ty�*��߉w���Ţ�[پ�I�k����F�Ia���li��m�C
��x���/�/~#5�	�'���l\yr1p6Mϳ�f��$�ԙ��p���-g�᳗#��J7��w$K�>�o5y@p�4��ΑĎ�!"%���C���s!Dh϶15UNf�gM���8QQEf�� w]H��܀�۟o�������'(�-j����E鏖�8ǟ�j�j���E��ѳ>�7��7�~���ϒ�"�W��՟,J�O�ߓ;w�X 9����r)�H�?�0���X-����!�2�{�](o� ����X6�����G���'������|9�UA{r�in�p���y�����10�mp�7�U��lJ����z�/���N �Y��:���Ѓ֡�m�`8���L �a��Z@����_���\�+��X�kI�������x&��F�����9~�|�P6�q�`耴7�d�l�-9�&��@�ŋ/���id��0���6�RV`8X��>���l6�X�u�[[̯/1�a0<�Y�_�8���s��}*��������Ń�� X��òѣ����$�=�1�D�F��$4ѱY�����	� mW���U���!�1�X�t��t�e ~��7n跐?��Ai�~�t��%y���o u@��>�H5�iK-VAI� �x� .�r�6����k=����|��c����Q�����sC] l�µZǘ4���w[���*0�1ߛ,} �b~��T:Ĵ	��V4~�������rzz"	�E�L1t����6���F�!�u���=曥,.3B6�����f%���� ?ǺG���� ��06���K�ק{Q�痸���7+��`�d��$��������(2Iq�ߙ<�/��1h������ځn�j�V	�5�@9ǀ)�(��;������zl�4o��~��W�,	�!�Nom�X)�(֊@�� �ȋ���c��(�
ᶕ�D��,
5@h.`�2���dA/�i�#-Y�#4������<�3U9DV���y�b �� t6�z��X�r�Y�׳s/uB�@:������Z��*��-��
`ص��
	��F���&H��M�$(�`�uK�f�`zM�' ��J��]?�7I�z~:V�[ݩ`�������X��l���)�	(��s,�cy� ���Ú��� ��4�����b�������aê��!`6����+�?O�(
��`PS�+�`恒����	,�D����Yv6^�v�1�Y�gO��].7�w2`	��Dύ��Ջ�6 B5>h�������:�G�aY����dg*xnY'k>���	C���3,ÃX�#eq}R��Y��R�)L:`�@uA�լ"�����{������Vo��m_�ڲ��>��ϸ藛�a���T��%���y��r~T�����:I�A\���詑�B�!d�B�o�ВB�e���K���=:�鼄5 ��˃�� �R d��I��%�_�|��|/ ��BX΁��%�s�%�K�f���rV���Ee�����%X��A�o���hE��g�h�ƽ&  )`'
$�w|(s+Hj_EP�^� i3Hop��ήx�K��K&�\����PHs)�	z�u*m�	� ��P Y�q� /�s �w$$�*;[./���t���֏ ��)�ײZ0���?a
]  4�u>z����!�.�1Z�g�2�M�N=�Ge��g����3�~	�kς��q���ǘ�7���܋���\���5��2>�ɵ��h�� �u���sA�����+���� l)�4�s�nl|�H�k���J��U5�8�҅�)A������h�V�9!�3ηU���[*f\
W��˂�E<�����`�ץ�O�[�{��?�u�zmƑb��4Qʃ?Յ�{����JP���U�z�=�VЋ���|��+�~!�=#���
^tN{�&h{{z.��{������c^�b���{����}�`�r���K��Ç2] c)@[�?�X��+�}���C�@P�>Ѓx����8����&Wj�� W�S0^:/�F>;�_P��4�y�]��U�q K:�`����-�֋~2�F���9���J#��Lvw���Aۃ��:X���^Aն㩤��ϼ�-��liI�h7`��" 2��[�=��G����J�j�K�q�؝MO0@Z�.��iߗ2�S��/y]H�6��6 �+r~<�;��@w���v`*���0���b����
k�b-m�{���/��?�ie-\�MK�P�<^��G}�jA[ d9x%�,���<s|����;�L C�0���u���c<a���	���yX�Q��z k�m�����I�/fk��;Ćah��:��HR�͝��&�?K t�n1��lV+x�\td,�^���;tFC�-���N� ��$�eSd.�����6-	zz���/4טb,����\�ox�
�ú�d����~�E�*X�	,��J�R��G��<y�޻wְc(ꃃ=�Z_i��)���~�����w?�� �d������Cx�2l���;X� �h����\� �C���݀��td6B5�%JbSd��l@�KX�T/�ۡl*���\����*Ɂ�wp�]z6Ɣ*@ɠ��	¾�K�BAe[�z��{r��*B��0/^<���7�y�!x`ι�xZ�US���hCo�� ��qsb<. ��C���.�X� ���� �����d<ѱ`8����ыõ	!X��H�O�W��k���
06&:�XB�#�g�2�C9[a�ٜ��(�0V��
�%�c�7�;ZM
�JP�(^�6&�e��e]��-��{T$��&9*d*=f�����������g���ű�z�kD��]/�0�ؑ��4����|����ޜ��B��!�k���� jR� 	e��=�g��m����N%�#���d�~7�8�(��T�5� 7���9o�Rٶ�̧���
�z�'�^�kG࿱�H�a�V$1�@ Wf� �T�S��y��s8���F}�c�kvz&�/eqr.�C� �[����L?����ٟN �p�����L��|.ǟ|"S51�Y�����Kzf�a�)�s	�PX�����z�������\6� �5ĳ��:9lл�V0��" [�����,|n�^�h�vJIiZ�W0���]���ćw$9������t�֤���%�O� �I���_�� �U�c��f�P��o0�<72�x�F���FX2������߇<������%��鍥���aMK���Gc�)�aD�1Pz|�wk�m��zjq-�H>�"W��CY�nq." =А��	��A&���ex_��>ˊ�;�
 fi�� KiRX��j0ߎ������9�r���qz�w�S�8����]^��t��.��S��#���K:���pf�7�K=�Xk=��2�`l9x,R�q�4q�ƌ�I<�����z�P��$Y˪H�6�z���S� �-������g��F��Ƿ� qx�! �b���s�?�9v�3n:�+����<x�X�w�P��;*�i�*2.5� ���:�O���L/y���R��^<�T拙*��^0�t<TF'b�JD?�ه���/d4�@��X��G�����,��`�����a���s�W習��c19=��FV ]Q��6����5ߌ�2�c���� �!�&�<{�~�2�ߕ���`\��TY�U�y��p�|9�:�eI���j�B�ߓ���)0R�q� �a������޾��?�de��e�5��O�2��&���ف����(t�s��C�Gϓ��z��r��z^X�	Ab� ��sӵMAixt!u�c�Zzi� �Q�r�%�ű��p�h~�zu4��{�;y�gT6��qN@�DLnz\z�sZn�>H-
5��f���j�=��Uk���\Cc�&R8��tkU&7�� T6v͐#��,��re+4�3��+�w� |)��e<¼����Po�|����T������0�̇�A������ ���lv�a�hK �v����|�艀��bћD�@��	J�4\W�*$��9Ǣ����@F=���W *� ��܍�ܻ#�q$�P���3(�L��(�$�P8t4Tp�.�Kߦ3�U�2�dL��ͩ�K��K�C@?�xR?W:�y�E�oz7B�K���Q�Y���i��U�hK�T�OLP �����(�l��窠�yZ663�k�bR���nB%��T*(1��֠ﬢ�C�jh� 	B@,�t���Ω�#�S'�z��&�"�ùn5��$`�]�2�s�o�r�k���~v5p�L z�&ߕ�c�-%A�c+]E0R*��z�ʓBi+P�x�^j����2C��h�cſ <�Q���d2.�ڔ �Wꭤ;�<��&Y����U+�>ڝ*��&�{�0���=�u�� �0�}<o������¸��%%A���ϔ�~`<��5n 4j��w4����� 0
W[��69�������X9 2�ۈO�B`�����xc�h*���!�O�V��������봽����rYſz}/���7�L�A(O�{*��=�=�R��X�Lb�
4P�P��8ԭ&
�U��O ��d!Wg���\���}�UҲ�+#���+r������T��`(p�	,(��p=)�n��1�(w
Z6P:����j%� } �/�/T���L�&!�Ok��k28�旭����ă��)��! T '�#� &
jN��%��q�y��syT&E�3I�|����A�������Co��������?�2�S0t�&�}�^�Рާ��'���������l��;`Ͼ|�^.��.�3�ng�Ka����c^�T�L����.י �˻!pP#��$֠�����<�J������e1�%�sLxln�y����x�*,~iU�]�"��8���c>k|��}����kBQL���B�!.�&g�|X����{�� �h{������\fJ��$� �Ihsl �L߬(���v���g�*'ڋl�y�^�� �K��֤����2�?����ІH���ל++�1����
�x[���ܖk�ZP&0,,�.=C{� �!��Di���HP1�+�!@�oAѻ�_񤇹c( z��Z��D��hV=��B�s..����5cg h�z�Y0�h��u��3��g�Wt<�W�Z8���KY��o%��{�.hoW.s�����e�sD%�5�./�Kq�l%���{w������3�����\R����*۪0<��=3�4����Ǐ� 4�a�
�����kr����E�K9QФ�:d�'����D�?x$�G����,+53��#�De>(�Q�����@��H�\/_�xVk�|)}.��p�֣IO��5�k' /`��6��0e����M�1=���T�'*�'� 3ڧ �u^!{ �\�?���C�&�N#	s� �|v)�� =\�v(y�2��!CdPs��ХDi�|ȶT��e��a"0�u��³Ԙ���[��3^9Љ�24�K��0���P�!��_�;{�����aM���O?�����	��#H�+3�`�ڍ�`�J,6)��}��!1[��Ѻ	�.1�>Ծ>+��7�B����2�����ۀ��	X+x`��9�a����҃e�\5�T�J�x�M<@�*jU2/�1c&N2���d�{�ߕ��L��o�=9��'5��.�@�0�3�+�m�gZ�Z�R-V�L!�\�x�����Lv�ñ, d����T�F�ՆnO�Y�󋫥
���x��rl'*&)2��g� *(8\�JV�i���t���DW.m8*��V���i1��9�3eX�qm�;e�����@�HT��%ǹKXo!�Fx�c��V1]���4
Z�V�]䖮}<K��-F��6SV)C@8F��9&ߑ��OOϷ���)��8������������F4u�iN�	K�Zv!
h�BE7��I�Ck�~�@��\� cD��i�®\z\4|!!s�  <��վ���XNc��µ�|� ��
|�Q�����#}l�X��^V��b��T��)TK�KQ�  H x(S�O0�@�nq�S�c���uc�j��3tDEϵ�h` $Ը.=��yQsi�WPt�U� �˅,�������d2��Z& .��c�d�aB Z��ƨuu��)��=�ޕ�P�#���!�#!>z%���������h(�Z�!7�� 8OR(=v/�����Ǵ�LJ��� 8�㍬륌�ԪA@�*��(��`-��:F����y>����O������G�zi�[m��9$L��=K(x�	>s�I�|b�"1	�P�9u1��ũHz����j�O��3z�Kp� =+z� �b7T:%�m-����(�|04�<���W��i^�ȸ鳚g ����A�%jW~1���Eg�����T�C��d~�iJ-d #@��&�AłX*�f� �L�VO*�!�+��i�ѐ���%�=���������YI{dҖ^�5���U�1��<��?ԧ���+���h
��/�zM��۳1�J�D�lԓ]k��O ؋���e�e�3S�ިG��eQ��v2�[����ߚ�����w�.�ÿj��1��C�F+�b��8��F*h��k0-7Z"L��)a������J�R�l�^����<��)p� �`J���I)�E�ۓ�ҥ�
����9 4��#c%�Z�.�I�EH���
�ʃ�dJ\#`��h*����!�g)>-:�}���,vn*�\
��.�ڈ����� `���\z�5�e:ȸ,M��61��QA9T *(���!	�����]q{#q��$���z�2��ߣ�u2 EO��Ru�Rp������`���Iv�W�t�g��mU0n+�ԛ��/ݾ�0�2cr�9��Z�+�F&�嚻Q8��x�B(��İ� �J&Gb"M�%P� �G���i���'��a	�e)W���*��z�������}v�Y�=-�i��߯�2Z�ժ'�nmU&���Zuӿz�V�8�ߢa&s�>���ꚏi)��g/0W�=!跆��La����1)F�~�S�}���5Qjb���ߖ8�m�Q��.���	��<	�a\�(K���5�(iL�WE��U`R/��)�4Y�������j��M�e�6��z8�jӵ��������d�8�+��RO &��de�U�&w��y5���4�4�|��{2��D�y��|�ƪ��{ގ�֙�B�8�X-i��،i��z�
&P@~�1��̭��;̛��6�����xg�&�HOFW�
Y��pM ��b����Mz�w�`�a�|��,3�_�����
�	�⹪�J���\sO�VA�K������2�P<>��L4�XLC�5s\�-����1d���)�"��� ���Åu���ԭIVH��)_�'�H�|m��',���[(hs���K��fJ�`mI
�=?����G�[^�h8���#�商i�G���i2��|O#�y�. �
����+)1�
 ���F�C@��}~�ϼĵ	��*)�X$� ����l���f���p^jpz� '��{��j�rMȋ����	hw�������V�ROAR(t]xj|� 2��Y�������C9�5���\-�$���	_Y�<�]ʹ�y�S�I����l�N���PvL�ru��?cڊ2�N�������H��	 T�\S-e[+V��ε����hh�;S��<��`�!C?eJ0�21��}�ƍ^e�Zb�L��ݣ�J"5��^Yj.?2�X6���t	�( 5�"����o x��a���P	A1����e����Rݔ��SyM΃IL3njEaT@6�>s���!$(B�t�w���� tT�����1�a
����ju
X� �f.B�9��HD�>�����$;Z����6CU�
�րy>����5Sw��8�t�K�Mo�a��8	V��$O+�<٥Uf�Y�lPʵ��M�K�ʟ��h}��bBQ�^ZRz�2��\sE,�04dI�P-�FC���i{_��a��,B����e�1�1�)��70w��-�0+��GïI���\sc�9@P�;�*+��I���U�� P����Վ0�6زZ��ϕd ̿��2}��
���á��*K=K�;�<E ��1��2�B@;y�
J�Pe:��d��\f�	��݄��JZmjbU��n���I����?��D�����b����cc����C|o�{��l�&T f1��!�
�)XTj8�Cù���#������r���#�͓m�u�u�0f��h�3'���k�p��!퐹�A&����F��[�LRR�	��#:"8!o1ə>��cx����s=U����a�X wv���:c��)�^OF R@���G��Oz����T��� #%����?�U*�߼�� �fg"%� �����aps|���Ђ�������	��s��񺘭5?��aߴ�#�Y�ytv�UQ��`��V�T��2�zp�X+���.�_���^��a@E��{�C��� ��H^g���ü��k?��Q�@�R�0&sQ,������o͕�iB2CsZ�
ټ��Uwq/o�=�1@���Ltg�[ߔM�{Vs!狼���:�|�J�����m/2���j��l5����.�v��baBfe==(D��n�hB�&���`S����вK+ A
��ZO���eՍ27K>�F/��r#>в��^W�B���M�k؄�G*DW3�MX�
�b�!c�N(�
B�v�W��V
��7I���P�8�������X���Z�Ҧ�ӲH�j��kZc��Y���j.���\-\�\�fZ�OF�胥f�|-IW�[juC��0�;�Zv-�G��!�9.1�x���"MƱ&����)p���;9������M�/@�4Y�_L�^Z0�3R˅UR�L5�v%ӄ5������V�����U���.V�t@``�xB4�GA�II�te>�e�ں�`@h�q#x���U�RW�ޖ�s�+Gkr�o�m�33����m���30\��-���4�qh�����ҴƓ��<�<�y�4E�0��'&�]+�SA��5������l�:�`�:�M��6tq7V(�Y� ��ys	�������Z�˙i`�)bU]Wg�i�8�����<���+6��'P��[��X��g�����XT���#��X�ؖ�ٕ�������#��tS�`�9,�c�&�!����b�(�i�i��S/����̟/?� | �� ;m`���s<��
���ؚ���2��0�i�݄�zh����^)��PQ ��)�>˕HL�!M����9��<�������3 @M�`��\����}v"���5��W���8&Ѽ�a$�����\��!_����r�ņM�*�L}���,�)��dG/�X\H��a�+��O (Nf�OC����y����J���L|�V�X:NH��*�*����r.�h(��x8ּ�r�y�ڲ� sp�����"��#��)��FF��xD<�޻�/�I~���=��)ڀ1�d67�K~f(�!��S�#+F-��H�Ҡa�8�u�m��3���"���\�m7����h��]�{87�1�EϹ��#6�,S0`�{�9��T���i�]��V��к����m/�`������ۖvqy�	�UK��U�-b[sl-��'C�5����2ƖՃ��.�Ulf��bc����(+/ػ�]aC͙����/��BBx@�+,$�d�X�W�!hڍ@<X�O���^j=��hy���r�8L_�J3ٴH�
XqB��ˇ`�]�,Z�Zq���x&Zጣ�u&bʿ��*�,����7 L�����ҋ0U��VE���~T��%D��M�5q�@��9�zi:��DȔ����Z��
PiJN}mrGO-��)ȧ:/�_k^J��]S9���U��
P�s�M���ƫ�U/�G����AC�M �6_�Chqv�__��[b2yo �-8i:@��c�w��s:����b�ٺ��"4�9��E�鶼G
����G�Gu�;�I�5	N�h���d�F�(o��*p�����PI��Tk;V�a+-MV/�6�5I����H:m��Ԏ&^Z>i�T�,a��ܙ�1�2O�([(d}~ѭ5dK�����2�\�"��&zL�B�L���g�6����z�ք�8>zY�K�X����Z2Ϧu@��6��+(�s }w��>����#A�
���WP�-G��� 	�P�B@��b%8U��d&G'���u�{���wž�ˇ��~~$��ە��P���i��HŽ
X	S���l��hK���5L��/��Ď� D���S��腜(0I��~�cك"�Ħ�ZZ�\��ə<��T|V��������Cpx~._~"��R�@X&4b�L=�B�MF�1�(�G��CO�l.��_��'J��K	٣ �t��CcLV=�D|\`|,_N���phcJMͶ~��'g2�L�u��Tb��b��J�&�����(��/��k6,�|�󾳳'�;O4����A��j��§|�X��e��S�b���� [��x�]��a�T��1|^V喖L3�����S�ZӃ�\,��m��S�c�c\g�uP��I�u,?ϗK������!V��:MŉLE��iG�7I����m/�_h$o���W�r&��5N��d�XD����ب�A���ʝ�#������&�8��Y����+Y��  7�3MC2Z���:b<�!&�Ҋ �)��rHkͩa6���NiY�O(�j�j>�)O�5q�U����!$Nώ`���e�2E��3?�IveY��+�� VxdP"��^�f�' ��3Ǥ��ˎ�,�\]��,�����C/	�ڂ ����Q�J5ϵTIE�0,Ш��yg��,�PT�v��aTt۳:�E�}��Z7�zX!�gFa�T7*w(6�d=fܳ�4�
1`�݂��sA�mo���FVm�U���"�[s�����"�Rn�Ok�^��ι~�3~��gb������������ߐ|�;��{w�3�'w���&!XO4�T0��v�
x��;:���	�w�u@����L�V�[����=M2����z�!CO�1��!X��|�R���a���ٖ��P�Ky�����m�[f�{؟jȘV8�����賕���r��E���l��}�y"��R筩~ ����^���X�Oz�|����!Cl��w��q}iX���\�x�&�L�ldv6�v�a_�`4|�[�����sq���Oށlj"�Ò/�1�y�3i�g���W������
L�k�J>�"m������P�G��OG���k��L���� �V
�X�|z|&*Y7<���}��(�J֡x���I�T��;�?��,ծ���ںao��~ۨaA�� ]�Z` ژ���\8�j�\K �M1ƶ��Ƌ�i�:&�*�l�31!�Y��UUЬx��Lx�ҒovP�1��V	���lj�0�+}f���*kn5D�j���a�d�@��={S�C�-GuA�<C��W�Ģ�T#�Q�H��Ѡ������~�J�"��l����2dB7�I�N@'od�9��M>�h�k�Л��H�-���u��1C00G*4���7��w��V��Z[<�V��^\^��o~��
�����~�].�J�a)1dÌ�����4�
eZ�L�e��ׯ�ӏ?����ruy��B]������d��1�����0��!��2޽'��|_&{�+F�5���7E����B�Y[����3�0	���q��*_^ɗ�>�\`�b�:��7�
o���2��PY���Ժ�6����- H6`�
�*�M���.f�0��Npm�֫��Ʋ�L�5

��k��A�c��;gK` ���a�b�f=���ZsK80R�����`ƩY}�>�eJ����Kj�7Z�O�V��X����Bm��ĄU4��2y-ֵ��3�$�-�0e;���tA���Z�������(��&��Gzl��|�|u��mΓn���z�H�
�������7N���oM�n����/�X܅69]I.�G~چ��2Ep�8[ό�I�M34�6T&��=_��҄O�&c�pL��t:�����������{���mtc�I�4>bV�Ԛ3E�� J tԚ�u�-U����Ţ��1�"�z}���L�\숝�-/�8�l-�ٕ,�O�>z.��CU�Zn���T0ׁɞ���JݼReh���	�'��{�����#��c�&.�	�g��I 0�׎���`%�@���'�j-��5��d�q��v\�T ]5�����JT���Y"TU�$��3vl�9+��ˋ3�w_����}�����O>Ԝ��>�k�𧥞j	�Rso!�׼� fKɘU�r	 u�Xh%$�fl�����Ō ��M��� ^�ɦa�k�7+�J�b�9G�e��Пj�f��c�!wٹ[��k����a���@�$�c�-�j�Z��+��~��	��#G�w�|M�e(���a|&GG��G�%�d�#�x�ބ%�z��]����}yr!�NO�SٻwO�{;�<�}��6B52��2��b�0��y�s�V�Ҡ�\���n�7�6�dn��*��vk�S)m����ܡ,د��VF���M|��&��ݞY�b�K�&f+��婺�+އ bäJ�M��&�V�(��'��S'���
���7r��9sL
X�=���k�h^H�<_ͮ�F�%=�]%Q��l d��?�ݻ��|���5�k]C%S�c�J�+M����@@���:y��j���Z"��H,{�4���( u�2:#���4��}6+���Ñ�.WsXk��ɍk�m�}�(��v��sKs*��(ZL��}A,Uc�Zr}`�N�M���� �л~�yL��� 2@�w�d4{���Zi�a�N�N�]?��Kbi1t`��[o�t���K��h��6�y}�m�]mmb�I逌9�����7�k�W��@K���-�����sl=-���r�g�+D]w=&��
�l7��~�͛��:��n��9<�I<�m�g�u��z��I̦���/��o7��5/\C�kE��K=x����nAiXy�a�-¼���`l*�+{�+'I+�d������l�]N-�W��V�(_����\�W3�F9*6�sF�L��ZJ��-��G��l�� �{;��@�w��8>��щ���8W%�X�Ȁ��]�	�8��n��]��J@��io�M!��%K������P�H
�@1�F<�/%�L&z �4V +���l�G��i���\\?~p ��]]�/���Vf�_ߋuMR�/�5ݬ�:�c�g����lt>3����ǭP4L�I����9�Z���`��7e���F"��
��Z�Ų]v�.m�b�*x�p���RnS�0=�]R9=m�p��^d�/�~@`��I ��h��ZM/�ْ�V�����.%N�o�V���B/��L��3��޴3�I�_�~#o`�.�?������lcʖRS��ǖ���ƥ�c�k�I�y�]��# �a${ai�	���]a���gG��1�g����G$ӧO���z�-�߄���eX�r�L�����K�Mf߬�ˉ�XI_K�5*]vmL�"�O�َ��J�F�p|�!�I�z����'�;||���Eޫ���> ��� ��d�y�V���˓�1i
nq&�ӂ##,!�^�|��F��SB�>܃ d�!P}�����Y�Xv�L��O��39=z�-�i��D7ݿ뮯���ez�h{x�s���"�8��W���]�`�̳�5��8<��
��9> ��i�ƴ�'�1��UB�<�EϾ/���h6#����2��2��|����.�k
Ǿ@~�ĸ��J���`v���̓h��]��W�$�� S���@�f!�ezK�Z`Y��V*(�`O���G��UmU�O�*�t�S��m��6�xF���]_�.WF�k�/�t�>��Ϙ�P��sy��hn\���D8`���ў5����%[�b@ĶW�u��#o�5b�<��׊I�i�e�6��h��۟��^$*%�tb����J����寶�yT:�u��wMg�v��4]�k�{>[���=ͯj�^Z[D�Q�F�Ϲn��GL��i��r9o�a��[�c���t�=n�eq��vc�S�{-%���9�F��({eHW��4��w��������K�>����{��D��;�t�=�BଥŽ��ѓT���	Z�^�J�Ds��笺�]zikWx�Q��ɦT��0�!�A��'�#�pK��.�5#=��v�.���v|�P��"��E�#�������j3�F�{�ޫ�2=�W��hO%n�g���Y�
�Y�-=B�m�Y��+-;��̛����3k��<7�ˊ�|a�h K��C�0���҄1ޟhވ�K݆�$��i�e�w�%�t3AI0s�Sy���TN��E���w��b��~2���N5D�t����v�0O����T����do_+v�._��^>ۼbG�Lޙ�WQv��"_i�5+;�ӊN��!~���2d}�h�]��6�
s�N���Y%�� �h�Ho�'O�_��'���I��iG��W
&�*н�.N.��9tϋ�2�L�╤�+Ky��L ��B����6��̯.Ħ'�6	��O������nSnR&���8��w�҈Ƿ���b6�!�2ɠT�,�Ӎ� 8(/���T�lOm6��*"XA�;=>���SY�g�����P��X����R7.dH�[:��h����$E�k@��x,�^���|������J�����7(3.l2"�.y� ���hs�N�0!����K���2����?���ky�7#���!{%�$�~�ɹT&��8w՚`윱UZ)�d�u��l�+m�E}��\���}�A����LE��cMr��b�P]f����M|T� ��x��1�W�#��5ļ��U��1�VP�@ �a�ګK�����cgGd��tKn2�s��m��H����5�ح6&-�.䡽Y�y3Z*�ǊV����V�� n���Rꮍm6<,�n�Fyw�6n�/T"Z��%�X�W�|f��u1�~K�m�Gi;O��*&>v}=4�e����t��� l�����ZS�mr��G��h0�xg�-���Kb�u����
����]o�y�5`�,�"�/Kd�a_��}�4gk��%x�X���
q$;�C� o��}y����0�Z!V}�-v�e�6��)؜�5
X�Q�)7�o����rCU&����`ʉ"���n����
���=�?���U����ikˮ���~+�8�=��񳒪�w�g���>7Y"���P�;�'C�$�hY�RoL��}Kبq0�J=ّ`��&�P��e����ď���d�Wg	�zq�K�7�1<����N��p^��[�{�s/��P(J�?�x�#�ݩ��K�(��x$�`�j!�"̩�X����	|�ᦳ w숻��>��� 0��
r�H��'�#�M! `TvtM��Nː�N���]�ۣ�S�e+(��w���}~9��b�`
��&����fm����9F�����2��Ν3����a�=���G@���B�)��j,�Ȭ!C�I8����tUslG�P�3��;;r�%7Q\��E�B�r�{�9=����@~������ }�����/@�d��}�HO������:�������C���g ����; R������w�G�"wE�m�������k�>�Sx�/{�E��v�6�O�p��[��/��Ȇ��5煙������%���VE*M���%CLgG���+�İ��>}W&�P��@W�T���p�Gzt�i��i���=^S�A*
�a���?���
�p�|��o���X�wv���~!�M�����
���m^�Z�M�{��Q(���[܇��<�PۨHpLԄ�zN�lTƊu�_�G-�n���I�L���4]~>�\����͵�M8�^U>*-��h�Q�%�D����;�����Ũjf2�%��u84�]�8��������X����ӎ�f��S��γ%{�hu�\����醑7�b�����Ʃa�B��VW�Z��Ґ����i��t�
�5ٽ���D�0M�%��q�ۘ�����b��u�T��${Ⲻ�[�t��ƍ�����׹.��H��+�]K�P�$l���T�%���3Z+��	�A�μ�*�G1��gS�����Az������@O�j��t��Gc(򁆏�K�\^�x:PYAЃVO�W�������$;jӈ�����<[�u�	�M�Xi�I��0����-z� >�>��dh,���ҩ�~�o�=�p��/_�g�}!)��1��9�+�ܻ/��=6��ܫ��7�L�9 A%��!���ϔ��$K�H���?~_���������@� ��D�^��X��1�ԓ�'����	�rK�sM<zp[W�5ϏN�����Fi���z��/�d�2���9��ڳ��w� w������z!�t�j)��-��H�GOE0�1�n5ؕWgsɡ�/0� O�6!>��_ىJ6�܌d���49�����O��>�3�V��%�F��Nqk�tc��:כ�2w&c?[I|~������a�Io~%�H�e�J�l����~��۫5<�}��[y. +�������=l�g��O�ݻ0.�T�LOί��O>�_b<C�������>�:}uy�����W�_~�ew:���*;����\Hsr.����@������-ǟ~,;x�s�ļY����=� 8�3�:ۨ7s)#߄�t(�S�L�ܺ�U�_���z��� ̳���5&��b��{�`�].f6�b_��q	%?C&���ְܻ'�H� ,�C���34��$,s� �
�/�$��ϩ����DS��[�ݑ���� ����A��޹+�p
�7�4��fy�Uю���m��^4|���Wr|�Z���)��G.?.IVea�3V�:�|V�\X%T���홍'��1�%�	��d,w��ա X�Y!Ȃ�ں)���I�5e����<W"|��2ˮ��6}c��I��t!�an��]aC)&W��Y��R���,[u��s�6(d2+XZ���א�6��M�,t���S%ÐR׭U�1��>Va��S�y��쮯������s19o�VG�V�	Y����4]xɀ�N�7_���<����Tm�Mosi��:�y�?�n���Bi������|hH��i�{h��k��_kӰ�<��Ti�H��N�1]?i��b���g�8�e�峄,ll�n�ǔ3
R���h(�Mz42M���$g
}�h���F���r��P�ʟ]sylu�M$��mfϪ��ͳ�ܪ ݷ��MI���c2��R��K)���!�[���bM`lf���#��D��Zf ߥ,��6�U#6��|>�# �s�ؽ���Da�ϒp��s>�T֕��=(�;������WZ
��֕V��w�e�> �䎰W2��iÞ���+6�x2 py�?�T.������H=Z����W��	,yjW����²��WɀI�l/A�O�p�~<�H2(�Bwg�3 <6?��e��# �]��c)cX�XO�D����P-�X�H�\1ٟ��>�f��{��D�"/{��{�
��������/X�R�������b��M���؁���8�#S��V/���_�{���#�w�H~�ϫ�
P�ʆ�k���QI��U�0{���!�9N�h2�&��A��s�(ߠ{�Ț96 �fv����a_���W���sy����CL��B���&��b�-&���-Z���O���c���'?�� ߓ%�g��{Y4��WV�~1����3٘�����Cd���6&
�-J���;||k��;�<��Xū:O*ӱ�W����eko���X�İ�J�������rq�}����tG�@��4���x0#Kؒ�B;.�!�{1�M���`�f6f������n���p Ò�_|����'&`�D@� ���L�f�W��̪������B�'g���KTνzt�^�^˄[���RX���V�r�4�EK'5��4�#�V���	�o�0�M�fh簧�z^0ޭ�#�h���V!�9��B�΂����h
�-f��P�X��r4���52�u�d*H&U�� +�m�I�Qⶮ���)�
H	 yG��7U/�ez�Ѓ��y�b�˓���w�$��4��ϊ=v,�%�.\���p��AB����+PjT�/ֶ������,M�6��:i�f��>RV�U��]���uZ��=w���Xo�A��^?w��D��<LM�!�zh�m���lP�wMR�AZ��H"�1���04{qi$�xtl 	?`��Ht? �������A]oe����NA���/���|���˿����;��s{�Mu��iIWa�p��gYlA���z尖a��Wl�ry%� �M٫Ƶ4�C@�j5��+�;���;0��ƫ�$}SI]�H9�5��iX��ơL�����3���2��|�����ٛW�׍E¼n�A�0��TP�9�
s�a #���T���Pc��I�R� � Ɔ~�0��{O��?~�r�<�)d�	���G{R�w�x�/ON�׿�@泥��
F+^�8�����kه�gK���]y����{,w�{�|s&} �����������1A+��]����@�[��!�/(��熎 5}��WϤ��6��B��\���)�������dyv�X��!�*�'�ew�@墆����ǃ9�̵!�����˗/�� h�D��xn��]�Y��� l��s�YBN'X}n ��i4�������q��a�ke+��~N�n\�}y�䩸{���j.g�+ ڥ\�_(0g����|��gj�i����|߽w����N/Ӕa��kX� cy�� =���Pz���u�d��IC�����4�/ƣI]8�N� 3��Gc��m����s��]/�ܶ|7�.�a�(��7b4V�Ixd����R���{�������ݬ�2O�Z�B�F˕qq'�L���)����$m:zZZ������ىv%�Ɂ�M�U��O^���2� � (E��4��`�:�U�С�!	��}\��+�s9��'���?���L�za����f_���EZ���A��z���Aэ�p���ucB��V"����n̵���j ��|�j~)��c)� .weow���so���^�F[[kb�n��s�/��`>{�0F�RQ��f��.j���f�[h<��aB"��c ��lA�6�C�*"�x����ެ�Zf_ �	�'�3c<-����A����1I�bJ����:�ʶ�H���ѼM�տo��pn �����
�n���X�׾׶�!�� �������=�4H�Uti2�ֳ�jO��V���1�iVP���2�j�����v̞Qҵ:g/�F�:����=Y�Z达��w�=��%}m�y�������`y$��X��F��n�3�<.�"u_�6�n�����K(�퓔�g��$N[ﵲ
���U�����͑\I��ǒ��X(�v��f��n.ݳ���=���ge&���l�f4���&��W���D�[,�s�F�'}'i�1L5��DdĽ~��?G�ӡ���v���Ɗ3y�lO��^�8<M��+��o�5emmEj;79�>��_v�h�D�GT$1�?5~�#����u�A�o8�ވe��'�q�!�B���Y�<�l�=(ؾ�s!�D�oЖ��4t�^ɟ��Z={"�?�	��r�Q�K+(ɫˮ�'�<�i򓓍����duK6��lT[��kz�9���� �K��&LSY(0*�������Y����	��P�Ӹ�q���/�6��#��M��
q7X��+p���'�߃pkE��-���N� 1Ĵ�kU�"'/�m[O�k��l�ӚU�����9)���Q.�:�JS�&�F�� ci������+俀��=3kX.*�jk2z[D�﹂ۯ����3��G�42����p3���*�(��s�Z=Z�=B��d{����]�m	�m�v\��d��{�i�o�I�q<&���H�h�M�$��H5��cK�=~Z�x�ANgSͳ0~��,#c#�����<�پ�H�M�icc]�*5%@�8o$\�-@��g��ASP��"r��4Du�$�fm��G�`��k]��v�28@Lw��O?d�A��$]8�W �Ƒ6	3� ����(x7����Z����%�#(3�;c7M�JZ�;P<�ߣr�@��i�08_L)�1.�l!i �A�ʦ �Cr^P�\L5���n\D�yq�+���Qm"U�i��(ʱ�B�~R�^�ns�����F�(ͦr|��� �T��rc� %�["(�Usb<37?ܬ2xF�崎ӊ�4d20���K�,��:G���Ti3uZTZlT؍���Lf�)o]���z��\!K=��Z��ڟ��3���R��u��r��z����g����mY:`�����ԍ�9+� �N B��Ï	���֡j�4��X�lݼ��tU3�%���7��㵠����{z�u��gW1*��	�D}�]���'��/��4����"ӷAk�" ��sU*E*َ.�8+�"=� K���Sy�r_?_I�Q�jM��'�Ő^;C�>�[����53/˻��-2۫k���O���?�bSn��1���s���˻
�VjT�vƱ�2+[4� 0Q��̼&*PpE+���[7w��^��t!_?z"��T�{�\��͟���#=�Lۻ;�����AUhX�X��fG�����ʯ~���߸�$��jJ�Yոv*����&SL�L(O��y~L
B�
���%�9}�����%O��-�^C%�Xړ}M�
z�����`��nC���?����ޖ�,�׺�#ޟ�&��� �5�M�I�4��sK���C��7��x���{�d�5�Wй�{6	��Â|?�5������T|JA�j�5Zl���g����u�ђzkU�
 �����}�����]k)�jʝ;w���.��wO�c��(T�k�:-4�v��p�v���7L(O�+�	S�?��du���qv��'c�UJL,"E���*�~n�@^���<k�� �er �bB!�"*&=~K���ؒ[�����-���nzZaC�"RU^����� I(UZVkj�̖ w�u���E�_e<:�z�Fk��4�\�Xl�EN�:�i|��:�"�@���R7�xЗݵ-f4(�⠤��l���g���c�jł_N�������'�D�N��a�5DT86Mq8��F� g���ׁ�ĭNO�	^L�Hn��2��X�bbm�����R.Y�']�����R��qTXuI������6��KG���� %��ǛЩ�'�@y�Ղ�]A�<<��ŀ�*&\�9\�^I��o�c`X߆#�v��[jb��>��z.�#I�u�x4Y�Ǹ1�a F.��qvǌ�b�-{όL�dm��
�P�W2B�5p���$e��s���7��q@�o�!�K�,���"G��'������͍-�^�d��#�!�@�"X���d"�|�����g�ȃ;�2�^�A!��B��9�
|��C����G�׉���+�9ǠA��.�֪E"Q�=;���P�R�%5+�ȫ�'l�9i���X��v�����QQDV�{���^���~C���˷Ϟ*ؿ��e_VrE)�6�ILB�z}��EGb���F�lhqAt2�{�ZkJ�Vԃw /�<�~�+�+벱�)0b}���|��9��&��P�g�����+-��'.Q����C=X/��͡����buU*î��g�z�àn�y4�V
��sb'`��a`���GR��n�& &1j�,@�*����6���״��?����I`[,����rtp��+Q���������
M�^���M��������Ф-C������H�����N��'�o�t]���]�2��|�����������9��4��-
4K��}9<8���i+��s����xF�_� woݖ������T��P..�Y�#���>P�������A�Sk��$
z�,���V�B*�le��T����H
ƹ�G�������?W^~(�8��:���v@�pA�F��qc=h{��z ��K��'M��)�-���g���v	W���������XjDy���Z�+�b��g�oz�Ayu��,�(�S����'��!����PӍ5��G�H}
�x�a��R�n�r��K��䭤�q��3������wN'ݾf"}�	�c�C��ԃ��`����H.//eпd�Cp�N?�G��5$pB�&QIBT��zr�y-yN��ȁ��ЙZ�rĒ�G�&����3	}��9����gbtv��ms���ҫ�F�H�~VUIl�f���ת^��o� �GqE��kS/+¤��3���w�������^ME���:_���˸-��$P�G ��qs�{�﷓D���p�*��\2�c<B%&�ʦ�����l?z㊢kB~�qf�E�i�j���=HSi��!����O�?~����� �@�9���O9��9Q�|ّ�gϤ�ky5��ʟ[�-5_0��� ����k�N��'��![:��b"{A��b�jb1�ʚǊ������C��S���c����[ȿ�ۿ�~H2ZH���}�ʳ�/�Yi��'�^�sp ���PU��hȇa ��j�J�̳���Z�jb�C
�*�
��y��;�b��bE���B�+���c����ֶ9����v�"Z,�}C�������{��T���R�p��//�w��}��g��V)0�@��T�gc�K��U�+g
�rU���H��kGA�R��Q_��J��o�����KC����o���w�{_n����(�X�`,FK��`e>�KU��J�-5�]h-�������r��k$�k�8M�+�鐬�<�/t�F��XV�8�ȳ�/��IJ�Z�ޖ��}*�������!c9S ���Y������ɑ\(� 﫠 ������Ahk��\3o^PT�\���D�J�k~��-(�M�����~M�}��H8�9����j*�I)��mCJ�R.�d'���1�O|`�E���Dبv��. ��)E�����.��ʸ���{H�,��п��bF�F����v:����S'�	���*T�(\ll�q����J�B�\��g��Ӄ���9=�8�y�Xt^L/��n��t��&���k�M'x��Hlaʘ�m�٤n: �؉�!���1��lȊ~?2���ʨ��,��5�w�1`�j�#p���������M�T�Uz(a�%�V�*���\!To�%�l�d��B�w;��H�Y/x4�L<#���Xtb��>+P���9&��Xe��#ٷ��p�\ߘ��xA���G�]�"MR7W������R%�F�}��D�甕S����z.LN�%gr��L��x` j�λ�.�󬵷H^N�G,f[̹Q��p+U�R\��d�NW���>��dfǧI�~�
3e�"� ,ؾ#��=�o�<[�X��p��]��jP����
�x�j��o��8�C0ƿ�z)}͆�Q1)��Zp4�� �kZ��0KOi_��V����	��)Z#��tC��s��RY�a0���H�g.�M��w%�������U�}pe*aQ�A�{��rG���GO�
�Iںo�ַ%�HiУ�x^����,|pB�&&^���q�Iگp��'&s���*�0�7�ȷO^ʗ�<�H�k��	F�?��Sr�"g��������zyyd����=��"Ji��H.56k%����@Y�����sʵ�Y��/Hӣ ^��� C%�0�'�@Ц)�4����b6���8rjV[����F����s����eumSnݾ'�����k��}�5������j��P^ojS�V��.�G�]MR��߯_��Z�^)���J`�u��H۳�lVbhl%&J؂��R/�)���ݞ/HYAR��"/���⍌|���,Ȟ���t~~������������H�L�qmNI(�|�����&��g�BG�* (CfC�T�Ş��"�l��W6]4���
��Ґ�O~.
�!~¯xA�ճ��d��@�Л����A�E1Jt(B�5��&*�5���.���# �t�E��?�SIq�p�u��}x��pH6�����#Yf�*Ҩ�@�yp��at3�D82��+Cn���	�UT(l�$%艡�9d��� �r�F]3�����������D�k���+�^�}�3ь	S��"��c�#�G���l�_��!Pa��
 8�5P  � )r4��-H���7w7��Ͷ����驔��h�f�
�J��F�-� V�^F�M,+D��u���R#�Z�)�X_��G�D�����k�d�$�Z2@��*D֧wc�$�&ɒ���+�qUdH9��"0��&�sL��!��]�[��k��1-{�80��6���	��*-oOe-� #�-�'�H×*q�1�T�U1<�*ZZ"�0tad����.�o�s���.�҄��Z	z*%����W���y���$J���秚�N��Y��T�"swU*��4_жM���Ja
��:�J
��Y�z@ih�<$�5Q�-�T� ����W�|*�۲�~C��Ky��;F�W(�W����!��Ufǃi_��)��}�IN�M�w�X�?B�G��2(F�Ѯ" �͹nC m>����z����L�d�h-XL%&YN�����ӧ�)���*��}���;�w��߲EDizzح�C�z ��%�$�o��R��#]texv�k+�'lOz}��au�4��t<]�F�a�K�|6�4L�dP��x�qH��.�]�6u��Ŷw��kr��.Ƕ�����1���~.k�5�=�&��Vca��/е:TP�6Z}u���E��;��Fk����k�jb6|�'#�\a�:�����L5C�h����`,�[�겱uK�ךRW�u���WO_I;
�����_|��e*=�w��S�o+�s��8�����[=�zSܾ� -�D*���^�APO���ZEP�@��Z�8g�w!��(���@�?	=riv�ޑ2�k$<ҴP����Cy�'��f������!x��R���
Z��"���'�"�!!+���s鵠���×#�a0׍
�{(Z��=�I�>ؖ��H�`,�x$�O���wO�T7>�[s� _��W��ĬJ']�*c��@�����h ��<�!*8� ��q�'�#����M=Z�1n�yK��87O:�e��9�G:�#�"y�&G(�.�Vy�`��0諥*��M}�gN�T�I� �5���ʇ$����w�n^͊��I䛏g�$����9r%f0�t�4 �"��f/��^�gF(s��	q40�Bj��� |p�lBȞ}fH�������[V0�u�G�ru`�2��kϸ��D�T����M�8�UQ�z��, P�8&�d�M2�f�`F�Z���ƭ��W|���Gs�������o��C��&֊,��b�2����p�ͩ	ϻ,�\��'�<b�-������t\�n�G�9����C�8��4��� �������{r�ؒ�U���⚧��Tˬl�E�R�^�	���u��*X���!_���U�dY����qm�@~̻��?O��>�f#����`,[+�u/��Zzg2�_�b�����&��=��i_�PҽR�������t��Z�҉�l�n��y���sv���u0��<��2;�x!'�V��j�\��D�h��A1d��&�M�^��Ն��&z�b�5с�~k�%?��|���P����������1���"u���
�{��Vܿ�S�n��+y���M��{!��P�P9!�*�G_�����_CM�����>#�j�h�L�����^�{_R`7b�	�Lc��l�ܐ�[w�� �܏Vަ�l�sC���80V1v[�}@{,�{��F��jI咕��U�*��|����A�KQ��&dUT\��8-7	�n<���T��}��y�������o^ɿ|�'�>���(��6C �
6H8�>�������8����k��m&�_��Ri�Y],�y��aSQ�	6�!�I��!������a�2X��+�].@�޻�g�Dψ*㆞�"j?���K7^�_J�3� ��,����R9/�\������R�`6��DR��V�����2
!���@��5X-E��(����;����e��W{�9?��Ֆ��pph�O1z�>IM_�dB0��j��,�An���?d�y"�s�_��-���	��� �Q����P��*��³�j��r�+dc.(�b� ���m��@����L5�A�ej��G����wn�������O��4���z�w�s=@.40%���9H�̦��E)����`Z(&Q�F��Ȣ�Ӗ��k�*J,3��d܏+_�ￒk5∶,Fe�	7��`�C�'�I����+{/j���>����������dd�G�����O��ZY�)`5�-4qc��s������֕dCV��]��U��]�xV��f(o�9m?\Vex��s�Uk��L��J����p��fΘ:�rJ0d٦\�|"L��q�wL�0�@e��Z��(h�ר��7�4z���Lt�Zvv�ʨߣwX	~E�
�]�dPT��G�i:����ʉ9�W�,�GN�H � p|���as)�v�>���w䣏~%��u(ܗӑ2�>o��i@h�T5��O�\%���0��g����Sy	���ē�X� �?�����G��*d�aP��$b�'tf�՚���{r睇�_���Mvn�f�<�o�R�W擱.�=$o c�kP�=?:���]y�����~����Bj��L� .��P����uσ7�)�2���������;�`@[��+h�Ft�~��C���~+s�b9~q)�{�_>4QO*ɱM�aډ�<A=��偊1����^v�~	��PB�x�>��ڐT�^�������e��o�|�-%�E=z��+�����R[ݐ��l�}������@&����U��������\��h}nck�*�E�nݒ���l�:99����\ir���N߀"E�=G�9J�~��n��2G�Gq�U繮)NR)@,�k)��i������^?*�B򧾘Q�1��T ������� ��3�xFr^^3������1މ�wT 7�ըh�R�wrH)���Y�\����SZ�_K�7�E�B��rŦK��[n� ��0����Jj@�<�cf�lG��!�9��Fo������x�"(� AEF%U�T��:�<�"<�NN�7@�K�����UٽuS>��s����K���ުJ�;ge�jP�P�o�Y{X!2 �D
]�e����,72��F��ȼ���jmF�%�5qc��Rv/�W6�#� ��4o�����À쥮���R�߽52'�7NZ��\����$�qlk��o����T�s���s�����Ʒ�_@B��$��Q��&
��u^Gj��6[k�B�nN9ǭ�Pʦ�� ������%��bQ}�qw��o}�w�bQ����E��w!��&
r�77�ԥ�h�����7߲*��'�������鷜���~�ip� E�`81o#D�$=R-:�;RwLU�8�� >w�����@i[���/�2�DๅzP�k��8~�/N��p	�4�x$�C�;�R��h³.���|Ր��3V�0P�.%F��_�>O��z�L1Y�b�d��`H�#�B�oݖ��[��o�RA�G�&�Dj�>�(;#�#��� 8תy�F�ѩ�E��zS:��/��ٟ�C����h����"h�@$;
F��̌���P�u�=BG�8eWT8�9b���j�{�˻�<���|'o���z�� �����F`�Y�p n١Q�U �a��ж�g{�Т*:�%U�������f�����-.N�}�1�=����}���	��~�o6�������;�廧/�?����3у�Z\ۻ[
��g��KN�Et��y���r��=M��<�`����hVaBM�>�ur��k�;��d,�x# �q^7���"3܇�2�
�"�����}�����ĩ>@P5�ZxF�L��`eϱd¬�R!�9�ug�PQ����b��-^%O����^Ѝ��~Oi��4��d#n�o�6��B��Qu�+q8dv����,<�V@����9&�f�׊`щV�#�h�fK��sKA�e�\�D��Z�k���ZP�͍�,*6I��U��fl����?>f�%ԑnp���wv�|�	3����w���$>�7_|� �,��P�1#ŵ��gT��	NhS�g��8䬒(볏��旌��6x��z]'��e#�&`�e�N�����.(fO6y�&,���\�`���F��r/�d}�G C)���'�\/��\����[dU1�>f�Tf�M;%#L���Ϧ6�Mn�\Ue|������C��4h���� 9W�:.�m�'I0��tn}�J�29y����*@����~7z�I��&\.ezz)��b�a`��r}}��3��عqS����Z���[���Z�!�zE��8A�ǁ-�� �C<�X�����f�5�+y�<-����|�|TX+�Zkʽ�`j����8��H�+QHׇ�g�:^�I�oвAƵc]��:�D2�O ��W�
�<�O/�՝��wd��>�q�����U(�Ӊ��v�0I�l���*ʲ��&����ܻ/���z���wيX�٢�^p�i*1!��IS(-�#�?�i�P�y�l�<>|GN��B���\Fo^��q�>�8���1� ���<�=@n5W�/U8�=�d���Q��gԮ���Օہ��x��(
^*�<����1�D��{M)Ty����
��`aݷ�e�f��Zh��u$�����~�1L���������آM��A�Ug<�cT@Vz�ϸ��&�ol�O�_������`�٨�����s4�ѣG�_���pgg��0 i�q���woS�DxzlN� �2¥�4|��~_e�qt�z��
���[,�b����g���+�}ڛM��ɔYzHƊ��^L�!T2RzF��)3]�l�Ĭ�1$��ߒ"��8 4b=9�ߓ�ϞI�ޒ�f%;��R�Z;�q�|�#�`�#�S.��X9U
=.T�=ԚR��	-���#�l��g��+2,��,��(�J��U[�7��i�/�M�@s�~}�L��c0�$�k;%���l��Hu��wwn�_�������Y~�ɯdE3峳y���|�ſ����l45+��$K�΢��i��)8\���'��h:l7��b��s ��
�3I�S��+�q�+Y�@�㬘\���Ov��n���M�a��.n,ت��a�8���vcO�Q�� �2�ߞk%M�����Y}���(�gP���r�iPL\��4�Wua*���0b2_�/��Z���=�.���yQ�C�
4�,�{cd��ܶF8a���KF�N	���#oF��42� ����a����'�.�2w(�c�z ~�`^82C9d�k�7��@�����m�o��޾sG�����3��_�*3{�
�%�d �ԩ�wX��f<�P��r��b9iR�����)p ��>e�g��YDu���;�l�(f��������H�(�k$���b1e�C�"i��d���x4w�!��l�]�a2a��t�BVT�%pA�� �;7����R�6���T���t�0�@خ�n�5��)��*^P���sM��2ˀ� ��&,��];�K���%F�uͣ�[C���ϭ�p�O���� �uBzJ=C򣋞��
tqQq��-��gg��|.o0��������LW~�*�\SS�z��J4bȍ�l�v�\^!!�e��l���t}����랙��`7Kdb��z���;p} �$a�ܗ�R�5e6i�$7��ƍMYk7��R')J�7on�G���-�u[�{�=�����P��\A�b0e���f�9Ϧ� Ȋ\vN�z>�xQFe�3��������	�~��\*M���Ϝ�ʫR�O��	 <�p��أ��[�i��Co�V�wyj=_���*yN3��l�9�e�%N7�ˮ�:'�Qd=W��1������^k`hQ��꩐(��#G�
v�x>�e/#L&3��]ȣǏ��h��v ����'��'O��3�Ȍ��ߞk�� � �ϚMR�6���n��\�c�R����
������!,]�0\��#_O�4�M�o���nR\�ݻ��������������Jy�)��S��~!_���|"�`!�Հ�IT0ՕG�M��4�T��m��E �a��� ~�Wb�r���R���+kW|�u��^&so� �����%���K���;�|bKm������J�ϸ?x�H�x�D�oP�l���G���w	�@>�G^��Zۼlg?�ɮq~(h)<��p��<��-��ȑ@�'c�'� ��bB�NM�����-!d�B�{������w�ԕY<dV )V��8`3�&n�ʈ�����8��,+@�\�=
w��/_�8�g gE�d[����Ζ��7���Ǧ̄鳢�|@gSAp�$8�|flՁ�r���{0Z��`�>�7�?���i�
K�u�`�����d�f�N}G�&����t�&
�&��
���u��Z�debk����7_m�{�mg2~����� (�	�%��јн����T򕦜赞�/)U �.۸��I�� \��l�t�4NQ}�rS�kN����59�T�F�.%<g���V]f
6˺nQ.5AK̉ӓ�c	��1�-X}�
8�j�NA�`2@KI�>�q�'O}+�O�����lߔ���o���wɉ���ɣ�?��O�q#��?�W��e7 lwoJSA�t8���I�g��+��4�R��6��X���da���M�hc�@U���o��ܲ5ޭOv��ڔWgG�O��o��wO��]����|�4i+R*b_�]������O壏>�8�yN�C��уR��lP:�c��#)�ʬ�a�"������m,��Ta��&�c��.EYm���ű�J����B+���P^��K-��|�qJ"�r_�=�݄(�O�ygR+A�$�4ܨX`�9��&{�!��3f���A��[7����)��ʓ'O�����{w�Ro����
�p� �0�v�ׂq6�yWqxh 
sf��g�2d�Ю_7�Kp4��b]k��)�&� �D��(u��oI��V�������Of2Pp���1�[�j����ȧ�}&���mp~NR�G߰�Ki�J���B¶�8�4>h�W�C�h@�q<�AI�#W�W(Ǿ��Cꪢ�} �������}FTda_�Mp��B�Bi�up��]q"gfs�����Q2��p�7\ޗJ�DM
�7�8��z���6a���/Ae�%��J<N�K�7mm�u�`�\�:E�ڜ^-���uϓЪ������w��2F�#��{Y+nَs
��l���p��$��8}�	
�`�)�K�]�����G)1:5H��O��
���騄>�]rz�����������j6�B�	�/����{�o��� �+�݅���f�0�=v����R���:H��I���i���>?���	lCʲv���L�����$�~i��҃�W��[��&QE*�}��5����ޥ~��_�7�AE6��4'�HJ�c����zd/�sMM�`\�A(SX��'̺i�@?0��W��,-Û7V��(q��<Ez�D?�&>I^�"�o�MB�K��)��Y�}���ZEH�O/��$�~���F�5��W ],�K�s�uYY]U��r*���86���&h��A|��S`%=ȱ��z�N�,d�� e�A_��KM�Z�(UM2...8�I��4"0@b
��OY�^m�d�����1���췛��d~q��D�^l(��o01�f�3�C�3O��(���(+����ٱ���˻R�e�9�~�Tnn��� k��=���shE6x�FPi��u1!���9����>y�#��Ŭ�҅�'�ܡ��0�M���US|��^ٍpn�	b��;)� @{KA��g��Cy!�!�c����/�0e`
��a��l:���0�����$�B�,�;x�Q��e��?.+$��i4Z�^�����Y�c����MY�EwP #�?1]�l47ӣ��f���+�cxj`t�`7+��lf�81�T ���"�S�u��-]�t=�x�Md�I�8��<լ���<��F���2~�O�����͛72t�]�����֦f�S��1��ĵ���Rj.�t�m�e�""�/�&%�h�*I�:�����"���W����k�>�#��|�9�5���y%Φ �C�$�q�,q���=#r�׎�����TdQh@�5q�@|H��`���v����O�������H��g	x
s#�t�?�Z?6!�,ɝFh�l�@���+E�� m�D9�����7���82�iԸ�:eݥ`��	�9҉����<�Ѵ/�$l��A�+�(K��՞�w��VѠ�k�#p�X#xAk4�C%y ���=9FR*�$�`��JP�+b:E��H3Z�3͝a_A�`�vK�z����}xx��Љ�-�{{����W
(W\�?e�si�ng9I�6'd���!G⿏
E�#�=�G�Gr�7�w�V5Nݤ��{�C���BҵMN �4VM�fAJl�kp)�b�9?���S���j����t��J���Y�8$ZE��9��Ip+�G����
^&z���ܑ3T�0�yz$�X�K��n4�J�	Jl c�^jF�y��M�G�މ��"�UH���%M5����{�BV�WYQXS@Z��d��R��~�a?��v{���*X8���과ԘR���D$c}�Y�5ֵ �U_ �"�8
~��Q4���t��#��mU��0��=�tl���,+�\�3z�=��Kٹ{C��39�{)���}�}��{��F��f�E�#ri�)�Nl_��#���u�Mdcs����U0h�K�<|��ـJVe���U���W�
��U5WU�=o0�ji��o8�'��q�����]X|�8hFJ	�9��7j�	�bA�!�ud��`��k8��Z$�.bhIx���j-f��
l M~9��X����zH5�MHUn�0�-���g�g�6�)�
��z`a�6WV�P�2����Kv�gdU.�T(�l�������C��6@<�pc��i���K"'�������wԟҭ��ھ���[;��߁M��� ��&��B���c�H?c�`%�����ĉ�EVW0�Y�9[#� �6I0��`��a���z��G0��Z0�A�M}���/�	(�-<Q��!�C4(m���?�9�U�X2���I��Fo��9��?��[L�a��<>'�
&�B�Ǔ�^�����!U��i���u	�V�����"��r���2�m����C��B�mb�.�@F�L�ypD��6l�?@ڜ�b���Q��	\e��,Vcl�������
H������< ��t���Ú�ѩ,SmW�3�wo��ߥ�V��<r<�7��0md�Ȥ7�6�����.�u�.��F�=kѢ$?e�� :eMp�
\#3X��D��b� �@;����|��k��ޑ�;���r��]= �|&�v�C�'�������lB%*o�Q�� |��B^>�V���Tvo�G��D�����w���ַu���3��ldC �f��}��7G���6��.(�v��my����(ˡ�;�
�&T��2ە =�_8Q)�����dPAP�{����r��Fn�������������_��L���0�Q�7�K]�b��M�PA-�s����5�r^轿�쒏����EY��nٺ�^={�I4�����lm���!�<U��U$0�Ե;�5�����7�]P�+ب��l��Hk�%����{^N��IK�kO�A9\a�8�R"s��A}YA6$'����O�wn�W�Wy�͟t������Q��>�T��nK�U��ـ{������	U����,�J����CT���y[��&*އ�O_�rE�<T��g6�����B|J��E�B����������d���Y=sR�/Ʌ��_?*�H��?u�����Ӭ� ���걤�i0�{1�fcU]$���~rP����9�~���BߡP�z{]
0��"%�5K�CA�Xa�@�Y'"N�MBw�ɂ�j�4�J3 �ƹ��>L�h�/��e��4�P%�8r.+�d��\pN��jqSH�]�%�Td�����̲s�8YQRЖ�ĆG�{I�@�c}P�$��E��j���Z)'�q_��=�h��	���"W}��80��N��G�0�$q�
�-�_kIF���Bjݾ�It6������>�  �pS[s�h��"0�RµIk�dٿg�|NdX�Fp��_��`�-�Z1^�dj�:��ߓx�P�����xxv8�Pq��+��*^�xK@�i�-��lT/���9>(IxAU&�X7A�+g�Ez�����VkF�̴c��&2H��k�Ѭ���-{#���P�����P)���ήGS�XP���U����H�wXI��;���ஔ4{�n�u�)�����ZjW)p���8�V%���L�p��s*m�!���nO�E�\V�䷿/���_��_�J�i����ߐ>&gF#V]H6�"b�;+�4�n���\>G���
 N�����TN� ��{����Ł<���L�����y>�}�2@�E�{0���ϡҚʹ��@؅��`��������֭��<�<=��t:�� ܲ���Ә��l=/)apUj���\��ƾޓ���V[�G׍��WG
^R��!Mr��=z�����D|Ĥ�j��@�v���h:6:��嘭��K+m#�+���ޒ�+
p���oI5M�n�ܕw��u�9c���;���J;�����&hnb��nCFo!=��-�xJ�ZiB ���M�EzL�uZ�s�U�bA�<�=��y6I�Y��ޕ���:�QK
Z�UV�w�ޜ�I���>�̶-TP �oH���[(���-)�����K(�2���T� �a ��K��
�u�1ɿ.��VrW��8I#������_?*�υ�}*��a�e���GIm�&�f+�� 9����4H�p�#���k����$9
!M��\���f�%�IT��%���i���`�M���#˘�}��Cq��f��fUu�<\F�Cc�IN2��L��K�C��x&R�6>���nڄ��xo����Z��V���B),[�oi�@�����/>�P���
Յ���D�|��C�J�'Y^�$���-�Sv��ρIh���00���B>��k*e�/�]pN�f��J����kMA׾8�{�p�&&X��&�Kٸ)� 0��9V�-p�0IdR�Ȍ ^9��Iq��E$�I��J��t���r��a1[F�SF���ӄv�s�cKm�J��E�`	�,�*��,���[�e�c�M&e���z�Q�ȼiL��]����2��T�3�$M'�	����<�cK� !�+`&r΀<�������װb���>�'fRhmԹ��
�}w�ݕ��+�~!��	�AWA�y��5�^ia\��l���&ep�P�� ���1��p@2>����[�d�880�-4�;��>[G9�yX�p%�����ϔ�=(f�
�����(0�ɋ���T������>��qG��?�,U��L�����
�!���;�T�SnUR���/�aQ�{�շ/^.۬���U��=~���@�3���������zP��sq�`W�C�,�����#k�1�˒��DO�7׌�Q��c%�V"�^�5y�=�H���h�fk� ��@�iRW[i�z�33�l��rsk[�j�m{����� �^s��S�v"�(K}��7��YIC|�f�EP��몯�$ 	ƹ�X�( �����H4����Vrs�z�ۚ�U�/����s�ru��V*� �<m�Py��~������ۂρgFݰ\h*�
�QY��\�/2�H8�g�XxNHO�4�>L������ӟ�����tsu�b�L���L�m�g���#ѯ���pM�4pY)���8u�^�������T��2���=�ATH�4�?|��Z��4�}�H�\�����.��Z�J-�E��j�,ݯh��{����آ�
@J�>��G�7"n��u�`/~f|6TeR�1وuXe1N�e�`��6��$���D�,�ż����.h)z���A�J���|�s��^d�h#+�h�p\##h�o�~iT���Q��
:'ˊ�u�NVq��g34i�t9�J�\w �%SUK\�eʩ� [��B�\�����R���9�4�jF���A�vlFy�/�q&w�zĊ��&���T��VYE�]����� �
=���y�`~��A�?��T8��qZ��߫e���o'��t`�:���|�l����`v�r��lmŶV��m�kT!�Ј���\\�-��E�w�|�����xε�)�\�V��Xtc�
�n�H��y������H����p`���ڡ�:���/"�D���J� vF�J8��u�7VV�ݬk�ߑ��~�jت��t/�l�e1�S0h��*LPp[� @����mi����/?҃S��ɾ�{��X��������QD2gG>�{:Q�����5�I^�y=�sz�e�ƚ�������}W��Y���� ��N�T O�C���7�v�)�;�lq������kNA�)\����_��������5���M�M�^$ ��W�0�>x-�
��`��C�xj���~W��B��X��L��e�/=Lk�[��9������>�������)�M��39<;>�ϟ+XKk�-�x��(����4���]�Jv��K�P `��o�]C#4��7��H��d�+�R�g���Za
H�X<�YB�E;-^�0s
6��-�ښ�K[������kQ�Ilg^*HNͬwF���@��|�.��45�DKVq��w0n��:��O���/�%���3jX�ct�tJ�@1���S"�vS7yK�����XQ(6��L�,��h��v(:���bJ��MP�J!Ug�;�L���W`��
���<Wb���Uжn�J�ݖidY�iw������d��Y7s;�� [Jk��.�KX�H��j��d��	�!�^)1f���9�R�/�����/� ����$̵�q	|A�@����y�A /�̤�Aܧ:����q#7m�p�&(5���h��'�Xi��&�%�RV�
�,[Fת1Yo	�#�@�"B��9'R��B��ǲ�ńx���b�e����9�#� ���l:'eU&s��}��8. �O��^�$�}��C�G��V��p�!��4K��s Gn���J�W��,B���\�� �;�C�!���e[�ek�,�ȳ{�x�+�o �����U�I7��:Oz�s&a^��r���!8�E�yH�iշ�`�S ���hV�a���o|� h����ݤ �ΈcȂ���Ɔ��%>�6ױ�K��}�Pz��	��.�4�묈e� θi�6Ė�� Si��ߏ�ܞ�;;��O��c��d��TjTv�+p5źFP{�ӻ��ل�M#uA�yH��0�S��[ۺ>/e�P���X��D5��pg�n ^d�U<$ >��-����>w� ��0��ۄggN�6�����!�.�N��N��4&)�>u/�z1a���7�C쇲� b��Ͱ/G��.�@��wJum�
�UU�{{���]�P��X_9��%+6O�}��W�]�{wnʻ�o��l��X�z}�� 4<;�KM����Ar�פ3Dr�{��v���=�S4���F�w<7|����F
t�y@�@�Gp�b�/��9G0��I΅\ �\�VN1�l��"~/&6u�;��z�6��e�ky�w�(h��������P^AP ,U��HQ�@����h}(�(�ϫ��Bc��fTu�Q�۵�o��qcG��p���4�7''tL3%�@�M��l7�r�J����̹f6�G'һ����4��3HS&��1�~��~�)'"����bS���9��lz�T~�b%`�1V���	������F*����h��A|���r̖a^Y��Ֆ��-)h��1�7��C�2�F2,d�g�^�sfc}�R��xr��"W�1\'�k��*L���*�6�Hvjf�����#/);����F�Jq�_�`^l ��|�3x�Z�U�Ll�kF$��XC��HX݀�m��ߛ�|O��0u-����	'��R���ЫQ�bz���oE�mM�=�C��w�ā��=0���X[��H"vdU%�Kn\L��G��J����o*�8")��I�n�T��Wf+�g��W�����$6����8a��^A6�+&���T��(V������tPt;=��8�?��_6Q�7Q E_R�d(�OP=����[$W����3�G��N;2Ѹ?A��D=����;�L	;�qA�~KP�}ߙ�������+�}�/w��
h�(��Ñ����}����I�4_�� �eb㷩�?����^�p<у��C@Z.UI��d�����BL�ľg4~}�-��[}wؓ�ڊ�zS)b��p�|]�=Ƶ�F�Ǥ��yy�
�+��޳�S�l��椇�!6Ο_
hӂς�)�l�v���=�7z?��,�݈D�cڌh?}�����x��L����FB-�e�ߟ�+���/���kYqO�n�P��?�sT Q��9�{C�e�1��͑}~h���H�i��* ���V�&���_ƌص�}�.)�
�oL}��C�6��ˑ�up���@.xIp"�#3�d���c
��U�{S��"��P�v����sV��3x���8�މ+&<@��������&����A���4P4��ߗ�AO6o�Ԭ�%�Z�.�I0�´DĲ2�v�ω�$0��� ��
������LaI�f\��	�x�J��)`����wdm}��'�� (��"&@X&�L�n,H�ё�]�J,�3���qE��MG.���5�nvHg�RV��$����8�yA5FO bf���tN5 V��l��λ��"�"h�}d���ߓ@�� >�J6��g#ɮ-!��S��W��p�O�C�P�Z�gY���8�.�%17�,d�b���U�ȷ����<�P少.��`wvz��A�7�q�����pzj:[
)By��Y=�>L$�鬀��/�k'GW^~ب� ��}�����Eqǩш�
s��1cj���I��)����>��t�͋9t/�~~�tY��k����7;����Z��'�wi)4��3��PA] ��Wk�ƫu�d�^�����*��G�;{NX�߅ ����r����"
�QMä�@b�c��������?QmM��A�����j�;���$����b���X߭|n��p�,��]�R�B�;�yp�P�<����'��F�ጠՖ	@�^�z3ϔ��Ȧ�ʥ����x4`�O1��^�B���٩U�Ecȴo^F�&�\��5)����\�\����{5Yu��SOM��ݻ�Hk톆���/��`�k�C�h��PcӜ��اp�n`���F�[a��B 
�?�&@!���	Z��!+����<?<�������I�T+�{�*'�^�"�X:�
�0އ��-3��ʂI'<`4t�h�L�B��%��{�]X4x
��3�>{*��{�����=�
�I��\bqת�3V�P�j��x).�e�U^�-�z[��8џM�N�B(�����9+�*v�[�)ڍNSG���ޅ�Т�ߣ8��������a�3f*�f 9)����Y�����p����!��*X�{��3�n�*�u!y��t�B� �~�7P%t<���'H`��aUK�$���X��g��V[�����ܹ/u��S�g|J^/0)>z��Ț�w+��(6 rfp�/,�,�6΂�%�˃�by9sr��˟�Ȭ�9T?P��F7&:Ђ�����&��������=cS!)J��FS��&�Y�ߝs�9�q�����C�N�+H��I±���%�8��j�����O���(o� l��Bv�,�vh8P��s>E�k BU|�B�BJƓ��6��h ���� �$��[0Z��f�%�H�8D tq("��Mh�Y��AȊZC~�
� YSd��Ne �d���=xQ�9AX
X]����&KMz��9���1�ܥ��B�Q��(���Ń[����K;8V��g�f�$&F�M���V������<��{b�� IyL�D�|L�T#��
 �̶�TZp^d~��&��B��+Vi�)z:� ��US���&3��N��%k-U�J��:��m@.���U��P����A9�`�ZQ�x�c}�FQ�z(�H
���\�Tc��{���}$�X�h���$���VS�>7Ȝ7� ~�3���Xu���D���KM����u��kC7J��^oK�_�^<聛��$7d��\�N�yH��ԫ9:<���7r�ݔ8%�+X(�T��� ��X�Qe  �%��/�y�!.6�>U�<y6=X0Ơ�$���M윆>τC�l�#�N��X	NQZ6$~ ��S�n8Kco����x4�iȯ8Z�I@��gI�^h�̤�+���g�U��ѱ~)h��X���J�t>����NH�������m֞#�>/+�������]0y��&N�P�r+AC@|�k��{�ľL�L�wh���2[��p�V�aR�Q�?���k��</� �����t�Ci �h`�`ԟ@� ��BY��e�be}E��6�?��˗��;Nec���D�,�����&='�-؆X�@���'$�G�� 	��b����g�����Ku�����_�[�+�<d��h��+�L��	�L�g�6���'��˓3���.�غjr#y9��E�yaR7[��� )nf��`�R �ΰZ��P-ԏ�r�4�*�&�w�U�#Ͷ�GÎ�9a���rɪ	�ZE��d��������8��IҴo�)�0��4��c�A�%r7� ���93^x|/���-�2cG$ 4�A���4 a���^ hӅ8d���T���LVr8�<#�B!�hߐ��I΄UQZ���Xbr��#��1.�:d��lS�a�U�J�*~�F���MW��]�������/AUv ���<�<���c� f�Țg�@�SI �φJ���'� �� 8�L�fwЍ�����AT	Ŧ����^BL������"^ȼ�h�߳�Z(��A��c#�ET>gN&����ZU��J�0�S�����/$·B^E=�r5�Ы��.g�KI���:[D1\��/kR�C�hđf�:T���.f� P���&�*�%��i4k�G�<Lk�K$	cH �,2��edpp��pN�Y��H����L�|� �q�ٔ�ށ��ǃ��U)[46�zE[((�Y�8�]�(��^}y��w�+��@$�^��0�Un41у���)�'�9����$���ƊLr~�BVk9~UtA�z�T��s�� �HuA?W2�K�	��
6����w�lf㞄���µy4���'� �b�^A{kE�8r�[�z��d��n���js�d\T� �'N"%1xN�|�:XGP�և؀R5ܤ��F��,.���5� Y�\:O��ܲ�>TܔӘ�i�uM�XQ�KK�n^��p2��Q (�^�����z
�Zb�-�J�T�7`�Ǧ-�2u�$
��G]�%�X]�ΛC�V�,����mqz,���Y;uY���Eݗ/��L�MVg����g���z!,�N�}���y�P��7�8��"��D/x��I�e�D6o�KyuM���_�����;rs���!ބ�,�Lp8P��X��T�@��z��dtCNƘB��ՋW���K9�����!�w������^���YZ2Eb�,���T��9J�Nm�,&S�)-��fձ�.���X � 陲,�O�T]sNh��G�Q�	�gd��y�� e��ʂJz�h55
%��.���H��=a#Q��a����R7��@�h�+��V0S�xA�H�A�iO�O�,�����c|�R(�kY��8]`�ۘ�zh��H\��� ���	�f��q��gQ�Ѓ��_�+6���_�N�� T�5m@�&0�vNL�� ��k-9��x$f#�$B�G��ac���x0�����Y*�,O��3u{#�rR-�Vɣp�NlRAq���6�s$w*g�XL��I��M�nKb$�^��E���$��3f�)fa����v����EV%�#r��y�ck��7�(J�h뭮o�W�0-��p���X�|��sf�`$���̤�f��<���¨���jS�$*!%����=1݋s����1����ʤ��l����\d�$p"0V�b<���4�M.���	U��Z���	*tDUF��L��!׃���K�7���4¤�ޛ<rz$V�X�5�9����S�P.�b��y�Q�A/$@���)�Z2�^/Ӻ�v*��
�
�}T z]�f��
�Q��Ց~�f2�<�x���I��P.�N������00�@�ɹM����K\��K��C��w���/:�  eM��<t����&�s�|(ȃҲ��f2L�[��
.1��&�&i����L�
Zp����gJ&#�Q]>��7�G��V�h�{�q���G۫d�7q��Y�٦IC��m(/��=���xS�T
�nE+u/ �����^��E��>�&���R}�E�3��X>?�׏
���0M4�c�D��~M3��pS�AA&��aߎ|D�#@�%�E36��v��s��������ʝ�]Z����Q�F��1h}D�����`@P���B 8|�O��~oD/��ʃ�>��Ɩf�%YpY��#�� ��cJ���Ȫb- ��f��n
e�I:1�{9��Ń�5�;#�<,dI&d�E�LX횸Q #��+�MRrj�؜ ��R��B S/�?���=���3����;��^�@����]��y�,���tT���W
U�����_�qhpm�;��̽9#���]���*
zm��K������m��YJĜ��R���y��<1Gi<�SD9jFx�f�C{��"ԃR�3���89Er]`  N���7�+��1cC��{p�̿�,Y�^�#��DnS �3g��6"m�?��=Lx�+5��{�^@��yreܩ#gƌP���W��xeܕ����ۺɦ�2o����8�4�rd`�o}��R9�|�Lٚ��θ'QM[��*�j��1Ί�.�U�.a�^?�Y0�6(?7���L
�#@5�� ��.�|.���C����Ԅ�0��!7WB��4���	�ͱvQ�ׯQy(�<�G1�/3��Od����J�h �
�b��ͱ��ӓ#99:�YM�"��1��Gb2��^�K��<�K2,"�P�3פJ���-���鐄v_|*�4�DMh��\<L����Va���M�{p�AE���:�к������9����R�>�n�!��29;IHBP%S�w��	���L?���鹌��zz�ӡ&Lz�|$h3��݁�ņ�g'�i� ����pJ�ا���o�od�� ��V��j�&�¾�{�Z?zĸ@Z�6�̅M�3����͡�7�8�:���E,S�5�v5�����s��q8��\/�N�lX�8�F4�G�a�� �ނ	�Me�P�)C'"� ]�#�1��C����)T�=�������wv֕��w2�;�K�}MZJۛ�����{xq���'��р���g_i☦8l1����
�jY�n�A;����|	b�9νX==l�Om�H�I�P���C���ы7��u�J��F�.�P��^v�dr��#|@Npp�_���}i�Zr��C�s��ܾ'��f@	�&�;�b���lR#Ƃ�"ŵi�f��6L1ދ�;]0H
��Ź\&�f#�P���:�đ}9�#��o#�aB-�%�!GS�ݙ�����d����a[q*;�o��qB
%R D��0f6ɍ��
!Di$a�� /^ȇ�����b�^%W�Q,�:)W�ؿ�lK����Y��0����'Ep;8m�V�m2��s��*&h�d�A��
+�:^0��!��#�ՠ_(g�6��	����aJ�>+VXCٳ��#���@�r�	�$TxQ2��_�޳I�4�μ.BG��,�]-�Gb g�h����,���4�/�ٮq)�%��,0�֥+3�Rg�p��Ϲ�GV�����&�r�;E���8��s�)S�B��6�ӫ��*	�Y�Z��aZ�ZZ����u�53A{�7RT��L�E;�qf)�5��2�l�jK�mAT]�˫
9k=���V͡Yc���D�/D-���6�v�r8DG�]��t���.!0����W˹�E�gN'`g ���%�6>I�����g<:<T��������@};�ٳ�w�� R��r�AD��K�s~u6!(bV��~MH�r�,	�b�'vgo_��(�Ζ��|��R�0�~P�0,Y�~��EJ7|A,��&P�-}M����u3��r!NxL$K��V���ҁT-S�N%Q�a/,,�����>:������a�_<��ť�ɴ��X��MW�:9w�qpu�����ϙ�3;�d%�������́���k�R���*�U�m6��s��O~�����?�x �pY�<z��%:����O�����_�g�}n�뙤' 4 ܥ���g�&�D�?gOV�xй�1����- ���r*@;�¯�,SK�L����j���I�v�|�n��aђ�����I\2��pgEV"Oܲ�I��,�{��.�|�T�$�����j�s8B���#��o��k^|rd�>�k��3�ٔ�s[�.}Qc,� �\ڌ�U�t��f~��=D=P�b9�ӓ�����s�wWīK�?~f������_��}p��o�=y�k;s��
K�)e�,�|�}{����;���=x걜aWK��E-��z���<�}��:uUj�u�i�Hg"�T)!�]3��d����[O�d�'"~A��v2ɝ�2�(qVk-��ǈ�*i�>�n%����M���o��x߷�d�$\%0P�����s�H��V��1�w����%��~F+�������C��1�@�fqĳ .��Wz�M�:�ZқBd8ܳ����/���}V	����,�kD��m��}�y.�f��;��OU�
���oǇz|�	�C��*e���XJ��LU�n(��U*�v�驇�WEWBVUhI�R�o�nn�MR�E(���J���s�����D�鑱)�\�*�$'gji��N6�Id�K��-@"���t<��e���@�~����>@ӟϝ��=�M��ϋ�0�p���
U�=�a�)'�,a����������!��o���/���T�S"�:{ñD�p�����بI`����,�L�k4���^�Bθv�߱C��!t���p Ȓ��P��Q����q�gE�3s��v >e���<���A�%G�pn��M�++��?g��m�tE��S��$��S��{��t5�W��v�����Ϭ99�����P�t�ߧ7����>UVe��ҍ��Y��k�_��-�|1��"����H��d�A0�%��zb,ZE�(+�m�c����>z����G���=�R5cɼ�w����7v��
��Z�+ ����hG�J�m��]~�2�\��Uhf�Z-�(�eC���ݎ��]N�\�ovs�8e.Yg�Q��BX��
sJu"��c��sʍ��m�6��絞'=��5�l�Jj�y���,���;&��z����~��<�ȕ�oYWL�̾ᯯx��h����W�x�ڎ�������"{eW�?�ًM~�#|J1r�d	$]z�psu��~<ڳ�d�6��P4}��^�ж����M<��I��ՙ��:I�g��Nl����o�y�-���'B�c1��&]Z���K&�M�f���Z��$���M�_����eWS���C�z��&<�+���P�U�8O�֍:�h��k�/��m��RʳNp]��~���`4�Z#����z�@����ͩ/��T�f�Z�Ķ�D��<��A$<�̵XY�+�\��4��li�m	��%H�K�ԩ�0�2M�J&\�o]?�v�mN�ΗN�:��h@<
�4��}����s�JXyY�<u\D��,2�Dp�Ots؈�C�Iߋn�����K%2�OJ1E����E*7��T��"��A���
�$�j9Υ�AYM
6<:l�o�*c�WD�9� Њ0Xu�����R�r�b߂�4��AM
��KpNL.�ke� �,�v����g_g�$�@ީ�})�~���m�J�.��V~XD��A"L�c���R)�܆B	g/_Z����珿�������Y�73e�JO��B��U*�e/JX�d
6I�C%ED�5늎�B�b�V�*%��$@��ǚ���5GU\�3t���v���d��{ :���F-���]XYVE-�_�e�7{E~U�Q��3��\j�i��ŗ_ڗ���zw����B����@º�A�LD���vq~Y�ϸ�L��Զ\�F��@���gk��nN�m��H�?S�*����L1huvn?�����������}��K{}v��3�+��|t���#�̦A0�{"c�~ɬ����P�����2��Gj�ῷY���0! ��Iݫ�#*B��4���)����'iW�Q��b?ZGY�ll��+X��o�ʒ�x/�4d��<�Zi�R��q��<P�̦� v�v�p���·&/6��o��k^�+��.��~yd/�<�����*���@�oV$U�I<�J��H~��ۮGDp_h=���m �����=��>�]�Xd�g��56޿o�ɁJ|S��]��GE_5VҕK6N2p,�N������h[��B�>W������������Omstj�<v�7����F0k��[��RȾrAf�P� ��b#e��RX<�z#D�]v�H�I��=���k�R�z�"^j�˛+;::R	�t�g���]{$�K�zQ����Ǣo������v�d[����E�H�y8��,��V�:	х�^j��O�M;�DꕑYt�(��xP�b���%[ ��@B�͂�?z�su��-��z}+��
�IG��6lu���D�n7y���^q͉���Y�D�T3Q11��)Ŗ��j߈x��x���d�[A¶�&��W��Ri�Z����%+0��2���M�Z���͂��s}�ã5SǗZ�����D٪	�@��u=M*9�_�5[��4� :���2@��sh�= ӺPm�lH�@٦�\�No�<)x=�.� ����čPYe^�C���ѱ�e?@w�]�YLT1w��8p6j���X���D�D[;�S$m�R⋬%�dh�44Z�)yP>��;jq�9���C!����ł/���a�Sr0�Y�0$ M| �`�`&�Q�CϲCW��Y*JF�R{E��݄*7YYp,�'�����ݨ�a�uY�ˉ���]j�j�k܁| ^�/m��k|=��*��d��d��sI��1"X[�*��r�8U�������x�ܞ=}l��v�@��(�A�ns���؟�nֵa'J6�s)���2AY/xH�*����M9r٩d�@�D�� J�]���5߄4�)���# D��8�%ڞ1a��$M�LF�'�p+�oPw���*D��s(�Hȗ�@(��c)�uB�w5�@�P�{Ii�l�Z݌=�!��ʸO�o2i�k^��h���&�v~z|�	%�/j�,�nG��:4|�o|�Qo�����D���}BB�R�	)�4���CM�H�a}Q~����&[s��O	[x�� ,��:	�1�;::h�8{S
����P�m�� x�����V/�m��1 �7�:B��*Xi����	��,e*(�D�"�B�M&�M���*<�|����<��!�p<]�Ɖ��7o��"έ�� ���9�;� �%��n�ÐC��<>,�=E=�/�ۖ�D2΂Xܪ�ٗ���E�y�hQ>J�%H��
d �q���� ��H�����l;���lO%r�J�5&���.��m�F��dp���{*W�"x�Q���YN4)�C��s���ϕI�u8I�I%�D�֓�'�islՈ�������г�@��kN�T�2�/-_g;*�*z�H�*�5��U�E�3q^ �B��qAK��'>��^��.d ^ ���M�.J���Db}�l8=e_"8 �? ���V�}�} �*���c_��Z�x��W��`�?�v-�f�77�s	w�uf��М߂*:y^d�8��r*J̓�{�����T"����v`2Üҿ���;B�ܤ��iӵ�0��6�+������L�2	:�Ƀ�ԳL�|�y˜�dQR*�<(�Ot�nŻ�=I�?�ߺS�V�6A5�sR�$ځ./�s4]B�5e�
�2��X�d���?\�t�t�к߀����1��*[J��ѻ��O���������yy���ym�a����}�P�!�C��� �w3(�E�ޓ?{) c��Y���J����u<io�n�Qd�Ȅ��+[����Y.m�Xx�֔�IY-�^�u�� �M�CQ_��n/�+��V�d��C���8���G�U�����@�6�K������ZTͦ���n�R����x�ͥA����/��uj9��=|(B�Q�9�u�Aj��4+�����k����(2>��U�3���߱˛Kuot�cy��{�7KtZ�����j�da�놡��T�A���Qt�pI��H�5�a��m��͑�/���al�7л*�ח�����h��!#��gQr�^m=.�6g�"�#/�mI&Wv ��H���t���h;=�Nҝsxx( ������OE&�uqv��vw�c�Ȱ�a��f
<�ȷ?A�pŭ�`�w�Ϋ���md޾t�%�~VYMBu��{��1-}C���\�SV+�Z�&V�K�k����?�r�Ju�&��Lt5���s���*R�T���\7-��g��-e��&��g׳��d���^��/ܣ�E�.�|ڔs��4�S��i� a�X����K�3�Y8[���|��׳-�j՟C�������3K��[RӶ�G�K��,߂A��+t�)˶��_,��%gAx��?ʙ��c�o)q96�ZBs����m�?)�#z�� &`.�J"q���ts}� �B��=?�G�6V�
��@�6k�]xwj�.�ʨm��-�f-o-�	����a��K�4�U����P�����������A���\���J^y�kTe���!��g�)8pi�o�1����>�d :�2p�6U����ލ�Uwر�y�X���G���=[�:�_�_���"��yo/@�˂N��%�Eқ�V����5[um�P�{����|���>J�+�je����NϮ|������_�������Ў��<��>�O?�������N^K�pxdE1=�|�F�=H�yZ�#���c�r�4�=hi~�m�ՈW�Ȳ�=��yU��\K���
f!�8����#y��H{�dob��{��`���b�Cg&���d.���<X�M�슜eV���C��Z}�>_��f�;��oӋ�Y��8�(�ַ����>�g���}��z�ήZ
�M,�B4v�D�{�16�\"��7���k�$7�����Q�-�I�$��b�D���US� 8�ÂI�<�����l���׶�Q���^+����Uc�_o�/�,er�]K:l�I�m�]�
ґdzRǋ�,���OHdӅ��&{-�;]��j�vs"Ft3��*K�H��L ;���(٭7�6�1j�^&�����If��,NO�o�9mwK�eԾ��;fa��h���:�4fAY���T�jt�d���>*y�I�	�?Z��\�gpAa��M� �g�z�����,�6����PM��.�*�=��̈$� 1\��R�U��N7���`�Մ�l׹
��@e?�u�jHgF%�R�*#&�+�,�y)٣L@��i5a���(%��p�<Sy,�4�;>�����k�5����܆~��e,�(��E�+�\�u|�L�p㵳F]�g�3�/�~�tj|��鳾���%d��O�6<<��c��[~b�<r�� ^~�;�ڡh�TK��4�[�CVm�xf�a���{���O��!I[B��(C�E��6��!u�v�!D�E�ǯ�Cy���E���0��� ��:\�	�����F�")����ܿo�L�lu��=��/��z�F�Y�,��:��V�/̖��y��:�> p��_�G�Df.[ݏ�M�^�x�\^���{%�d������ڷ��-���������'O������������5V�PIs����P�z��yf0�)���C�n)k YF�pr)�^-�5�d��4_��m�+���֧,���&��p����c������U��"��m��P銬�&e�U9��N�`d��󉐎{H=�%��'z�%sV��rzc����x)�)�r>���l�7ŋ/��_���d���<z��*��X��%*�Gz�̄��	�۔(>� �N~(��f;��_d�v�G�������kĤ�pV٣	Ѱ+�0(���0�[�+��	�%8P�����b��R�D����`�1ѕ��B}#��2��T[������Jǿ��h#��{��c�v���@��ԣ����d���� �����P�J"��l��+�s�� �:.��e�e"��6�ɵ�]�V�΂Ъ#�������&������-��O:[�H^{���fK\�\M��k�:��#����@�"����
�	�D&B���!����d"�H�@��$�.DQbn&7�ė���,*�UaN�a�)�߄^.�B�}_8�s�l��]�8�Z�
�$��f�h]�lQ��3i�e&���+%��n�����g�/�4I�]�����J�s�R���6�!NP����ʯ�NǛ��)�*�D��SW��HH�;PY��#��-D^>�*��|�u�oA����jۖ���D+��&A 5�}N-HE�L��ү�,g���*���J�Q��h�&�Cq ��rSrG�%kK�m� �J�hNі��=���9��|�(�ocY%�W}�p������x�2�e�*e�+�RQ�6�{
�j���~3��[k�bu�OH�#RV���i��<��o��>���G��?��=x�����=�W��_�O~�g������ǿ���s	��r�u�7]�ga��tos��cc�6ʸ0� @��5�)+Juv����!��k���$%,2�(�΢��g����,:ɜ���S���\�����|��GpA�'��9`���u�@���M���1��i~Iu��N����m=*K�F�|���0�?��O>��:J��պ��E�phߤ0�"�"��<��nH����`���PK� ߗ�%����IH>�0ңh����͊���U�����F��k�`��0��//m~|b������J���{ �S������Dy7I:�.nu�nS��u4U*���q�5u����&��͇A)�.�" K�*������^<V�8��V�����^��婻����������R��@�h�hTJ+���Y�t�R�l;������n�,i���L�m���Bb�
�Y(�h��\TGvfskd	y��̖xL�ΫhK-�j{�7)K�K>'��S�������Cd��&8R�my'�γh8J��v��� /�"體EwKznR)�C�< J��J�}�Md���*ȯG���������"O��U���h-����nw�f�ߖOx�;k	��Ý���O�9:��q!��<�����2�x�)�ѾZ2�����w�jig�ͨUn��>_�sA�䇝�ʛ�J'�|�x6������v���Kx�6aQ��D��v-R�)�F=�-E�}�J�~�_z���Y�*H�Ԕ1/��M�-�2x�(&/�?z@u �<�sY�|تZY��MJ�֢�'`v�E ܡ\��I �<�xYeT�����Ū	1D��ؙ�F�\�H-Ex$�W������፴d ���oyy|�2�����������������������}����{�g�ݾ�IW��������R�|� ��ͩ�.�m���ܮ?ڌ��X�x�al
_�5ϐ����2#����S� v"���6�o���g�$�$�� ��(���8t��H��st�Ҟ>}l�Wv�� ��w��ҍ�s����h�,(�I]4�o�5 ��xE^��ԃ^�H lгwh����mvtloH����f�A?�.�ƈO��o\�D:~�ܻo���`u4���C�c�擅�Nj����8d���`8�a��*���H��� ����"6���N�_��\^��v���e�]���L��FK6BӰ�%��6�P�j�A���d��-�j\;C��P E-���Og��Mr����Ïl��сp��C�>������~;�_+��F���`�׷n��8�p���]E�dL�	G���ߤC+���J2N�R3�wD��ۈ�L���a���n*T��:j� �e"~��"���0S�FF|U��KZS�[q6Ɛdl?��h^�_4�fn8D�"�&�J��~��K��]:|�*q~��t��ݨ��4m�XܶJ���Dj;�P�6.�]0}^* @$�_�Z��fN��wR����z��Ro���H5v�e���Ͱ��W3�Ļ
v�(x�������|���5��fƃΎ:i� ���r#Q�پ%���2l��3 �`���j�>?;�ڃ�f�?Y�NOm�Y]��o�ْ��{�n����ܤrYx:	pG:*��)����~��_������`JN�\$Je� �G�,�hU���Bk���8Ȩu���ݞ���*ES�B�k�1P�P����(�2G)�s_s4�|l�����T	���5��\����|���,��3r��U���\�5,�ԡ��t���$��HV�����:��恍���7������ڃw߱���9>i�?V�����������أw޳��S�:P-�t�5Q����f:w 5�YI���4}cI�e>H3?6<xz ,�({� /� b?�j�K�Ж����hD
����7;;>����E9���Zk��E�	�$�@�y&�"?�Zv�L�ܽk�g/l�]{V.�` ����g
6�&2Җ8;l4�n�;��[�*�:�S4U�����C:Z�G�N���u᭕��%�(u���S�������>f�
o|#����ёM�������
�]�>3J��nwd�?l��@P����I)�:��N7��p�҂<�?(��+|*^����Ϭ7]��L�R�L@��ei�k�V�u�nPk��M�݀��:�\6@��<�`x�4�+�=����Vc$JK���NO^��A�o��Jgw�����zf!Wok�l�m��F:�n��H��M���:���[�"O��"�[��&��+d��V��$��;�\����7�w�hH�/�Qs�*2��)���I7�C�zul��p�nKr��"T��j�����YK�*�5�����%��@D��%�\-K���G�P{l�jFi'���R�xCQN�T��\��"�H7:4N��0�D�����γ��o�)y�M�g��%#K�ώqѶ��7�={	�LcÜ�Nv�l�A�,&�j�\w�E��j���z;��>���T�d���'�i#[�?<fK��\.��'�Bơp=",qF(A�]��=�պ����ŤyӤ�������aXm�	��8�|��h���ŹU���rfBH��Sph�q`�����n(��{�j(Ŭ<�v�8B�2$�1U��yV��J[�����\�|���ךH�M�� n��q�����~l�_���b:���ɅTZ��*�j%D�F	�z-+��#X�i?�W���
e�����O���>G��z�ѻJ޵���ѩ���:���E�aR:��Wgϟ?�/^Z߯�����OM��Pk��r��i"_QFP�P������twцM�?��c��u���s��{��3d*�e b���jK�;�a�:H�w����|��ެ;���׾�����مo�|�̮gS6'��L���Haȴ���:��/4f�aU��˼�V�;}���e�J_8�G�&�o6I���M�t���ڑ��(΋��!��_���f=�����oǿ،�d(��W/�ɉ��jɾ�>|���ٽc���>��e�Ǘ�IAi�HƇ� /*� <&�^C 8�B�A��g��#�w8�먏��h.�27u�W'+v�m)ŪTwO��v�t�ے��Ȁ�qaaj��W�X��1�j5Z�t�Q��Q%���R�(Q	��AG6��-�Zz���N�m�S�Y�G�.D��L�x-�!�Ruh����M��e���i�GP���f{���d:��$P�q[p�oRHyĸs(s�����.��2�7ȃ�(�f��N��X�!�qNZ;y*�uR�t��d��>�$R�����5w�[��� 0U�JhHy'�H�Aω.�Ե%�%�I��Iٝ2�k���J�Wm6��8�۬D�V�w*���	Ls���=R)���*ܲe�8���ɛ7a�A֒�z���Y��M��
�)"�³�a���c�_
��x״�`c��&��0 ��^Ev�o	�-O��'�W������&ʥ���̃�^��b+P��J���e󙝡��Fa>1��0���~�EihC�Mca	�s�U�=��Ϟ"|}�=-i=�\$ne�6�,�1�� YO��y �����se�������}��eWO_xPU�ҁ����a�B;H�7���:�t����U^�������2��*4�����UY�;��<�O��|kU�Z�裏d�rvraϞ>_�9�3ٳ���\bKe%�C�`���=@-Dd�g��z��F�;\9��[�  C� ;�\������q����7u@V��]��#C9F�eY*� 3Vv���+<��������\�A?����}P��z ��������Dt��\5R�w�>0�I(�w��kD���Mg0����oӫ��`+� ���	BOL�upN0��`YM���\d��[ddm�R����&4��-��{��w����_hc�'��˽�\|����ٷ��{������,��EEK2%�Z)�80��PD�z�a���8"��$E6\����BX%�C��-�×������+���'7iޮ/�¨]񬚥Mo�	m��M�	pCf�9U�|�n�n�<ږY��;5�o�� G��X�=�}s`e�H���3�*�$ 
�җ�{#br{�h�K]ayʾ�����b�j#�� �3�y��Ȯ=9�}�N���Z):C�2L7�G�BI��>��g��K���5�s�ἲT*����A��d�� �����a�%"cѓ�J[�['�F� ��vqm��?X��M�}�۲S�r�:x��H~��sl�h.*��2�}H�j�u����]Yt�A�n3@m��榶�hU�'e�á3F��U'�䳮�MTƠ���EdCP	���%�t �%���� �R<ҡ��ZN�}��D���ul�R���$ ɼ*4l�c������&�j�6p�RP�R.��%��DF��,����
`�/Z��mt��<Q�T�T�����$�L�8��/����+�^���]��3h7Ҭ"x�Ě�1s]DP�t���]
���m�B����������gW�V���>|d���߳��m���2!���鰾�*Y�P��A�7��̕-Z��7tm5��J>@��|8P��S4w(�����^���W�������S�Q��t!
���'�_��_j�x����l9����Z �e�ȸ��9WI	�r=������ǒVq�?�tޥ�y��p+���Y�\]y K�i��|��l����ff�<:� �}��υ�K;˟N/��諳7��]��L�����-N����Idl�$QP�Z���ݟ���ڮ���|�=�e%O��p�t��+�V���׽���{�k��:�t;s�hh`���4���c�>ƿ҂����w�ks�v�7v~~aW	�U)���~)U��X�z|1^�����Ɯ�ѡ3�Uu��4Ġ�L�S�B^���IWH�L��$�Մ�-��oK�k]4��]-M�&i#^{��R�2����y�Q$��\ ��*Ekl���C��M����;�¶����Z�8��B�:��or��i�7S[��q3]��?�?�M�?6�1f�r��X�4�#W6v�E*�ۮ#8'p[��rsdAp�$��&2He� ?�uZ�BjO���un��[��|Z��
���\MC:����e�t�8���M�h�
�~o� a�a���ǯD�p��Ij��6p�ιV�H�x����"|uq��d�\p��K	�1G�SS������(K޻��M���=���36�:�^�'"~Ƞ��W��ad�P��v~��d���&���4���� DD��J��'SD��M�H��P�%CD盲d�ב ���(�*K�Iur��L�`�������؃�6�x џ�d�#8�s�y����M^��2����߯f0P"�<)	�C[�/�0l=�Ͼ�|<����g7�Hq0��B�ݦ�R}���8,��	���V�PƐ��P|���Hs#��+զM�0�J<���A�G�-���̿�Tvz"�i���;!���׵��J�~@޳���C�p`����Q9�?�L��U��G���YJ���WA �<ҿ��vC��k���Vw����1���#[|��.Ϯ��b~_ݮ�(WRyۈ#X�<�\�������hӕ��zu�r{��Ǥ����+Tb��xm+v ę'}�C&���x+s�������������~j/��5ݽ��|�+G�������:L��7	�����^�sz��͌�?�?�=__~���.L�:pX9H��W�z����4��;*`�U4T ������Mw0�q0x#QQ�N���봩�s���\�8#6G���bv-�v������ӏm�駶��U�a'��3tf�ϱyx�&|���ྜྷ��9����c�9t�*x~3__+�Roz>*?�ݯB�rN�4�E�R)D$S�Za#�:C�)�=��ቁ�꺶���Յ-ߜYņ[!�|���'G6�Q$���I��/i/}�=���xt_�9 2�tD9&�G�Q�C�
�)�t�'�u���rx�LW;i�7����m�s��Ԗ�$�*E��-�B��3��j3�ǁ�{<������=�S_��=��3b�)c��!P/>.�2%���G*�8<J��:�=����� eh�i_�N;ߨ�*��&�P��$�]$�5�6�q+���%���C$N�pi��V
"���)����L)Ux���N�mB˺@a�T�A��1CP�W��P�-[kI}<K
�������9Z��&D�Z�	��h���d�ȠHn��5}c\�&�Z���I0e���eQi��l�X���L;�O��X3r%ݾ��!�ŜJ٤��E/T��u�U�3�+�{ɂ��}5y���At��^��[��h��Q������=?h��~���{�:�d+0�ݨ�g�`��p������z ѯW*71�5��*��hV��q�`N�5�$����0�ԉ�e�,+��$i�&�M��d�6u 8Z����P�t��	�=ܳ��c;�����F����!���= �P[ù�e��3� k�D�1�p|�?����_���u#�y����y6e�:�R�o�s ۄF�\�i.������N�R�ݽ{�NP ���+3qSE6
+���~ciTJ�ю���-��د�����7S�� �_%"���e�����۩����+?��"�~����?�3���e�^�����o��������W��;�P�DAw!�r"��Jh]�;�穀3���Y����3Ŝ"?9�k�䁍���l=�?;����q���@ߠ�{���o���ߟ⍄6�������L��`(4Gh`}$��
��	���wh�Ll}t���#0�Al�ѻ���=[;h�|����u�����;�`8.�Uu+��}}��K��6��f�jH��O}c�2��g�r
/xEZ(��橝���G��ǯUo��!��Ftw$��9���Pi��N��w#��OO/��g�X�7fql� �0�mh,�)��z��[��J�A HpL⚛T�u+�����oIO�&qU��4ʡ�6n����k��2 I�h��re��O��w>��p�J ��D��\�&%b(�{+E�l����Y.Ri۩���k*�Ef%�"C�%B�T^���|�D\� SXd�*z�%��j��R�*@�J
�1f ��:��r�΢��LI�f�D94��	XJ�~�
� �F���[����{Q�p���ŵ�<*F���o�8��}h����F��H衤I��D��cmx�Q3
�2+S?�ӹ0��s�	|+>d=� 1M�*���g���ۃB��w[���Zg�B�ܙ�s��)iR-H�� B�4<�Zk�lA �\\���<�C�T��b�ך����U!�ؕ�NdW���?���W)`Pw��&6���n��r��x��؈�Q�s��2DVq�� h��նѫ�T �T��(��/�Do��4ƀ��Ύ�����7�,����s)i��5e�� I�R�I2�n����dץ- �?��qu3�ק���U����"��,�.�Y[٠W*��OC%ׂ��@D��=z�}ͳ�}�w宍s��?������y� \b�<|f�q ����A&���AU�tpng�S������L�9�)IuB0t`?J���B��_��m����:�$�;_~��}����umc�on�~i��2r G-W��a��B`�;q�����6�s_��i��r�+j�ʭ�!�'�O('��X%�IS`���P�?�/����������������wD�%����ߔ6�ȷ{ﾝ����~�i�t ��~:�G����`̟�ot�r���G��Π_VU��:��g^_��;��E�!�%�_e/���Hu��`gj�6E�)2qJ־�_��)Z��(�r_�m��AD�>!�R%j�5�������:��[�]�;��<m�M�a�hc/�C��M�̕�1O5�*I�n���9��V��V+�f)�6�.E�Eg+J�]q�(���8pd�j�v���Vٙ�|}��G6�"�[���{X��}W|�����Y�6M.|���J��fI��yks�lZ��[A��wZ^�V�6e����b��@Nu�t���}2�`�1��6�C_m�!�޲��m3����3� P�H�S6)%��GZ��&�א��{��JVj���ͥwS�|��Yڈ���qd���R�� 9���{Df�{;:�r����������e���PZ�e�ʹ��{��ĊJi��Ñ�˶�ٔ媤>�'�z(���xM2x-��$����ꪕ����]�EB���q[���&ä������9�MgI��Dɽ(m�((�@ݻ���?ܳ���byc����q,r t�:=���Ț�C��c��p��M�E�VLQsm�si��� ��ʏd	(�G���u������(I����Y=�Z~@�Ѯ����ͥ�8��8z������������g_|� �ٞ���]��6�vc�y]8@C!�p�L�����������2|�m{�{���5v������������?X��g''���g��P~���n9<��� �C���k��WO=Z�}..S��b�9�~!�)d�8^\�?���"���n�Wص��5��_�_�Ç(�WѮ��h"�������8�W����dh=����m��g�H���v��e�G���g�kiɖ6�������A��i��L��P���9�Dע�A�P7�����T�@�yB�����U�~N80Z���f(� O P��C�/n�$s��::1c,���we�ߦWwST���H7� ��a{���*(Ρy�&��V��� �ೋG�t@ll@����P�f��(�4C��w�E0��t�ruzf�7������CJ�p�,�_6�8kaE�Yt�0��F�G:�d�-�J�"�E���"�m��-�y�]S߯���9�6����[*��܇���|zio>�����=�P��1�^�6��-����%0�l8m[p��f�ϫR�P��S�k��f�1�r�!��KǅH�J��l�[�7� H��YD��=@���\ϯ�t����Hi�`_懀�&e]�6U^|.��iF)+�	N	 ,�ӊY)Ze-S���DH�K���+ʕ�A^^^�t�k*s�	�e��8� '�c�8���08U'R���{@&|F$-W�h{��๏"`}���1��VS�M��(l=y�ິ�@ʤ��-<kZ�u��,38�:Du��.�5Eݭ �-�;��Z����V#����� �oD�F�u�(ܔA"P���u�f�Je�j���yr�~��L���{F����;y�����6����S3 K<�\du�G�fc�U)����(ҎS �����v����JToN���l���/�09��X�����~��ȣ�5-��]Λ<ƽwx׮�}J�d��o���ث�_�ˋsۡDY�J��ӛ�{��E�Ym'���~�U�G�X)q�u~x��u��]��^�����������ܯ������к���u�>�-�.�^�����&ֽ��e�������"�.Ke)�W��M��W� `v~n�OO#:qLy���ܛ�˗G۬1눘
 ����j0�9>:
�"D�|M �G��;و�>D�[��p�ІwZ�]C7�[��c2Q��_�ʁ��M���o��!i,T�O��:������H�Vbu+�S�M������}Hl��cY���;�i�Nm��́�@O�����;6�*|~���\y�2���՘6�@�MX7�6�}��K�)���ZO|rѥ��X��n��$(�e�����Cd�f�/�
�*t5h����5I"�	�B:uj$V�H���V^r��=����l�$)u9|��4��X
��:�����r�����")�Q����Y���Z^y�\j�b��ʡPV�ba׎����l�H��Y�G�8�~/_=����L��ʬ�ݠ�1x�2��8� ֶ_��t��D�r8D�� 8������p@�^�VQS���ƸJ3JC~L])�ӧ�7e$��0[z}��wR�*�K�kJ���|�͡AĔ'EN�=�F���SF�1m;�Z��4av��x,�� 1��t:$���f���8��߹�g��\k|�\��
�G�����l�$aD�^�z���l;�R2�I���"S���ȸ��¹�:���6K��)���3���'}kɖYُ�d��V�ʗ���hW]���m�w��℔<��~&�����@(4�|� ����jze���oٱ  ��IDATm������lcW~x��ؙ��t.}���e�7���;%�+_1���t���Xࠗ��0K�k����&�F\J�����C�89��M���� {����Y�@�w���;��W�4�Űw����O�EW����::y-������TR��|vcoN/����Ǻo���4���(��VZa>� پ�u%��Mte��=����<�aO�wP\<yb3��F;��T���W6��q��T*gq8I++}��>�s���L���J$`��ؐ�������{@E��x<�R�E��b��� �%g�3�؞�/� q�O��~�e�����}��}.@հ��)ڙ��c7���#i+�E��r��v�t�(��R9ے��f2��/���f5Q�r;�r)���F��� /�
��� ��H3��]�ˉ>t���{7��߁�ߪ�G��g�,��'�Z-#�B>��D�����	]���ݑ�z��j#XϦB��iq^�l����F:�����sхA�.Sk�,J���#�\zUj�#��܍��i�g9A$l���C��%��e[	�V?#dг�,�݂�<��A����tR�$c���P,�8�#R)��J�1�����իجٌӵ"�Ni�^'������h 0*Y���ܔ������1ҽm�Yj�d�S���C*�B��=�Q~[.j#@)c#V*��Cԃ�Q�4-<�����PQͷ ����\���q����e<�zW���NLu��
-�!:��{[�Ƹv��F%�5��x��Q&��d��]��ǚ��N�f�0��`��X1�	�22`R�|��0]x�\F&1@ ��D�/h�'ϖj;��Ab,*�Ѣl���v���v��9c��DJ�<qy��B!KVғAs�W�� E�p��XpJ�~�m����%ƦݠV�0_�m�c�aǤDS���j\A�����67��x��[w&���H�� �.ײ!��k�`-s�ȪtZ��k�@���x@�f��!�v�2ќLve���Wǯ�m����<xh�xd���^��LYJ+k@5{%E�j[��:�ѫvr�Җ~���>��u��Zrd !�j��;>=u߱�ݑ�d8��-}�n.�ʼ��9�j�T��9��vFV:p�vwD��i�ڥ�qo�����)��Á�33��s�Q��Ad���;rVv� ��z��#{���"���uA�a��kc0��g7��\���ȇ�`���&��~�=�����@��D]�h�Y���}��O�7޷���=�^jv�Ee�����2��| �J2~C�gO݉�\�(#Ě�C�X��2>��
Yv[r�,�'��|Ji�ʦt�wſ���g� :�N �HY�Nr_(>��:�DV�u,�*��� �q�W�Pt����V�eX�iQ�J�QVPKr)��C�y�b�2RxY�w�^8���[/�)Dd_�l��AF����a�7�ArhޑAY�VF"*!jy�Cմ��5�8$������c��5���!N)z��Z�D�Ry�	���v��W�-x�z�����[�6=JeDh����*[U���k�^!y�I�Ttq~���f�p�V�i�&Q��#"�3�ntGی�a�A2_k�����\�.�,��bk*5Y�'�Ԃ�V�8��&|}ZEӭA^���C!E���Y(���=�����O:;�`M22lR�D�F��Rv�R���?����c�Z!�V`��e�~>�yo�ն��
�m�s�~5�"�|�� ��!��&e�r"��.O��y��g!�F �5����.�P� #,Z��8��.����@V)����i�s���']��wm�b1-�D�2����[��M0ܑ�Gx�mC��(�n��7�)�|og��H=[F	��;���~VH�ws�c��sܮ����|1�2�w��%�Vg�F|�v�1d�ѥwv~mw��S��LG[LϷ�~�ǯ��B�\��N:~�f�P�]�I�� �6��0�Ϧ�d���@y���}\'�{v����F.��eCܓ}��5��7�k�8��k8��ݱ]?���"���=I������1����W� B�SD�sLn�}�YtW�p�W�D�#y`�x0�r#�����c�?����>w3�s��ڷ~��>�P��/?��vv|l�]�=˖˫{���:������t(2K�~�;4D������� D�{k�y:���]�0�]G�
MHܜ���f(��"�9s0[��s��<d���Iw6])H"@��8XO���j&5wJN�����$�	Yn��%�\�:��m�,���e�y���J�P-�pf,��7���/��+ڟ[���'�@�,ώ��y��Pҁ�e����D���9�k�������M��:|%��W���B(X� ��6VD���P9u���Ԃ�A��[o��D'f}7ef�櫠��҃G:����	��:~�f�Ta�؊���lV+E� �˳s��+	�e�Z��y���2�����
<�E��Ѫ��24��},���ʣD4��.��i��=x¥�T���US6a�GـțMq�r�m�	���d'GK(���!���f���C�>U6��ߔ�;�9�:\x$�^f�j,y}$r�d]��/�_�2�7Y�m'��fN��-ѹ�~�Eb���^�,�~��f��U�1�{#o���,7���mT�i`�@���|z�	@K�lu3�d!ӭ�r�n��{��ݺU&.#��iۻ�(
`@�����%E�ZA���87鐬=��yD=��d�h�-�ky*?�׀���QTQ����B���l��/�"4]�.�:X�"q�z�wx��Z��`�2�(25w�%�?�5���]~J�C&`ó��V5�yŮ1��	UY�~�Q�Uy�E�+���cdD�I�X��j�	T�SxKTg�\_M���Fi��/l��ᕽz��A�e�.�^x�1P� }uQ�p��z4����(�m2���FhC�:8�3��w|�t8tR���T{}-Pf����:����3��q���>fI�O�o�j^9����ڟ�{?���?�k���?����Ս=���G���w���&}|� �D�H��.��>�?��?��O�P��Y��L�m��Ⱥ�w�yQ��O�����\�[��5���������@��d3�g�M��A:���N���x}jgg:S���< ����=NðAڃ�zI9?+�.ā!�T�<IJ��������z{���7�ų'��w�/��&���ql����
�ī�[�e�>�;M�ē�F^��X�t��(���q!q�$�/uT���<)�͹TwK&uW&y�U-ؔ��0TI<N�zZ-��uh�#2	��=��:ٖL2�-@N��f[i��F��ޖNxe��Wk4]1�*]���[i��*R�DC��fK���ޜ��P$��g�xtFg���]-N"9�1���zyd{���!��+Eʤ��y-�9� �ZR1S<�f�`t��g��,�~�Aiu�pr���M��!i y����$oY�<�V�7�G�`"��f=�8Z���g�JTd������0�9L*�zƛj�Ւ�[K�e(�r����g�T�]�32�֙��vyz�¯{�H���<� e*G�OV��NЖ[^R뵥�jE֪��g�E��c��.e#�����XHLܖ��Y��ȼ-���,IdQz�ĳ�C�듗>.��u�u����.�n8e\�\��UJ�D�5��	��
 |#�TT�~�N�>�s�q��Z���Qʻ[�\O�ɰt)2:Y�7o��0ڝþ�kԳG���{�2��@@}���<X:�+��zZ{��>�>|�6��4���{�����=b������h�ϸO		%�R��0�T��x�PI�5��r�7��0_�$��p�u��������J�>6x�&��^�|-����x�2BA������
P���|�K�y@w��?cF	0��|9��s�tr|��;H�ݩuR"�y�'��"�3��eutl㇯D�����[�ؕ�O?��.�o���d"@GC���W��3�ׯ���˧���^��?�e��<{����}�� ���ut���d��G�v��xt�S�yW�x��n�i�1d�2����M�3N%iec"/_������Ͽ��=>��c�{���ɟ��~�u;e~Ma ��?~�2*��W��̹;*g�@�J{��	n0N\����;l|�nB����Z��jݫ�/U�_�	iV$��,�\���d&io�%�%D9��	ȉp[��P�ah�K�G��L�a�}�$�_V��.�FY8�F��}t��Q��fO,U���	��'�D��Ԋ��������QU�W�sq;j����f;�Ĭ6۔=��c�lv<�$�p�ќ�|1���E�oB����Z��@yw�ƈ���a�ф�]d����;JM�%���,�%JXE�TtZmV������%u}�uw�u{�mfj�8'mYA&~څ*�q/d X�Y�9�z�
�� ���In�q�]����:��/K�><E���ÓA�����D$� �H%$2XHA6݃��l��f4���saܫd"H�Y�n^�ǧ�F_% RԛJύ���d��m፵z�d��@� kɸ �<X�݂8e$F��X�ͺȌ��	Lb#Y�#��!��Q*Q2��w���P��pgbo.���s����p"^τ. �k�d��7�hh��s&�4�dH�[�C
��y*ˮð��,��.�x����n�apz����v|�s]�ȣ�
!�*2�c�U?J�7�W�\�{�?�du�So^�VY���K{��g�K����o���_�_������Z�D�mKz�2��它�MݓK?�/u N 
�Kt�(}u�(�B���
#ر�ÎJ��|Sza���O����;�D�\|C|�䱽>z�@oe��ۄV��@�;S�RI�d� j�_uU���\��fog�6���3�M=��
��K����|>�����T6S��g��}����l~��^x�4��{w���]����u�u���wVE���4G�N�m�����ޜ��g���������g���9_�n�G����ڄҙ�'�5jx�$k��\ ̬�����D�6k8V���}=M�W��ё}��6��a]���p��ݷ?���= �Y��#���n���Ϯ�� K]XtYH��A�a{){ثD���e��:���^_�;Pd��i��<iY���I���pX%�'�-�Gn�2��K�H3��o=��m�N*Cp�U�ӤT��$�4��M.y�U��*n!=ɺC�#����uT6
���<~پ�r�o���b�P�J)��Q���|7�][ �a8�d���LT�B�a�9�"�J�~�s,2�ﾣE<��ao�@D��
���44ю�h�+r�E�4����,�'tt����������}�D�}�e:)��I]X����dH)s���f7�l�|�֋�S��Lc���E�v��o��%�W��J�W�!��JC� p�8` VN�z{m|��邢�2��[�X�s͡u����;�5�s|C��īr�o{�@!��b�:q���5q���v��1JI]f;JMYi���U��ؖg��+ٗ�U>d	�n��~��H��	-W�.m|��sN�Z�8����vx��������м�A���A���Z�F%�eJD��m�p�7�Ǌ��Ȕe�Y�s_�S�\G�:��i�߻�@�+Ͼxj��&ΦzV�R��]��1'����Ͼ:m��I�-D�������O�ڞ=��>�������G�<��^�D{a�G���mv�>�U����"~"��̮N3�E��zXC��׶�;��N��o�tm�s�������.��5m=��+�zqc�����)��G�o���+S��a������m�QF'kmy�U�J*��u�p����������S���*�;�D��ڟ{��Y���*�Ɓ���x"��=yb����k���>��}��''v��^��1�"��NY�+_|��!��$���y<�Я"+Id2�8$K��C���\h�åT�eB��ψ�Z�qreS��ןD��[��u��|�'1�zf_>~b�}�X�3�}��E���g>Ñ�)�C�����j�Ⱥ��?�����V�e5�V�ޗ�5l�z���U�	�!לh�{D?����W��J����ہ(�T1��Bm�!<W�7S�K�fC�Û/Hi�*	��I�kR MŨ8撔=9�Uj�,my'��R/u�4-�|�6��V�3r��m���A0��̑�`Y�Y+�VD?p���јUM��#�+�q��B��Ot	�����҉�`��蹞��ᡟ]�v~��`�	����,L��ؤ�@+�����ΰ9=[<���ƳHNڼb�xD�����,	�%XӖk���������>\Jz3!~��
ϥrE�:7D�N���0�����vUuR;�D�|S�EVFo�� 6s���3l�Nm��)�m�d10����ۡ����.���F
Or(�6ȶK�#7��|����E�u��[�i���+�H3�K�[��[�҂���c�^�^�8YYh��r�G	2���ǹ�/ ���v����*7^x�����|��X��,�G���K��/��8�K(8��1��s<�n���sqE ���{X�D7�&j;>�Ci:j2��g׳ٕ6㍝���_�G��n�ә�<7��冗ή�9���g�~lϟ<����9>� k$�&��ׯ^��ɱ=�����������_�Z@��w��?�Ⱥ'#C�ˎL����w����ϐ�G�i&�Zi��ٓ�V}�.$����lxM,=[@����;;���H^E�����ț�EԐ������T�)s��/�f��d;tZ]k%����5�v�LcT����������ni>�'o^���sk>���{�\��֪�����E�[	־������qp"1�'p�:��=���;�{��7�V�ϋ�{34����U����<�+������l�7������{�_�|�*�ɗ/�g�wzN�pc�PF���u4­Q#�J����P���S���'���{|h�� '��}]�w@V\�dD�r����l��j�@�����>�$f�C�o\y�����ѯ�����^f��r k�m�m���ؖ/l�Dfd��":$����2�՝Ѧg{��ֲ ���aYF۵��CCv�'���O��_
@S8��S(����JS�V��u! B���w���e#h��U8u��r�gi__�{i�����R�	P�V�K������u4FM���{�%^ t20>l �������$�������'�~���6�{h�i=�ϐo2Á@@|���h:� 0��%U�2 G��_K:��qkx��^��ROK��ZuW�z)ވ�I����I��gJ�"O�����Q�):���ͺ͘�IݹYU�D��;�ö�W�/,*�-J�R�e~0�my0u�,A��a2��F&'��s�p=�kiQñȹ���zYZW%ѹ%� �8���1|F���`�l�4g6Ɇ��A�ı�2�>�<�p,�IK�NQA�M��m˸�D�h����ť����=�����ٻ��Y�|ziO�>Uv,26];}s.-���Ɓ�Ji�5Ɖ�A�f����4���vU+?��bԳɞ�FG;��AGO��SJ�~8�;C���\�$"Gy���uq�F����v�<�m�����>�>x!n��\������=���v'{2�<�۱��yTT{>�6}�خ�/�P?�UfRG�?��?�>-�ʆ�^4�q޻c�+{��Ku��#͟���1~MK��a��a�m �D^�Lx=z�������O~�c���׳���۝����o� ��?穽�u}��ʥ*	�� ����p��,��\�*	WDǝ�%2K��A�{�>�{������چ�w��^�^ϝ6be7�P�F��bv),%,��&~YdK����#?�ڞ?�AohGO^��ٵ:�^<�����9!ɋZD��/M��
j��,-�l?���x׾��8P��O?��={~d�χ˩]�zz����ud/�{i��9rvy�2/6d_�r����s��w��r5��W�|b'��l�k����g�<|����-y_Ce5�T��F,�j|O_�����U6/��-m�sǆ��u�V���ă㣕G$G$9]�j)�v���W���7d;���.�a3O�dxI];�:~:�C�D�\!��0�pe��+:'�A�riḐ�YR���=�ي=�-`�J'J�Es�w���Z�jĤL]5��X�Vg#y�(��ڂ-鼼��1�	�&��Vb��JdM����т�Rj�,�އxXq �φ�	D���Qw��羙�%qvye�����wD�#)//����6�$2�G�zx?2/��G��m+2�Q�jK�m[��.07d>Em�Y�?S+��T뻇-����Iĭ��a�GM�Z����l�[�Q#�Y�I���[�/MH��q�7	��c�4�Nm���ͫ�kj���c�����:��TB{V�G�7�M�Sd��0���2�� �'�^)Pg��c��Z�[�bY�~�a���R˷*@Yz����,ֲ�:[{8��Ý��u�����z���K$M�RCqbD�����3yH�<H^�`$�[?0)G�lI�d��8H$�dO���Pw8��y�C����[-+@b�@7�C]Uw���������Z���g�x϶�Rq�!1���?B�`'(bSҝ ��r]�;w^�o�"����P8��-�(�,��z+��$�Ft3��m�ٌ�0�o��c��s-+ E�%�)��֬������m�L�4����j�^g;�r���r»@��O����	��6��l��k/ߖo��F�Xb����Ƶ�u0
��d����"  �W,���jn�
�W��@�L/m��%k+u�wN�=�IC��
����.�)��������4�������!����벧����/��٩t��*�|�+�x�Ϋ��]�A�R���M��j}�$�"��0 �nQ��
y~�X�_�N�Hñ/���bT����5�� ^Q0?���{N�Tpdn=��(ڱ��VPf�w4U xΑs�?�0}�'~Znܸ)} vw��wx���H�<>��w1vV�N�
��Xp�.9�	J5�πD�͝i?=���ߒb5�?}����o�ŷ�+}$�zMʰ��5�x�����u� �J��勳��k;��=�����
�Nu�?�����`�X� 8�כ-�,F�MQ���9lH0���J�V> m� U��谱��B���>V�%]�n+���R�nz��=C�Z���#�TWMdN7$�W�]S���x*X4���夿;Qt;�ე�|��zġZYa�.��JM��ֿ���9q�tvA�e��)#�V���b�"�%�]1�Kn<H��\{�M�$�XF��j\G̤#�c��;��J�,����CP�Ɔ2E�Z���Ǌ�	uN��c0��>	��=Z�-y��0�Ad�@��z-�͍�Ӳ �0%��Z	�:�_�9Ҟ��xD$��%�\��M9q��ç@(�>I 8��L����PSdNS�!�ڊ.�q9>��i�Q��O)|���1��T���FS�`[B�K9�cղ|��ҍ��΅R	W����*�*Jަ�ܽXq�Ǭt]��F ������Id����B
_`/�n	�q@����8�畫�Q����9]Lٖx03#S�s旉k��Xs��9�䅵$)^�_�ZɴZ�x<�P��b./zr]A���u��λ����#���3Zv��?�urF�;� �c"f�c��f�	?� ��Av�H���k�����>#y��
7L1a3ь�tGހ�!�Z]_�GNc�%�����xH	۱*��٪������īwd��s�~O��w%- �X3xx��Ӏ:�)�,��k���H�*��1%���܏8=ƪ��Mc�.��[r�����\�WW���*�Ofp����V׹�
�X��d/Ďx���8����}��H��c`��"<~��N>x$�\|]��\	�ڈ���Ecue9���3�pj\jCA �#z^P���)þ�(�*/�1
���e�Qo�y~��'�De.v�wkk�@���|v����
�Z
�j�[r}�&���޾�}����]L���.\؁4_о�}Ӡ�� �*1.h�>chyq�ST��~W����WA,oʲ�w��M<�h���"2�@ t}�� x �������&7n���{�Sb)4�
}e���D��h�+�ހ���<�Ц�>��qS�H��U�Ǒx�+?��F+�lͳB?����R����v�����ʔz.�hƼ���|UNQ
)��QyIW�3��$�}���P�t�� ��T]$"�4ڹ�e��'�Mi�R+2� @�s���4A(�l���'���-p�VA��i�0�8�s�/N��O��	=s�#3�^��t7��l�����#��'.�)�=��Q_i�H�08݂p�LcmsK��<x �]#��;ݖ�k��tٖ9=����T7�cy�7�[{�9�O�Y(#�Dz��F��`!��bΉp~�i��=+
�abl��80 &�FzF� (&�R��ۘ38��p�I��D'_��I�g�2���wV}�J?�J�+�X?�1U�,���Q�(~B����Ī�{�  �Ҳb��F�6�`�.����X�۶���C�	p�Y[f}�r�&�<���O�2��&����"T�<)�6M��Y&�*c�R�K�Z=�d�$OO#Sgf���z�B��̥�����w�6�d<&=�����Y	5��g��i[޽/��]9<���E��\��7��X��6跥T���@���>C�RŽ���)`�?��pY[J����u)5�h@���lf�<�tJ����#�f����g��>׻r[��Y�T]k��Z��l�n����~kmU^i`ʤ.��[��c���>)�Ͻ*�epٗ۷_R�����=j����B�ݡ\�ܦ9 �!�BiIbƃ��a����ʵuy��my���\lj�^5���D���k�B�ܝ�]A׍��R)�ɉ��������E�Qu����GJ����ܔ�K�p�[2/��g2�5�V�H�)Z-4���YSp�d%��8������	�^�
8Yz�+��I)d�}��e4Ѯ����z�%Y�ޑ�_zIv������� s���6& ���S*����BXoT������+����K/�(������k��O�.'�~CR�w�EO�ό�r�4_ �-����q��-���������X0�~IueM����n���xb/�}k�>�p"�#��jz�ˡ��W�k2���{[��q����l�g~��֝�����"��L&]]�C)�uHg
��+r��P��p������SW*u��z�3��KŇ���
���NV;s]P��TL�*�N@�>�ME��
\���Y ���.��mэ|�Ȅ����'����}�k��G��a��)�p�[L��r��Dgi6[ �R����N8q4ׇ���Փ��q� k�������;?�q(k�qU7	�>�o��_Gs�l5[r��F��^2�M�X�X��ʕ����!#]7lF�N����x��C�8ۻ��ꫯ����|(�N<�M����39:ڑ���q���=8*j���[��$Xp�c6Im͜]�����dBf~�Y��S7�	��T��Y��Ϝ&�鈴ld�ܗsދ<�	�s7���V	��9�%F8���y�\K&s#��,|Gvu�v����xK�*�z���Y��/���F�QFK󊎫(Q'5~���k��$�<5S7�"D&TH��G���qV��^�rL�h	�x��b�)�,���z����s��e�y�I���T���]s�;���t���˷��rpx)�y��1�R�%���[�u][�z��7U�rv|L�1�S� D4*���-�8A�8���,�q���B5�^�(x(���}	�e�����o�D��%Ȗz���6dcsW�n�$��H_�:+mh!�%L2A��,���z
��O%ƴް�U`�Ǩ �@����<�;}��t�p,eM�J��iG���u[@�"�Z�"��+��� $�Y8u��j�������r��<x���A#����e8�i�7����ۼ;���7��ߖϾ��������~�wem�&_|�sr��r[���w�B�u��7��$5
��.�Wd�ĩNbsG+���#xn�"��= �`d!z=��d��5y�'?+�_{M�K��~Z��)n"@6t]�A����)�z}�~0���{_���;��?���s]Z��o�������'�GP�I�\�%�r%��$�7p/�t@eUx]Sh��:I}>b52M��9�zCkQ�y ����u���c��H��������	���0�V��ں�R�9j��u^�{q��t�
&�B��m�u�$��U��!q��*��%��0@b?⯏x��Z!���gn����52��ZF����fI���~�Y ������b%~2�BY*� ��43���m_3��:�	���O�z�f�פ�S�|����_�r6��_�SrmcC�O�}v)z��C�y����w3k��6id�#��p2v���9p�v�p"y�抣@Y���!�6�R���#^��������Z��oj��	 �`<d��'��ѣG��^���7��_�H�rvtO&��ts�|���\"L�+��Q	܃"���dY�Z(!4f|Gv�&��<cz�����<4c5w�D���/jk���kه�b�e�ܿg�3N��:��#Վ�n���"lN�p�P��D\Kp���fT��q�CW��ظ['钺��+�ep�P�0q�v6�{j�
�T��&�(vVGP��3����6�M���4AM&Kb:�$ �yL�u�*�o��؋-�r��n���J�nZCA�l�R��L��c.����5��m�����^RS��H���,o�z���ݵ�x]����
��.��U�����C(�K�D�~�]��q�h A��6��j0[���_�N�� uϞ��κ��7������M9}�H��4+��A *9b ����j�I����@e���#V"��@~����?�I���oɁ^'�Q�~z�T�����w�#�
ZU�Do�����������#_��_��v���JS6�JxT0��!�u_`��s�M5���o�X�8_.��5 SQp�������Ip�
LW́�{��9�`(�i�Z�b��n�)bS;&��15�x���������c���#�u�|��-�����������\wh/z �b��5|��������';������h�X���� qw[�粈H�^���g���mgSAMK.��2��[Ja�>�`E����k[���S�����1�7*��fem*�O��n2��nߕ��k�B�j��;�ԩ}�ݟ����Mg��J�^/��مW���\�����7,���\���=l$����D�̌��w@ƅ��v�RC)�f:�M?Y`�^!J���f��^��b%��r`� ��{�?9!��I08kb�K�)Me⥌�)�Z��/��r1�=Qf���+�䐻&�NS�e�.'x�L���2h���3^�ag�����L=~�Xj���^s���t3ǟ0oCp���t��n����}S����d��I��2}�ݑ����z�8���L�͗Մةr��\��6b���mR�"q����@��� .���וr��1lvy�bɿ�8�?�����.�~�jZ��̉�΄�M*��{uтK����!�n>_ Z��6��H@��`c/��r���G�=~d�K�>���@��*^��8��=<g�� ��ԗ3�i9��M�a��ըP�� �65�lK����_H��R�
G*��k��q��֐�L8.ᏂT`�.&���Z�sM$4`6̃^`m7�yߪ\�bȠB�I�o|�:��Q���vw���ή><������vN��Lf��R�D�(����M��_�O~�����zK�JCꍚ�9^���̸KpV���=���Mޣ�鍇
�DN�2�)� ���T�~S�۫��|F^��䳋���~M^Q��o���>���J`����s�Zߠ���c��wߐ��~[��3��ׯ˶��O$  @��B����1>��6��:]�ך뺿�?OcV�ӹ.�2�����CL�A�01>�jkM^i5d�����T~�w~G=|(�������q=�p�E�K.�&P�OO�UDJ���{  �~F�����4�5�<��W���g����*5��u�P�}QJ��jl��C9���U�YZ�K�{3yԹ��&���9�^��벵���]Q��sNPbz>�����Ę�B�����ܹsG��m�����Q��;ߗ7��r}oW���w�=��RY��$ ]!*QU��(1�q)!?//id�}����,Ĩ�n�l�3P�6'���$ ���\�d'���+�� �`T�E����YB��E�e��[x�?����Z��h^hf>��^��=��Ά�f��ʵjك8�"*�2\$���և���Q�*vj4f� �Q�y%_nnV8~vT:˧o�_��ھ\�ۆN�O �)�J��R��ٔY����gA���-�K{�����[a׶v	TV�*�>|�@��Q�ċ
M]�ĥ�����@-�AU���@JÈc��fćw;ⴕ������i��)/�(�tO� �d����?�2k/�*y���9�'n�+��y��Wx���n�ӳP���~�r˰���ځ�Teƹa=Ǚ�yNW�d�BP�Q��	�Y���S��m�)q�.v�g-Nf9��,�X�尰�l�Z�\!�l��Z��8~�����e�Ƴfa�g���=Y���nb=�s���d����L�a#FF��Ԫ7��s D�h���o~O�^��H�{0�Ľ�Cu:@��5��6�O&��
+��E��t�t��'�Om�n�A�c�3>~r$��P���륬��H ,�?@!�h mA���r��}�W�U�X��Y��ɮ�S@
�-����b��bE+�d�}ÇhCk��6j|�{x�.�d��XE��z�~<�{�-��y>zr �+묌B�dk{Oϣ*���\�{p�yʩ���sN�@�;o�I^�]��'�_����j�RcʐZ+B��XA���$_A�W5��M�caЪ�}4�Jcc�*ih����k���P�� @�t��k��79�x|z������REk*��۲����i*?x�}���]���/�qV\�ޕh7������7�zU'C�~��VSMH������'�L�)�o��s'D	��1�0m@�oVX9	;�q���\�=@՜�`"�q_?c�A��8�Y�@X���z.��[_��d���:����+��|G�����8}�pM+R(7tM�T�E�H��Rs^o�����:�����|�^�	OuC]�Y���h�b�µJ�9yA��1|"��F`��1�f�E��r�BJA��l���Z�V����x{}{���;[�_�Z;��Y���|ܛ��Z�{��������v/�{�Y�٪��Uꋠ�=�E�R�=Kd�QIҹ�ѩK��".��9*�����/x����s�t�,G�*3���NT{�7�32�)�4z�u����3n<�م<y�X?ڗ��5}�j�qWZG��������ފ�Ƶ���&<��H�h���d�CL�P��*"�`C[8����3:Yz��
$a'$��m�r�/X=�2>�i@����k"�g��ƹt�N�+"��Wj���_���쉫H85Z��������vˊϳ��.۞�	�j�KT�L�gf,�s:ȷ�B��?|/H�����9���@�Us�]+�xE�PD�M�������uZ���ֆ��.��l$�~��^t�J�i���Af�&v����]XKA����LN���*��U��Nn뺬WKr��}�k��i��{
ѴɈ�
�.�E4���JM� �9~>F�t��h}*�Χ��O�2����pK5�߻w_��o���i�����ym�yaŜ�����
�}o������]}n���<��OO�|[F���{� D�ڤs�B��OM��M�E�`ʦ�h� j׳�k�]Cik��t/)� ^���e�9VX<?�OeE�T ��Z�ӳ���{LA}�[ߑ��{���<::8�8��� qgu]�z��ĔS�
�0 킯�Z���Vmr��%Y��B0*��l�b��@�A6�L����y(�u����݇˺��JU��7�s�]}zܖ��K�Cr����Vv8b٢ɷu�'��ݕhБ�^�u݃tו8 b�Mj&����WW�4��gc]�'<,���O<�R2��Z�ei��[��c���m���xvQ�	#����A�����=I�3Z0���B�z]pl���t! ���6�j�����]P�H
��%9_w$�<m��z�� ��ј�&L�az������n\(E�"k��h�x�́b�>օ7��.��,-U�������ӟ���?�����gvN>��_�E���w|���G��������ճ���H�psks=*Wk@��i}�,�����uc�={��=���u�⑍�a"e.�/b���c'�*��JH������~QZ��!��q�G�R*��z�0BC�����Mf�}�0���P��+�~~K�o�Ț~�?��>��Ύ�^����Jl:}��u���(����ss��|a-(x�x��bR/�������]8k�����j�b@�:^/=kߤn
)s���A�$��q���;�ɖ��i7����g�R���r��̩|�OȽ�	Y�* �e%�7�q���4��m�)o�Q�'v�B�./�D�,�&��+�.��ULpFpW��:D��w���!G,4^V�/R��w|�̬4|���v�ޏ�E�X8�ñFc�%��.C��4Cn_�sܺuS�|�Y�����sd����w�h0@b�鲌��]�:��Yp�9X6[	���пek�$�JS�AO�K��P�����x��|._��%�{{����dmk��k�4�\)�� `x��X��ƛ�����IS3�����L���]H�A��E�z�Hu/{��4<������^@���Hz�3#��0
����}�T.�mY( [[A+h�IH[^|�e)�r}����v9����`$?x�*���e��K���m�s���@�chޠ�W-V�U_��4��4ݧI�L�UA�[�?�U]��JՀ�^�@�{m~*�=_�=>?os�ju�>F����,�Aw�a��S�׵V�q�=��˨^wmQK� f�L��2��� �6R�7�����Z�d-G��D��u9ro��֍~��K�;��`&Y*�?�H�E�9OX8�"���;��  ���6jY��h�p��P�O�2Y�@��X��@�O��g]�'^M��&���д�Nd��t�n�
�^>Z�_����O��X�܄9d������b<��KGi�)�È�pL�+�&� (�ܺ��o|�K��;?�K����_��y^��v$����p���������ƃo����h�����K�b�giLC����9m���>hY0��Y�ˣe�wɥ[�^p��co���B u�4YN�䕄B)��W�q6f���/AJ�2�BT�v![+���E��>D4���z�~q�4�-��Mʞa����X����5[2���uyٜZO���,	�_Jp`��p|��]�L�"�𽬚��Ń�>##�� ���e (�V���*�����r��� ��sx����D�ý�.�2�Y��JY�Q��x�4+��R��� ���a�0�J85>�- a��'�2��#�$����jJ�P�e{�8�C,�������f0BD=��31��~�U�Rע�g���dK!`N���Q���-�2ɣ��T`I&�d�p�d�!W+y퓟���������2ǐ��@8R :��&���x���S�,3mL�� S�%'�gˊ��^P�U@	c�>���]��BaummE>~�*!tE�z-�ʚ��2F���29>9�Ǐ��Um����	~B�	/T���=�7�y�h�3^D�lUh9�Xۚ��}V��aY�37�<�܋���+��/_��?����\���3�����ߦ��=�>��%������oX;	EH�C�P �եTm�b�l���Ʈ�
I�z�h?�J��3$����M�V	�J�B+����y�UWW(9q6�#}��8;��z�զ�*��J��E�fXXk�<�y4�X�q:ҟnO
�7��J��Ǧ�o'��� h����k�$c�60�]�`���e��NxW��;�CSo%^P�H��A��!y
�����P�Qj��M��6�������Yo�L�N 4����==���YT�S����ہA�ׁ�������1�G�-F����nZ�"N/�vIjN��wU�ΝZ���q��)���d��Ť��~�������ſ��_����y�����>�˿<��{���������~����{���/���ʦ�g���`0r��JL��,.���Z� .3�Ǽ��g����5��Fs),���M,l}!%ޏ�ԍ���W�A&�7�V/��"�%��Q��ghEzu
��!�D���4K�X�j-2/�����0}P�K�h��8r�p�S(vf�t�ld@�V̂��8ȿ�A��@���J�����/^1���p�x��k��&	���ԁ�a��>�:'
^^��U~�3#�f`��S`v|%�jt;|fc�'b"7�Ό2����8��g�?%����tZJuXq"z<��]
�1R�d��@xų�1_!o�,0�`}
�e�� 8A!2��g���_�£���煮�J_A�e�/��LN���u/��W_[���ɝW�ȫ�xM����(�3؁H9�w�&A��ܯ�9�Q*��f�ܫܞ��AR�a�� �N�w�^(�<|$�R�k��䘎��;�����C�T2� ��R���=C[������{ѕ�u8�w./%���< ���cR ���]i�ZRS�U��HiW1�k<I��|k�y�����EGZAn?��>Ov���yF� �'
��������/�"P___���S#u���K�H]o*x��ڙCM�������S�$*רs"��_t�(C�(�Z5��F�-�ص���
����w ?�r���m�|�������<x�DVa���6�Xx�U?-�%IM�;*V�ư"��� *�zܗ����w���k��н:�p��R0w{ [��P��%& 3�&6��t�
�؎1�J(yt�X2+�b
 �! ��C&��轈i֚2UP���5^,U�����_M^�Ւ4"=/]/o���$�ܔ��-��i�XQ͂R���Z����`�@[�W��w�D��J��G���/�����/O�8���4D�a5vɵ_���R[��N��i��5��d0��~��O���/������֯=�������K��������_��8�w��`�[��f`�f#��ĖM�wR�}O��Fj�%�q[���č���e�6MbA9���g�z���
����d �G�R�ɗ>9x Q���6�G$sz���J�{)�fs�&�N3k3�xғ�����c��1��+�왷N^N�w��?M(�n�b�FԘ#�cKL��fy��G�w�ט&f��I�jW�g@$�z�`Y���rc� N��U%��YK`�?���,��}��c���(�\��$?�}�ЦIl��CU��'ȹ�9q;�:9�oCf���VCq3��e�)5�2�<��"�����av�N�(P��<6�P��UP����Z�j/4@`�	º�[��`I�P�ՀX��v"�g�
Z.5+o�+
V�+p��g>-/�|��*���aCNŌz�Q���O%�V
�s
'�pG�4H��Osʔ7��� U-�m�6}W� .I�����Z���7�y�����k@[�>N�� �TM�KS3h?�Ct�q��J��LY;�@Z���3ᶌ�	�'�Y�%r� �:Iu�ãZ n'Q=��BQ�GO�X��$�ֻoqr�_���F��ݐ�"$% 2P��gcZ�R��E��$ղ�us^C��/RK2b�Æ�"���.�d6��F�V�L�Q��JR2�`h�����+�I��"_��7���yC����_C7�R�����>�@�-R�1�F'P�]L�?�@b�������,�&�{�T}�P��$ vg�5JbW�L]�Tݠ�k6OM]WO\pTp.hs�F
���=�^o@�c�
��E�E	�.�z�Ge��C����	8=���#T�'���R�S|x֖3]��΅T4Y@{����RUk3rjݹ�H9��چ*�E��F=�_��y�Y�c� ���>/��;�ݐx�C&���s�_�> �d�8����������7��_=���Ա����v>����������_��^�p}sc�z����|)��~'�m\��}�<8�x9'���u���<�g��3�!+F�'�(3#y�Z`���*:�Q�%�Ӈ���Y׌->�D��K��B��O�	l��ZQ��n$��)��ͱy ЕYB�a�*%n�8?h���IlQ��9���m�To�gtY0<+m?��r��j�?��a��x��[?s@��^hc.1�[.�敔�Ut�|�)��ߍ,3�G�Y�D����pI�s�`��H5+�����1�����3����-���*��R#������{���3�]g�����9�9u���x~��i�_��Ʀ�f���x��({f;��&�l�llmi@X�����;wdsg[���2P��>�1�Y5ľ��&��N�?���9��b����˜��м�X
n�|��\C/i �5˞b"e��B3�J�*[�&�����48��x���1�uX��^R���3��X�ވ�?����8#�&���9y���L)D611��#w��_��Q�T�U.�J���Ӂ���K��P�E��A`��ݣ�޵�{��@m2��h�����4�.TG�'>н)���?��@F���/5�Y�EB]�m	��P�mL�r1dU��Y1�R4����	���e0�1�V��VZ��'_��Ύ����Z�SOG'O�}zQݭ��w�k��Ȍ�.)����S����� ���˪͢^{�W�IQ��E_:c��T���'�Ĉ��|\[�i�բ���d8���jgh��8�x�� Tc�ݠ�T��K����Mh��PA�x��I���"�!��}ep�� =�{���̱_+ �=(�[���\�5\g3�z����x	�������;�R�����D7�(T����T�Ă�jք�	2�4�2ݼ'[�ko�y����G��{�?�cs���K?���o2�7��Q��ܔ���
"ƒ�f��,�U�2{ڳ�X�ɒ��=3�Lʃ�m<"6�vS��H�U%�6*-��~���s��y��4Y8_��us�F$��*LM�l|(M_^�)ڔvb��t��.��*[�T��Oxq�!��{�C�`�m 1�4�
����3���0�Ř�����m�Y7��x!3+ƶx�q>��Н?����̲��S�dT��Z*���c֗gF�3�2�i0>3ψ%]��$f��9 �7���#�՟�����\�Y��-W�o��qDf7u�1�\Iȳ)&�-���O� �-���Z�?��@ڨ�fs�{�h��AF�6)8G�����{!J(=�U��^�}��u}���S?��t�)���5�C}��P�4�{�A�q=rcKk
9ϔuc�U��������*�^sN���<P3Up[�q��uZZ�U�4��F�APg ���uL��v�7�Y��X��T��d��g4�� ���b��P
<��`���v
%aA t��� 0�o���v��`�P	�C���s^�Z1~�vT�|�$T���x$gg�|N�=+��O��-�m+C�O��rQF����kŪ\߽.M��'�H�vPd�"�^[z�s��Nj�_��Z<�:4���d�**�����n�S?����W(��r~r�=��l�g>�Ii5�������o�!���Sp7�נ����R����l����ܐ���S/ܑ�w���=y�k"��z���tҚDiE�wNx�3 ��m�	�-@Dƌ�;��L�3N���������z.PEn(�:��	�\,�Y&*yz������5��K)����ql]�5Mڂ�JE�J�';�e,��L���� JFE�xC�J �D��P��PtA�kX��b�C�Ə��c^�I���〨���,��V��
�(��+|j�	`��,��ꫯ��Ͼz�W}��]�����[����� �|8��1���
�G�ZyF4�+�F��e��C!ld6Ib�}榀�.�/���z�af �">Y^ G��kF���'O��D3�/`��F�l�j�@�S-h�>�c�3B"�o��]m6x�S�;�!�z����s�N�~ς5��_S��zNc�{��y�,#�����U5�v�\�Qr��ʕ#7��c����%��]g75����������,T�`�HXG[���t��!W�*���k�q!d滔� �k&?G{�ȜUb\�Ź3����6"	�b�ȸ0��̞A
tW�5O\^ߌ$�l��8#վ0LX�Aۑ]>Tۂ�ԛ�E���%�l
��4��������[�k,FU�@s����!��8��th`�����������@1 �)[�APw*�Ƞ1L� �J����ES/2X	���M��g
L4�-��}G���(��L��=���U���3�s ���vɇ�y ��NN�T[���(�����ZE�
J*�<���3k�W�;�@�ݶ��D��8S?������N��{Aٜ~OxB�P1�פ���u��j \k�'kͦd��L�2S�V+������x�ƃ�X�oi�#��}[�Υ��=NԤ�Y�9�k8K-������i_ʨ,��h��L�'͖�D�u��D�)��az��S5�\FC���zC�?�Y�����ں��~ֻ�Gѹ��[�~>�q�&�QMVo^���u�����-���#�w���
t�i4cE���XNB�+��mU<G
��|�a;�Zk�2չ�ˣ��X	[ս�>��Oesg_J�
�� @��~b}�f�����X`2���5�� >+XH�9�sV邢x,H�P���4�������&�����e�>��KSQ �})YE?v����Ƴ�?�b�`2d]a�sE���9�a�f&�S3������R��+���ʯ������Ǹ�������w��g�����ѡw~q�4��is`E��Žrb�M��>K�������1I�S�K�!�BG��?@F:BeƇ�\�emuCZ
Lc��2���M��h9U�E���W3��JM:����kN�x^g�� �ͦ
V�-P�(P#���p#���UM�0�ɒz*�6;��H�b�����NFd���6���UJpa�ty��[�ڌs���Sκ�$�	I��2@���9^K$��3N[uLL2�#���9��x2�'�e@��?*�x��\����+�M��1"���g'&2
����~��N��ؚa��pLs�'��ZH�f���Q$*������-sǛ��kN�7�'�3��CX+,V�����r���\3���B��hJ;Fq1]��I�вZm�8��0ʢ�z.UR�-�%�!&D�Je�3��(�����ƈ	,%�5�B�3Vg *�1�VSj�����|F�$ �x 0�翵�A.�71��c���`�4�B��@m�@�q��HY�Ki<���z��-ݿfg'�\�k�/K�\#Y�P��J���7�ʬ�������>�a��׻�w]N�;�6֘�p��R�(\��麬�Q7�fP�)�YY���ܞlի�ӐTq1���x������{��W���4p+ I/�Jܻ��R �r����mm������@���spDjz����)��8z"U��F���I�
Bf
 "(�����J�'k{{S>��g�9=�/ܔ*<}�s)�Z�^[�p�<���1+'�(d;ȴ�2&S]��
�R4�(S�Ҍ�s�+S>Op��"*k���>��j��^��µ.�/	�(_Ͽ�=X�\A�()u]� ��0��gA�y����T�^oIa4�� �y��������E]� ������lI*����K�g�3�?���xI5�� =��%�����hl�jD>��`V��X�������.�2E���<+��W�������{��{���Q��ʗ �A�����]�eޖ��NqS�$�k�kAX�%o1��4�a ɮ*�eM(DKK'c�r���y�����U"�8�1����A�D5^���	��l"�>��F����r�i<ai|�R7#F��! �&�Go�r�W@�}X���E��G�ync�d�Y`#� ��Q���E�3F��l�lI����)d�bU�l#�yVD�w���!~�l����u05��
`���=+-���rp �(�^Pqb�N_}�.˞�`z��rY~ɬ��ߧ��{2�.cSj���$o*/Xo�����)�>5�	�9�=�K|�/9%��Ў�[j�5�	��2�zt�.�&�㨢 a4��Br��U�M&y Sz�5d�-��ӡ\>������F��J�eNą2ԥ70��oղ(0�TNlzϞ�����SFA�u��F�&���
:P���٩�w�i�i yr`O�Ǥq'�\��{�^��FS�j-ߕRC�1}�bd���V���Am6�l�M�bJ�}!�Ǉ�`[���c5L�5����29=��f�u���'�r ��Є����ն�����*+*mPԝ��o����y��\B5"*U�F�ޞ�V���?9��q�9�*�%x�0�vj�R.ߓ�fE��>���\��ezq����UXh��;VXi)��Qq����1r=��&@��yG�|B�28 8ONd]��5��'�$ӂ�3н ��於��m��)p����{��$�d���Kb���%
���������J�x@����`a�A�uO>�+]��4���R�W9i�\�x)�N[棈c�Pt�����$�l�J?@q��m&U]�M=�|��1[C�������!]��8#�� ��^R�RC��S�E%�-���.c���c^�����s6���59�)�g��d�9t�!��Oi��Y�F=��k�XL+�J�d
���]���nj��4�b������bGF2G��Gh9Wd��=9���Jʪ�2�w��,<WT�ԍ�qd Bd���pȅ	,���°2�
���Ǉ�D�����^ 	���bȱh�ONϥ��J����[a<gV\��K� ��L��5�5�л�	��j���%V
4H��ʔ8���S.���=��t�#�.+/��ꅈ|!�g�;�V��fh�U����+�U�#4�s~N�k�9�Xd)0G ��A�.�c>ed����|����s��qze�ȎS�u�9<H�U�L#�4�k��<�YC[�zoL��B��Z�X+��rX�tQŊU�*y�2��P7����I��n��Q�|�r� S�
�	��u�э����'6%�vkse��u��hs��m1����m�H7n�\^����[o���V�4�k��x���s]Ѣ3��'��H�\�r�L��M�Ig��F�y=P	)/Dͦ#�e1îB�D�����x���1f;O8�]�ҵ��3ӿ����]O.@\���������7j"qv&���4�{���{���� �=�ދ�o�'�tG�\�ݰ0M�D�,
@0��c�g�Oezy!0�h�d�6WB�@��	F����4$J�p4�{ӄ�0�HRİchV���#w ��ciUr�^��Gr��������J
��.��$g6��t"+�V�:��Gn�~V�~�=/fE���ߖ�&6u�5 ��:���� � VY�kZa��z}*z�0�=@)i�9Oe�����I	���Vץ}�X��(b�������u?-VLs������N�
�zl�����#&m�٧�BL��[�)HAN1�{s���*����ʶ�b{�=��X4Bw��=*_?/�W�5\Di�TW��,��1�
j��%u%(nB�A=��2����&��/?�W/
��< "�)2A/U@ձ,���]A��T�|TWL��O]��f�p���Y�~�gs��c�@]DY }H��䮙K�B�⌛tBx��g"�%x�uӋ�	]�i�2� ��~Hx��f�<�~��'ǲZ/����y2��8e9�X��(��@7K��#GB����$6	Ϸ1wji���5�0I��$I�V���&�|Z�:�Aj[�Mr�%�x���]rZ
!��µ�����s�y�8p��eEǁ�@�L'Ʌ	�*� ��0~�xr���q�ظ4��?��s�.�����ϨF�hQ��dD9q�>�)a�V�ؙB�z.��E7�eS�=Y����\���F=�T��PvG�ߟ�ܝsҨ�2������2�� �p�v8V���ߔ�5	������sSQ5cn�4%�@�
]�/�GRjV!��A/ŏ�@�Ƚ_�?��~��"G���B��pq.?{{����f��:����̾��s�x��T5`Lg#�\P�ǵ�z�T��+LcC�H=���2���
>�u�`O���ZLu?C+
DL=�>ך��N4��� �L�m�X��c�����{2�+xr@��Seb�X{����pzpD�3�m�g|Hm}�X�X��;YR
$IFU��{W*�zKl뾣�Yk������]�������hS�����P���G��R��n�3ӓ1+v�F�%ZF�Z�{�4��*$��ewuUzz��RI���la��}�<�~����&M����Wu�����WC���`�}xA;�!��D�i�
?;0
8F�,U�zO��_������=Y;=�v���]+�t��L���Ic�� l"�} GO�S*�9��Z-�[k=���m�i|y���esg�U��Z�.� ��u�^RKi�MK?���/ ������: 44�0ɦM�^�Ͱ�c��Q{M����u�0�D0I��	�*d�(?���T]�@��1_z�@E2�<�����������ti&�GO��L}x�V��	Y�ǒ_���Z�NH�a]",�9�l㮄/)��<ON�2q�3�-�����ZAxa>��V�yQ3�#�9��^KdBȄ9�:����Y~F޼i�$h�@�?�7�N�Є���x4���74�x���b/0��#Wr�E��d��6�K��v�͘-�|P1-�TX6a�;b�����$�idN�ٳ?�W^Q�[$بrnR�	2+[[��\k�Y7�gA�����*��$�nl�͹K��*A�r*�Xyɖ�S�g�	J�
^��A6M�E����>ҵT[[�w���G`�+)�KNIqhɧ )����*"0�`��Zfɔ�u���|�C����T@��)�=���g�`���j ��f���.�ќ%��/�j�%
7r�)3)w��\jp�0i��������5��:UOHj�<�м��
�f٣�'rv�L�
�ucr*�n�²�
�����h�*��^�r�̉�"��'�4X{�J ���C���y�}�乐������k<�˺&�nj�B�v��	��J�����| �j����v/�B�7��^�V�r���D�`R�p�|3z8a�+��4wU�Dƨp)8cb@k]�eԁ�M	 ��Fn���VJ�+e)�~��w����0��%��{���� ;��)��,T�Yb�l��/�HJ����ǃ����4��� ßMG<�u�{��$���S��Ӄ�G�S��yPY��H2�������L0+��z
t��gB��J1:��1^_Ĕ���2�Pa7u 0�ڝ��������L6/�P����w��n��C�L�Fߋ��,�Q�|�B)�F�F�1�>�)G�5�ߓ�_���y��\$����)��j
5!j�e�����b_A�ϻ>C�ԡu[�8m��*g��g�7;~(]����c^�Q�C�M�3�J�#s�
����+[[[z�=y|r���ͽ~���^.�=�_t��s�";�n�z��ņ��9�%|#��3�c�NL�2���	�b�5��`�5+��@�lK@�uX��42T!�~	d�'���b�$`���J|�V,B�	/���*Z�d��ŐK��+�ش+B<`�9���������1�f��A� �8s�G!g}��`��y����v��ь�eQl�E��"*V�:�4	�!'�P�F/|��NG�Y�;���5��)���Xu�F-��I����
�0��������e	b���5_���s; 75Mދ8}�ef��k�\�/Efb85�ZT��܋�2�l�H�+8MH�u��^dR����ZĈ&>��A�:�� ��P�� t�5��$�A�8x��d8�@���8i`�Ik�$�Jb�fv���V �h�G��T0�4�ߙ��!�F4�f���'�l*+���k�L�Im�`����L���y���IW�YLb�z�ڒ�f˂pw"Ͱ([��Rn�(�w��ryѓ��4�4��q��i���W�|�t�cJ5s]��0�h��>���,���Uֵ\U�AO��+���L���������L,��{��߁f��� ����׊4��D��\���j֨֜*���m�Z����I��3�q09�����D�ߕ�[��AW��'p�0�K'�	C�j\��H�h�)�����S�H�ao0��b����Ǧx@��.Us�W�/to8O�N,a�X�$*�,aۧ�Y =wԵ��8<�%��^ ]!T5�4�pҮ��*��8\���UH)%�=E�a����Ș���L��A�X?K�RE�k�TjJy���������r0������FU�5�l�7���=�F�P��I�w[�4�g�~��V� J���)����+z�uPF�K��w���H�c���p-��g\���1x�(�t��}L�=�j�O )(�q\�!�'�dCcC{N�X��NO���7��V����W����_��]���n��BTҍ\�U�@z\8�J�l#�`��� ��6�(� 陶������Цk�x���Z�SА�Ā����#��Ĕ���AB�	��ϜN�17s�)�w�BFSB�\`zۡ�-Efzx��}��`��P,V!^AA�E�Fʞ�쎊�<����J��NTL\�&p�{E�V�TohC�=���� t����X7�)���Z��;�FB�u���Y2�T�,��������e10|��hp��B��,wO����9��58��°��x���:sfs�KPĦ`f�(<���v~��<�� �4(VS]KeY[ݑ��B.��h5��W��_�4��-��|3����rCp'�Zi��R�6-�@ t�Zb���~X�d_�Ϛf�(����NR����1u@�ρ��o�^��/��qB��i���xH�2��yB@�S��2��z_F��Գ��ȝ���EQ�<:k���\��\��X��6��	m&�e�����7��g~BZ��4�-Js�[��ɡ�h��z/*�h����q�VU�E&'�O�����?I�up�4�hT$֌��7�-rt"ŋ����7@�@z}SI�L�C ǥ`H!�����0%D%������%V����.�[�z�J��?ϊ3����r��yl�nh�_���R\<=���G�G)0X�>Մa ����ZI U�Û���[��M����m��"
�)h�B-dfz��lD��S$
&�z_E&U���]�{Q?��٩�ߧ����ME�G��*F����:�X蚫��gI��!D�<V�1^��V娬��I�9z/J����:���"/Z+s�e���C�dћ)�LeC�L)Y�K��t���Idђ�l�h�(<��VK	��86��Z/��
��{�.��ab�dm�G�A2!ƹ>
Tga8�1x�(�r�^�� ���`I�Def���L�fi�M�ݵ{��sG���g������_�j�����]��0�
+ͺ����|�H�?�����Ǹ9)���,88Tro�<R�f���o�'�6p��H�,�)���D� E�Cs\Z��ĲN��Z�A�a��ή Ƈ$���Vqj����F��w��U�_7���5yE=�70��f5�M�>�Pa���J��E��`�0sm��"`K�=]�Qa��~o.MF�
�6<Kp �Y� � 9 �40Q��
�PС��P��<Ϭ-�u�C���0z�����:,!�UNW�o(����-yƓ|�;�^'�+��8rvN���+ 1�&�*s�|p3_��Y���k��vU�-�	2�U�j��8��#4�̮m���.��z!�K�9�~GU����r`�9��p��i�<+8`
"n����=�� Ģ�,&К�i�+A~E����L��Fи ��7 b����u���1i�)�L����2l_���\*�U�k�N)�X�)V�뾡���ƶ�������;R�ؒB�)Fw��X������V�ym��
��ɱ���P�Xƥ�U�ʂ��t(��yz.�7�y�D��S�3��6�����zOo���y�����
�Z�m��e���T�����;k��T p�'ɧ� %�����X�xU}?F�#�v�q��?���L/_�h:���#9����}b]�D]�d30�X��b��^ߑ�aY ���X�f��	$��Y�������w�u��#9��9C�J�� �h��z	�
�gϷ�%���F��}�
2��B��	<;�BE�
��1m)�c�{])T��i(��S@V��Zg[u��"c�-�7/Cb��3c��ZE��N(��:�8�&���{cMȺ��3SJ��*))�(k�juL�Q����&�Z�z��҂u��;��r�@�[p/�q�u �t�U�(�_�Jjj���i�ǜ���+,�zް��e�\��w
�>8&(	�ws�2Pd|�nKrͺ4jUO���p���o~�O~���������N���w�R�>P��?��;���/i渡���S�NW��$l�e*�F�C@c�ŷ��tac���y�Z��-2\0i@�b0k��xг�L�� �E%KLk���Z��
��M�c�M1���!]�B������1�2�	�C?��ϱC�1�1�uN`$�D��9��R�cƑ�%by+�M�t�k&�A$Q���2�)��B����E�ad捸�
��$g���!dn��������g1�a���_y	L��Ge_ψ�࢘�J����3���^ߟ8���+���&���tr�>,�趦�ѨΡ����.��FC�^�� 2�ʴ�jN�Ԕ��I�@��  �g�en�!�	�٫�� ��p�U�`L�u�Q	*H���p����=���9����B3^�Q�Q�qgT�0�=���ʆ�kʪh?z`j��4(�{;�,X�GK��eL¸ɫ�	1H�يL�hK�A<]W�¡ =V>C�=�A�S�~��[����؍���Os�)���PwD�?��3��@q�ۺ�S�Uk�B��m ��V�m���+'O�(@��CLiAZ�@{	�U�lS?\�$dĊB;�Ր����K/I���k��c�-Fe�)0?�!����핰�������-AhemH�f=������|0$�m�B��V4b��]�~O�s��x&��!�W9�H�_��^���p(u��}*���	(!G���P�홴،��O5�l����d��{P�\�5� C?g��5�3����o�ƚ��yB���P��J�^����8�=b}K|�d��ө� ��z�u�(3�PRH" 虉������3׽��1�P� j4������]��͝�Bgr��9���e��;I��uX��f�ˀD1,�dl_Mg�ui��.>��=/���|T^;����~D�U��2=����Q�#aK���<�PQ:M05�?�z��޻o~�������/����.�7�\!���������/�w������l֊u#��m>�����K1���F�ω�e,ͲL:MmLVLB��\��_�M�x$��!_ �V�����p�K{@!8l0CͲJ����en��}��'�#cj������4D`0W�gG�TZQ����b�v���st6�0p}�f��Z ��@.��>#�z���?�zO�1L�c)��-R��t\L�]��1#H�Fච�Q���hiX3g	B�Yc��7��T��$b%�\g�ϝ��*�q7hk�$O� ���	�wC"p��&�ud�eu��X���ɘ"�ē7g���83�<Ch�A3����t��6dk�A�h�ӟ��С��lq=! ��"��esG7�r�`
�7�j��d8���� �GQ���K#"Ӆ�y���%����G�!���a}���Z@ ?�WRmT�tt�k�-�S3�3����5���64���]����d~�ɨ�VL��"�!~�A�0tǘ��Q�1'q#����P��� 
��}�x��J���	�#���H,GE�Ah��(��6��B V�F>g�Vg"հ�g|�0�]�i���Q[�.l��(�K��1fb�L�fR2K�����$rh1[hO�u�ǁ�����YH�'6���2�ϐ>�%�(=���q�J\ gj�{����˲��-�9y��|�����0=�ڢ��hؓ�ŉ��Ƌ�k�Ж��t���[�uE����zzJ@MQ��5e���J�a���R-�����ޛ�J��W~�1G�9ǚ��HJbKvC�'5,À0<�x������?0��K?�pÍnx�eI�	-�`�5�,�XY���w�s���o}��M���S�PA\f��{#��g�o\�Z����˭������s��TX��t��+5��x�6���lb�oἵ.�=_<�x��� �MB����5�� u�X���eX�5S���bU���l?���A� ��K�K����{l=*���=a��o�����fu�>��<w���D'CƳC,��;&f����6�
�	���Q�gy�+�����?L������ܛ�?���#������/~��U��n�Jj�)7c �7��D��S^���!�h���,~��v��}��*u�m�J�*�9&��! .3dB�p.�Af�ד����/�n��w�!��ϲC5�h0rU\q^�(oA����ca�05P$�Lj�>k-���1�d{�%���k�\x�(8�V�88��ZJ�pK4flO�@�Ga��=�<��@�/�;����UB*Q�"2;9��'�n�`:U^*���$�օ=���:�����5k]��u��k4���H�2�=P�D*����܈z�H��c�MXC9)�ڍLճ�$�R���El���X���|r|l�?w%�f�����8<~�X��ޞ��ׯ��م4k&�ʮ#Wƾ��iR��BK�.EQ�D�&�p48ƃ'c?C&��(���h�09E�"2�x���RU ��Y����Y�����}ֶ�3[�5��F��$Nkd�9��4R9�J��u���͛��(����u�^�ry6(!۵��,�*��A]� E [��2*|d�v/8�@�#�
��
Rٚ��_lwD��w�
�!gs��}Z�B�6a����y8a��2��1m��{�C���}6:�Fe�V���q��v/��?S3Knm?�	��}��ɏC1�������X�ځ����!��҃N��W���'fsN쫵���Y�<y�����l��!�=���(�-��p�u�g[��he�k��ѯ��m{.��LnwL7:���t	��3�+�ձ�1IȎ�a��z[ҵd�܂]�K}� ܋'b��h|rrA�u��Q�Sk�'��;�K�J�q�9��:�֨��i<�^m��۰�_��\Җ{|R��+��w�m������#K`�=������Mڤl�����~�^f���婜b$�*b��H�+�������=qO�9)=��9@��.��o�������������)S���m�����������>�ɏ���,~`����/ H��/��+˔�HO�(��Y�( �+mx���׫�W�ʲ0D�D&Y�CRU\�6����Ei�)d�]�<��{8��}�{ᝏ>+��3w�(^u� 01�{���xU��^�?f]���{������<x�2�:�ױ?4�Np�K1��de>��52����C�<W�jRzik2 �z�d��N%�@�ES��h�\��$�J��F{+����:v���f}}#��\�(��%�ʓ�S�s?���#�>����G'c�F��a�~���o��Y�+����;���;{�U��*��UE�GfO�ev3줡ӈM�0� ��qU��g#�0k0�-�s�TC�-�E����Z�����9m5��v�m��Z�[�IM��'���X��D
�m7s��EH��x(�l�|�Osn�S�����~�g
�z��gd�=[ˁ�#��
!��ز��d6j��T9 ;����m$:i��{�#�����ة�;�۫�&���=;?�Y�&�ym�b=��B�ô�'������K���a�ŧas}��:X�U�h�3���Z{b4�ʢ���ȾN��UX��g��?���<��y�J����.]���ւ�/, XK� r|v�s)��[�#��s�C;���>��N�������8��>�"_�Uち�{s���K��;{��ԞY���_X 5��k���k��.s�X�2=o ��!>Ԙ��(M,Y*S����<�l�1�LUI*���|u-��Tg��T0����R�� ��Y:0��=�S8O�y8�GR(���흰8$���!���,��$���	��NՖ� ��h�1�SW� /�Zp{ws+R���±%c��H,L1�`�K�ь����%S҈����/��7�ݯګ׿K��m�IddI%��������U81����w�`G����!t|�U���������d4�����{���o��o��n \���w�����������A�M���}��r� ���K-&zNN��0��pR����TL� ��V�� �\��L���h`��%�^�����2�0���<|�[�?��gB�d����=��'/>Ʊ�؏��.�W�Dҝ��>2e�s�[]�����8�9�� ɍ���(�pbN�q��șZ���(�;H*T ���P��q��m�?Ae�
ۄ��P�w��Y�H���*1{�"'�6^�W�����ե���"�����#�&���7㟪�@�q�(�����}����ߋ쵎�C�U�7�_����ֈ���߻��tIg�W���Ap묗ays�Of!3���e}/�a���	�s.��B������H%�Io����u��q�%YleϬ�7
@��坰*k�mꡂ&�2s�T���vp�9��	��Yh����yu��g�´7�IXn� �w���E�r��Ʈ%�U�b����Ԃ�ks��7�«�yh��(YF	�
�p�oNCa	̨|�=ɚ֮�_|7{���:��o	T-G/,��}H��pe�8bJ���˭��W���d����/�m���1O�v�7�P�z�Ջ��5�fa5�9JŴ��*j��~��P��2����a�1�R;��%Ȁ�o�,g�m��Y��L��%��V�P��jc��ve�n����̂ 0Ggr�����2�m�x�|��(i?3o��b݂�חΠl϶��]ZPfA
���<W�xA�a&��N4n��!�}���ְ*l��u��pB�0��$WE2���H�l�F}os�'@^2�j�;dA`{sc���{8;�	��Uk�O�7v^��+�CM��b ȴք6��mX~�E�������/��Z��Y�x�Y8{�q8癗[K?�'�\綧H�?Qp,mu�)����_��%�[�TU3��T�a�%�E��J��3�=�r��g$������(�q �~?�����������"��_����_��������}�/��Dgggӿ�{����?������_��gf�SJ�����U�\�j��P?P���xB��s �f��8�K0�f�w��J�ˌ C�"\ u���V�Q���3fp�ui�1�,�a�2������d[�eѨ���.3l0_�B�Y�:�V����WJ������aL:w0���,@��o�l���h��� �}�I
ʸ��$�v����Y8��JŤ�/��T�M���LI�n�*s���iq:w�8��=L���8;�� ���и�@vh=���_GR�,<;il#�x������I^�:qݘa��'-Y��gR�%H�f�lk_�նf����P<},3��va����j�AƓgO��2vF�C���i��#�Ys��ҹo�>0����BXp��-�X�����>�WPiJ��lHW�q/d��@WT ����XoO���>o��:�g�fk�7�3=�:L�ah�EX�������� l�W�J����_J���ؓ�g��밓\S��Y�*l�t�{a^��P��)F�)y_3Y�o%g�y�N� U�D�؂�;sHw���eQ��J���`E��U2�|oY�]�Hd�T6a��Rm=�� �*`��[�v�8ǐ�Q ���^�O�d�8�+��ߎ�rB@WJ�
�m=�_�cMYY��R9��U&*9T���"ۺ�ba��^Y��[j ��)�y����[(G��[���w�ľ�{5���(��N2��߆-U'0K�B>s�Xl,�XK{��+��Y�"�e1��8������f�prv����:�������{ZSbgg���\�ѽ�ޝ��#�ΰXɧ�JJh1����~_^Z@y�77���g�勰��i(�қ��fN��b�U�F����qe�<��İL�B��"��ן����.x#�V�2� L�d��K3b�T�1�&�d��+����!!%��x|����o��������o~�?�����������]��y��v׳M;�����>{�緿�����Liaqfp�2O�=���h�Ъv����O��"��4�"30�M���.���V	z��m<��tO!�+�Ԓ�P���
@A�y����h��c��&,�g3��(Z��f��Z�C�p$�j~�̳�B�G%+�@㶳�_Η�rT�$%O�9�e��l��O�#��������X��d��4�A6V];)[M�%�a��'�w'��qH�3��i8/��~�Ru�.�������pi����T��2Rz��z_��}�ޕ����c����Ox������+.>n��e��:6ݎ�G���I����o�6�hW\KM�b��-� e�ud[�O������N���h�+a����FQjv�jВ! Y�j'!�&�u}�;x�)M,'�&�07�|�����W�>U] j�^��@L�=�d�HH�C�n֚���]�+sVh�{;S�}��s�£!H��k�_[f��$�-�ZNjh��:��'�)2e�7�F?Ҩu_@;���P�u���t��}Op�26�7p���l�KF�{�xp?҃g�ZQC��s5-�b�ak��H=Ϙ9 �^��	���nZ�Fh<���ϝ�\�@����N��V���YޢH2M�@��6���ގ\)����!�"�*�>�]7r��gak�sl�oj��L3��v˭��u777z�GO.B��܂�Ԃjʭ��B쵷щM-���{mz"E�%K��k%^�|=�p�z� �����|n7KmT��]��8�V�=M�ۅ�7lw�˰��`�)a-hZ�G�|�D׹��$�Vu�ֳ����E�Y��v<֙�t���$��'�bę�]���h0��}V=��Ă��k��,���B~6�]��l����ׂ���4l�ݙy9��#	��!� �Q�-�����.x���t�ZR�4ɁL��D�PkW.|Fj|ۍ��KG5O�6E���~J&��g����S�X~�ŧ����/>yi;��K�I�[���U9[.6���|��O/NN`��pQ�mޕ�p���i�}�X�`D��^�S?`�;�i�&��0Z~�{I���'сR݀��+�?:7�4;�O�����������㟆����[�z[Psa���W_��g0�Hl7��������}i���خ�a:pY�Rg{-���9���[X֊0"y⠰�{{u%"9��2ouQ�&�!�ǘ��>'v�f�)H�>�l��ހ6X*�o�@�t)s�)k�Y$�k��M��?�'��	�������S�ⶤ*�KBr��������9��{���8�F�jT�]��$c�x��Q��|K4�3�2�7��4���-܏�a��cϜg��f��H$�G��7r"ǖ��m�/7������*x�ᠧ��[�z]+s��7z����r�m�:�8�]Aq��̱9�fз/_�	�Q���@UgkA��~a��9'Q���zc�9f�'�4�����&dT=����XL�h`�V��KF\#M�!@�sk����Ѹ?�}���4-f�$y�#�'2��,m���.��6�k�ǅv�F��w�p<T�P��nN��Y���+���^�]cA��십*U�%ǉ��L����[�3ڮlǑ�-�{�r�9�ڨ��!Y���8��$��so�Ck�fR��=0n�qL��W �n���f���sm���O�=���!#c׼�[8�B�b�`�7ǡ�&�]-4�-��ނ��w7"���t�����[h��+���>��Y/�j�Pq���z��n�珟�'����Mby��Fx��%�Rغ�k(h���%ac��-�� �I���l�*b�ԑF��&	Qg-H���u%��ħ�9�Jۗ�����x{��8u�-6��V�tK�����P��6�W(uM.\���6���_��eZ�>�[)F�"��E!bt���� ��CF�%[Y��[!��a	<��kW����|n��Ss ���<� !����ERo�	cm�g��@;q6 l0ɞء�*�(&H��q~	ܡ����Z�A �m��}D��j9`�Ϩ(��iR!��5X6�,ÖQZv��������?�o^� ���9�A8�������w�Y=���<� cy���W��Y�� 蹹�V&N��<����^��=�51L�����~+p����ޢ�_o׺�N���K�,=��X�x��{�>+�T�6�قw@ۄJZ�*�SZP�T�dֵ������FMTPǔ�Y'�虜lt����f����gJKfYi���T�dd���+<R`�����Y�)|��| ��[����D��(���*�t�~p�����?�+��
�i���&\���Y�r��<)c��Wka�zd���uY�����_�u�pP������p&i����L-��|m� ��d�h��؏�A�3R���OT��"�$	�&>�n�5��j+�n3�l���܎Ӟtiz���$*��G�@� ��q4� � �ܪ�>�+��sTu� F>����0*��c˟z��'Dy��ht�RK' �aϞ �A[��X!}k�N��;*q(
�;+�y*�`�8@��جO��צU�N���u��A�8�Mb;iG��^�>L--ZK�-��
-�F�S���{�҈���ъ%â��,д)�����X������z�i7�a�q�)���tlI�.�~V�^�R%Un�!C�M�ݚ]�߇
�A�E 4���l�1 _���b��;�T���a�7�Wc�a9��z|r���AZ��K��CZ��4�4ާ�,�^�N����B�U3�v*��^��n���4S�>ȏ$������TI�+���}�n1jNk�)�KE����S2��ԙ�8fM_L�0cL�L4���s�'��1�m�����*��z��f#ph�=AJ���H/l��ۛ���K�,���͑��Ys�e��6���R�F{�$��/�t�ʂ��ڡ�Wo?�(��**��V��vW��J�z)G=�4Fr3��[���3��J�4��<N��{:Qv�xj+�j�P���$���
��Γg��L��ҜY��x�2'k����l��EuE)q:xkW����DY'Fcq7��[��ת���'c���/̀f�i4����Nj�����>�H�q'*�~m3����P[����TRve\[S'a`�{̌q��>j^G��FՖ�>N�7+�V�-m#��6#:Y"�=(�3���r��r�o����drTr<L5e�����`���6V���I�$8\gq���������\T�Ж���=w'��F�����ֲ���R�0D�z'fe����co�ݷ�ǆ�
�v[�7��	�)�3�[/�b�o����Wr�`.�^����-Ñ����@	�5���P��C���ܦĉ��&���S��Co���q�V��jY�~o��H�Ȝ��s�6:��r'�	�}�$5m���k}D7��v�H2i�[a&��ko�Hg�	�l=$Y`F�W������Ω�iܴN��@�Q�5ڙ=��4�9��1)���I��K*�*�t������W����%Қ��qЋ|;�����8��"�[b�NB�hPI���������?��!��#Հ��9�]Ӝ�6�意�}�R��
�ak����{��ْ~p-�S�N����2��3-��LK&��W!5�:�=3��C AE��I9�.�yXٽ�^���,���f���m���VÙ�Mg�m����{^Ak
Τ>������l�6��j
x�O6��OP�x8(����ׅ��!84|T�.����$�(� ��k�\��]�շ��\^(M	C�yG�?��Q�����I>��At�k���^�G��W���k�CBLN���'- ��	P��.//����y靬���(�)���ļP��S}V�m�KH\�'��� ���>�@wD0�E�g%QT�2#[02����бӿmr�h�J"0S���(�_$h�;Dz����Ӱ�{X؆��1C�}���N ��;�r~��b�m� ���/B�Z���f��K;�w�۰[-���Kaw��LU#+��،��������x��0u�QE��/�a�����`v�n��y߮���w������f�U�A�u����O,�8;�����|f�0$d��ٙ�gm�p bu����d�bL�j��d��D`2���y �#���o��)T��������;����J�DT֩��1`jDX�zW�q舴	���h19F�Ϛ̍}�x��N+E�R t�>�J�(]v��������e�9��:����oo�3�R$g��W�+����ե��u`	`O�����o�D 5���i] �*-�ֈ�9�珞����-�����ŋ�~x�x���̾�9 z{{�^_���}><k<�g�ؘ}j�v~w޼y��;~�T���$j�e���9o�HvH�*8�}�z���Ʊ�k�<��K��~lJ1F$+�i��$����$V�GO�H`���i!m�FU�<^�n�W˴ږJvfv�8���=����)��%qĞpY׉���z@��^oe�H&VU�P[ϕ��kz�ח�D3QGPv'A��y��lhᰖ��b�*�ZK8�>-3��$?��س�-V�$��hroICr��U7��;E���%p�{�NBp���7�f���ŋӣpzr,������ �� 	S	]��ٯ"�&�~ǧ01�a���~n��[n�!i5����h:��(�/�I�=��,�xծuP��pE�K�?t ��c	����U�({�-b��j&��$Q������v[�=~�����tE�؇�(�������ګ����f��'5��. k3cQ�V�hpf�s��/��?�I�� ��eipl�q�{��OADg��, ^�������4���Qeo5Ek^;
�	�$㱜}�|��?�4Ի����F���DތQ�Z;zC��Ğ����2^j�@gΘ��j1H����D�_�߅kz�vHӓ�����6���W�������ga��B�#8ԑ�#3h�t�4X/���UXZ�B�w2*C ��C����&gg�(���(�h��ؕ�Ȍl_m����K�e��y��١�!�43T��kh����'O޷�t���b�
�7/Ý9a�i��qh�!��Z�g�8��4�� Y��{�{�%�$Q4�ZZJD	�b
A?�	�&2(�;LP�b�I]��q�|%���#����A�*� �3K�:�r��� ���Xw�\��ٽ�B�=��5�{�I/1��uQ���I��g��J���>@ms�����H�o������=g��ɣ��q���g*.�/�Ά��x[4id�#H����n�p��  �`܎�k��'��6�٣s�����YGp;��2��W��r`�ޟ�ȫz�c����s�X,������̂����5�J+klkzd�n����V��v�@H�I��ğ�Z=88J��:v�N̴̝aC��!�D_�J����:�qmQ@{�:j����*v~-@L�"Ac��^����0�=9:NK6l�j�D��%Q׭�<k�)2�}i�8�dU���"��7�@�ڻ֙��8ar��!8� ^±u���J��Y�g��� %� �#���"�5g�Zg�K���r�h��H�"h	�����$�,�Z�ѿB�`���Z�`ی:����sڙ�9�­��j3� N�������'�6$(Ma��X�B�q" �
�UL9����*�@mBO��&�LEZ�UU�H�޲?P4NU�@��d4����+�����U���5B$��3w|U ��[�1h�6�������H
�g`ᦙԪߟ~�|�^�崙d���5yRMQp���L�M z��aH&���5G�?:O�?��jz��Ob��Ha�֫�*��C�UǾo����Dn�4Rt;-e]o?Zf�����)t΢�7��456��ۦ�u�TM���CUt�ޚ�
f�o���m���m�W��ٺ\��:{�n�\<�Ӣ��fM����,<=��@���z��T*��|��\��`=_��L/���C�v��8)���;�������2͉���&aG3��9 2�~����Yvc�p䜯�j�������$R���0�,;y��G{�Y��GI�LO��q���q�ǜ�q#d�Y���?����$� ���9ZR�����!����6���Ce�r:�H����yФ�m#`��P0=Qŝ�O�Q1P0M��!��H�M*�;cZ�8+ ư�ZP��>z,��]�� ��ZY��tq�ߙ؞xtv��V�@�~�����`b{�J@_�jj�s<���\<�9�l�2�մ41,�&����}6UG4�����md�&�����;@��Y;�M�
ZoTVF��N�	�u�`)�{L�W�S�K¶��Y��E�>Ϥ�S�@�s��VYxe܏&�E��z�QW��v.�j��6�[��F�0]�:��͝����qA�Ğ]f���>a�:r� c�O�\D��t��JKe6��$���5�$8tL�.��54����'Ǫ ���rT��, �&���Ҷr"��w�p�'�X֠v
�<N�\�&��6�=�(l�p`�%�30�;&��T�))�F{���v]����X���W����H�'��KF~f{��j������%�58���*��<�M��rq#\�jU�˥���	����,��aU�¨�*�!�T�[���O�c����T\�ݙCe�}�f!�� ���jj�)����pF�⊶���A-�{x9�_�8�[I�h��u���:����%T�|�6���>|w��~V�-��5�	�Ţ��9��T�M����{�Yxtl���d㇚v�	�`7F9�u�����"�Ch�n�ǵppp�-�Qu&Fݬ& 598�#�0�ͱn,s�( 4� U����p������M��I�M���1�Z����`�1�NQ�M��y�b��d���,������U�A���`�MĿqt�<��=;2\Z �!�V����š7���G攦�pQeDޜJ�d����9��9ݍe�4Kִm/�W^���	 �:f�Dz��.H7�$�F�bFo4�` }~(�S9E�l����a\]�01A��jq/��{��9�cF��	��8T@dJٵ��E�G� �++�4�@���h][�5��gE��k(1C\E��Z����ȵ�?IV�����r�`#�{�ȬT����6:D9p���W J)��'�T\`1���0FIEvn�;���g�M,f����:Rs�]E=�*eӔO��R;���{?��!mŢ�~פJ��n�a��V�%�!t�wLJ��³��<0M����?�d� ��ɫ}ڢL�@Ըc�Qv˼	^�t�s���F{�~����1;�j�Uv M����~�H��`�Q${9ڻ�gdgbZ����%
�v!�9%|&��9?jW��1��ڵ�ʭ�2Q��{�͌,Æ��|�O����i���ًh��@�z+/�t�`_�b1ؙ�Fyy���%9��=�D��w�H��ue��b����2�#��@xvr�i���#�&��C��]��;�� Ba�O`���
����>�
yn�>�����_����.V��8���l�TM�I�Y�4-R�u�pN�8/�gҰ^��O��anv�����s���^�nW�R�	3�?��`���IrUe9��!������ʕ��+I]�^D�mz��tXƎJ��7�O�AJ��s)�����X�m��/_��'?	a��s�-��z&h����t�`������,,1�p�̙�����w�O,�9�{W��,�W/R���&j,hjz�}	��%��O�Xc���]�ꕨ�9$)^S?�E#,���2e_�
��F31�fNQx�����$�Z �~��9R��w�/����ѷOS��nQB� �ۭ9̞�ӫG*~ǈ�}a���}�}�FT���>��+�p�e�C�*u	���FI}�W� ���b�zo��z�ADy}�����Zz���#�	J�"�A�7��<m"�Ib����rI5Cl�&#�q��C�Pٶ�c�Ty�j#���VS/�1 @���q�k��-΄��{6���JDlbЋ�*�II�;J'd�Q�i�B�k�_S��,�9�,?��L@��ܯ��im��u^�~[��Oi��*U��ֻ�+E�9��v��c�>���-�܁�#%��:�84t��?�����p\d�FE<I���M�W�*�<~O$\�f����W�Jp?���^��3�B@���0����ݙ��t~&�#�&o��u5��e�k�5�3*F9�e�`K���0N`z�Q�H��n�������_SDn�*sY�F�w{��*{�!�i�u��g�Q.,�����p�[��0�G-#Բ�9>R�Fd?_)�M���ɉ�]��4Y��i������1<=�9��$��Q�+�js�X�SO���*�j)�~�	�����/ʜ�%�KR�gϮ����Ղe����3�M�n��]�8��L�h� %b7�P��X��m4*��<iqa�g�f���V��+%�6'�j�/�v;��Y���
?��?	?{���i?>7���a�Om�����vQئ�tt�$��D\7i�h�v�!���lF���C	!�ջ,�3l�{��t�"۴#�S��+EA���Z\��5�X���Ї��!���}�|3m�U{�7I��{b7���5z��B�ӧ\j�l��]&jvwk���c����q��N��*�'"֔J��oc�.#��%�F�7
m�,FЕFV��3Zʪ�PGf�@-���l�ᢏ����N��a�ݤC���Qݖ@���f��dP�pNΟ�����z�Jp�O����kν�_9Q����1�<��fun�a;w�U��ႀ�B��+Z�l��IHfG*t�����n0Ny�Au�v�����J�!�����O\� \A�:�Z���}+��Tϒ�O��qi�%���]H:�~e�P�C���3τ�$M�ht��QUq^��8�%P��^�ы�6j��"�K4>��n@���ul-/�ٱ��û8�8���[%��ڙM�8����g��	��ꋗ�[Z|� ��t�+�A�J��.������c� ��ۮ���q��F�c����P���4v�:4p�{hZI���d������@Ր"!���~(h�Jc��4���m�*P~5_J��(��h50�Y{+�g	�f�=���&�����Ȃ���ӓi�����DO�sT�wwz�p��#O�DSs@4ag�~��ן�U����;!SZ��}"�����b@Zı������Κ�9a��|��P]_*���ӟMb�@匠H4��0��="�F-�`|ܧ)o�Q���x��/��N-���:�l+�TZ�_J]�	pf�%0V��"�-Hc�aOBВ8����"�0-|��
}Zu�bq���x��	6Ȑ:F���L�hek�1��<[{��zJ,�a8a�٪�6�GT'��]� Mwd�5>	s{γ>��w������Oj�8�.���7q���>�X"�AWxi�4�lw���R��eH�7#�T�5�pL��Y�4XW�i�Z�&q��	5`g��yMu�
AK]Gv�0�ߐ�}%_v8��p�p&G�pb��Z�8�7c�;`�9��v�R�F�7@C�6��#{��>���IŜ������	j�nW%ј��/�n-��Ĳ�dɮ���'}M�e#��˴1��C6�srhN���Npj�Q��8�>����p��C��<�2rrf�܌����rL]m�̌i���/u=�_;}��<�.`]^-�B9>����'*%T\0�dz���2��0M�5�Шr�ڬ-Q�@ʲ8�sY��O�@I�:O�;^2�8$k����Zy5�̀��^��|$x�B4pJv�6�U�*B����+1e�'�
w���@@f�^*JM�L��%�q�Ld}W��G��p_i����`80Q �����)��&�28�5�E#�#�g�O����;P��g��`�&H�t��Q�橯ݺtL/*� ��k��,FVK�t-�9�5²u�"A�pZU�jL�IĹ����p$e�e� �h%���\`Z�Um�J���}�
&v�mX �����>2�Ь�#����#$�N��AEU8#s����ϥ��Z�mI��٭ծd�����[�y�hjks�TS������9�������(MuM5$[�c����W����p�Z�=H��ő��FǈY|��%T	bw�^�v�����H���9�i���j��V�.����pb��`R�8�RFձck��M)(��6�4��\��h�P��{����d��ڠ����=������9�3n�DSo7v�W���^�=x�<��;���R����cI6�lo�X���A�GTp |!v���0�Q��O��&���"�]�����w~�����ٙd�bO�\�t���9���*5Sq�4��Q��39
�>
���QX�W�ǿ�����]����O����`��i�� �z�����耹��Q�����7�-o��"">�[P�x��J����A쒠���\�}/\�>/Jo%Hc�������خ�����Hs�WI�K�g��^���	���f-m%��'#�"b��5m��{�}�c`�D�?E�z6<@]���n`1*�	�������؁(���ZL��	7�^Dy�Z&�e�Q&?�<L?�v0��QODcu>	�v�>�0�۾�_�*�P�S��s^�����2�]]��x��G��9�<\�����&ЁC%b�DJw�=l���*A������w�*��Z09ޣٷ��K9v^��;ܴ�tR�����<����M���E�G�������8c�~a~��Lu~{/�>�������̉��8idPGf�c���FY�{���S�j�b�ڀ�"M|<���Ƃ!��b��hΚ�/Y[�:q�$�C�vd���Lnd"p�E��R��F{��zON�A�V윕�܊��,%�WZi�f x��7��,��O�n���{��Z�g����7�� �	X[a�l�n���-�Y��3��4��c����:W�m���Udp��Wە�#s1 n�4(+���=�s��э�w`g��X��ꨨ�̇�5�g��a�Q�Ͽ�`w�U�S�TjT� 3��l�a�q�\��γ�ߺ�E�+���
�ҭ���Ғ���ԭ�+�O�C����U�kI��9=>�^��� NaMډ������r�#��[�~Ǿ�n���L`}��oiHf*�j����5����	�z��o�|��u�KkrNOO��"bW�&����� �ɦ�?�8���;�!ڙ-X��<Zo9<~�$|p�	&-�۴7�y���u0��Pp�
���m�����S~GA�{����ٹ1��@
`�
'�g჏-��?s1������{��-� ����ff�fjA[`m�E%'��Z�=����%���p�ǷamghIk��� Yg]�8$����1*� qLJA����r��:X;��Vj�y[m�$V\����[PN��m�,
�z�����w�(`ǉ2�&�L"�NK���aƯ��]��{W�\��F�e%��*�'��@��i�'0Sb�����UҧT(���0�˿�ĭ�S���iIdTL���t�)��Ӡ��p��H
���HKy����XBp0lȆ���fȓ�h���.�'r���F뢸�� �s;��O�ftP�7�+s<+�.˘�^��7oJ�3��&�^Y����? �S��j���N���2�ji�a���:u��P�S
�>���"|y�F%s��+��=��-���xؽk��2��L-��:ƔlM@?qX��a}�ǁ�[Y��b̡̆��#�P��2
�G�(��F�΀���ŕ�/<���sF*�3�a?�\�������	��ƌ�z��2
�g`��x���Nv�p��w�e�T+��%��xg�Տ�J��5�s3�%&� H�Lc����ފ�3�5����Qm��B8U��b�9�٫u�Ύ�J�8�T;ɹ�p���;��0P������#'~�k��oEj�9f��X�Ɓ�Ρ��|�J渓Q_�˷�7v]�p=��M�����u��J��_l�0�µr�Il拁��L�I��q��ֹ:V���T,)���6^Y Ĉ6���e���0��}�]����NAƠ��GL�v��v��� y>�l癲��-�8�
=#���Ó�~�����N�^������FqQ�C4v���'�E������ҵ�8[�˫}x�����6�s��n� ���f��طஏĩ�SV��]����
��%=�ϛ�ͭ֔�٭6
��y�w��pk��d�r��Bt��V{� �B�:?�|i�'��_XP���e%��Ιa~��&|r��ֈj��lo��~�٩x�����{�'?�����p���P�sG���ztd�����Q�$��oz;H��0F��Z`��;f�9Ѹ��-Q:��@�I-��;λ��Q�ŵ�|���\Au�iop�4jc��V�L���A��	��Ep7"˚���_�+��Vi�ԽoF����&I���J��Q�c��tS��
����	�"Fjf�u�F�׮~{�q�&�K�rjE��"��l��P��7q%�ܹ��_�v:�l�^�E%�oFukG����{�:����M��IK��>XGn��d�
G�q��_���?_\_*(�8�ݏ�����]��o���Z�j2�u�a��t�*�f��[�5�ņ 2(��B~f�6vΏe�� i���rW:Z�m*�)*�Ս�Y� �`��N�����8q)���am��a�G��1�|��U�Z��д�]�Ǵ��\�3z���[������gZ!��#�9oo	fo���c=V�Pq��U���yڈ0���_�z����J�� �0OT�Pۢp�q�j�¤���	pm�d�.ˈ���u,�i;�����vcho�0
�k�������k}�	�)���@����E�z�ӳ�K�ɡ}�:_��2�xz!��N��D o 0%�əP�))�!y�����Q�*x�/���f�%�P��\�sTZ�ӁcoO�M+@=�4���-&m��r�d�'~l��[ 3�z[��ϸ�}��0���!�T�
��7��esx�\�biA�ʫjgm6@,���=������I�<;����`��%੼�B0*\�Ƭ;])�sP�� ��oOվ���ؽ-_���ݛ��7�$y�HҒ���}�#�W�F-�g�W7�§7_���]T�`b�?/��o^����^���{��7ՙ��@�~��Ia� ���S�)�x��j���&	:�o���>��	���w�~p���}ʯ�g��ax�)��������}f����| Y�F�@e�o 4�D�Q�>��$���W`���i|�=�U��A�U�t�WvGڄ�>v�ǣe�����c�I��p```tr�<��Bςv_����Km�%J���ә���vܯ����i���+��$�`;�ÜIY�+N|Z��H� 4ᅘj+rF��⃁��,-��h�-� ������=`x��<J��,�%�A#�N��Ne��N"�[�#��@/�'��dG.D9T�ksj�+W���(�ڵ_��ajӫ���������Ϟ���G'� 	WAHm��0#O)]�6�z@MԉY'�[S��
Z�RC���		��_�գ�o�yР�ϤR2� �Rf���#�Ժ7Ld3-��_��R�K�:�����ڽt:�=�H�A��!�kZ'N��ȴs��L��Щ�(n�����\��E�A���[����/|�h����ĔѩՑ�<�sxd2� s=��BG!�F�uCB-����4�}�	T�Ҽ�\�� �ѫ�G����R�g�(ܸ��wLӬq����H��OF��\����c�Y���u ����<�B�x��s��g��췍F�qby�`r�˹Ɇ:K7�,���Z��y 5HGj��y�
W&HИ/�h�,םSM��v�VZ��o�dd���dj��ԩ����h�ٺ����N@ןz�`Y���qn��낼M*���k-3o�M���
��[�Q5�%\t�PM�ӳcC�n,!�5NkgAt��I%�-ි����@�aZR�;�|u���=�$YpK��@���EU�b@�W�Y�m��]�ܲȻ�}����\s�-`����6�;�=�^E�"O����-��.�"`�>lv��_�{��&fW���?.6�:���%,w�_ؾ�W�v�U�ڳx��(<��A|a��p�P	�Z�Q�;'�k�(@�=��h��~K�ݭ��2/1p�p���	G�3o�t�.>֜�Mt �����I*�Y_�2��
Y�<B�`/r�0����L���Q�FS^m��׫���|�^��y�f�%�H�Z ��*Z��"w�J���-�M0u�[����!��Xy["�(-��nD����h N&*Bgj_���9Ү�⤊�W��2$_��0��ʸ�U�h}�<��r�ss�s3��<�E�H���*-{�5��s��߄��kɴ�6��󻹜�m� I�a^4�q�d+�G��E�{~4*��'���&��a'z���`�n�8^߅����]�K���Sw�P���N���>���5ylh�c��TQ(��{Q�lY�^7fܖtY+ϣ�Ō>0^�׺;�ylJA�/'�3/T�hP'�J�����{⣓u�P�	��)͢�����!q��	aO���ŕ
�;�Q&�b���ؖD��_�4?P]�E�_�w Nz@��h��Jt?���.8Q,NU`%3�y/�?"���J��"h�g��F���b�Kճ�9�vk�a�i��4����8؍y�>�����E`"�Gi�����[�qjLS`�*�՗8`"}%�^��q�.��K��ݝf6����S�RqE3i��g���ɩTuE����"6�9�oW�u����;�a<�x%��G���<k���Py�_U(��\D�;T[�X���D`���=�+�LW1�r��{σ�}�xvA�>���� w�	��!���"��:��e�C@�g�.4�4R����`l&i9?;	��p���!�&�H��k��6�v�{�g��c�H�Z�ӟ���p��+��f�0fac���Q~��?�f�<=	�fi�|�o���2<��+gB=2;S#��#k[������������q�(v.��MG;4Rv�Ѥ��U�}�Jmu�3� ;�)���V�Y]�tYσ7�+�
 %衂��Um����%W��ĥ�"�wRe����W�݌��]��jC(��;��!��g�����P��ȩ�H�г)�($t���W �����[�C� K�0��T��O����퓸�p��*�UA; č̈�m�]��N���k��{�٣�;���co����W���8Ϟ_���Z��m��c��@���;�ؽ�"�#U�\n�p�}��f�*�/yo"N���$��I�fb��="ǅT�'�����������K�d0k˘J~�#}�hV�9P �!.���U�\�U~Ƈ�Q�.�0ā
���N�g�����ǒ:3��U���M�$�8��յI��m�Z�������=�S��0V����Y㣢>��q58���އ=�ek�[j_��&��M�|�g�dc|k���׼׏l����<Hl��X��q�0�=��*<M�r@��o����qx��Bg�'�L�'/u�����t��4�9e�����7��g��H�D����7[��6b}�#�,uW9�����1��3���0�cwN�������rv�5�L���W��<�́#;Bńi�'N0����,������F���Pm�086��
^tyt^h�����qT
�-x9�Luц���ҟ����`@�+E�mC�]�����x�Y��g�t�"s>�J�&ޚKBd��NO���Ž�f����;����N�̯�<�:q�2\�l8Ӵ���&xA�\0dL�?� ������0���g>����5� �2�p6�H|������f��/o��mi��u��u���� �vX��0�ж��f��j��Ĺv�.���ҭ��{%q�'֊�@�����7�)%g]�d�c��X
U3ق.7�Pr�xT3�L�����!�d �pc�} !o���2K�"��֮�gմe=U�k���^�3{f��$)L9TK(o�ن����dL�I]؎M��%�L�`�lPe�Zt,e�]���
g	�9�|�x`R����a98�����ĊM�[=`��T������E�(����:����4����mS��2��i�g�!���$<���x�[���k��,��l�w<gO���"���YSgS>�@�g*՗��O�Q���2X�@�хc�Y9y�6����f0���NYF�7;\�mT��#z�+c�D*��&X�(�}��Z2/���H�Шݐŀ�+cw��=B�1פSU�	��P�b��8��"v c+�<?pt��w|�%�Fx��U��
�u�u�y�W4ƃ��݃�E�܎�/Db1��꬛�I�c,�*c�p�o�h�q�Y!7I|�^� "�%I�2v���> ;�:i$��c�*f�]{�k{�����	�X�/P�H���8��`g;E~����p�U�C�܀;�=դ�����ܶ�C
U\�s� &s�&9�����S}@�~��(�Z��mҁ����E�w�E¿�/���+0�����F�"��:�X� N��;���p��Pmj��YGO��"ڷHH9{L��]$0 ��X0�ĂE@�y|&�~���svd%^5�E/R��w{��y���}غL�뼥��U�r�&�8+��T�:G>��TvZ���*�)��G�7m��^I��Ȅ+���5��4�����������>
��5=����0�~����N��G?
����?cᩒpf��,����l�.�X0���px|*���т��̂��؃�,�i�
�����g��^Ciۉo/�+�y�"	h�Z��?���R'�|�DUh���%��); �Ci �B�Vv8��.�6�����ek������/x	�<$:�d��C�FF��0od�
A�Y�������Q��"C������(a2���Z%�4�v�'Ü1��tJ80�v8��}p��d�Cl�q�\��i���3��Ӽv,���� ����쥢@�-̉&vM�$\[�E�1������3˂��_\�	�8;\���?�8|�{�W�V�J���o��6"kK2�
U7ݐ:>���@O�t�/���Vl����Ǥ	�s��z������{�ؖ�~:��* �a,���kٹ$A�����+�V"��C���t���wK��-z~Q9>�Օ.@�^�LT�>�����{ɹg�C��<������C[���"�pȈ%�ޣ�����p��CQ��$�MG�"}��h]6�)a]h�����;3*[R�� ����(��F`A�K1,�²K��{�(2�A��kmt��LJ��9tU�N��k�YAY]ؚ�^
'�)�.HMC�`���}M-Ŗ�n�F���Ֆ���&���Ր���G���+q��{	��q^i���jC!'%�B��y�[K�x�n�O�LFg����\���sg�ڗ�X)N\
D8�(TI���v��݈Uy{�u�����;E�?�~L�}yF�,IW�t��A�6�ABT�ǹ����8�A$�N)��#&�R�lv�5��D`Z�5�r����q]e�$���lz�O��-O%��6lw�#�k��w�V����}QT� Xf��yH� .%M鉇�S�I-���]��臋�Up K�E�k��� ����\��C�j���a"�1�����=Ɂ.A	�8�*�D�7����[,uL E���0)��/�3�mg,������'� �ؙC������W�U�6˳e�7��� f��äE�잞,Y�90u��|�AP~��N0A�RZ0 ��X�&�2	Z��DSL��W!���ZJ�2Ǎ�T�8��3q8�4��DMǪq�d�
b���Bޗ�iU����z߷���!(�	�ۅ��7��*˯-�xs{�A/��;�
��[�f��?��O�"��������_����]��?�@��Ed(��̉(W�����4NR'0��)�� �r��R>5'���)#SV�^�eO���n��핍�
�u�r�* @W��QE��� �Z�I�$�M�^�6�L��Į��}���������`ieD�_����S�ht�o��Ut���Cu���肭 �	!���D��+��0Z��#�|�*@��$
6��qrR�j���
'ϣ�Bߜ�׵�o����x�l�`�&�4��;<7T��Ǩ6�As����b�`e��U紩t1~���ձ��g��N2���8�]*�&�*A�WcZ�$��#3�M�\'m�:p>ꆅȝ�6�b��db�NUi�`/���'�C@�j!���A�Y:r]�(�	�,�]��f��=������TS;(�z=��Cz�̜�T6��e%K��9bۘ��t2
�I?V{��]����i����n�*��>Z�yԋMb�RA
�$��y�_�N��Gl����JP'arM���C�]��L�ejo�yKӁZL�74�^�)�ť5�4�F�oS��3��Ϝ�������ql??Ӛ~���J��?�Qxq}&��������g�6T�+9z�w�0=uQX02���z*�b�T����q���l�j���yJT]
�z;��|r�j��|>��Ae;aȠ(����ȧ�4�0�iKޣ}�|s�̞��l�նH����u��/������k�lJ3�m�$]t�eـ��Q*�R4+#��a<�l=
�"��� Ϗ`���2�|�*�����Q���h���:,�o����V�������p�K��c<,0)��F��2�:[Q^��d�#a�`�,}||jF�/��s�Үi4�FG'�Y���
w����g/U6�蝏B�NC�V�o�&C��9ۦ� g�*�*�J���k&�6Yg�(qbqT�6����1A^ߜ
Y8$m��I���uR'i��I9t6�d����Q��Y!G����V����QN���k��� �D��aba�[���8�}���3옍c̻����nz���]v��v��C��>�E;��6Y�QnV���DХr�d�����h�'��d���Bq�Þڕ]{��9&P�Ҵ��}�ȲJZ����Q��F�@U��1�7�>��C֖:�W�-���G-C�| ժ^�I�7g�r��Xv�T�Tq,%.�@5� ��8� e��J��	� ��qG��~q'�g�x:t�D�fz�jk��������P�R����o'��Ǜ(�ՓՆ�b[���L"�`҇�&�7����_��;m�p	�K������v�*��A_�#�b�v� ix�vF������}�f'��{��DQ�J�x�|���i�W�@еw; �ߝ4x-O�\ĕ��l61��c����"S�=UϜ�����z�Ha˸����y��e�=;��}�}s>��i���Ex��Q���£'�ó�g�������_������x��kC�+q޺��b��&U�?;��[F���2��9�]��pY`�D�;n���1z�}�g�Zًv�����rd�	&�����l�A�J�Y�m�htdK`�n�֭��Y��qn BJ=;�n��̡��w�ݽ��}=_�p�����M���mo0,��Q�+�D�(Z1�ҜV_U��z��BzŠLJ����I, !�yUa�|d��xN��F�arv&v�*t�Tf���׵��Ͱ:9
�)����P^_���c����L ��C��� ?�Y���.f����iEdԸd �`d�n�՗o����%ѿ��g/����c�?�4_\�U���O���?��k�p|t�h#��1�CA�3 �!���J6�Y3A���eK��0�#���vL�{��隐0C@ej�Y	�v�k��vc������N��R���ѻ�5�E���¢Px8p���I��Ә�'Ӱ�Gഭi��i�ޜҿO�c_:���<�S3u�3���4>{uL����a(�E��#�%;EEZ��̵l�I�L�q~h���# �P��E�- �݌�Id����p6�����٨|��b���J��#M:�R��΍9�3 �Y�g��2�̢v8yP?E�,y������Ck��)sPc�})�۪�cP����zg׌� ���a�Z���S��k	�֚�Y�*h/��A�i��Y=U��Zڄ��)RQ��e�yxn8�z��Idt��Q��g�8���ȫr�w2��5�4:M U�C�;)�-}zONM�X����|�9��ŽM��w/��՗3��D"���'vVk��C����Ϟ-�ıd��<�T�N�JR�fE�ԫ�a
�=��v����vp�8"�CL�uo;е:>DU��w��u�<�Q��S���D���t�R�f�{�?�4��>~�o�����?��?S 7���w��������v�xt��i�����Ă�e��yV%Ә}%O��y������d�iߘ]�d�D��\P�F�a6Tio6i|�(���)�� :�|� W�D��-U�`��z��F߮z�M�"J 79���`,v�$�Kg��Y�KʤA�����.6��ϒi�&)�Ѹ6�vx�z��0_��/\����߭���� ),`i1�C�
�Q�'��ש�;�\,[O`���c�JA�hy:�Pg�����qX�/�,Wan��"�m&6;A ���Ix<�n�~���MQ�x9�	��r���e~��[k��G�k��ڈ��%�Z�b���x/fP�C�]���+U���+���,s��G��o݇��v&�{O�f�a�v,e���;3n� s}�ٹ�z�=�/��$Ikqb4�5�| ��2�7v� �C?�R
$�b��zYӬ�?D�F�jHɿ�5�|UI�O�g3T6"�I��e ��Nړ�e�j��Rw�_��g��zc����o�ao�Q� �R���g��F`��9f���Ϋ�x퉦�2�Ĕ��Q�>41k�Y>x�﹯G+1�pl�K�@�q�
GC�L~B-�����
m��T��[�T0#�trF85�huh�>���y� O|M��^�D�/�GU��/�5*�D�쟏�fO�r|��Uӣ�w��dvN��1v�K���t�Y�|��>�$�iA+��7K�?w�O#mTLy.��	kX���iw�CK��?l�bj�|O�}4q��&�� ӉW\I����z�ժ�U�����L���c�wm�*�I�v��L, v;��ڬ^���8��8�6�9��\hOg�LaU*���^iU�S�j�
BG��y���\��k���󊙟G��kl�-�಍8��k����h�����,�k��վ��9U&���~��$[h��=����,�M����pk����X����G��/��{�{�����|���"���W��iv��T��{﹩s��Ɂ3���M�"H�9  X�dȀ?�� @�m� ��{��`X"i�EM�LO��o�N�S�O�k���U�94$qL����9u����/����k��фVx �x�ń9��L��������eƟ������
^4�=�#�������T��{��P����K`T���� �qG�ʻCr� �@~m�e	rrl=Z0�:`c-��1��W����[i����|�k$ ��9��$�O2/?n�(z�z���'s=��o�=B)!--����Z��c�KN�\f�C�G�{��dCBdPtr �q��5�=>b�qO'����^�TP�v�������j��f�Ϟ��76��_��#YBHm�H��)��N@��H�C/"��+�\�s�4� �؎G4��a������R�ѦF{x;:��t�T���ͤbn֕�ƶ\~�1.�F��g���%��c���+�9��6!OȢiKQ�� ��p�V��� �yk+"c�� �jWf鬪���X�^�4ż,4KX2�u���S��)�V�b!iµ�*FR����R&�mm�T�[���و�������ځ0����4]j�1�U�8>�E�tN��"�\	��+�2T7ixk��C�J���h܎�i���Y�Ġ��wx�`Σ}�e�@�������#��8D$\��Vdj�8�Т���(�ϒ��Ȏ�#m�r � Y2���P���--����> �V��ˌ�D�uhJ,3t�P^2 ,o�d֡3�.4(q�Ԃ�)f��w&�e$I.�gQ�-�9���|��Vu�𱘹A���F�y�yYPV�'��)�ž��ֲ!X37K#�g�1;-�ߒP�	�0|.�,��c�F��2N���1j�^ چ2]p���*�:6q{r�
�L�������L®,���sXv1y�8��2�(���
�f�/;�,@r˼��Ѿ�������S�>./>��<��K���hC.*`��l��/�',���ϓ���S�~�����V��-M���i��X��zt�/hD�� ^Rd�޿A�O��ya�G��G�0��4Zug� �g��Ьqr,;[�$c� '��B��ށ�\�ޖ?� �VƷ��B�~��s��҈µN�I}j���9��G��Ӳ(��rY�s��"���GZXc�c�bi9�ؙd=��Þd0�R\:rk:��n��ܽ+�ܻW�so���������ɢ������wo{s�`0����գ���L�ڷ�l���N)nF��m�|=a����c���%�)c;��d,�:��ZQ�DVJ�"��P�h�?�[�����
�vY�z�>"p�E+�B���d!�G'�<��?��#rywW.n�6����'�W_���$��t"�\���<��n����07:n^�:Ȁ `�BӄY�*��H&��i\��"`��g�j�k$D�KVi�&�&"A�6�U}���:p2��B�{oaD]5��Ff|��>H�Ce-��!$�܈�B�Im�m�"i��p|��
&����d�CG	���>���:x��ی��p�@���)�x2߮;ChFx�D�+#"�Q�T;ZO�T��' ��E��P;h�![�.KMwl�uy� �E���Ef&a����sv81� R�n�8�n7|6j#�5��¸�s���\ �igOV�iܣp�P$�S=C���Q�8T�&�)+��f�b�:Q7�	�曆�H  &�����)רʺ�
��h�j��0JL�`�3���q���+�F��)���t�́��;���OEO0����Z��#D�(�@w%kw�Wb��p�b�A>a�~(7����@f.M?������<�{f{12s.�͍F���':���T�E+�w%0���g֖s?&���?/g/���^���<�#?��$�þƞ��QP�üB6R_@&�� �k�;ؗ��lw�>�O�9�$fG�1�����X��vw��߸ʌ7�WFXK��X�t+e=�!�lOC��9s�7��b�&	K}���_����2;ˍw�к���/�E7���76d�!���<7�9�)���1��_R�q4������sGQ�.�Rϕ�0g�A�]���te.�u*p�G]ګ�Ṇ���{{rs�P�tB]��W�:<���խ��'�����s������'��Q{�휫�eպw�����~�㯿��S7�^��a+}����Y��G:Y�Kj$��u7��{j�-���H�H��dvKf QME[/8%���6L��], l p~EV�wp(/�������s4�>��D:�7���(��}W�0��ר�;@�j6�b�p+/��~��K���f`��$�Cr��=�AԌi��M�n5zd��¦�d��٬�y��e	�D��6"M��C�]:(�@H]kƛP�d:�[�$�>���p�B�5ҿ'?�@  �m��[�A���:q����J{�:��3"�^�b�:��?�t'���f�U�H�5V ��8gG7-=M,;|�=�f�~b ���nlY�FI6:Y�e�jf^�!;x��@v�j	���HǬM)�H�2G���pF:��§��2�Y��SQ��	[�#L�G8��8K( ��XDU�	��B)"��Yڐ�4K�5ߟ�!W2�E�5��H��� Vd�9/+�uL�ٯŞ������
A&H�7�B�yy�;��(�$�n']=z�f ��a	�H?�h��.?��#3�b��ARF��� �mh�fu1�zo��Ib�z)vF� ��<��+��Qqى��$��&�O�O�(�F&d�*���S�H��kټ`Z�'O=�؉y��v3A#��tY.�ٔ���g�C����r2�e�K�NE�kgЗ��y��62�UF�dQ�eYCxk!˘6h�2/`����y�l���J��ö�4����=x�eqµ4[Tr�ܮLu`4���4�畑�7|\�pA�ݹK��Z�����������K��L4 =�sh9��� �y�b.Gӹ�q�9O��u�U�)F24��N�F�e��Q�ӳE����=	^L��U�ApH��P֮�Z��_h�,u��P��(&遻�)�N����ܼw �^�*�(���r�6�;���ŏ|�s�K��O_����۹N�&�s��^x�������g���|�?{����]�v{�<��tcE�u"}�e�o��k3xqH�aKi���Q"�@�W�=:�E| �]hh�\���܀�iD�R���|Hn���������N�m��+}�~���X_���SCM��S�ᣍ0&���n������ kC�UL�"����ې��DE�BB�����H�pb+�֑�$jJRE��1QγѦ��ђ�L%�~?8�9�]�"v4�.�T�<7�'d$P�a4|㥙�D���q����(����[(M�&����8���8Ն��86Bj�B�*��V�2tj-��X�R�6q�*�&�S��l8��A���-�d�k��Y�����Z�^M�����<C��2�x<�P�Vٔ1��8x��(�����9
�J���	}��<�4K�lh�nKIޑyk%�i�
=��62��e<P@���1ޅh团� �$"�%	��Y/���7�k�`] �^Z�,��{8��Ԣ)#�{-����,ovK����#���Φ�m���X#p�nyf��Y�"i�� J2�
��� W�V��C������
�kF����D��,�uL������ƌ������4�̼��o���EA����,�p��}n�k`1����+oK1ݒ3xT�x��F}��9T3=�#g���ps(ÍM9<�'h{�L,#�^�|���90I"�\h��w\�<g�:;��2�V�C�������|��|��ے�*�c�S����#;��ek笜�xIz�A�����Us��m�9\�vM^�M��59�q&��)6����<e����;�ԟ��f�H���tj<N�͙X��L
|E�������=	^�"�t�-ZIZ�@�!V�	�|qYfAyE���t.���ߓ[G��N���ߔ��o�ͣV�;���g�����o|���w����G�J��^��O?�`��/~�o�����g��O���\�u>���@':J:m��s+{��Ɇ6Ln�u�]�HQM�m�P�E��X_7Uzy���BL�O�����"����9sF�66��_`jRs��k��eS�v� ��ͭJ��Ia��I�dm�y�FO��}�8du�S�3�f�),�D���28���hG.�H��pl~��w��"lx�,��##G#��*@S�0�$�!�]*0Aj�n�s�F�)I���u�JF�A��>7u�
�5�7Α\X[C�(��!��%����n�ύ����"��Zc�qXo�^�F��j�l�Ӆ��9'@�h�<�k����q}�,*x����Ш+oE�sH��O<�mF?&;\�Z0C��s�A\Cj�]B��ںQ�je���z3₃��Q��\�J~~�M�α�DЄ���r�e���JJsP|���E�l�c���R����N��PV��F\�u�����U21��lTm��\m�s<�ڜ}X:ԥ7i2H4nhc����+��7�+�q��.��jx������Hp�"����h���(Y�C��E�%�t(���?��`�a�l�l<�������(:X�!�@Z�	^���A�*��ʺ�h���M�̂�Ѵ�t͢ub3:带P)��٬8��S�*C���s	��>u-���� ֞�n;�_0��5�흮�te>�dz(���l�~��Wur���X#�Ya`	�h�����˒��t�.�����)��{�k��`(]}^��#��酡���S�����Gr����3��ʇ?�)��OV���G��}��lk��fs16(k����/������Y98<a�4tu䓣���A�2��)����H�Ƽ�����ͪ�������L����ˏ�J��	��D�[wvd�/���~�Kkc ��ɮ7����#������n�������ß�:�˿͵|��/��pp4��/~�k�Gu�k�^gWc�x b��,L)X
�6���tk�CG�u�e4p�B���-`��n!q'�A�b����k��Q��֖��-/#�B��6��0$��LD���K��G�����Q%�n'5@̸u���u�����C!��nײ�?V,51��K#�U,��im�س+����9�����uB��H�V�IEv��}� �:&�gy0'fK.27̂k���sc�C��h� (rҷyU�ɓ��)6;�J���?F�5{P�?�5�d�J�li���W�Iɺy�0p���J���K��#m�t	�`���~i@�qץe��ܱ�E�~KL3\�w@Dt�E�'����L�����m�K?B�hNJ�A2+���cb��p��,����IIܑ:��C'�����!���ʵl��1��� J�z���TZf!�kg��\���آp��[��еv��5�<���`K���9'��6�)u�[n��M�v��V���<���v�`�-!��=����K묶���"+������RL���#u�캀��Yf�Yݘ�c�o���U&���*��`^Yd&;/�TF��K�LV��g����^����`�^�\r������ ;�6�f�bʳb���آp��+	]{e1�V{ Ћ���z���"K6%�@Ĵ,��U���l;{nC��|�����0s�kx$������A� #rQ&
4fǇ�Id��Nx������[G���z�''S�(�Y�F.^�$��k?���g��X.\~��Ͳ�0�욊9�0{��0�K���Ͼ�e����g<{ܧXv� 4ƸN�2���t&}Tt�]�  ��IDAT�|(d��	���U7u����=	^�\�8���T���Kg�Ƃ�%Jȭ�P�z�/:�u,t�Ci���2�A��UGyq������������gN�]� �g�ym����׿���,Me��g�D�"�Kh�FU��&wn��$�!��}؈
7���Kd���d"�Z�]"�2���t
��$�95F;���@�G�ty(��v$����|r0�0	��1p�� ���f�d�o%Tj�+���?":X��G	
�p�e�:K,��l�P��:ݾ�Y�-"�wA�
�G���Є�h�f'��) ��c��g��*^��)��,�`8Ȏ�[��#٨����o���Ja�Y�Z-���w�T�L�LLaU�,�F+u��[u3���zKqĶ]�J���M�.f��Ȫ���3�gD���W#��Y~H��80+����v���>@���
��jE�q���<���x�СV��$����Qe]>� �ݼ�[׍�#�&;|�bC�Ɖ�ٵ���=���:�j/G�9��t��(1W�����@��nQb��)��+K�Y�,q.5�ȥ��Df&��8]�n��-7p�4|%��@�t�u�9S<\�1SY�,t�YƣlJp��!
o�w�Z�v�?���3�n�H�>':I۳��4�c*��[���[�#4jf|J�F�$���}A�u��vb?��᳢�̥��1T[G(���p) p��� ƌ�hu:}f@�Zx�yD!:��v'������T�A�hl��2@�B�BKAA�~_C�9��)#�\��S�Y.ˉ_� ��kD���}Y(x�6� z:0��'�W���>�1�����/k:���hBsP)��(��?4������#���/ʝ;7%9�-��m������hHЂ���{}�j���n0�G{	�O�E��{�o��/��R�Щ���Yd1R[� )�]ή���h ��F͙N�cy��-����8r�������'���~�W������;_����_�·{���;��������F�uN��>�,5��ڑ�%PH����j���`j�ԅ?�v�D¢�.]#��F�n��,�@?+2�h-�yz�u�,�L+D�̪@����[����Q�F�3C��M��шPa�K\%���l!n�������X�r�N&<���R�L}$!�y|���'׈$Tn�qBmb���d.�Lƛ��F.塀)��."~��ƹ�����!�@�Ė�������\�LG]Y�1�7�J&3Bf�Y7ddD� gt�������XU�[��]��Mm��;��d�KQ��)�,��t��@,]�ޗЦ-~�Xs���_���s���Bc��'��aWU���=�K䔰:�C���ce�x�{�Y����	}��|���g��U�񑕣/�b�(v����"�^��զo�k�d��#�ԦilP�q~�Q�9鬒��P���u�y#����s���� ���ڭv��������z�m s�}��w$�{P7%��U�W���2^<0̘�x�P��w�k/"�E���Ҡ,��u$�-T�n�Ȳ��9I \3����2t��% Ĭ\��>�}#��-�,��3����W���6�z�>����������� A������=�]����i^�: y:��e�¸^(��^����<tz�r�{�A�'?�i��_�婧?&�M��,lb���cX�^YG-����ϦV2|���Xn���lv�Z�=�'�Ҡ'�`mN�Թ��+UɃ 7��C�V�����=	^����R�)=;z���#�I͟��7>�ܔ#� �f3�?�g�"�����x���[����>�����]8�w~'����?���_y�_�;:��N�Po�WGWy@��?K�m�(aԑ�[Yr�,��G�r�<hL ^F���y8Oh<W�`8R���w8��`"�L�])����\g�c�;"��}c���O���fIp��a��A��\�ڝiY�s0�t%O��Y��r���̶��P�:GgC���+���4;7>\��p�M����ɔ��9@ -�\��0"*����M�6����$"�`%��
��J r&��V`�3�q��*P{z�<��� 3��!u��ˑzF�_�VP�e�-�NZ�g�GjJ��eu,q��yr��*v�E&���2��_i5�-�@�{��ƣhzm��m��b���N���q'QS,+``-����Y8��M��� ��=�/����O��{W-�Ak���"��i�l-ˉ��@H��5��2`��Bנe�|Xj��TVB���,��l$J�Ⱥ�c��ׄ�C�YA�w�)�Y�s���d�E�)E��he��G���W<��];�9Q��ŬQ-kG`8T ��F�V���e�
�������y}5IJQls�2�%�94��ݔ;y�ՠ1��z�6��k<��$ΐ�`&��&�p��r�+�}�{E��hqAc��\m@�\�*�C�TfH��$�{QU'�ڥ���26B5�r]6�O��>(���M>񙟑�ً�Y3��i��½�,�űL-(�t����?h�e<9�����C�J�ld��[r�����C�#:F��[m�x�8ɲ��//�M�ҫ�N��r��v�4�;ۙ�bw�D!�J�:|���X���#����b��s�O?��~�O*��Q]���{o���/������1ϗ;���LH5/�M�-���v>���7��88������$�c�O��P��sK�c�u�+e�iT��˲0}�������+?C����u��Җ̼�A޺"6��&;m��m��o��FOm3Ģ�lY5�%؀h��pb�d�v����SG��
l���	3��q�z�c\I�,�O| �K����ƪZu��$-�h�~H����;Rg��ƶ1���u�я%"���X�b�]:X���z�%��N�C3B����(2uR� �A��J<�P{+kMB�����,n�P�f!1��j��Z0�j[^��8��^EBC�J%ZE�.���$d�Ox�%BO'X������ߐ^F��T��l6�v~XV]9��9,���+�.�u�A��Y(w��"k�����6�Iӑ��R���BIГ	�B��7�/�aݼg�g���筋>�߷���\����� ���������؁	�� ���5�T+��u����W�I��}!F�V�~az�9��b�D�B��+(lH�������,ϲ�O*�!+o�D�������Ǆ��+f�j\��Τ�7�j蹜��;=?��?���ONFg�Qh���eY��)�=-�<{Ef��y��k��e���~N^y�%�
!>�%O&���R�R:��s���I��Zpu���dH�V��y��|���ce�TS��2�Ȳ�m��-��I'co���e������L���E~�}��[�KO������O^�u��f�XHԙ�$����b�[�P�f�x��QO��-V�R'nE�X����Љ<�3Pt����۷eo�.5=,�̹Ic���E
߀�Y�6�Z�Ji]8ش ���oZq3�errpե��a�bD�YF�(�&�è+2}:��(17��%�)M�`��� D�a��؁�2O�_��י9�����[��ȣ֞���8L <`���l77��bņ���G��ua���g\L�W<�Ԛ�~����Y&�6X{uj�`OI�@�rV�{Z)ɢjK�G�_7 TqC�
7�$&�R�pVԁ�b.�ֶ+��Bto�D넓��iҠC�&�����!��#R���è6�mܤ]��� 	�i�|����
��k�+��uX�̩�r�?09��z��xA�������1���C X�+pRնFM%��I�Z��g�<��<j�sh��Ƽ��Q�-�| T#��J+��K(Ve3����qX��@H�S t]m�T�A�|�2"y���uA�����W"��aޑ+g�]; �z���x(3D�'A|o�R�ţf�� T�5�u�'�%j#�S�?2��NP�՟!#��/�}�*��2-��H��~�U,f�R���` �nc���N~t��©]"�Bu7�u����>�!ٽ�-H�"fIZ�n����N��pٲo.�h\x���剧?$��z]��ǲ=��t�dsF^I���E����/s۟(��b^��4����8>��n�v0����$]�ٗ�z�ԝ��ua��&r�Q��(����{�o��o��\��я��˛���i6Z�X��:���itvĦ�.���Vl��<��m;�H�7�^w J/��;�	���xP�%!�-ƥ������XzP�!��uߑL�P�\�T�5U��fߴ��]��5ZfQ"[l���[��t.  ���n�쮁
R�b�]D�,�2���4t!�π���v �p��[:��t�C5��)oa��,��Ӂ����z�ת�$����n MmpŲ<,�P�Y���H�LMɵ�<�,-"e&£y<�M���dM6�*�]�iYw��R��0Т0`@��q/���@ *��.!�6�ԟoQ�ŔSW{X��!���X5�3F��͵,�d�Pn��d��[�:��e�>vU�LϜ�i���0�v�t���|.�(����)���v7� j'�G���g�S�D�*��˔P/(h��gT,���@���[��-�6.n�c�ZgC	׉�!���x�b��*��>����:���k��?1�Q�9��!��*�c�vȠ�|�L%�����ǅYUM��t0�~1;�*������T����HЦ	�){|�� 5G(���0�U�묨��;��vWy�s	��!�����*9�тV0��0[G.��}|D�Y8���ΐ���Ζ�n_��`Cbݏ�������5�(T����vhL�-����eΠw��h�hߗ��/�}H��/t��쉡�.qas�ք�M1�K眳	"�fC��;_���~��Е�����am�P ��1;X��unYK�3d����2)O�����G\�UzHT��!_2<.M%���i��d��6�xǈ|�p[Y�k�\�t�U�#}<U7��ܫ�9�5*֤�J,�+k�N�������V�s�`,F�F�MBY�$˽���RԊM.�-�s/�䬋�؎�-e�唄_.+�s���LȆ����� �t�[��&T�!׺��"^#9 bY�*�躈�XW�v��8I�ND4_��2y��IW{J�����s��|����}[�,�97T��d>aZ��������M�-֥�%lǮ��`::�v^�Od���iG4v�O�7�Hl-M�TS��1R`T^.�!;1qx�)�GAHX�s���:0m���)k6�e-Q��&BdnD��S�B���.��c�mV����@��ݚM�[1ۗ��\[��x	�y��ȣ̆b�x]V.�%M��u?��R�g�ME\�/��]À����tV�kӶ��&#�N�����a����ٜ���M/� ��4`�k�b\)+�ȭ<S�C����q�ct)�v?�!"��uo��K�XD�Z��½�?�nA/)��4QZ�1�g�]���{C�i�S'��S��ܢre�f>�\"���X	�4�*��_(�W�+X�楕o�͌*/�X�g��g>�s8��D$�w��OqJ���rN�,��QD���X���m�;Խ�=��,�������K#РQZM��׉!��P�Me�<lCz�t�}�9V�{�!9w�,Mk��eZ=]���р�ۊN��L�!ۣ{D'I��>�<�ؓ��W��/�7�����D�Yny��|-��F�<5�*LS�6���'��ׇu��+r)�d�������4��铹���&�ûB^�=ѝt�Wu}���i�Gu?�s9�xn�(���s���={��r	���~�N�49%��@]z��-��F�	�˜)��d*�r�t՘N���
��������B_���\A�f2��Hۻ<P׆�W�@͢d�]��iqSV �w�ϝ���vdsЕ^^-Ӊ��w�n�L�ES�����  �}�E ��4�sƓ	7��Ɛ�s��x~s�Z"����$��v��ԏ��i>��RU�X<;a�gZ-F5�&�H�����i���N�*26��:�I�^��ׁg��̶�p݊��k� ګ-be�-2�iVo����iv���٣�K$�
��&A��I~Е�+-�#V
��8���צ��m7����Fx$��Vd�>���K�W%0�uY'�Fi�*"�H2�8(v��~8���H �\��g5K������eSK\?(��,$j�.%�d��2Ui�b��^� �uH�Ӂ/F�n���Vr��u�ū2˪a���ee�'�Gk��3�5nI�ժ�v�cY����/�/>��u�Wn��+>�oie�P��s����՜i_�2g��SI��rv]6�D^�^2��� ��� j����A'&�d�#U������t��t��;�`ٙ�V�)(m���L�x�`i_Դ���@a��KG6�wd��yk��w��͒�+�: � �bguW���b�9���{���&�����|8����M��Y���6_8��g��������I���l�~��v"��[���A"��T8}.0���p4�z���#iml��i�(�Qg_Ξ}1:Y�Sx|�Q���u��L�'0؊���|Su���	�L���n"�a[N�BN�aSl+H�:k���\��Xj,�.��k����9��'����'弖�l��e���ԺI��})��uc=��p��) �.,�Հ bJ���M��}���e�+�t�+��F�lQ�$��l`�Z Ϛpk�(��6�)������0��}eoOR��u�뽝�����с����qG7[K9#�Ԩ�����<�Q���&��JC�<H��lAL<�D�C��� 
�A����qA9��٠셱B��%/'�b�Ħ[���?D����*��FצL�Ö]/K�¨؂��t��%��`/�M�Z�a�37����Jv���!:�6x�Z��q���"��*��0$�*d����Ȋ$J���<���(�=[��7^����,��$<��̒���h��<�H����7D�9���C��_���ʴh���
�1uEVh����1"��y�e�����ٳ]�i;��,�Ē�y�2Z/�)roh��2�8!�gmޡ��8:,׭�p�<ɒ���3o��%�< �K��}Rji�F�<p���R�R �`U��YU�VB�Y���1���Ԃi���>�L��ͬkM��?/�8(��H�g7w�_�
k\4�_'M�ɼ}��-�.>N�H�;�Ao(mAń��붨�Fy�9������Y��@DUx�}}��K)��S,�M��^�P`LM�\�w/&|�+��/�u��u)�%�<*�є�{NΔ݋�f�/���+s:e�[A���߷��$x�[i���	�YJ��6����!�Z��cy���������$k��i]y�F���ν���53�n��/�$�邆by���j7�J3�Ԁ��뵤A������ �ӂMRĦ�(�l�d�ٕtgCA�i��)M�[v8T�S� ��m�~7��BlC�A����P������aK�c�����M�� Z���c��L3��kԏ���rE_KCz<A]$:�H��C��ߝ��"�`r���~���6[:Fq�)�H{]nH'��}�!���q�FhY�1����c���J�"3
�%��e]��ӯ)�S+�Hq����Px��vP�%����l�-l�v|ؒ�a@�H*��);��:��z��n6Dd��S��򬆕_�Zx&h�8�2H����/ԧ������-�m������C�����y���p�ALYΥ����Mߤ^��D"�kɈ���$p�u.�Am$]�{�I����mR�f�@,|c�r�1N�
����S�2���2t�."�E|qqԔ���d�L\.dfc'����#�
M����j�~�����KA5�>=���2���;-�~�Y������K��ˉ�Ą����v,V*L"Z+ɒ�� '_��l{�deda4E��%t$�ڐ�����g��2f��2���M����Gy���M�2���X[A��ӎ��S<T߷����� ��<����r�h��g���	�*'�s=�Flߗ�e�?M@��3�}��;����yVf9�a�vϩ��W==�f��'R`oʬ$Gb2��3��G�'U�Σ4IN��ߗ��,x�kc�2�K�Q8��J+�\����_�n�Mo6K��e�sr������������b1�u*9۷�KY�B��x��=���Q~�AI��2�V����d��ς&c�tQF�@S1�j���Rɸ�Ij�zx�J�x�ߕ���d�ăһW��!�j:�e�ZiQG4{3�u�Xv��V���]yG���e�{�ˠ�m۬��� �M�J/o Q_'v�P���T��.����t7�R����dqt(�_Az�Q��)�����pS�n��lYq�ZM
`��d�9��UuC/&.8 ,R1�UD�L!Ǯ�L"�F�5D������V�����A#߰-�ݏDTp�ύ1�SQ(�CQ{����a��̉vO(YT�ɘ�K��8苔$4oջ`��D�C�(����a�4Z�:�����G�5x�ݻM�&k"�:]W�ۡd�#���1�c%q��$R{�?Zu3A�0r�5�_�2;�uR5�2��z�� qS�ɧ���@A��� ��i�����_+�ó�A��B�T�Xمߓ��x�]�j�h������8�Oe��6~'�D��%T�db������sE�����Q�Ց�#kb7]���fa�ƱO`~��Y�;iJY�EYAF{@@3;+�Je{s���(�,͉G2ں���6�ܹ����7dz|�H2�yJ��s�yQ^�|Z�&��֥E ]9��s��֖��7�b)G��rr<f�{D�k��X��;���BZY�+��c�A�ݻ,#��#��Xn޾�f����R#֔��c�Ot�2|�{�p-G��V����G�����D�nd�~;2f:P5�m�펌��ѝ̑ڟG��<w������/w𣼶;oO6���a��ݤ�#�JI5��eXB:���`���Y�@�r0���3�*�)#���U��3��E�Z����SI3t2NI��"/ى5���]7�;2��>����"��;H���4�{W^�����gO�rF?#p{�p�m|7���wnȞF�ށsI��ql`���	P��J�a���ߍ�|B�|���~�1�������-��c����nf��hv�ӏ˹��֨/s�hf�1�}�U�����}����%C&&nIc���x(��5�@J^��΄)�ާ�0x��G���r�Y�u�P������j�z;!Ӄ^.N�e�� ����� \Y��b#2.��}�"��h��k�r�q$�g!�x��/=��`�5�@�݇b�	�xSTh��k(r_!v�T�kɻ"j�i�8p%3�*j�$��j��]5qSC%�-,ZeVE`Sx���|��#ym��Q$�>��y?����epj�xm��$T~(�����%+f-��$p��s�Z�)�"��仕y׿���RN�j���א�<��Q��v?fUu�+��g�紭� :h��jy���M�u�?�����ݛ����p�癑X���=����n�(1�O�Z���);;��"�����'���(��C�$����\_Yi�r�� �� �#��a&�f ���[w�p��y�e�.#���tN�3v��I�2Y��Ef:�Nk+O���_�ί0�!��kt��:��	�Jȶ7{��]��[TsLv^~<�����,��%�ƙ�
����':q���Q�HV(8�hzt���k������'?���P�3�<�_����|��v��jO���B����Ƒo������C/V����v��L⍾؟�^E�Ī�J:;�#=��꬟?Ob�~ZM5�IIՌzJ3��y"�V&ݡ��݋"�
8 u�V�9��P�)��D�%7F�Pj1��}��A�Y��	��
0���[ץԍj�V�]5TMcsA�,�P�k�K��.W�ߕ~������'6�eu��s�Q������R�r��9���Ge���";2T�2}�mNS9~�-�-X"۸tY�\�,����l,�;
�n���;�*2;�F#�A6FW�r&sȖ�g�g�)��5����@Vvrc:s<�e�$�ŲVp�h����(I*�J7�����$6I :�Uj�h�D�]�\�Ä�j��b��c�5Y�p(���_/����%t��+?��ȗOb��=t��m%��Wo8z�8^���t���|D�[Ѷ�&�SZ�l��0q"���DZ�b�C>�;X/�51��tFj=Ä�lMh%��j,��$�j,�ru�;�%u���u��pMֲe��[?�V�^���+���~f,�2k��.�5 ��|��j#��Cυ�@���t���{���ҏ9J�f� :�  �W�֖,z��^_Z��^��~��"aќ����������p_ap���i1��p4>���X6a8��چ�烉Yb�ZNu�M�sY�D"F `�PL'���[��{���,���= i���w��s/1bn�r\r�@�@���
��y�ܺu�kן�_�zP�^��� ��pǠ�!#1��XY�qvA�O�I����)Eyeu~�)��n����!^�	�+h=tp��������:�ͧ�>��˿��P�e�k����n���aY<��Z�@ߏt.�j�4�p�?��Z�I��4�=�H�
�
�M�4���i-ݪLIv�Z$��D���ԧ��\��ؔ5rh�6�����?�sE�@
C6���ϰҸ@�1K��Ԯ�)�9Ķ�sg��m�pr����;�~�$���2'�b4T��z��`���N4�9��+�'> r�y��n� "�E���e����}K�͡��O��?(r�� ��@_�������=9�{M�vG��|R�}�"g��h�P���.o|�[r�n�����}�lo�&�����-_�B��vb�#��YJ��zEstr�͡�n���b�c8����򬟙~e��Ee�P3�; t��7F�F5Mv�GV��Y�c��)� ��AX�k3ڏPŵz�pH�6O�W�����,�I���f�,Z�(7���cQPO�h|�$k_���Y][�ƕ+��ԣxY�H �JZ�J!�H(ӹ ���t(k����m뇺E��o�˲��h�绀�����2R̴M�Ƥɪ�-(;���
H�����e�P���@�\9\@ƠIN]�)®��u��͵N�!|-��J�dF`�����LAB��d�� 
�i�\��=�{��V�̎�/]���z����w�����JO� J/݁��1��j%�]_��� ��}9�{K�NiJ3��21�8/2�G��n��,4`Y@�V�����7ޔ?��W��2Ԁ����?_�i��:�VY'������Ƌ%%��7�xM���w���]~*�CxA�8e �L5v������_R�|��L��J�}�xO��G��e�@@d$a��|�0�5�1i@(���ݮln�d����Չ����������?���"���|�/`��o��ٯ~��#+��d��:�*������B׃���8V�Q��rmڪ�*jt�|�H�&g�nȩ�ȅ���(���M���ZG���PQ܍��.�i�n�@Alʭ`�ŕ���e6^Z'�Q"P�Y�A�ķ*	�ú��և�&3����%aC�|���}�\���.�̜���8}�	�=�aS���J�'Lع$�f��FI�}
���lh�fL�& wl*�џ��x<����|H_[�"�h`�I�����7e�K�>(;���d�]��:�����_�����,�Q99JV_b��)�ں�<��ZL������1;�� �/kؿ���I��)�K�AD�;��wuc����<2�zZ�q�C�t,�#��0x/a�� ^�~.��y/���e-�\ˢ�0���R�"�E�����"9�]��>���F��^�]X)��="O��?׍����h%i�b#3�S�l�>.�J�.k����y���`�̔T�AP�H�ʤW���f�c��>u'6>F.>�� Q ���Q3�^BZ{�U�O��$k\�pH�^&C��+�_I���<.f�*�)"�Y�\ǔq��>P,b=w2ܑ��Y,�O�L���Kۊ:ශ�mI_c�ml�a�F�˒�����c��?o�~�g���K���\r��%aw���=����,ْ_��_�ls�<3�g��ƌ��i�(�$(֔��8��nܼ._��o�9�I��a�3�=�]���Ȣ�Q���$�[�,��D���>�"���K�SY����u�����'��Bج"o�v��ԳR�Mt[��;���ɯ|��_*&���_��K��o�u��9�o~��7���crp�7��|bSC�}�~^�!W8�մ*���C��U5�-;)���#耀Ke���ŀL'���C�@�#9l���8�Hw/���Ǎ���PV�h(�N�@R�A���� .�t�r�i�
D9��$�Í�Ί)-u����ٔ�ӏ��m�粗��d|Ob���ċ�-�-�r��;m���[g8��n��+��f6''�!qC虞[E��� _��F�	�5��^�th��v�F�,}A�;�md�"����H��#"�Ήh�5T0���)�k7d>��$���pӢ,�L�6ƈ�9̽:�n���Ϡ�z��A�\/��1.��e��̣�Hv���:wc��W�@3qE����2,�[���J�<،�ȿ/X�����'�ip�n���~~8L����>^��g!�.���;�o��{��G�y�f�?�.'����q|��OL��~���vl�=6���հ�qX�w���l\@�5:H�Py׎�l�|�ܚ�L���U>vA��C\�^���x0��U��$��z���+;e|�������4/}���������/tB6e��z1a4��X+rD�]�EI�^Z���1��p]Y��k�帪���J��v�kn<9f���9�ww�3���h�2�"�i;aV*(�M�9y��4�3�|b �r�˫��*��O�D�������d�.˸���ݥkS�6I�(2;p~Zz�s�my�_��~��r��m}�5��t_h@�L�i�Ӏb>�����Q+���e�b��ٓ��������X��z���ۢ�T*�X�l�d&�A[�:���o��r������A�7ƽVk�֍���F���x��~�_���?����u<�����/��}_�W��׫��߾�1|�U׽TcAdz&I�׸I�mվDA֜����Z�H"�@ݞ����`��ʶF�n
P�Fž��'	V>���`c�7����Otq���Œ�f	J��t� ��*l�n��ϲZ�^��1���ٌ`%���^{�?� #�������:��L�r��B�Jv��d�%��L�C[�Z?���N���b.G��!h���]enֺ�H~�\׍$�Me�����o��7���lرC�ށ�ܸ&�сl�*�9�q]6.�
Y��u���G�qZ7��d̬�D ��тy��D�H��� U]�2f�A�ʺ�. �W?���L��F�=���6�E �9�Ƞl�$Qp�z�<��t{L���A(�!;f�nS�"��;Fߦ�;"M_]��\�ͲC��ۘ蕧��U�ÿJ���»W���U0��􋮞"ᰫNevl�X��<�"/�Ќ�0E��.V|��2x�8��ש)�Sk��늽L>�-��=�a���WJ��]Ϧ�6��Bk(�U�����|T�k,Q�vGk�h�G�v_xA����]߲{~���黻�LU1�n%��H��j 1 �e#JJM��3�^˾���B�h��H�(�0���fw�>:[�)˗�g}X�/W&�ȸ@�2���2�2R�N �s0hD��Dpd�(mw��ݡAfq2Ǳ6�Q�U�ee�X�����W��C�5�*�q_��F�@�?
�jP����T�����x������A� d_����Q}�#����ZiKU qKɬ]�y}��My�o�w��My����g�O��e�dK�3�g������G~ �%ĸtؓZ�z���LON��=���{���'rҨo8hCE4�э}�s~��D*0�����Nt�]��'o���l�9'_���3�n]��l�8������}�k���w��/���y&��J����7_{����_;��]���-��F dAe�1��,��&mL���<X�:^��b'uYD�X�7��2zq�<�M೯��3@�j��Rs	�Đ���ˈ��5�$q%�X��Y��� ��F^<F�r��e	᭜�Q=��dk�S�/LV�� `둇��ܮ�?~�MY�:��qwz�\��=�f���(@��{ݽuK��-�)r��ȇe���l�nݐ���})��B�q9�vS�|�{�?:���KS��;r����Τ��tt�����Qݜ�yD�����r�/Ik�@P#��+7e�����W7�W��=�����ɯ^���d����RZJ<b��o����� ��\�5�&��.q�lJ���|����xD6���v	Z
vә�UY4s��ˎ.�a~7:A�,�d���>"u��1Ta�.o����P�*q0�q]4�Md�u}u .ѩC^�ȯ��q�%�wR�+��S��]��Q�<��q�<~��A���F�q� �ZY�A��ʠ@a�Έ��ڻ��ږu���N@S @0�B6�0���-D"lj�ULh�GRY� ���eq�C��v�(��l����"{>�:�A�6+��2m#wW�a�S�w󥕇Z�Z��iV�2�~��ג:ed>E6c�%J
31Tif����YO4�^�xAy{%�U���tS�V�e_����]�c�̺��1,ȳ*k3���<��%��ˆ��J�$�TP��e_�����D��O~�3�яR���Sr��9.OX��,���AB��kW�ȟ����{�yN����,��G�.G�F��ܢnWWf�����{���	�,y2MAJ���xO�<`k"L�q&���L���uT!W@��@�.��P���(~���Rp;:�N�$ڿ��s�����|�;[W�z��|���|�������'/.���}�E|o�Nz-_���7��|���?���o���O���쎆�껐u���l�z%"�
)ۈFl�;60�Z�-h�[�D�zn�9)��j���pHrk�2Tx0mJ�ѕ��QZ�v}'��ꊙ�.�X
������"FlqddǠ��&8���Y����ЊH��G���RtaW.�9���#{���h*IW�ㄵ�v�H��b;/�ޯ�+o�����p��[��xG�|�������6�����ܻ{(ë�X�4Z�&
�nߓ�x,۽7˫�}_�
p����h,�/�-NhTW)�:��k��L��מ#�]�%��#�]�20T0���<d2�T�-�Ga��=��h^.���w�2�)��{}ٺ�>���S�z�~I�(��UBX*�4�Y����2M�Ȁ�u�XiIߧ�QGN%�<���#�~f�i��p��k��ELH�tlb:6M�P���g ��j�g:6<w�bۅҜ�Zy��}�.`ڋ���z�ͪ:
:�M�4&K��	��W��b����gw�}��$��1W�\l�G]{�%� s��I�'hޔ�Kx0�%��p���1-����((���-�\�~�L�\\;ر=�<���������P��_�J��hL11tH/#�V%�����d��!3 ��3&�Ҷ�zD���L�������l�ƃ���nSB7��������t�a/N�py���� L;�Q2�N���J^A-���i���ؐ]����s
J�ɫ��(�����>�itm�8�����nݾ-�?��������_���=��AY\3jE��Ƙ�L��9էA2�8��JC}��bo�.�?ɼ�8>�C�Lt73���,ttt��QE�à�H�DO���)�2��,�H��Ҿ���t&w4r>�q]7�L���FQ�������?�}�����'��n����Z��b'���;?����^�un��NG�N4�������C��,�ɾ�-�-�w����%{�+z�@�626l�����%�͙�$ŭ��� ��/�Q�k��w��+D�W1m^O[��w8��%	�0H�S3�J�0)�+�#�k)r�o�c�9�Υ���\��Oɨ�-7�r�;/���{�����u���4���z�׽�%ȯ o��X����
7�4,�
"�,�y�Q�\r���f��&@�^ح�#ٻqWf{2�̥}8���@AQ�%�j��W��}y��M��]|@2}�#ݬ��pFߣ�;��d�rY2�L�ɧ̼X���J��I�����>��c�k��}qWzO<"��C�$���#t2 �Ng���pN�s��x�š46�ְ��� ʮ��+�aC&�����Q�"�E�=���Le�4+��&RQ��O�����w�XfR��Y�r��y�M�G~4���qE~������ْ�O滒�w#�x_��U��tHˌ�!��e>v��#}���r���O��<H�|�M���ZG��>{���n����"���ݦ�r�[��Z9f�̉,˝4[�}$M-3P����Fj=c̊�k㣄�)�AQ;�+�-����	�W��̧R��'l�U1`"�N���Yfܻ��^ۺ$������o�wG&+�2��³+r6�$�����佢�5�@h/�BA����̑e�MF�z�y�ߖW��-��G>��4^�ϝ;w��7ߐW_]�鞲\ ۢ��Ɛ�K��T߫�]K��sφ��R���2�|Y�I����� �l�9׉R���;ֺ ��'� jU&�\�����%Y椲L�r4�G�2��j�Q�ng˪��+�Ţ=����(�'5Uku�+4�����ҙ]ϧzF2����DںQ�e�H��-�`e��-;�(�W[*�G�G�I��/�Q�l&ɲo�y6+q�ߪ&�*��	EekʼhDi��jЁA-�A�LEG���Y���)�
�E��ĥ`�����\�����ka�"��yY�����:#��3�h
0
���5��_�{P����y����l��G���I�чe��#=��wve����o}On�ٗ~�/g�H������%}��LN��@7��+���sJ�|'z���x\�\�QO������Wez����O���)�e��#�r4�t6�Aw�ܪ��{2P�
-�Qú���`&�&a��g/�&�o[C���B��R�$;�%��3"�ω�l��h�\x��m�Z��Ĩ���b���F�@����;
:C�5n����sr�Ɲ�ʯ^&�}�DZ4ˋU�p��|���\Ȯ�XuݘR�&8x�l�A�ٙPv���o��38�tu� ?�J��$�ML����$�]�_s�"�!�[+��v�5�.6�u��8T+�b�����ߖ��Y����w��5��]z���1^Y����,� +��j��D���%�'�@�)!9�`��gbMp�L���~C�F1B85MĮ��� �4}��y.� n���+��5[iڸ��Zk6�j��P���X�C���v�7 qf�MCd6𕻓<8.���/N�޽=9�:����M0��V���^����\�[�*�"֪�`��Y~p�ү��P�z�5e��u����K/����Cvy��2����9��6xw�"�ߗ������S��ʒ�y{��������w�4��T.��/y����W�{�c�xς�X�0��Dà�Y���Ct��d�"������R/5b�*��$�U�wC�DW�x��D~��~~���� E'F
��"�}2�ā�r�� �:�}CK �E)��f')�=�N�E�".��c�L�r��&yX*���[��$�������d7Di���:P
eTK��]�QC�R���!��#���em�Щ�!��>�(="��u<��g1��c�l���r� �?�`�Dv<��B�a�q�u�Q�#����s��̮_�}d&�o��ND6dw{K.>񨴟���E�-]� �mt�#��t�y�K��M�-g�_.=��D����6�\z�>�����oʍ�#��|����OJA¦�np7������d�wd����<��������X���7����IFD[$�#�%5m�U���s"�Ĉ�S >��gXꦶ`��dp���xD�~P����T�
� 0��. `�4���KE'ފ*�U�:�W	Z4n��5��Ӹ&���x0�F�,�|�/n��ݯW��
0���X�����'�L=ب$�!�	����>B G5���bW,�kL`4��	щqY����k���]�-9��K�"j�I|?wSN��5I|@p;h�7#�+��0B~ȃ �V�
|� ��O�ݻu�-��kĄ9h�/"�FK�++˒4|()���J���{��.��AJD�R��5�@��\�Q��Ў���SLR���O+�/�VW�5������hH�j����PE�b�A 24̪����L�11�ɚ�hi��(���#/��^��1���������4���;��cC��;u[[,#/����cu�����Q�����n��G��ڵ���k�!���"�6�F�A 8m�|�u�������/O�ם$�B��^����:� (�dV���R΍����2�Xk0�3�[��'�w|,�XhW�Zb	TF��D�B�F��v�D�  ��|�u��hA�7�Y�=̏]�K�'�/���bmyl�(d�t����F�ы�@���B�lSke���A�ti<  �N0O���g%����<#R�6f���C��#�2�C�p!����qݒ�S1��P߅��V���z=�Pl�TԒP���j���C�ْ�=%��{�����+�ؗ��]9������{�w<#����}J��(��/���e����N�������轖Rn�H��������r&\�OF 	x�a��1t���5���#�������D6�қ��!����^��7%^LeW���"��M�A?4 m�ץ�	3��ȁ�yA-�R#phZ��,�~J�> 2����K��cgW� �)���2#J�<��Q����>�X-B4_xT������o�f��3qr%��0ۂ� ޣ��p^E�.JßX;p�d����t����p�v\�=����^��I�-����JmS�"�2΅ī��2�֦Krfm%���P�k����I8����;^du��"�$QG���)�a��Y����e���1�"�"v��)��JV"}"HbI,�E�̢�@-�n�w�;����c�Y�(vN[�����A��ǕX�{�WW���ϻy�1� �4K4 �%�`hC
Ůb�c-~J�-"�Iw7H� �]�� `���y۾��_�<'��UoHI��������n]��̓�'O�cЧo���llg�� p7e:�(K�%P���E~In���u̲�s��7�ñ`��l?M�Σj /A�
�~~в�1�"�ffP��@�UX���"�*S�{�^����1�E�8�"����¼>�);%�/j 0
� ����x+b��ФJ���VM�]�%�	j����].�~��[�s�}�hn@��$7&�����.o;i�M��!��m,sD��� 9bG�Xo�H��.�*��H����Q�g�|��g��.�}�e��ڜ1�£.ܕ9�����@�3CQ�P\���0TA��%;��G)�h� ���|p\��!��+c�341���Jೈ��-�m����Oŭ���L��AP��F=}��Fm�'�ԴG"$r��
���1�sߢ�����{�7��)�bid�A���@��xDUC޳�,-ɑ�cĶ�y[v6n�)���!��=�$�!��	���ٖ�/h����P5eY^x2��jzε��Q�ZȖ�"��6�R�0�~���x��0���VG�[C��P&{rd�e�[dbP���J����dG�5��<��u|���M5{sR9�&��G,�����i�~`��y8�J=����!����ϔq2F��Hr���42�pS�jĸO�Yh�$1��"�"ٖ��24���c���B�,��uN��1���yy/A�f�p�=��3�`�-۠#�e���y��1�s�6)&$�F��U���cŲ�Q �I䜜�����(���9
���M�w�.�p�T`ÿ)�$���T�u�s�X.w_��z��6a ��lmԜ���4v�p���ږ���^�t�n�����:(gۨ��M�R7�L��<.�T�A!�F|H����ih�T̎95ɏ���3Q��l�%�#S�c�Ƕn����/�δdJ�.3�z�!j� �>�Qd��gDV	Zؒ�� 
���Ik�r�I��8-|<6�bC��>9�H!���gv�b�Pֿי��T:
���ZL�>{7�$��ػV�vË��'�o��<�?�0=�!����'�����'�S��7�o���ֻ:��c��SѨ��{R��H{iQ����"���<��#;[�%�&���ǀHA?s��Q�z*#-�!4�ID�X�EH�3�D�� ����2H�\�]v����:�]T�E���ܐ�:�b{�Y&8�j� ���C=�Lc�<��W��P#���/K9����p������F\ �����Ad �7PJ�UgT��J���j2��qB��J`NOF����έP�7����M��*C~�òq���	� �-HG�)[�eq^"��B�a.{��R�����W����ăe=�Ӳ�Aj��3i�}ھ�%�o��'�uG��=�n����o����M���m?��沂!i���^��ss�� �%Ḁf� �}�yEz��  �5d:3�
�Μ`���#L��l��].wN �12ށs�H�ڋ<��p�J��H�#RD�<,;� w9�ш �Z1C�h6eO&`�e���$��$�,OgG�M <ޘ�l�ʒ�rKA)�-��<�O���٘��Y��9I�W��ZBt�S��*U�ц�`�%Q}6�5L��x���ƬXb��2�I���̠q�
rNj��l�S��1��g��z�ifP��$3ۣ8-�8Ш�\#���e��z�(A�H�&�G�0X5/1� 6I�xx]�Z��c[p�ֆs�j���-����,��`�H�f�N��� d�B�0(4�~�^����1�b�
��zL�@H.=�L���Ԇl&����A����՗�yNUH����OkG
�3??��Ž���G}~�|gޮ�~mll0���2:
����0=��0M=�^:J��@F�����J�˒#��#/��4��}M��%�g�d���]�X�mZP��jV�8�?R�V]\�_�L���Ot�=�P�uBޣX�@�%+52��h����es�?P^z�moH���ٝ��S�z���l�J0�``J2�X�6�b�w5D�h!a��cX/� %C)�9�c2�伋E�#2���#�L���t��)���9 #	M��Z)�μ+��dtBi��8�x���!6���{�j����,��[M5nʨ`m�4f�&�x}�aP8�U���\D��Hڡ� 1����C��r����2#!�!]�B��=�֞�8Bj��]Aˆ��]+��hn����Ӳz����r�۷��������(ZX␶u��-�^�.�;ے�=���om��g��U�6�:zܾ#�+�%��W𦟧@���/��ʲ4�����o}Snݒ�^˞��݋We�g���*#M�^Rp�IC��	��qQp�GqT��Q)���܊8��A��S� �����G��vH�vCA�e�<b�������8�&Eʒ�l���$e��8t\`=����+$��#���Q��r9��.�r��tl�V� �	�vF��#8,�Z�W���Dbw��\w� :��s8�<�d��턥 �@��W�,^W�5�yq8� W�`@:��;z��=+��a�b]f�-�1mܦГL�[��?0�Z�sM�p�	:g!f$و�އR�`l�!���2m����8w�3~�6
�
2z<�$�	��Z���L�/5+�p����Y����5������n��G	 ��{�1�t���V�V�@a�\���2���g�Ǒ��-)Up�EV���!��u6�Z��L�ú�T#����]�xN8?L���(��5�lF'��1�v�LC"1�	?���A!���_u}�V�=M�$a�P��1��Y�Vj�3�W��K(E��Ɉ�ֲݚ&(hM�$ram���]_�|�� K���,!��L�{݂�R4P9�T�ZL�8gM�M��!�6�Ke T
�e��>�vJ)hDXQa���	KP��9��k43��E���:�z�'���]OiC�-����?�T3�<-��[����R�L[1}���~����`# ���/�ÃRR$hL)�|RD�W����8EF�0�̜�k0���N��
��xʟ������=be)���{95�KX���:]��l���Ӂ����uFd~N>"��֥wm���{o_�-O<)���e�T��ۍ��Ƌ�Q}w^�}C�Y��5yA��s����dY��Mm�H� 'R�uT�9o<�uپs�k��^�&�������r���e{����A4wkCVGy���Gjt��7�6b�GUe����M��bS�-8��ʒxB����8sV���Q���'��4�/ᚋ�e�����-��܋(*��V]�Lg�w� �8O���E�  ��1N��9�Z�J�� ��5j���Q?�j��cmOB�1���,A�_#t��{����<�z�Zm���A_��k�ʹ+�ھ ���C�+K�6ɘC�	�e ?
8���#F�: #Ga8,��%B��4���x�Gf�8��wp�������O&`�5���'>ΑC�t�ݽ.�� W:w8Q����H��z9��L���c[\\,�����D�;"�l�Z�kT��T�vn�$���9��'�r斁Q�Mpm%uS�f@����f՛��8W ���.A�<⾴ -ڕAj���z�h�/lq�s�T��w�sd��:Y�i���yc (�ȤE��1�����'���i���#3�P�3���hI���yQ� ��YP��T{/�]ٻxE��GzD {����B���gHaU+d7����x{Â�8f�5J!H�UIP��ĀZn=2�V��TAR���e�Ψ���Я3Ң�~��e3�i��(�먂tk6%�*��K�׌`	�T��v�<s2[�J��`��):�8�F�?Z��A�u��8u4��Ń1��b��QL���p��	uJHt�FMEɑ�˚?����K���̊x��T'��C,=y�,�0�Ri2�GN���&9 ��e�ZkN�$��D����ݐ;W��hiE&���&A{,7.]���*��YE���i��FX�`�"��V�lmK��!5��r[#���j2VC����l5� @dOҼ�Sb����`ZA�F<�fAw"B��o�\(��3����"�k�2��8g��� ��.���*�W�� ��FWt����U�b�mM~�
�A�y8�v�S:+�c��͙�hg�8D�|�F$M�.�g�/8S|w�$����u��UG��׷�xP�DJά�9���2�L�0��\\Z�~�Tp��2�K����:2� ���k�?dg��8v��_�������\g8N���pK/�8q`�`׃�õ�ﳥ%��C���'�����ɰ<FSҮ������%����?��,����<\��u���2�`80AF ����hv��S>�m��S�By@��L�6x/3�@/���X�F�.I�}֙���y��Q	+p�_î"˒E�tH֊>�=�@� �Lj�h��O��f�Rg�(��&A���𻃊�[�֙���a���6�L6	�w�զ�A�`\!v�/���wv$�d�<"�a�%����pmq�� �-��A \���������y*p���&��CRaK3r.(a�i_?X�>Ҟ�6�R�齀/��31@u�(�+�5G�=���@��d  �L��� e�X��&Lc�[w��o�ۇD�0�������1�h�5C]����T�JR��PPS��0��8Kˈ��`��F���>�5Kl�mZ�����Ad�msf|�R��]�pf�hX�8v��]q@1��V�qP��q��H�#��]:v�Z?,GO��5�j��P�7��d�uK���P����o������$�oɸ ݫ�������.���h��~�y�A)�eW�>��l�|A&;]YZ���<"�����j{/�&�ϝgD��DI����IP#��[\��n���H B�,��ˉ�����F�s�.:�b�C�+���p�4S�5�o�CW��.xEg +6�4�c���w=8��^{M�߄N���;K���ERc��)"=���`����CC�'��!����NN�֭[�:t���`�m���`~���مr��U�_�=*Ǐ�`tm�F��v/Q]]{��ܼu�\�����}��.�0���&�'�����g�M8o\�� F�%R��
<�s��l6f�$���l���֌�AzWG� �?��Y"��7���rr��M<��� ��,�QE]����x����{)����v��+	�+)�OM@y��tb��<�ך�)BK�L�K(}�c���a��M������7�~�?�-y�����i�u�e�w@��x��h�,��{�{Szt������p��� 泀��6��bt�����w��Jg^mmU�=�_%�� ���I
k��<4�E�;�a6���W�E�U��T��T��2��kB�e2�ŉ��Q���ܞ�FD��H�7�0&�{a$& tH�������4�k0�U*�1Ȯԛ�"�$AZw���&k5��'���ˎ���#��ɓ�a�3��iL�g�s�&5A,��(#S��� ���"	v�ϋ�a� �(W��F�%�(OI]�L)EJ����GS���-b5�((��#��m���y�3m�e���rk%% ,�n%�B��H��g'W�v��B��>�2H�-;*���9򮷋�s��;﹥��)�yY?��3�|��q����9u\d��l���u���MW6w���!y�co��w<*�4/��RWg����Ɲm��X��t���t�6ԭږ�;=ٺ|�@uA��	�6$2�d@�7H��[ͱ��
x-�$�H��Dv�4;�`d�1̓PR�,�����*���������Ǧ��J������w�w'���zǆ�C�N�����=��=�������?g�9$A���ǋ/����߲܁��g |�d��� \��^~. �M��σ}���_��\�|YΝ;'����+����N�1������:�����җ�${Q?����}��}1I&\ �(�y��@D�q]p�VVVdM��,��A��Gφx�q�<�䓼Fx���\x� �3ǎ�����.�;��N���8v|�����-�ǎcėg�(��=��#rZן�I/a�g�#���^��Qf;s�����ـi:�A��L^��d7Yl�u_�.�7ͤ�!�rU^U�NG����C����6;^j�%�ܺ)@����Tw=��ڟ��g�F x�76�YD>t�Y�C�Pl#Q
IK{yxa�ۈ�6��G�u}��lo�0� ��(H�C�
��F�Aa�Y�~:q~R�)�EQ���V8z������{��$#8��.���Z�0=�tb%��Il
�0�ј�o�ٕ�%Wkjx��WTٽ��I�X|��Շ�u0��Fx�  � �O'�z'Z�˖��Z5Aڝ0�)��G�Ϙ�Աe�ru���EH����#6� >���Y����0��ll�RBC��K}���zi��Q��wN�%�0�jH`+���M���J.F	ڈ�,�"�7r
#�zh�Wmv,P|)�'��������t֎�ɑ�ܧ���l�uC����?��}���x�Ei$u��ѵ���"�f]�Ϟ��K����Yj5d�ѷ�뎐{#�rL�{��u�v�l��;K"�+6��7kR[8$��v�k�%(�B�*�Ŷ�	���9�6T��s�8�.�#Gض��PC�F��$YY���W�H�R5�Ea���̶�bs��QH+L4Gd��/|A����XU|G��[�RE.'O%��ܽg��2J�r̈́eT��r�]f�����3�zJ����$alpī���f�w��@/����=�G���aI�l�E9�Yk�l;�m�sϞ��}�/��矗�zH��ɻ��vD�#�v]�`D�1a#���_������\# .�O�Q�t�����m�"�t�5����D~�w~����_cl�#2 v������������.��&�@F'�k�(���?�#�˿�Kf;p����k�g������ʐ��(FL7�ux ���{.�vQ������ѳ7�7~o��'���?���K��K
�;�K��Cg �+��"���!.\������/������& �e� be��� |�� 8�46X�Zn�ѡe:/˞��}���l�VЀ����sP��:�H���E8o���>��������I���
|C���6��6�I���m�i�1�B�����#ݨUlLd�E��[k8��Ȫ ��'f�Ui��qO��N��A�_sV��{�>@�}�=`��	e�������}2�݊�6�oX��_��aO0�&��|�WԦR,�mD�,5$&Q�y��;��C����h���W�R#�+Q'f
���ʬm�|�6>tX`52Xbj�&0�Y|8Y���ȺQ���z��b��$4�q�Ր0;$��
�A� N����g86�#�
!Jec�;(Id�C�,;��;&wރ�xB9���#)952�/��fz���K�Cj�y�1��Q)w���U>�(i!��{��εlD3�T���2�..Iga�m����,c3�l� ��cFZ�w4�����9��<�p]y 嬭�Ikn��=��u�������EQҐ|,�k�?���ET��h&���k��6�jd�W/h�Ր#�ze��T�´�	�w;U���g!��)s�O�]���;w��,0K�(^Z`-]�JK�ZGÒ�i�&�l�&$D��֠�s�}�ɫ��ʌ�����?� �0�x�������5��x��s9? (
$�F�z��6#!�V��c�}�{�5�!�H:����>ǇL@~F���R��p	���� �� � 3���؟g]��=��\��^�8py�t�k�lL��x��}�l�L��L����L[�"�}^q-q�L ��~��r�0ދc@�u�����vk�x,!�R��U26�u�,��~�,K�� k�%���9?*.�Z�6M䜭�k�e�Uڕ�}��<�~(�~50(r�D� '�� ��/�jsZ���$������k�63���G��C�0�n�@&յ�����@�Q��� 9C�(���1#���S5�9��XYH@�O�۫��5p�i0j9G��p^��'��
�5eږ���V�N>�C)�%�@]�p
Щ@Y��T�X�z�bB�W�A�M���'���x[��D�*�5a�FÚZD��:n� ;�W�9(�<
 �Ήu��wBu�I��Z��0� E65�[�>2�6��Y���/�2�v�`@X�[>�������dZ+v%a�M$�F�Ǖ������ar��n��җ��*�
��1���`�MD��m<��D���9Aز ���zaT����hD�Ƙ�i]����&���=ٿzK�ΎH�f�"�5{�Rj��ɲ����j��Y����a��_xY�W��|�(n([^��jr��e��/{�\��K�jZ��k>
5�@�c���]N���~�� �b��rupJ�xQC�t� ��X����}qy/�h��+s�h��YpL�~HhݍC9�|����g�gIᥗ^��W�ʣo{�����s:�K�.щ:!����ӂC���?��r�8'N�(ɠ tdY^��>��< ���7䉯|������g��>�y'K
^��1;��k�� f-t� X*mL���vK������� ~~�aY;r��^��%�� ,�oL�ű�)hd�^H�c��?��s� �]�~�@������<g\#'��9r2��;�	\��x��Gy��sK[ >m��_���?��Ǆr����Ϙ�k ���o������\q8&\{��� �.<�8W%?���v��r�����'~��-y�[�ȿ���H�	� ������{cfI�׎0�am��p�w���G<pJl�S����I$(��&	Ӿ#K�Ru�e)�״�0�ٰ��\�0D��,O6�&[[;�{gK�X��
�nx搭�����fM@�<��l��N+E�0�֫��Y��kX�K�5T5Dm4�	6��l���*���>��@?@�¢fۓF /
Zr�9Ѵ{�M��!��<���"�C�����;ބPZ�e�Fe{8R�Ĥ�f��|�[��:*�`�5�lE�q��b�i��6O<CR��XksD��4�c�Hr�A*6��$<(q`�c��s��R#�B���$8y8�@D�"�~�.�e+�@��wŢ=�5��Tύd����~5Q���C��]��H���!�2�հ,�]9"��E1-JX$�3�2��S���>Y����6��G�<����k�s�&�By���a��//˺~�,)�-�WoJ_�j�2Md��Kru�iY��}|��U{
Jn<���nm+�i&r��<����2���3����MY ph��F�p6_~U�}�o�K[��C.6�Y�K(0�U�Q�Fļ+Eרsу�k��@ϫrhEZG���	��5���,�����8�f�TS�6�=�Xx$�6w �1����
8����}��\V�V�z8X����I�I x�����ȟ�ٟѹ����8����J��KE?2
oy�[��19{������.3>��������G��8�u�Й�+�`�/y*��L~�l�%�u����O�?��_~Y����� <90��R�3~��g>�������g��A�oN�uN�P�����������ɯ�����?�o��Ń��@e�����x&ųIޥ��\/������{\�{�`���R9��+^�����o��y���������lg�������~���/��/�����k�Ar�3K��5�u�2tG���L��߻�f���w�N�d񐝍-k��){�X�%̚2��aM@��*hP�[G2�{b��h��E	��@K��v��A�@a�Ó�cBEl��5EM��(LbB�b3y��<8{~�+Ȁ���M�P�&g�ɐ$���hp�yP?F���?�3� !f�2$�nڅ~���Ө6�mqo��	^��W|���v-���Ҡ��-}<�A�;�#7 
2�c�����N�j�%�E�,R��S�~k����|���)|��Ng� 2�3/��ft�Z�~nG���}`�é������������\l|j�����4�+L��]m�yv�!�;�v��O�S
�O�j��H:-� gT��63/3Q~\1.JZY[�O�
�H���ˠӱ&&�d�X�*�$�<l	�X���#�U��{]K9�I��t�L77��/?��I#��$sm���o���4�>�qyE�Wnȥ�k���-��N�ZȆ:���_��nW��[��[�]���w$AIC����m9����ޫnO�~��u{W��Z����Ci�`@m������#R��N��~�ת<�h�%z�������xź�����Y�x�cS��ʹH�n��˳-�&ܦF��.��":Gۇ>�!F�^�)3n"e�>��v��������zV��䭏��_�����[w� �Q�y�8�^�@����l�Fv�xa��-�;��7���|� ��B�<���t������A��m��ҕ���?�'��<P��WIZ�;X��λ|�|�Uf]��{���gN��9
)y'�:������_�"p�����/���^� D��mo�ӧO�}z�Y����4��:�yP�Cv���l���
�_~�efB?�*py\�9w��A'�z��|��s;s�����<��3�����?ο�

z��t<�t��k����,��Ϡbl*̡+���Oo�gY	�d���[�g��s<�P^�=����'�.���/(%V����rmE��Q :��<#QB���`��2=�9	Ԋ+A���@�'0��Cnc��V��Nl��G��hcz<?�LTV�c8�1g9�C�D�29��� ^E�����'�� F�����7$x�V�U�Y\�$P �	�p�� ¤�>ػ��$��5�*�G�3E����fT���`%��|`�q�e�;��S��U��0�W�0�2h�)�fD56�DV˭��dO$/�gI���F��1ZegI�x��p�,��� ����q�d����%ȉ�0"�cPAE�Yg�xF�1*�I���(�8qVQl��@�V5Ù��,�$L�)�c��4��0�jDR_E��D
�#��;����`l�#Muu�0
��7e���RU�q8�����HA�H��(��`O��1���m��*c"s��@Gd�#�F�wvt]���˄����u�;�.�}�i�w6%��)��m^hU)oI�"�<���#�: �� �VS4��zh=,kgϘ��^������d<J�mA�cgQ1.��ԑ������ɻ0�dW�
����h�[�g5I�w؏s��@T.��,��9؝%Jb��4��o(�N��Ƶ@��zVF�
�"X�����Y�9��!�@�uِY�s�6?��_�� ��T�͵K@dwҪg�?</~�e�! ��J��� �@�@�����3��c��goS��F28�����׻� VP���+痰g�e��s�|�;�
4qк:��}�/'�ߑ��~q�(�����Y���:?�.�[�^O��]O��ސ���ܴh��jKyq�~��6��ն�2�����7��D���?��X��α�ۋ�@�U8�����g��&k��ȂȻ �k�CP#�K��-0�Y2�i�0#���HdhFC�4,]��bZv�^!�]U�J�!��V.�5O��0��3��šԏ8�;"u߶�:��<{�_�Ʃ���h(�M�%���Q�4����И���rY	X� .�b"}D����5�Dvz#r9�A-�����F
<��\��&>���ij�����. `*�h��G�e�j���p�L7"���*J.IbN���3�g�gjh�u��D��4dS�ig �`00��A��1�[�jk!� `a:�L�=��b+�a+��� u^<��R��#n�P���a�*�64k��Z�Hgu�����@�ZE�ʁٹ���Y��q�Y���S𲿲({��y[Fc��y����ʒ��x�8� מ�wwG��,��ɉ�Y=$�Td��%y�K_��7��L��P�l@�sq�)�L'C��2W�u�p隁���Q_gO���$�b=Ba��z"D�ֲ>��[vt��l�%��7άK���V�Ċ�yVٖ��Y{�_F��t��UQ����!������d�VM�3�9��x[���]+�v�T�u�H�����R�}��@	�Ķ�ʌ���"�"��w��ЇeQ�ح�;,�}��$9��g��/���  ���'�;�*nb-�AY҆륖A�y�<@�O���A�� �5i�F����(l������_�qP��N$��dB�YB�m�8W����8�ʌ)�q�5ǀ�$��6yϼ೰�/|�$�"��������u����3N�{��,�J_�&�W��o� �C��n62�)ʤ/�{�[�8U��Π隵H���
�^c٨F/�~�@P��z���7w��NK% R��)w�zpL��aDWb-���Z�!|�s }�,d��uC��p@ �����s�S�@M|����,ԞE�"��"����N��tB�Y�%%`�Md�Lk�����|�����"�K�Lv���W�/Tح��R�ð��r�	j����s.�6גH�`\�?�䲸�2Dtw�Dôa�/Aa�Fhk�B;��LqV�Be�fsT�P��D�p>@�le�fL�%�Ç�c��bF�$rb�:��*t��!��d�@�2�������	�l�F#ɘ�iT�n�0z ��I���T�a���A�#jh��{J�����I@Bn1�J�9�l�Ȇ�U0ٕ#+e�В,�9#'}H�_�W�4�j�rC����.J�җS��o}Hԋ�t�
�ʛ7��p,�mn�θ+G�˱��]��i�smyA5�_yB�޾���/+�֌�H�*]�?�$+�-#��el�P�p�8S&2Eݾ����@v�l:wF��9̹�G]���JQ/x�&�1k�a$2;¸�%.�G�
s����ؚ���с䉌�k��r\�����k=�=[��o�rm�MT�)\�t����̇+��yMl��X�jp��L�e
���]�z[��t����?-����ʿ�O����R�&�s��X�Z��>�`V�[��E�y8f��q�؀2����[˥�] �;��ٻJ��/��"��|6�'�x���S#�5����Z�ol��8��	�zL���X�����~��������,�����o�:6���|fy-F��.�NO3+Vr1�K�����R	�Q��ց�XOgE�H�vwy^ ��Ӟ��Uv�")��:��B���p&"w=CDsSAG��˄�%7:��s�d�ef�\����c���y��Ah@�2I��n��u��QA��kB��P����:�.fC���Jp�ω7Y�Fo�3ooH��w��H�ՈE���˝71��w%��v����]S�k�2���4#��b�#m�В�N[:�,�`�"f��]ٗ���H6)��8�QC4��5#��p�!�3E��M5�:�``^Fy:�>k�Sɲ��p�f��J�VE|>�ʁ�����ssT�zK�Q4*�c�^�!zĂp�CÍ�N��,��v��������R>`p��B�:I(������&胖Ed����@��sޛDL=�ֱCr�o��G�9}��n�YT ڨ�$�ݺq[�����
8��ׁ���H�H��]�!r��m���RG�U�G���0:��]>"�m����!��g[�����YgY��xX�hztvMpR��Z�a�Y*	�c���ʑ��I������45Wc�6�P����i0��"����YIy�4���z�S��G�e����U��MwŁ�*Ȯ�Yqgr���98�s��uU�l)��w��=�V����P�2��VU���<��R�Ƭ���0[jepj�d;~\����,�X�l��������� ,Pa��F�L�����Px��� ���g�f��zl�!�k!|�
���k�z�ϔ���@J c��?>W	_Ȏx�S�=pXf<k���3����q� 3c��8��n�ח���{G��}p@{7P���(�S���tKp�Exm���+�F��Ra7�}��:��ڣL`��n_m������0�W �P�G��vc�Y[	YI>&����sT>O6Wβ-&�s�AL�&����3���)2���a�b�#dT��V{0��LE�`]`����}�ʈ�{�ʴ��bEQ��ø�X�� s��D�bY�{SooH�"�y c���!0C"<�hh��b�c@�c�Lx�P/�g��Y�����V��5I�X�4���8c�b������"�}�;��ޥz/x2htąi�8��f��� �0[�!������#��H��3f#�(�6��I��$ѣ l��H7���@M��q��g��E�h�npvl}7+	:^˂�5v��z2&����pX�)��'�L���lVAa6����N��@�F�~%����A`��^�CP\7#c����� �XY���'D�VD�-w�9ߒƱ��zB��D�K
Hl�C;����Z[?C�/�ɇj�G�{R�#lK�}�9��}��59|�:S5��;j���X"*�@-A6"��S���� y��z�$*��?vD��Qc�6o�+5\���]Q��}x�'�
���Lb�"�!rt�>��HO�>Mb)�h}^_?B��	�#��V8B�e�w����c	��)d�.�94�(�)��ꍰl"y�T!C8v�z]�XWآ���yz�������������k���	�^`2�{�s94���9��	�X8�/��<>���x�� ���PW� �2Z����H��n%��Y�9����YR.����
@�:?�?@ �.%8e|6��̡��p���q�b��B�iW���pOA�9o��(�S8�����ǻ�fe|�w��õ[2̔P.B�Y�"��<}�@��8���w;��w/og���$�{[�0{������&���F�d�Q?�f~\B	r�0��i���c����QNuQ�8cH�՟�j�z���^���0	\�Xbx(�g����r�D��
;�"]�M�m�O�`(��]9P�6�d�`f.��@�efӷQ�h�Ŷk�T�#���2ԜY6sL�7���@]0�a��q��x�X;2�zLfʇT�5Q6�D�[�HUX�����yM0\��7�ٙ���:vX��07�`w�uq�V���@�����(֖5R�rg]�����J=Js4�{��:���k�	v���׈�� jd��H	y���^�(�Z�K]\��IїF�Y(�;�yNrdi�������o���d�7�@�_-�Pך�y��.�X�C1�� �#0�h�e
�����m>���F�
�>��u�s���Cu�y�xe�ZmʌQM#����b�;����F��A�5��S���d���ܚ��0-�P����@b����ӎ���k7da�FA��p[�A�Ƹe� �Y_���.�q��79�hUׁ(0R+�S�\�$˂H�+�k����/�'�*�h���Ioސ
FN�L�r	S���r��3����5!�1v��T�V��#H�2/Ү���H��B��I�3��\;H��e�'׹#�-�g���qU:���4px�<�tG��Z{�,��� |���yD�/�3��
ۇ��A׃�;O�s&q=piXr���0"����0����C���ka�ӏ���=�����ןV����%1�m��>��$u|0�- !����?��?����ߗO~� $.��%d0�����s�������' ���AS8��D��E5� �F!K]���O�n, �>��_��'h�,�u�?��oLvA��
R�!��n)d�c��Ե�s������=G���O�|p����x�P�E�
��N�v����f7\o_c�hD֍�g�C� I fh��)ۡ_V���(�Ĳ�T�m�ƛ3[��xG c�FS^y�yY���>��רGUjt�n)@����蚊Z��{ ��[
hR}��;��N�Xgid���b��Y��S�0Q  ��P@�~z/O���/�F� ����{;�
>��R�W鞮�7
,w�t F�6GU܃��
���>%�2ÞLl �0L���G5͢DQ[
��&�ސ'����/�]?����[����i�z�$0�w��H�E��5%��( YTGr��Q*��+z�����'eW�8/0�`���0�������I;͹\�S���(n���j��N��"��ؐ������y]#|c�[#q��p2r�r��[
 ����D5��(j��|��>��4X����.{���9D�}H0����jJ��W��arM�������� �������u�b��i�B@Y
N*S�Y�B;������v�%UHJ�+CQ�& F�c�L{��8P����܈r�21��3�bA�	m���d��0�W�ykK:+U��KGD���
���'Ѡ/mԂ���y�U�{�I���H��JTv�l^xQҭ۲�F������HC�w`!�p{[��We	�T��w�F�=�_���OAXw,5�u�?uUj	��� o*���_��� �=���,?
�5A��z@q�`��I�J!:�i����t��]m�����{�o1�y�i��CB�8��88g�X`_�.�y.�[��J%ڒ�2�m�!����^��񴛍�k�M<ӑ2�(*�pyB��g0|�b�O2I��+'�{�<�dʥ`�"p�B�͛��}�,�g\�$�����z�|��$��/�I�I@ϻ1��r��6�y龐]y�/���F�}�o������|�+_&������!�ָr.�V�Z`�26�&��8��w�xg}߹{	�p��{�urG�%��s�mp:��i ��K�R������ kFp毫羾���� @�����n�ȍ[Wd��fYWT�=ֹV[�Rk���۲��%G#�אaぉ�"�;�~��7T۽;�I-3��rO�{��`cyAZ�5��&E�)��{8�e[��5�5=�Gπ@���61��Ϝ�S�O�j�>}.�ҽ}C�����d��`�����]��՟z�P�E��2d_��q,B��ױ����ĕԨ<o��	^�E��		��	�MZ��8(b�_W���AW���e�Hj�4�<��F�FI}}(n)*��xCA��=��'�8��w�z���������K
d�9�YQz��A�a"oYh�X��_nh�߆a�E7��fM�{d�������Xw����ԥ������� �j��Ƣ�@���{'S�0"UY�j��voc���x(Y�i��xOf��2eK=���+p��}ٿ�/�w�hD�\A%r�5OR4�JM�а ���4���k07�&/D�`��5E[22&���h�� G	�1��ٕjĴi�Tˤ����7���Z
�*2��ʵ�^��q"�4�HVV��
�ve����/Ik�lQUF���ӟ�9�أ�td]���۷�w��,�/Jz0��k�ȵ��"�H�p
:��97-|��HO�'iO�mT�U��A�-�Ҽ��2�b����2�.�=�jPc����c'���D�����% )��1���k,�'޺���"l��ڇ����w��ѳ�����# yl>+�z�}�^FkxGIA钸��%�@h�c����EzV�l��<Y*�M���b�`
k ���@6���̖�pp�p�8_�᠌��Dp�,����q�*� �����Z9[�?cV��K@$E����vw�=�)	��+��0��.�W$�>�����:h� ����A#�C/e#ދ�y�tic#k�vB�ϰ�,��Cf��5��Rٙƫ�<g5�`n��>3��#�r��w�&O�hi5oC1q�(Q&[��F�T�C�"�}�6�/.�K��u�  !�F���q�&W�+	�m5�HW_�RoM�]U��9|HAKM2��Wo��׮˶�{�!Ǹ@�#h ����sg<������ܑ���r�겜}�Q�Y�!��Io�׸ݡ
� Kow �q�d$�&q��_�i)ֈ�B�X��q:���m���[$��k�?����؉:1�xk���V@R��Ψ�ؖt�%�'O�"ɥ����֦��u`���륺�1<�n�~����y���d�Don���C�l�?�<��7�n_�qtwo���6n�p�R����|'�c�|$�4�tĨ2��#�u�a)�2#�!���Rpw����T���'1����45@F)�?걔��52#���'��$5kq�l�j41��l�[��Ðtո*���ؒW/�*�._��$2.�3Y[]���'d��)i,,jd1���u�뵜Wg}���ʂ>���A�2�hO#Q5<�������HH�_�.W_8/=}�!���8/'��CGV�F�E,��Kl�Ɔ\W�����15�� m�Q:�y].}�kҿ��F��J{^�
4��ܐ[�T�H���]�~W�۲�j�h:d�߼-�0�YK0�-�Rcg����yO4���eA�[U�b���ժ�%�Jp�*əF�	�
�]�z'�0��9+2�D02�4���KX���LA��LK��KB+��!@F�K�5TX�`��\/��e�Q�l>�S@d�*�����Rّ"�Vl�pq��e-��]���"G?�,��Z8��Rj�*�{�2�qg����3��r?O���]�Q��
`0�N����+3���O��3�~��|�k_�O}�S<G}�d�� ��S��L85���P#FF���aNy�uE�2�����8�� q�\�%�B}�+_�1r�~�����A�� ����� ��4lϤx���K|w � ���q~�g��lT��־�T��7�.�`�X��x��~��\]���KJ]��~ܪ��XTl`("ëE�� ��v�8eG�D��H�FnT�JN�e��+,d_�4�#�zS�ǃj#r��M���3�=��GRi4Y�6�	3%ˋR�ޑ=l;�#ά����srjqI˺��e���|�� ]b(O%B^d)y��atv��'a������'i����%�a���)E��[�.�>��	ՉV��CԿ�"=u�]]��7��u|C}��^tgxe���g�y��߻��|~8lv?�O���ǃ�[�;����_��S������Z�-���㢈��V@���P��8����
ۢH�� 3�3��C?�4D[���M���ܦ��|�K���M��iV�2�x�C[v2!����%R��0�w�ƣ�rM^�h��F;[�
J�t0�2�㹥�x��eyW�.'�Ʃ`��+���W.��C�rZ�i��(;��&�;[2�ڗ���Ζ4�uYC�PRS��+/����^�a2T�#Ӵ	�4�P#�B��.��mm�p�AB�rQ6 -�{rD�,dq��DV��s{GF�6`5���]��~Z�P���$���Z75�B�A��n�5�P�\����WI��FF&�F������>� ����Y��� "ةK�Њ�;AP���Juc�@m��Nʮ�(�f\��XN����9��ݡ�Cp�����yPR�pûJ:Y�9��p䐏����-��W����/��/P�e��KB�L�D�i���߻�$�E���p�yyӻڮQZȧ��8 (� �HP'��W�n��6� '�Z-�ؑ9�� d�01��~��(�?{Mq�|(���[�|�w�@�Y��h�K6U�E��A�s��?]Q����϶os�kJ�5�:!�q=� 0qX��(�)�P"�l��>�g�C���7��G��]�пf���3yނ���;�8�f�c�fF���e)*�Eqh[��ҕJB�g�f�Y��y� _s~�qmP�'��}#������������U�0��D���d@3� �?���v]r��������R�g�5�݃]�g}�����{d��a�_�(�����@ǭ��ܸ�a�O�$ݗ���GΜQ{z\�t5�ە#G`�q^�	�{���(q���1	��ma���8���yu�e��v{Â�Lj
���d��� 0`���G'X��^!%�k+�]��/�*�B��ِ]5
�(�����c���w�}������;�ſ����� ����_��Ϝ�kW_y�|�R[~_u2^�6���S]68����t���P�Ў�ӫ5
��*Ǭ�	�����j���H'4Ε$�Ar<���Qi��)���2�"%ɓ�w��t~h'��E1Pc��9���/��{b��=$[\Q ���#i5���;�6:L��s��l����Q����ټzC���RW@k�1�s[�2�gTǽ�-��2�zU����r��c���뱌G2�}��Ii�1n�Шv�Ӳ#�����vgM���
���������=��`'�CWWQX�a��$�VP��}�Hf����WL�N�������5����/J
��\I.Sh�`l7h=`���1Y8��E�^Dk93X�<1A$f�e�Y����tc̖Rf����y	�KB����Bg� �5�n��[��m P�>f�V|�U�-����p0��3�<�ׅ(���E��,��Z����R�(� �.'�T���}&�Jz��\8:�
���%ߧ?C�H}?Gt��G��o~�� �G���I��S�jp\(�<{��?q\����yf] 4���5Af  �j��?{����(���ȹ8d� �P"�ǉ�~O ����ش�~y~���ﱗ���C{�뉃UCVh����=����lZrݗ,�Ͱ6d����^X��ϩ-��-1��%$�0�l���];�Ӈ�3�!�8�㌶(9���?�e��@�dzu����Y�����H	�}���U���SgenyE������o}�
ǧϜT�:��y��<�yC����+���t5��'�����"����h����@Yv?�(<gЯ�@ ��4]E&3"UQ�R��o��^�pP��TH�D�,
�����\���|G���䊀'��7Ց]ܼ#�=f���S����X\=�������O|�?�����������������\�����:��؆��p�h�5����f�Դ���a��A����A����WWt�}��=����ae���c�Q�"���!9gT��W�0��1�����-Y\X�'Z�uF&
��w�f����,��yA�<��9{5�
��.�(���J]��71�O�����-��ʭ;2�4h
v����W���,'T~�;��ѩ( E7W���H��l_�������5��YU���*�`T?�łm�U�.����ި����� 9$g��%a.	�y5��� ����#�z��HbD�?�ُ���[=w��a֌����/1a҈Di�G��G �LC˩��9���;��8����:��v�<۱�Ѽgq�Q ĻMf��l��f����Q�p1;����f���+A:��yY3�J�W1vN2tƀ�k]6S���υgi��6	�t>9@��Yp6K��>X��-��g���ձMBD�]$�� 8�_Y3��A`����g:j
Z�w>�ڕo�囎:d���C� �7�s�6�!���!9aw�|g:��u��Y��9Q������[n�x]v�>�+6�s�Wq<U4�k�\>����ˌ�85e�Y���z��ՠdU��
J�K�.�p�)�T�fDM40CWj%�\ϯ��E:�s�}l�/ʦ0�j���n������A�d]̓��������^9~��,Z�z ��=?���J��zN/W ��g>+�~���+�����)9�l�R�Vm�9P/܃"�)�~� �hc]�i>Ѩ~�@ߤ��T4�Ԋ�iTK�F$=����ǔ_uhl��ˠ˰ɍ�-�s��ο1�,����~Qy��?�) ��1�ȏ��ӿ���ǧvn�N����*0&<�Eৈ��Fe�$�:ᗬ+�6�ٙ���PZ��ҘPQ�f���������H��_��e���R��M�vٺ2rv��#��yp֬ f�@&m�d�*���N�{�ON�5e<ג��a�;s�}���oo�@AK��@�KAK�w�=���=�5��,�%��%5I�1��@u&)������it����R��F!�#�w��R>��%��(�zL�
�nv�r��r~Ƹ^�P����#u�}�g[�DZs�R��]��D�h�R��?���X^P�8&yB���)�L���
R�@�P#�BhU�az,� �FL�e���(�[:uJ�G�����L�~�m�-i�T}tV���ms@P:�@��m��sgdT��#��&�Y��Y�5�!!��*A��,�3,�4����tޒ���G�P*l^VQ�=�,A̔������"6n�<�V���@h�=7?v^������%�=���r�������lǳ^��2�0>���;Y��P����=����%�_h��C�Y��༱8^/�U���8�,�1��̙3� �~;P�엷R�����f\|:(���TT%�p��u��Y>��Ŵ�i��ivf�T�Q?/�_�`ڎ+����Q3`Ya�2���8K�R�٢ �.%t����1_�� ��&C��H�ȖŒ*���Z�!��܂H�>�]��cd�#y�{�!?���w��}���&�y�q�Q14�L�X8����і����u�=zP��S��מ��ԯ�d��{e]A��i�[f�kU͊� ddsc�u�M�b�'�w�˷�VM�ա�BY}�`#��n�%Ӈ��Y�	d�]�b���:n� V��ݽr�ĩ��o������ן����������g�������{;{Gڕ:�<"�b��Ğ�;��9F�ıd�=�#
w�p�������� 7)���t2n@=ꅁ�oosQ{�
6 ����3���#�C!�F�ŌJ���ڊ�זe����ܞ�d=Ie!�H��qi��Z!�2�_  9�jR{Eo��B�Tv1 M�I|U�J��%}���ݸ#�����-f���e��2�p��Ӳ��N���ҫ��u}]_w��QY=��yH�~"��4b�;�刾o��Y9t����w�e��5�������m9�tH�Q�Z=$c]#G�8�-.QȮ?�˅�Jt0�������v�d��%I7nɖ~-���\�j�ݾtj��ej�d�����L��F0�%�k�".Fk�w&���8t�9���Ƹ�k��7�/�x���/}�Kl����4a�=�2��ْ�����gy�i�쎈m�����lF���!���Deɢ�2@<�X�A��Yb�4ܸv$��ch����:��q �� 
Y�j8/�����0��\�YH��:)wV ��c�2_ �(5a��/��;�N�O;�p�fɳ.�����{o�S?�S�?84�.�c xB�	��������;��y�/�1��M"S���E�"&�_�v�����<)&e���<1e[�_����a�=C�����>���pN�s�J~K%bIƞ�F�K?p�P�G�晷��-Y���5�W��+��ch���2�L�`%��f�累6����P�������G���g���y�ڊz�5>�IP����ωjw��+���2����y����'�����R]�)���>e$j�����\�2�0z!rE̺��S6�v�X��h*���@��V��  T�k���*��zrG���O�����j�ſ~��}�o�g�l ���O|�7W���'�����u���kpSP�X{h`L�%�V׀a5a�n!>�3 %�"�M��!�6��#�8D3t
��k��j4-fPZ�ҨsE�{��}-�4�:�{��ۼ&��MY�:)���rZE2��R��^@�eqA�;s��+zR:&���o0�0v�ӕݗ/�޻�!�����;j<��-�a�(!���$k��(�Z�A����r�����I�j�oݑ�����</����)8@��Ⱥ~�9��C"k�Ywe��M�'M�8~V�+hz��!9��c�YY�����*/dG����cA+��nvtM5��{G�[�=/��nI� �3�. 	����e'�H��*��U�A�]  ¢%ҧ<�b�-�iF��)�2�u�}���90�p�� �8��3:b��s���(���G��!�c��+���Tvl�n��p@v�APN't�L��r�L%�鴠2�8��\M[k�n� ��'*y1\yf�啠���\J~�45[>�����|~�����׈�ϙ���e��H��w_���y�|�eeZ2����21��:yi�s�O�d��� �kb�$� �����5\xl3�<S^:���a�%Ӗw�,I�ʂ�[��5��*��R��%!'��$$�'a&���	5_X�)�wu����>���0�f�Y*]������{k��R��fG�z��RG'��B�����T��+(��m��?�������rh�0�-�������
�6@J�e=��<D�W_yI���?g+���s
���E�8YZ�x������Le&ǽ��7,x��LAzq�E�S����p�QGF$W�� auAެ5�'Y�����|�#W�����;��ُ��w��S�"���5h�4!�Ғj���UwL��� ª%�i4�_���D(G�N���a����@c��>w��T�+�0]�T��9[%���`�u�B���|N��EI���$����on�֋/���l�ܒ���ʉ��H�����������8�Gh�����P[՝;�r����ȡ�2���C���"{�n��j1R�`����ډ�"H���ɍ^��˗D.ޖ�{ ���\��-y=�k;r��+#�PνM����/��c�늴��@��M=�g��-YW�v��%9u�4������e�idf힢 M�/�!�����|�eIzꠇ�%���=*��5��Bd��(��#"K��m���u��5>tXDRr^,��O���(��J��i:�ۈ�)��d�A܄���+���0���3�z��2��:86� �	e�Yq�0Cf!�HB�	�_��<!t�8I�E� ���q�x�6�q��+ɴ�߽-�7��L5B��D�l� �怅���{�������0��t��:�ƅ�P�A��}/���@&��5d]����"d^�lc_�0����q�$q@�k�͵#�)���c�q��㠌�c�tG���Ҏs)��YΒ����Z�#�)6��rB�H����7���sp�����A�]W��:���ޜ3+k��4��l�`�쇱�1?�& ~���h��?�h�tt�yģ���c6��؍1�$c�e˚U�U�*�\9������^��L����I���H��s��g�}�����4�I��Nb��������P�z���D��z�L�EO ��Ia��^y�ԁ�{�����J���I3�pR��H/��}���Bյna��rq0SkZ�A�z�U�j��n�����P�����7�(����ɢ�/*G��~�U��scK6g<�x>c�9_���\u�M�����9~L^z�Ay��+2{�e��D��J<�g>/�0^�����rϋ		��x݂���V8��4�,�샰�P��"��T���&���Q&���r�/��]�����^:�r���S�xe[�I���t���*��)�ς�����ӂND�>�E\/K�3����2�b�����c�����,K�����m�+�A̎����	�t��|�@�VK��z��������WN��O>#O=���~�l�mKw�/3��*�&A�RzQ��. ȬQ�aU_թY�sPC/�G���f�)���?�O_�e9�ۖ���r�De�^�@�՞�����W��}�46֥�����=^.�6���u�r�\����]��q9s����p�!�+�����T6?��%[��H����sr�ŗdc{M�r�Z����e�<�&�T��X`����})�zA��k�3:k(�9���J�0�ן�;��[��7�4���*�v�n�V��'�y*V��VUX� ֹ�K_��5UA	���5�������Њk�ǔ�}Ǽ�.���+�k%�y0&P�?���ƛ�"{U��	�I-" a�.T��l.���
�����x���1�� �K�}{'�]@������~��,)���}��G�\ㇲcwjV���V�^J�|���\�ǽ�N��|�c�����r`5��W�*_��W�0�y���� LX~�
��_��_d����w�������O~��k#<���$����Qpe�.�3`���/��/��̇�|7$$�8�;��bh̉9�Geu�m����hdX���P���s@ɟ�j"��|~L�C�΅BoB0�7��hNr_�1$���4�
��������z����~y�+�8/�w(��iۿ	J5������YQ�S�������+���^:�O�yϻeY�o�;`�����UM�9?��.�%ۺw|O
lT�|�]r��wˉ���ТD?[PP:�;��e����w�p��HE��T�:��
�7��/9��n�X\�/�U��
B�[��%S�7j���R��eߊ�Eg���9tx��wzl7-,d�<�Z?}�x��`�_6��X7,�u�B7���c��Ȼñ�A�L|���y�N�5��e�W��;cӳ�tZ��߃+2.M���ė�3��/^�t+����<s3ο����%��d��,�/�4���"ׇ�<p~K���*�M�8�[�<4��K�і�l�.��Pa��_�
J���9��eF����M}�>��	��c�+�I�z�0�����g%Ckk
�L�X��)E�'/�xј��f�諢ݳ(��<�Х��c
v~�9���2�0#�NK_y���r9�ʵuǜ��Z�k�/ȳ�<&۽-ٻ� # �>�ؼ��2ؾQn��M�:�Y��Fg����#W�)��Pa��9^Z��%����b]�S�+������ݨ#�&����&���υ�E��k����E�� ÔB �gP�P8P��X�γƖ�i���N ���ї�����Pw�(q �����;i����ya�#k�g�m|넲��^cS�'���;�.��疕�3BNC�qװ�X��.�B�6�Z wPrO?�4�X,���0B7��liq� ɱS
F�����(�P�x����S�7�EC����Y�h��g~��Hr�H.[����93@~D�6�1�q$m(��w��7����!������6  �rp�Ҙ�׆�׵�ZȀ�����O� w��~��C��h��$R�!p�T�l���cd�u6a7�V����ꚅ�R�=�gF�Z߇�H�G$�0rs}�� oD��`�ā��M��mw�)���=R��I�Ij.�+�h�Z��t�\i?<S���cm��=Cn �0^݃��Bt�<��˩�5Y]���
��6��@p.*&JIG�z�P��� ����I	��%��p��t��v��sI�5��`#C�P_i�]u�UO��e�;=>0��<����i:�O�$S�Ӧ��A]ѱTY^[c(a�D���V�&�o��<�������[�#J�-+/��8,����x+TU}U�E�Eta�UЗ�w�X��� �q��+�����ؐ�o�Q�z�M2?���Ҭ��2��X�
%������g&d��M�@����C�{qF��[��퓧i����{nV�3C��j��Ϩ�&Co�L�6�dfZZ-ݹ)9����%V@p��W�A�ƩL�;#=�,�`�߈�]X[�5�ԓ�ȕW���r����nKG�����x ���j��HK1Q�>��*�'�ɋϿ�� �f:G���^�$F�l�$!��\�қj������Vwev��6f��+%QM&a��>���~76��3���bL��8P�P�PvPf��R���(sw(_+�5o�%��*��(yS|N�U&��������_T�T��%[��%{�m�����zQ{�pa�I�=N�|����d�H�X�㓉� �<`np=�H���	+�8v(0_d��M�rr˅��!�(|M_�V�z�]uҵ�^+S�3��C��[�.=5�P�q��BHX�G}������tђR�s��� /�33�|Y	9��B��< .K��[@�~�ںupW l[[_�l�H@p�a� wD~��3��G�:;��YV�Dl|���uв��+�{쓥���<�A|�e�U1�x}�-�jGL'����n��6۽�����ʀC���_N����4J	`��H8G	5��=���P�$|��/��G��,+�������AO�on�4O��`&���V���iȥD�8z��b(,!�|�.����8�{���B!r����
�B-�� ��q%�i�z����©{��	a��L�juL!��urϥ���!�	Y�:�0$%&gU���U��q]\�糨*��Y L���M�o����K��b�\��a��y��刷���������/Hc�/�[c����d�5���0�aa�>}�Kkf^_h��ј���a<;�TV�}Y�9�RE�� �l�=��1U���Jh�f�IŞ�{�*�B-�jK��Z�g�J:أ��Cr��qYU��E)�e��k�1=%�S'�؉3��1%�K����TgB�Z���X�ҍG2���9@5���y�z�@ZU�I�Vl���I{��)�)F��U5��lǬB�W!����e��a��S��$�B�RRq�.9�c����t;�o#�jF	>1q���ZX�ao�7�
�b4xaBn�!)��*r��'S���-a��;5�����r�-���aء���݁kA	 \A�Z>���ń��閛ɣ��]��$���`䫓"G)��,����_y������r������^_���♠���C�@lχ��N�Q�t�+e��wm�yc��0���s��EE��[o��|�#�FE�c`��0	��7��ɳ�["(�A���T 0��m|�ǔ�q��ȁ��*��{bόg�� ��=a9:�e�-�[� s����Z������R j.�伐nON�(*�}eƙ�HIx!�9�(.��y�~�;�wx�؛}�ڥg�y��`mӘ�a��Դ��C9�^{���}��V�� �Qob��B�8�|.��w"5F꼃������a9� �RcT�*Cu��פ�rC�D�A�$oz^^Ӈ.x��RA�6BXnp$ɐ�H����U�_�(�!�Nt�d��YF�*�"�=d|��r���]��D��s��)�T檘��Y%j�1��'��t�~��QX�x�"G�����UIP�EU�T�_p��3�(��6�BOǍ�7g���r�WKoS�ǅUy�ge�̆Z}ی�6�eny���
i#7d�,���$}� C_�fkJ��9�/-JE-^������	*���� ��rA�9��٧J��d������R\q����\�jY���e��*��j��_AO�4�S�r���ϝ��b&s�M���k��nɾ�9���B��V��--4��{W�=��ѩV0E��i��7k27Ւ�NSZ��=+(��Ut)GH��V���Hs����k��7J4�r��-��&�������7�uL�s	O)+G�*��� �,Q�r) �M�X2�%�Z�*��y	,aҪ�����V�%X��7v�g��"#3w7�Ag��ʜ�a�w9�e�P����k��i�7|I.�Ed9AH�ƥq��cI�	!/�'R�<V
]���]���}7�zH��b
�J����b����N �cN189D�C1�`({<7�1�-�N<��aI�\_6��Ocgӝ)���ɽx�D�a=����Z�2ƈg`��	ဧ�C�PI�g�����<�;�����S��'���w����XɤB��R�(y}�����)
<�e�J�)!bY�9��A�}@,������|g����ltY�\�s��/�^5$���B k5��7ٳWf��\�z \��H�5}�]���~gH{$�!��ٌ���?H�Y\���E��uF����c����;0bL����8��<�,"��E�o��u^�,GE4�� 82Uk�X�Ϲ@ܴڮ�ʠ+#&��g��b�F=��q����S����$|��%�8�6:
��3��4�ƞuRhe�*.	M�@��dE����4@;�{!�V��$e�媬U�F��Y����,�z�9,�qO��zc皇e�����
�QW6�U�QPD�:xHn��Kmn��~���P��&{��C�eq�~�͕L�M���\��Q_�7��ᒹKK<;��?/��I�Y��H���\��d���j�^q�ޜ��9�D���G�s��|��*(����Z-�
���=[:xY_ݒ��{A�D�
wI���m�� g�%�֊uP��l���|D��}Q.��2�V���!(t��~��nI�	@ڧ�*CU�`[j�Z�����#���eϴ
��!ki!
�:H������G%�:�N�	B��%e��J�'�nyٿ��t�iY	�9�� ɄI�a®�3�C9�F��`�ǹP@Pjf�B���0n�jLjE�(U\�9-B�!ı�꧐���-�Ej�Ǹ��c`ށ�{:��CE����p��h:,�V�GP�g�wڞ{����|.�=��U��3o'�]s��e>Gn��$�A�Œ�̰�6K��8l^�=���w0\f�����۔?䁕�[���u3��s��Vw��kf�a8H�*4���1�'XpG
��3gΔ�1lAa �xC&\�'��i���򪺎ϦQ�<{���<Ǯ/�*��a�*��^_%�;_%�?���l�mo�aq<Dun�ICI֢|������L�+2����sk% /���b�C�9{^���X�LB}���	șK6'��'�k�<�Q��0@BuR�`0�aH2��}��a�~HMT�mٶ`9l*7���5�^���P�T�(�yio��u^�\�"s�}t�9�U���E1t/�*��*�j�w7ח^x����}���WW��c[:r$ZY?�Rk��T����� h���~�p}v�Y���{w��M�y6��w����x5Ȼ�8,���e&p��^9��ԅnd2wB�����/��ű��5@���N��3��c��v�Z����ɤ
�FM�Ŵ��fTs�ʊZԒ�n�A.�ޕZ²��om�M�77djZ��="�i�<����]D�$�\~��2��IWIT�Eƫ�d��Y9� ����}P�´�gZRo�W���P��9����{����̓Oʥ
���_F�ځ����sly�G����s"GO��W���*s
Xf�\|n~��Pf��,)xl�m��rN��Z�bixU�^O糯��[oJ��Y��j��� jB٥V[5u�A�v�]G}���{��G�j�!�����6��b�JenT>�Sc�%d�574���V�0�����pJ29o%#��A_�d°kaQ>�����Q��dcS�J ��!5�8_j��[�˞)��.#=+�l���]Ob��I�#.��xR�>�yC;aRo8�5�.Z�%�|- GL0Vens�����sN�xG���@T��@dB2}�C���|(�_�5�u�<&+o6�[s�6�����s����T�F��e���^'�c�0^7s ���uA�w�������i�j�E#��p̂����7=� �)�*��/�̫C3V a$��Ҝ�%�8�Z���:;��,}�R��ϝ=���Y2Nl���I�=�"oo�s��� �)�ŵ����r����[���g��5@��*�,Q����������)�R2��䯵�u^�;!^$�h2&>7@7dnI0��F���)"-E^�}��;�<�П�3�����?��}�_N��EYn�[S#�%��j�8T$�TOG�l�a���$ߊ]/�"W���Ev;ʆ���
fÏ�64��P���47س��8��/�v֓�L�H���Br� V���lw�dc�*�
�>_�� y��<HvSFɓs�2q�ڔ��C
����`]���0Zd�8�+@�eR]�ȁ楬 ����){g�l
�<)۲v��&c�ܸ �}Xj뫲xp����G�_�������r�e�eOw�^W�ǟ����˧α!g}u�k'�ș����K�dO?���9�>&�X-/K�8����@(?y�Ϸgu ��*�W�K�xI���d�=�F=���
�eϭ�Ⱦ[nٷDA:�@���<Hlt���\����b�$���K���凄	��=SH8L�J��[�+e%��"q�?��AZL�H7���.�6NG +Z�3�9�� �}wh�������-s���`5�**�:\���Ť��}��I|�H�� �6Q4&\;��΀[�vl`}.Ԕ��q�y3�W���~������eK?�F�?�@Ӽ,��{Y��oaC���4�1��I�5&��l���"Ŭбy4�F�n{&��h0c\Ze���7謤;�_�gY��o��0�:��c���C�P��ڀ4	�T��ו���}ES��XV�W�P�'��^U�sZ��s'O������`�rEd1�P��g�Mb�p��p�G"���<��Sr��12O#����Gژ�-�*I���2��ńL��B�FVT�ov�~�I%���]8I�8�n����2�bӿ�t3N7Z����f6�'�Q�5jQtݑ'����yhE_���w���oٻ�ս�9�U�FY�ưU��p����k��4��A`	��C��a}�1�rQ9E}�&����6R���Z��v�$�U�*�cP��8�*ڮ����&rx�tL�����s�J��I��%R��% �"�q_�w�4�=�p<yteR�w��
K̲p�t����ƒd*��%��k��^�C��6d����K�ʼ6^;/+���}I33R���[��ecCz.��5����ZR"gU����cr��ȡ�P����ʚl�;'u��=�32x��U S�]��'EON>�8�a���;��k��)y�4�:�=���uX9�t�2�w���6Y��f�K�3�w{�'�N\�Q(3�ח����ڱ�Q�+J�/:,W濘'#;=1ab��S�f��-B!��j���N�X�Tv�tBb9���{��J�-/&L6�S˭�m�m�3v����桁���X`�//�ͫd�	�YLa����%)qm	l���=Q�����Md����Q��
���P}�	'�	���p�=ˮ듦��e¶&6�歲� ����\��C��ŷC<����5'��}���́���1v�1+.]9z(-F��s�H}a�c��YO��0�&���d=PP��2�u� dq��^ �c�E�-�  20�&d���Qy�[�;f�dzz����4ὬB�CEU
�k�&L��%w��lD��sG��G�����43'U�ԑ<?�q�� !E�0��K�vY�N!�vB�t�n����*p��إ�d����숰꤭ `u{C�Þt�S��=K�g��~�G=��?��?��@��7������>w�B�[�4�%`�e+w����Ao�X_��3;t	;�8a����o��u�{�υ�"�]I5�.q(:��I�9�%ژ�A��K�q3Tgc,۫k�r�96$�/� �/a�v�Y���������̢#���9�`���q_�������?�Ʈ䴂�˰N��:#Vɸ'�3���3O˱���)Y��U
pH#�7�,l�;K/TL�:O5s��a���E署�Uhiܕ��:�K���iN����x7�]E�,�탿%��l�}P%B���Yi���R��]۔u����m!jaA�_*��V��Ad�^�N���~6"��K@L�t�a�8w4�q��\By�G����	��wæ����w��X�'�a�������Й?��?�����}���>�ZzA�|���+��+��<�0xQ�N8�wcW�2�=���������	�U8����sZ�� in�
L2�r����%r����k��*��й��w���;뗔�����`��BI[��-r���M*\�j9l��dk�����ɶ�A�Z�����T�/�5����BJ�Ls�w�Ĺ����xT��<���d r����<-���Z�x򤬟=�`��# hb�~X�y��������și*��hM�����s/�#~Cn��V���C^�kM�w4v�2siT���ݦ�g|[ u۫�r���弎o^�4��0Z���nҪb4��!�JT-Q��o��^�G��5��p/��sǡ����ח��=�� Hc�b����[�F�%��>q�G����^z�?��/��O�����g>�|�ӿ}���Xj4/i�;I'�a�/ +�W���,�
��r^xA9��5HG/���:`��UT������ܦ �[V2���]")xO�e��Z >��t��7n�K�P����\��i����]�!_��L��y���̵�8^�)�>��@�!�*!�.�|��![!�Ď�"	^�H��i�$��T�l�>)�UY���6h��������+ �Cc4�mZ/�/�L��iLw�,��`с�̗*��4rJ��$��k�	/k*�ªp�������_��}9�xEj㙖4�+�C�_}%�tZ��2�'`5#Ȅ@Fh�)���pE��j��}`<�)w����9��׌_�v��a�!U�0/�%��I��b�;�B�u��IX&TBa�*7�sA1�������$�s[U�X��	�q۸�I>Pxb���(�rQ�D�>AA2k8vc����]��C���{�~0f�"XO�y�	�I������H�u�Xwy�J�X�:����&B�RhK�k�`��{*����^�6+��*�^�]�I)}�K����v��@ ����Ҳ1��,8vǎ'�\(�ח�Uf�ϝ�9߃��,��4V �9�O5H[�M�R��UT�{�BU���SV��o<(w�}��ݳ,��c���»��5���R�G�j����yꑇ��ѣ�"/��a���ڀ�$��0UCtR�
+�G������/&�ҽ�[x����r��!,j݈md��曪�λ�x*[�*����&����w}㟿�?�j|�~��?���ÿ�u��{�����ۿs��<�1EF�*�V�Z�Z����Pz���#gu�c���E�ٽƱ�{�9��"�V*�H0c</�n�$��(���.���t��ݪI]��HiI���IT�'����H�*rVlmm0צU��u�������\8G����.A�3C�GΉZÁ��g�7���|���c]�m�8*�8���Z�������X��_BG��ԱWFT@To�pԗT�
I�d����V
ke;w 6�����k��W��A�8���K�ݒ|�#��r遽�:�_���L��_ZT`X����sV�#G��-D2mƩ3����T�]�>���-�l�����Ę�o��EU�v�j�J�7�tp��@C�GS�L,)�[�,΁�wJ�+T7@z�ޣc^�����������oދkӲ/A�/\⭰��R���?L���a�p���b�I)�/���n�TX�{�P����t<a�5�A�����64+���N�������9���h~/ �T��^	�
���Ћ�J��H�[�/��_�d�w�(�=U9�OA��3���� >6V ��+��I�X�-�q��h{@)��"�A�N	$jihD"���{g�2�>�v�%IS�  ���Ûz��ǎ�?�9i���;�ٙ!���U��$�ۉ�_į�e��)y���募�9�כ�k-u��	��Ɔ4�3�ykG>|#D��/�ʽS�U �7��/y5-*I��ebB)"}�.�n2��AORP��B�����Z�弾�����ʼ����˯����~�?���f>�}������_B�̧>��?��������D#/~`���vG����q@�1�*W%/k�A��s���t̳��rk ��X����x`v2�"�]�Df��d���e�3-���DY�rlx*j���@E\��f�}<�������)�A�<0xY����C!΁઼�����V �òZd��kTۻ��G=�2�<�<�n_�ѡx8"8�%J�S
�X&V|O�!��tG�
N�;mg�bB����|�&d
f��y�� ��hȮ�L����ݙ����R��ֹd������,�����܆>I��?t�
�ns&���;@2_Ɛ�N��/=B��{�QV���}πJZ��m��0���A%�7��c"�`�>4�]��?Kܼ�P�o.z�^v�(�ɶv<.|�-���C{���0sΒ����&#�"�{1|ļ%)=v�	��Z�ǚ^��r>IN�J���vO+60'����`&�������3�;�	���ޣ�Cf-_$�d�4��{ظa�<�>pi�I��� pQ��Ȣ;�U69p����n�]�SĐl�<"˭B8{�=K���`�f�1/�� �v��{Pܮפ���oWj�D��O�U��ޔ����Ҩ���eW]'�3s:愆P���f>����u��˱���_��+�m�ˡ�iY��Ȟ�i)���mS��Q9O1�JJ*����*��M�����!�J��i�����vO�N����D�E�ӭ�tC����ҿ��M�"���b����o>8��������ɿ9���9��x��ƀ0�}�����������N��ѥf��f+����%����S���/@�ʬ�b����#�	��Vi�u*}d����=7 
5���I���2^:(�c�"-U�W��N�ӞS��^Xg��j�y �ci�bG�6F�9;��H^Y�������%V����
���M�ᖰL
l�HIfd%��aJ�^��w @�g��^#��m�%��]�Z$� $�xb}�n� t s9��/��s%q� ��lH���7{`�ёר�3EWm�� bvu}�2�R8��@,%�8��Bzi�%'z6<ؕ�,�Z.�D�r^쑌q� ����"�%zRBPb
�`ջ٣@	�y|���P�a���'j�L'H��gh�}QZ�g�62���3��&��Tخc4z��+�I)�n��je��ٳ��U�x�3�!#&�&�j��Y����%���a�r���,��=a�������D��7��<����F.g��u�ӛ*|�6�q(7����k	v}	��iX9e���R����g��8v��{[\��׷�N@�L�C����y�N�N��04F�X�@L��<|ޙ��5X9`^�ˤ��vܶ���}���񅳥���TC@�9�Q&`Q��0=�U5���p`kS�Gu��T������?+XO�=�}��|�m�Væ95��6������#��i<����sO��}E������s����\�wI/,���HݫWWdJ�ќ�b�(��������4�F���n��7��/i1�U�'|���:xR(~$8��2�ږ���n�Y���5�,?A\�
�[�zSf:�h�U�u�w^8y�������/}�w~����K��g�7�����}]�X{����/���������~��q�b�vpyj�5�@B��`Q�<�Y���Y�������k��5�f�@�T����* z���v(Ȝ+�/��@��$U��I�f�»%�R�}{d��˥��W\�5�1�,�n��]?�^���/!���IM6�+d�e�X�2���|�o����tJ�͕L�끖�n�m��G��|<+\��
(\��i�eX���v���X"�G���[���9~���1� ��5�yi:�b/!|Gµ��~�<@�K���$S��9�Vf��W�j�5�E�1 ��h�9e�Ҥ�:�\�f��T�\wwIRv[߻��m�$w� �w-�Ѭ���v.)s��q���o�Ae�-dV���q��N��nе�k�1<�<08 �c�T�o����$�@��U1W�N������[��m������T��� ��w(�I~��Ǭ���'V�{0v1�H8_�ڕ��x�#�;׃���r�����ڝ�^��PF�ƪ�Q�� 	��œ5@o�Z�Q΢:���,/�1���_!y$��X�B��憴X�0ݬ��۔���}��!�Re���9YW���ޔo}�9��iy�����ny�����y����\[���xJ�|�9�ط��G��
���2���2/w]w�4zy��J�ݕ��pE�Q�����v���Aʝ��\�5������V�b0�diN���벊�f�`�m��U7ʆ��`M��M�B2���B��X-�,1-�
 �
��2e���uWμ��p��3����lv�M�[�Vj�t8j�on�no���ڼ������N3��6�9Rp2�g��>^QyE�S�(���� ��E�Jv��B���|�a��䏕B�]�R$$�&>�=���pϊ�ڨ��>�d�TT��؍�=?�8�jC`�謦�5��ʅ�c  9��I&$�A�A��D4G,��H���Y^M����<*�MB����  º�c��e�K��yʇLLK(��@9��=��תȼkV0a^I����\c�S?�ñ;`L?/ ^�xQ�Dk�˩��$f���Ξ��(���ʅ����:D�lF"E=k�<���Z���@�ӻ21���]��7>ߋ@!Y	iX�b�+a��]+Tڜ� ���*��q^ͣP�;n�|^J昜M��·\�P������\`���q�g2O�����y�/����`L�9�����Rd�.���y�a��%<��Wq�@v�D��@!|�_Y��=/0�j���w��|ވ�3;�U�-�D����",^�����W�b�1�i>w�r�ʿMO����(�yg0�	I.q)�	˺�OK0caO|�*�F~|c5*�n�Y|�B;TCik傴���7Ԡ)d�)��W���P����G�j�����#���S'؉�������Z��,Pv�������r�<��y��#��q�-��jʥ��r���\:7+�ƆtW�UG��NY9��i0|ƙca�ܭ3���
�����26�����^Ծ�dY��Y�)�<���
Rt"QT����S�ټ$��L#�
L�m�\�P=3$�X�&҂�V���p��>�i���+�"��{T��e��9n7[�Y�^�bS�j4]�KC�t�냥1�$����E�cD�?�݀S ?UV���quG���5�}�r��J!'�
�/#Z����H��L���ry5xQ�S���}=�i��-���ΐJ����C��:��r�S/�gS�Y���})���%��$c�Nn`u�a��76vY&�s��\��8���2d<�B���z��K�J0b&\K:�� 3*�=�U�刅���	'�*-C��AbA�Xj�y;e`��e�@]�EA�P-��
���,c�MA���yw�{�O�R�W��6s�|#Z������ĜW˅��l�N1L��첒MY�
��J,	֔�������N;<�$=�J׼+�L�&��Ƌ|4��|�O	����#�H���Y+�㕵�4�qY�F{��:'��]*�7E�	q[~+���I�h�|�a�0�e�ż1�+���Q ��kXޏzBV�U��%��9d��@ī=/�CD��k����&��\��@x���<�1�ݞ��8'�����"�K9��$�C��]��t�>Wg�7a�-��ؠ���ݬa�@�����X��S�L���PM�ސX������ E�m�u�� ��F��rN��ڐ��?"G.�T�g:zOU��l����w{mni����nȬ������kd|T�N�4��	����q�.�r{��	D+�d
�Ë���`���ڳ M��c����n$���g�֐a�'� 0��ҙjK[Rg�"��.k
pV7����j��ǉn�NR�u�b��C�w{|1[����@Hg6�J}Yꠔ�����B�KI�������G�ϑ�p�1得ۭ��AL3�ݘ� �	�*m�<�C8)�I���M�@����x���fSK�i�}��a淨b���5E�s���yH\cGrG��ʿ*N��A2�r*&�R dL.�}
 :OKQ�%���̨�`���>��
�4r���e�RƲK�7��7���d8N�'\���	�o(����a���=CǺ�m��h��"�֨q.�ft�V��'�����̅Pz�*��Q��<��O���)1�p�2�"�L�<#NqN�w)�%亘T����f��0��2� H�w)N��`�N`݇���5�b����^��*ܳ��*U���2�;�z2h�����O";@}������f��$�˼W�\��������xr���u�2e=6�!hu�%8)�nw�ˢ��/*�����Vab1���·�LZQ��x��f>��O]�jT��b���L�M���ؽ���W����f���ڣ��z�*�Z0��'GE_�ZuR�Eo�����s�S���#�iA�z}Y��6�ff�%��80=�b4SA����xcC��5��D���!�'�;�&�Y:fu��ࡍ����,7[2�����: �����;#[�����s�Ǯsuf��pRs{5g�L�	�/�,���/�V�`���$u}�(34ǠsN�gH![H@�@����[]���R���]kl����)]4Eӗ��H9�������@�G��`ߐ���)�F�� H��G,-��#R�#$��$r%vd�/> c�d�عX����^��%��~�dT� - %N��7TJ�ո�K��9D^�-��H�qZ�*&*q�NJ���_׳��X�p	.���O��ܱ���3�ɘax!��
`�a9:��M�U8m�C��aV:2��S��/L�̭�b�+�mM�� �(�1v�D��8uU՚��/�f���s�ș[�bt��p��1QiHP6a�h�b���+�9j�:QŤ��Ue �u�oRD*�ȷ�d�L����e����G��˕ �T��3��w��B����-d�5b�(T(�^jɓ�֮30"y�i`^���� �ru����b�ply0�+��μB7���|8��0�����;�w�	��ݓ 
�o��(���d�;�Y6��!���x>?�;�>�d��͆�*!���X���PZ	��e����}�;����0,�do��`=/�E��[h(�y	�p2�]:���i��3�.vG@������N�8����|z�*Du��_�t��H��&grK{���YYhM�F:TY�';nT0�<tH�F+JjjT�RR*��a_uT�����;���n����������3�q���H�UPS�� V���RgD%!��}�\�4&�Q��7��/q�d��d���/���3RK�8-E��B��P�M���֥�������շ�dZQ��O2��*�>�Ut3�R�L#iwZ2��]l�n�����������NS3�!�ݚ��"L`%殳�������X\��o<M�*�O�ȸ;����j䛒#�OFE��W�S8�
ֺ*jd� ,��'�B�����6 #�.�?a6��`�S5u�'��QUa��Yqc�k�7Rc��ʜ��;J|
�ԱE�(X���[Pa�����,Y��K�kE����7�\�2�_�Va+E��=�X�b�a�K'������o�� *X2^h�M�(�9�n�K�; ��`���a�sW�WE� �+�T�����I����zN�ʤ���L[��v6K��l�c�
�����-�q�3S�f��������#��X���ݚ���qn�7fS:�H�|���J��|Mc��vn��1?����gw�-W �Bz;r����%�f�_�R�o%0��t\60sUJV\�x&L-���-��ͭr,�,�6����$��P�T� H5߳&xn���W�>������LbT�`��n�12�2LU��l	f}�4dֶ�0&�L������a��*w����i��C��9��A|�.�q���ҍnި6�|�5��4��s���L�(�<����
�$�����Ԕ�>���rN��L��j��j�\~���n��f_V66ek�Rw@f��	�Z�^L)H�s��̫��恹�vy����H�R��������+RS=���H'ql��&<.����#-����׳���z�n��.T���L�������]�2Sd���&��X�����Tt�GSME�m���ږ)U�}��.��!������"�R�k��F�o�0in��-��X��MAN��R�!1 4���K��n8G�Ao���\	Z*<s߻)(�,C �����(;9;H��N -��D��ZG%<5.m�I����"]�
��Q��A���K��L���4����#��=����Pިj�'�ݜ���a����W�9::u5f���dтnZq�wG�=���`�@�#N�,�����[�KҏgM�cᔖ
��V��58�u6rUF ���� �L,���YL�t��p}� �pω�d��Э��
!p_�J3��y1Bk�l��c�XL���G��a��m�Z>A�	<>e��>�2��)��cz'v犔y+':# �K ����Y����Q��ت�����d�����Г��
��|�s�$�\5j}�>�'
)��I��hI�@@����I�^�����^9=`���C�a���X���w>��7P�iR���y��Rڢ2��=���	=7&�\�{gy������<"����֏�%�;�(s�K23������*A�+U""����W�0/m�g2�ӫ�2$��aVe[��MT������O)�XR���zۍ�웙�T﹡���!��#����Z�S�GA־=K2�2䐎yZA|U����I�6���r`�33�Ώ�c���"0��c�瓡]��|ez���/�գ�f4Y�&c��*2��6�� .��4��h�u��2.��W��*��n����)�RQĞ(���e�<�L*�jv* �:�HF W����g�}?��4ﬨrc�ۚs��b��]*l����Qx"��a$J �s���	f����b3��i�x��ޒM3W>�	��!�c2���ƈxdV[N�^��i�A�ۖZ�j!N�%���I�8A��o�x�
ѹ�a� �Z�	_\����R)Z�*$x�%��* ���f}k�J���FV��h�<�F�Y�Hƞ���y��_�����H��h����`�'H��x���i4�M:�.r�z��s�;���y����T8�X�B����BH⪒X�Y�x8p�n�t�E�14Ԣ�~�TVĬVj4ZNq�ݒÄV��+�}ו���ye��eK�|�x�֜� �q]<�u���.���G�'�MK�Uq��h6�w\��=��}|�j9
����5m\7ε1
��V���{y �='wt��MمX��{Sn���� =0^�b|R0'xn\�3sc�K�Ֆ�ԅ=1WM}7�Ã�܅xb�J���Ƚ���H8����϶>k{���3�ˆw���̀E��q�}��Õz&_}5��諆֑���]�N�}���I�kt���Oݬ�����C�=j�1٢9vIȨ��d��\��r!a�,R.��&!�S�B��RV"Wlb9����]��L��/���}�dy���Q驒߿��N�U���S��XX`��������pnA�q����vq�;R��oy�}�ή��+V$ۮ�yK'v�h���Z��-�cl�j�w�.�l��.sě���<�+d�_ֻ�u��?-��mi�\~��LCf�.�T�y� k��#�1���<^��|�Mz��*/��p�&xy��a��$��$�Ĺ�� w�p�d��Y����*ȯЗy�ѕ�
�і
�fW�
�Z�a$�6uSd�P�Dt�,M_"��"�����]`���Op�̪$���L�+|#;��}\�g�[���gI�%�ƃ��J�tҕ�"yAP�9k*�</Ej�x_vJ����õ	��
 �SǏS����=q�	 ������W%\s��ZUN�9M%E� N�]x��ju(�766�̙3� ��9B`��u�X��	us|eEs�W�����,-p��)y�W(8!�17P�x�Ç��	ם��]R[n�0��-I\6�[Q�	ϼ�J�֧
M�!�}��IK�
< `���f���~$�ϟ�Wt�Cc;p���]���k��o��^.�ʚ'a/P���vH���<�ك9{���������bJ�<���-�����y3OG�̈�p����y����~��I�6@����%���@L�k�Y^�K/��
�#<��/��G��3��Y]]���%�馛x=;��u�3���|Wr�[�c\\\���p���:���<an0�sj	c���TΞ=˽�=iݬ�놱b=��Xɧ��rx6f�^�<Wx�lb�`���y>p�X�Vc�=g@��	�s��Y���#*������wcC�T���%��~X���_��9:�r��ā��٩�9�1���UD��%����Jڅ�����BQ��(z4�`�8W6��f��ʞt\8o��g���g�T�j�Z<�ֻn�	C;�NgH�EC\������/t=n��M����6�a����F@��}�#h�2�ﭫ|,x]T�Vu��:��fW.;%ٹUI׷���|N�Y��r�4Y�Y]�A{콖	�̔�0R$���c��:��W��^_����㱮[�YB]�D�H�H�X�O�!v�s�Ӱ��z�&F�Qo��H_�J�⟺9+�𑯐�� ue���4�@N*I�0,Lp���c�p�ڰ!9��N�-.^��  ��IDATX|9LD�v����O�ĽnI�8� �0��$����[]y��'���B�K�*��.=$����{�-3*�x�g��_�:��{��^���'�����_�/}�K����/��]�����?���ٟ�)6 �o���k@��r�-�3?�3r�W���J�k_��l�^��K>��ORɘ���IX���GO&U�e�9KP"�G$_��^
l��!���������Z�����p���C�g����^뻿���������]旖��c(���/~Q��^}�s�&�c��� �䮷�-�x�;�mo{[��q�o|����\3(e<���O|�J:�O��K/ɟ�ɟ�������p/�̰�����8?�s`��<���)�)��'��뷧���߯{��%q��\��?-O=�T����G~D.��*u����/� ��ԧ���8����'�'�{��{	^�M�Y��
�~�w~G���or��9���(�EX��}�s?���r�b.-�������Ϲ&���O��p-���<���<`a�4�u?��/�r�ؾ{�ᇹ��կ� �����?���}��b�c�X���� � �"��H	6�>xwp����-
��汧W�_�G}T>�����zĘ��{�G���wq� ��w�+G��/���ñ�S�m�H|��Oq`Y�+,�ޝT��}'�-a��	�춂>��ju���ݚR�1-���C50�Q�4`�,-.ˠrT����A�"$e�o��W������t`E�թ<�9X`�ㅵu�\�b�Fe�-���ࣽ
��g[q�F��	s/PkSR��BAK�?tDxզ���Q��/��].I_U�Ǫτ�X�MG�灧���͜��GŘ��}���]#�/xa�Z�<��`����E:��ں�GՂ-ϑ)���TD?��"�NrIȋV��B����@묷�=�D�91�{#vO��������p	���2F#|ʲ	V��@
1{4��d�\��P�����O��yR.��r�3�ɽ;�\�P���@AaiB��c�=&����H���n�r�UE
a���sx	�LP��e�,x s�'�A��߸7�1�cܻw/A\}���ypa�C͡I�j�|��q�9�1;=CA�t쥣��s�ɵ�^+Ksv�ء<1�O=���y���ʁ9(�v{J1�1�:O�"�E�-WŅ1�1OP��j��b�&<< ����q��Pp�����@ ���s�ߖ�5�"�| �0$X>���
�x��Y���X;���s�e�8���q/�'��<��C�����?��r�UW�`�� ��Y��k�߸�)n������;�c�Z�Ł{� �o}�[	��=x�F�&�@	?�q��  H�����}�}k����e���t�c,//s��{	 �}�c�8߀@�	��������>�vr�����: ( wXCz�<�,��Ï=*��ַ8�V���:v���pF��
a"xu��3b �aMa�1Q<r�:��w�Q��_��w���<0;vT��&2���ae���mH�ڦ@�Ņ����v��\�;^'T���7mSeL�恲[g׋͓�k�Aft�b
zY`�����#��;lȶ���[�i����_ �E�x��@ˁi����Vu\s� �X\��gn��a�b�d<���������X�/���7Ջ8��d52��.C@�d�7/��Q"��� .��u�ő���}w�>�Yӧ��.��y��!d�y��u�-��s��.?��	��LV����x�.��n�	?�n�s1�,.+�F�4@�P���R������~�G���g\扵,��B�����],^�s��WS��ʇ� �����[��n?�?@Ai�x6�@��> #�ʩw�#�~ŕW҂��8¼@P� ��0�y��,�ē�A�mmu��g�����{�M��穧�$���{�c�y��vG�,B���%�����^�/�% �U
�r� �>�����*��/}�˼��>p`S �`�~H���z���]���,�,w�y������1�(̷��� q���|�<^���Ūi���'u�����u����u�1\��`?���(��J!/x�>����|<�!�.P��;P�?�?�糤c�����������3��qO��-��}i xN�>xư� Ζ$�#�	��S?�S�� @�F��]w�Bew��]������gcu�φq`��o����؏q��#��`�qb���1^<�%�b�q�χ{�{��Ç����& 	B��g W0@���=��/<��O=�g(r��½����ˆ��{���#Gx=�B�oܿZo�����y`��9�����U�dwb1���o��a�xX�_�|��!8�yCjզ��}:���ʹ��_�d��!��"&��,{���2�+��V�>�єe�I�r�=���� ���
�N��f�r*H_�3껫�lƪ�>�KL2�Ե��?�w�9�|Q��+����
@�0&����@Τ�kJ'�[$*�JQ�}�Ͱ�k��Y�%���^\��p%���Q���c;�K����u_�T�@r�ܑUKx>@U-�ޏ�<�x>!��e���RHȀ�H'T����J]&%��waތ#�{�#bմ΃���x�}���yW�('(9X(p�CHA9�Ӳ�Ь||?�p+[��L_<(�� F`�B�C2��������{`,8�e��>,BP�� ��7� ��z+=!����.hS~�?��%tBV>��3�%�q�{�}T$P�����esA*s}>�=(*�%`�=�&�ʁ����c³�~8��:�Z�����:6<���P4#�%�i!E<#�Ɖ����o�u��x^z�<7XZ�j]�aɻ���1������#�����waC)#�	����|��I�����x��X����O�� �CY��?Pο�ۿ-��˽���Þ��?�c�$|�<G�(qoxP�����!�K &<' ���>�5�� -�L0G?��?K`�5 ������q 0a_ �����8C��ѩ��,��?� & ��	9��o��oɟ�ٟq� ��<�/�X����v���g�c��{���%�7��W�W�A�kaO>��B� ���αbQ~���� 돰��V��'�olN1V�ǭ��N~{^���0Mט�����Sza���9�~k��²�H^x�9ٺ�N��w��[�B�*�`
�ޛ�䒭:�.
�p�E�)�&��A���Q/L�4\�JN����qߢ�xV��
� C�h�`�N\��]���)�"��,䉫0͜�K|�ޔI�5��7�F��#�UUoG>����TTV���(o���
m��5<$�<�t�W�n�r�yx��آ� =*��S�V�O̕�"p G��S)�W�'�4_$O��O.N�%�;����wI�e�F�$�R�}�����>�ot���Q�`!��*V�xK�B�5�.�a��`5Û K�
B�����	\ϒK��Pk��	���ɔ֛������b\�P�޸.�K_�aI�`tAYZH��wPI����\��i�Jo��R�fݍ����P݄��;�Kff��<T�����en��=���<B�:g�a�����:��#j�bN �0� 
�; 
  �8������< 9PV�+Æn>��='\siU1���|\3,� ³�~ k 
7�|3Âv���r`*�zXU�B��7������\�;��僑�M�
�/���<sP�P��* �X(�bϫ��/<� A� ��G�Bx,ٖ�����8��ާ)�>Y��=Y̧��^�k������ )̱yH�~nW�s�����|c��,��V�`�	C����P ��C�����!A��c��)T1ṱ�����X(��\��L��w��15;#�/9�u����dϾ}R򲨁�����c>q�$|�<_a��n�b�6��ᵜ�����`S�k��k�$��{��Josk�{
�(,���1^K|�A4i��꭪�+� {�طp��1� ���T�W*�<�iI���­��x/z2/�3�=�m�Kq`[��/q�acD
P�I"N����֬7s��I�U��/��Cl�����$OU������n]\�Rg�:!�d��qK�cϫ��H�92')C�9�z�4��4e��rs�$�J�bV����ºd^�lᙑ;�g̗����+/`e��1_
Հgǫ@�E</� XZ�Ji�CY��2n��Y<�|T0^��߰z!�! !h� d�>�P�K�,t�JcU��)V��N�uQ��u�� +�/� 8-� ����WY�;t��9�C# ��� ��jŸay�VM`�����{�Z� ́\ 9(M<��O�d,�����1�z������aٵ'2���
����(�� �x&�P�� 1K��2X�F���a���mX��<%����	�x��L�;8�Ə55�RߗZCAS �����E���O'b���@�(�p��C,��B3����o9+FP��@4���+΅2�K����2�S&$o��Ϫ�G�+o$��\��A³�� �w���\3��g|�3�xq}۷�gc���u`�,����A�>���=���Ǽ���X���i �r����"�]���
� �9���3N6���i��"3NxXΝ�0q��9�[ޟ�)�aҮ;��� w�-�[���nwX�C"n��o0q�^T�����
�r
�O*����b'ߋ�Մ��H՘ �c�*h]ז�����^x�a��(d;�fzv��5w�Q"�a�(�BG��PPTa�R& ���qFXN����ē��^X�}��V��V�x\e%r�ȑ.�L97�����|)�H����qI���< �
�%���#���Hp&�g��]
]=�KH749* ���z�=1oE�����'�Ȼ<B�$�*d��c��E��f!�,e��ka���J&Lh�1�I^_�g�s9�	�!�)��?�g�'DB��Ä?·u�� ���ׅ
J �6���yV<�9�m��P�uF� \�x(,�6�@B�9�I]��ȇ�ª��|I���Z���Y��a?|�e��@�vX�N��
����u�����$E���j��Q�J���q�`^�@�-�sw'+��$ C(��C� ��ax.�&Pv�*�7emJ��-���
Fh�`�3�j�`�(�߰�r3vZ��XY�%�b��x��Ȃ��=�T�=���u��
 +6��{�J���n�o� '�?P�P��iб�</�H �~�w�^S3�+���
[#x�-�!tϑ%�b~�N�݁gϳ��c��a8}^\c��0��K>
A8�p�d ��y��� � >x7\c���� %���Da�����4���<����p��l�<#�g������� �������2��2q��q�{���_p�}��9G���܃#�6���±V��扇��a�.�c!C��|^[�1�ːF@�ĝ�u��[������+��=��oVe�hЗ:BfC��1y���c�l��4s����p��rV��j���TW�;9��5�~}�F0{�ҁ���� I�ț��˜�=��@&"
0.BR$���kE��{��6�o��u^F���n�Q0���
�R@`F0!��3)��o�+@A#��G�8��PQ4fϱ�����$�l�(OK�< NoDVX�a�'bJ��8
�q<�K�Ď��{J�xnRzx.*FD�r4���:a�����W@���Z6e����sÒڐ����}�,S|na���H�;9������h�_��!ؠ\��p@����5
?��u
���ml\f�YhȪr�Sc�//����|��
*o\�]�uT�  �P�|FN��E���?��^(v���h�=`�B�A����i݇H�֋��V�(�?��?�������}���@Y�m��sA�!G�5q?��"��Ǹu�m���Xi�� kHօ�D�*�8ڞ�7o��a�~��}�^����k���yY<�5�x0/�|����_�5����*oS�V�c{��@��������z�'�/��/0�����6��rl0��<6⫾���q���������|�J�:�G �=�S��oȉ��� ���3̙��bO!��e� f��"3<pM���ʯ�
A�����~�x���D��=�q�؃(��/}��
�0����b���,��4b�E�p-/ $	�>�9I�X0ȅB�6�]���\��3.�܍V ������=���ӹ�W�i`�K��{���������5���êfTV����R�z8�
e�p�����T�ɻ�>q��d��E�����5Qu�˘_ICr4.=c��b�n����F�{6:�CG�����z�qL�}��Q�ϵ�$��U���q�4�7��k���c�I*�rӓ:/�\r�a8�^���)���h��Q��M��/0JD��ƀ��(j��,X�V#�C�]��>��J'ё��y��B|3;߀�$qރb@�5L���&����ޛGKvUg���oΗs*%���,1�r�m�$��L���^���v��r/�rv��6 �qUA`$@ � 	���&$4fJ9���q���9ߍ��^�Q�E���b�|/"�=��s������۪b�f1@F�E0 ڈǰ�`���L뿤���i���en�Bj��΅j�QKX���Ҍ��* "���"�vf�($���#�ߥ|9`w4�A��Կ��Q�S,>/��Q:)/y!T�<�6�w�`BDK��|[�s���_�z����c^���b�N\ƿm�N+(7FފÇ��o|�[V_B��0">?�i��������bބ��|�)�2< ���'�P@�%^�9�J���"GY�:�2�D�f��?f��7�h]���3�q�<�)�6P8�X��z����M��7�z%M�8�+u�=�рO"~	�F��~x0 sB"�z��k�f�,w<�X����Ƌ@p뭷ye�݈��^-k?�-<�*�	��;����@E�T�Ay�fP�xo Z�
�C9��O "���y�;��� p�XCɳ6�����/۞�Ns��=�Y�;��s����g�j�x�xH���g���8z�V�����<2V 󡢐�ϔ�����3��e/���{�+9��02�qM��
0d�ꍪ��97 �sp]���K�N&��SI�LO嗾�-�G=����9�7���À�ԙ+<�n~.�É^�r �V���� ����5i%��O&+̨�p�8�g#K�?Y��vbX�kkl�	����8�MebvW�<2xj��j�F��2'?َ���^��]�QsL��%�h)�;�zJ�q�,�'�qʂ��(Rg�� JP�s�Y�7J��`[�Ph�E�a	F�k��gF�mÝ1��W�'�-�n��Ю��Σ��B�F�����q�n�P6l(3Ha%s_����s�z/2��2��,�Q�*�7E��"(��.ţan�0h��(X.�_���W��E^g��ƴ�,ȴ���/�h])�5����{8\�Ɨ����!��n������Z0~��R�_�V�Qy����
��h�,�#y6�X�X� ,2k8dbݾ���67<���E�2�D�����w����-E*�<>׼� ��=����w�\�(9DT���q���?h�EpPxω\��GR�|y����s���}�u`=����<Xi�C�iPz�A^�k��o���c�y���?����k�2VRͩ#�}6Tj_�d�/���XX�0�
֚y (#R��ݯ1�G2|� ��g=+`�+"�R�9 7 %֚s\q���T���7������PaR�ky��'��{O��u?<x�HG�0F �\'�?��x���}���H�@/�[���W�1�$�B��b��h��b��6�Ye2����",��-r�;��Z �YS��?�B^	�N2Ec�>M=1z�U��d�n���V���;��olyFU�ݪ cy�E�]�, �v����/3�&�|�����z�e�v����G��^�!W�1�Р�
�6V����괭q!��L5��p�\��ؑ5ε�Z�ڬ�g$t��y���%��Gr
�
^~R8/~�eN�&��'�Hઘ�F��/��a�.������hX/�A,`�]K��P�6EVwp�A���nz�,��H]�\����nwC&O�aZ�Gzo��|i&����.�Ҕ���IGQ���.��4p4��͓)�������z�eؘgg�72s��Z�L�Z=��l\�w�8t�T�WI��M�Q.(E�C�&bf)���{�S��Ac7���傠��M��i�A(
79J��jx�а��`���Ro�#k�_���5�1�k�%ro 1BJ��91>�8��Q�(`<���}g���a^pVb��"�^��hS�؎YT�J^������B(*<��������b^�B�U�; `#�f��mn0Uև��Um�b�[�'���o�/����?u��G�[��V#�*�@E���,�^�V#.{��M��������>xY �DD����>�S�e�a�.��B?���c�ϱV(x#3���x��Q�y������TƑ�zytxp�,�cUdnD����a�'�>������}��/{���� j�{*XC��Zx8�_�����7�6�P���@q͗��^�җ������S�<��b� 6�9w�]c~v��[)�xo�Vx�b�2�=@='�<;�����=Sr_=����9�3.�[�`���Z1��
UJ~��L��,3�6<���(U�M�@��܂����z,�P)(��۹e�}�9(5��1^�e#b{]0��1�g���k��V�0A}�a%d��9(D �N��7���En^��:�����yQ/iϮ�� J94�d��x6�si�?ʃ�4l��z���o�BS9��͛�(v�WS���s:��j�Mw����{��Ro��XG�]���U�>�i�*�{W�AՄ(F���mmXC�!E���:͐I��I�o����p�1	��E p�D�4xK��3V+�Z���s�p��G��ǅ�����(���oNZ]ׄI" �P�&��%�w�	d����DܔpRz�B9�H�jMt^]��k��OK�f�� 
�XA7�h���9U�T�|Nq�|�8 ( ���.�܊����HCp�H���
���n)j]K]�9��FȺ��w�f�j�'����؍L;ƥ{A��}5B�ܩB�B9�BZ�#x�(�Hs����4� h�xg�3,u�Ax��JY�<L�1dͨ/ ��� ʺ1�)k�=�`r!Z�x>�GBb�+���B�%���G�0c����H�-Rd���LX��"l�0a%��"m
�Z��ɚ��G����#��,�O��e|#��r �ӱ��
�c.��� \�14��gH���]���	pi�����~y��y�Z�[[#B��s�c�ߌ���!{��t�y�e��V. �BL��B������Cs3'��S9$�f�W
��H�C2�(���0,��"��b ���7Ts7��3՟ȋ<��@5��BG�m�[aԞ?g�߱еnۍ)xJH�u9[�w� ��b*�;��;μq��;Y��*^!]�(R��$=�M�Z�uSY�	da�L�CY�ȁ4C˼F�ܝ��~�㔾E��s����-�Rf�K¦�`���m���Z�tp�U�n}�uS^�S�q�[j��9㽴�PAw�iq�@��s#R�)4��������q;:�N]hG�t�9
r��ڃ3��d/(������{+��+汉�hk�->	
)L��d�ᘔ��EZ j@��Ye�;a\�Jk���e.�"�.!���)� %iY��?���p�".qx#�P�H�cq�<d��@���XE�*�.i�}*\ "0�p1�k�+�K��t�J�H�y^ayn��n��n�y�	�ӄj�z(�'x������'<�9�m\L[�(9�G�~;���ƈu��%����%.a�����Ӑ �S6�#"%���@E�rJ/�;tV�S煽�reb(HM�P��3�g�K������ZP �f�g����F���jspNq6�mP�P�S�!�j�TJ�Oף����kAt�~�Wq�8���87����#E�\>�'�
_Ɗ��5�
�`�������̑zK��� �8�]Cgq��$/^�BX�� �ג7�ҲgB�"H�߿�w��d�[�"R���Ut���w�W�jע,@@�Z�+!�L�fɅ 'F ٔ����J��H��]�+E��ixY������݉c��!��	���m�u[9z��m��=�� �换��1vc��� ��+T`o;^�t���1^������C5��F�zMM7Cv�7t^g���дw<�d���:ꎃ�ju��ݎ21��?�`�C�����E}ࢼ��,�S�g�`�)^��j^){�S�᝔�%㻄���)p��*Z�hyŃ��Qϵ=��=���L��[�\}~�M�	�o�u�U��[��u��CۀzIT��p�U�믹�?��U�Y]���L��Vؤ~�6�*b%x����ܩ��}4��R���1mڬ���KH�bFμI�
�b�ݔb��h/�b��{��M�L�
A̡��pPFn2�eA�`\�J�E�b�@� Lj�+�A-��B!:�1���:�Tp�1����Z�������-3k�sdPv|VJٺW�4K�����������%��j�x����F�,a� �֠����r�v���%e�^���g�}�Y�c�&�O��c��~��[햋�p��p��gy�T4���C�u�<O�E5K�#���8G��)�z5�A8��{�.�<�����>��-�nCnl��6�T_eN��"�{�$���~� ��9�#����\nl��# �ς���3 �yŌ�a���^ ,�y�L�%��Г�R?*9qP�,8�҈�>P�G��MA>@���y�aw�7�e�&nϲZ����WJ�yaS�fέ��<��p�=�!2o��
�j�j<.���CVUٯ��H0�K+���Ȟgn���a�|��P�v�a���ǖ�3^-��R�����뭰���ɡ��΋�-����{ӌ򪅳�f.W�֪�Q���V��Q�o�&@�V���_277�Z^��<]��2|�e bzf�u[�I���j��]���;H X�x��ٿ��1�̔��^�b����2U��q��7�W��]o��o�'}�AM���H�U�j�k/Mk�e�7E��v0F����M��Jɟ7���^���e����>NY�2��;4 @��2~�1�A���p�<pY�,D䥍�߹��l_t��y�{%�៧�K��z�[�Vy��w�HM��3ͩ�u�J�z�4?=��ھ����H��6��<x�ES�p!�+�+�zf�  `k�Ǳ���Y�pO��S��WlUoQ��뱿	-T6��hl
F.�I*l��	9x��7�&{Q3�ba�qk�K�k���8aV�S.��,^�����<����U�C���n��s�� uS�ۊ19�w�#v��k��N��3O?�]p�y���u_���q~qKѮ �f��\����o�'�ȇǎ�o��7;?g@�1@�C�X�~Ș����%k�P]%aP����X�p5�Q��Q�PR2�<�L;�_��_���>Ad��q�^7���_��Y=��k�c���7 7��=y�����g��*��Yae�c�cU0���Ç܇��#&����9�,���h�t�Xsŀ��	a�j�u�%{ N�V2�ؘ���P߃�u�W�(����}�T��˺$����7�����n@��2|/�ȵ�6��N+I﯅�~����]Sf�Ra��;��/��/n��*⫼�U�
��c�κq=�P���þ��N�Q��T>��7S�;�q<۶,��ls;������/!>���T��,�V�#��I{O�g}ʃ�Y����.����C �by6'#1���^Cc�Ǻ��	���y� �ʲ�|���8R����^<�x���満y�N����]VȔ������%@E�1N'm<�o�f��Pr�VV@�,�,�	��2w��c^�zPX�յc��[w3u�Y�Z���p�H���h�����
@4�e����+����>@%=�ڄ>�#�+��ۀ�}���]�����Զn�ǵ���)������i/�s7m$���5v��0��suW�v�z����Y�F����P�u*#I��o#<hu�56���V���{��c�����8e�KcX�+��8[�U5��B�ne��\�����}��z��>;�7�7�k����5�k��ѕ%���ᵖkyl��:��h����Fm	cw<�M�ϴ�����ΖG���޳wf�iW����/K��5$�Z��z�a5"�W�US�Ⱥ\�޲>� �+�2YO^ yK���J�!��0rTBh`R�E1ay�p����1�kc)�ÄЖd%!`��w�>-���0�*�������I��N��K]��� �+1��G��o�e���hH![//dķPsD����s 
�d	F����H���1cZ�B$�(P,d,v��Z��([>���x���c!��N �ba���=���}�h�P �Ҭ
�$��{�b�y�]!\ԟ����+��zjr�<��L  7�E�6ˤ�����' p%�� XQ�p�Pޓ^��ߙ<�y�,��?֐'��VYُ���3�|q=�LTP���2�1��p�ҭӢz�#�;p]x&:���B��+� �������� �l!�f��~��w���N�~�Gb�gU�,Y��.,j��<��כ���y�3�g�=�x�����kG��qA���2��12 :�yVVMֹ�#��+���]"΋+�s%Y2J�j���{�S@</|F�e�t=)^9I�^V8��k������nt(��[潡سq����=8i��h�z%wk��K�^����8�V�����,�'��ʱ�餯%/� �-W���-�3fg��.?ϳMW�p����5������w��F�Vu���*yC�Y.����vn�gf�$���W[�����B��F��n�r�KQϏ?Q�#���x@��8�4f̂�>�~
^~b��`�{dL	aC������/b�w�ldh��� `ۂ��q��N������n�?�H�#r��:�ro����(��P��������:3}t4�[^؍=����6Zg��,_r���\u<>{�937��ˍr�Ӱ�.ѝ:TC,#nJf|ۀY [$�~Ss�,TH��5�+#����#!�6p)rl�m�V��|�=���	���a�p���)�(DP�)�@xm�55�����{��p0n���2MP�(
�QY0V���A�R�cJ�����B!ܦ<ql�	J��u�\	�S�(�| �!��.��ܨ��U9}�6^��jq�0�,.2�S����9*Z0��R�ʠ ��D 
��Ov�k�� ��YGyg��$�Q�c���
��� kH]�YX�P/�`!m��߸. M
�^���'��\�e��fe��\���>���}��
�IP�
Ӱ~̙2��7q32Y?�NB�rnUF9Ãa��-�b���R�y�h�۹����o����Y�yo��7�n�XXN%���1�kr�!�s�}���H��m�]��3f��<�۲m��E$ն��n�>fn�ݚu&��q��#�����\�!��|�'�*�5M���S���"� �����B*��bY
�}���2��CGvq\B��Ղ�o�6�!�j &ؚyh'0�u����ghݡ{�cn��K�|��X1���7�f�z��W�2�F]�����n�ˁ�v7_�h��:��?���^�U%ˇM΃kk�{��7��m�uѶ�խӍ�ig�u�v��=w��2O,�"KF(��Ä�k<ǖq��;2B�g���'�qʂ�z)� L��AΤ��ih8t���ʾW�O�t�5�̹�����'ګ){Kg�7�5\yjf�>/o�n7����K�{�%�{l˅����7��QH���>�����ܼx�׿��>���O}�|�~Ʈ����Lf�iX0%��g� Z�#8&Xb�;�ly�)�-X�M�JA�Fݍ7Bj�)47a�K!�@�~����`E�qྨc����7�"[���$�XJ--X7�Y�}#�QB��&�Ҫ���@ؐbk�V0���rM�2�R_�q
�Ge]�eW�[���8��ى;��؞�
J�)T~Gh�h�m�Z.�c|�h�s�1^���$�%�E�Tmeg	xA;�?����R�~W��ʪQq7S�(�D�d�㺠Tc];���{D�:m-������5�e9Ph|7M�nĢg'P�
*o�@��n�+�#��9�d)�D�R<'eYi=P�x:P��<��lB�N�G� ���-t�e/�����V��:$x�, �I�'u�f��,59L�^��}��y�u�v;��W΀B�:���ڰ�����}�H����k2�q��17�k��֢�	2��~�m��#�ՃM�>��m{�mN�<��Mo��ypq�	�k��em��LL�f�+5�\S�Z_���8��~�@m�[*Ɨ�=8��w?�x��s�n�Vrk���@�{���p~l�=n�re�����=��ڽ��~p����WF��2��������΃�N���O9|��Y�9���3�j������q+��w�.-�-^o5�ѝ18�1DD�j��P?&��՚����.�)^����s@�q\;�T���j��x�+���<��O7]���^H��}���;�q��?Q����K���/�ٟ��������7��n1*\p��+���M_��mw����������<?��uX�K�Υx]H�#N낇d��V�!���)���M!�yx�����j��l��Q�"��0��	�H�K����$��W���qP.� J(�T��~T�4�� �F�ƑD�i��͝��xAH�c���	���$l��X�&,�����\���$m[�tR2m�H��Ga�����.�`QHU"MӽUa�C
A &��#³2�Ҟ0�.��1)�qI1��&U����q���XӼ+�{�oF�&�7�%)��˗�p��׺�{I K�j�i�̫�=J)��|�����Ջ��l��\Hq�}���B�ZK���Eq3Pƃa*��h�4���� ����)�$p++�8�a�Y��;A6����3�V�m��z��y��ɖ���Z�] ���Z@��=��.ʱ�t9֤�7�m�YQ�������pԟ��{I$��	 ��E�R؏�ʔL�a��oIH�G��z���W}���"[�����\��cں��I�<֎4w�8#��r��[�hH����L�1|��i���V�c�K��nmy�NL-4����>��?�w�>�I�^8��3~u(���믨;6W}���?���s�����t����W*��u�3Oڳ������Ԭ[t]��f���(��V��R�äYe�Y�9sr�'�qʂ�^u@�r�##@R"���H����EQ��,�3����U�n�F������ޒ9��q�A������}����9Oy�����ou~�q\~��#��=����>��/~�|��G�5ϟ/U~t��.RL��8�4
uXj�<�u�I� �s�a�b�2:?�촎Qd��R�����,�X@��g)T�tyc�� ��2O�x�7I
N�G`B���	��@��4a]���[]B͔�pPheO�����%p`�V
�%��\�J���(MM+��Y�j ORY� ���Hw��%�J�j�����H��\�s��'�
�a�ԛ�zX�u�P�ݫyG�uQ��,��Z�i��O�1�V~M��_�)�����!j�uL�z��y�K�>�|̖�FOH
�*,�' ��w�v]��N��t��3�c�a����J&�.�����W K����AD��AM,M ���W��s�\A�%�]`Pi�z��[J`H���>p�'�#oJ����릵9����Z΂3��f���8� �(8Yʭg����k�����%�8~�89�32��2t��Xe�}d�����~o覑�P\�>GpX-LJmT���п�#~L�^�<�|�=�q��-wg����v~�����3����^/�'Z�=��^��+�ļ:�Їni�~�c7����~߽o)M�<c�����]���[;�Xh�h}�F�Ց��mN��a��<�����)^��.AH%���B�h6�s[���+�X���s�.[�wnf֭-/�G���K+���Y�����]������������G�{�'��qu�����J>�`�Q���=� j㡅��OL�cҠ)O�L�\臔�E`�* �hK0��G�.%�G!��2yhQP���G�BJ����,
aY�c;W(z!l{��4�R����l�T����46������Z�B��9$ދ��q��n���+!i��A��y�BOآ�H��-�A��bV/��%�'�)Ӫ�z)l%�C�)�ԣ#e&��{IT�;,�C 0%0����k�P	� FJV�rS,����Q(�U�&�3�F��K�X{G
&U6Z�F�s�z�8d&<�	��TH.(�!��r�D�֘R �*��a;zFa7�g��=@�^
�*q�=XI�zy�6 �"��q������6�Ѱ�vI!��)����<..���i8*�Y��RCόR�9�c�0��?���v���)X����}-��<_�a=�%}&�=A.L�s�7��x<(�dF�Z��y�#�(��i�2s|{0V�	V��_iuɵ:-��Cݔ4|�<أ�twn��K]+6W�涑w��r���#�z[͆q&7�5W:��ꊻ��Aw�����3�[?}�s_��������ܟ����Y���?��?��k�]��wo��c'����׾�~�X�\�%�'�n�ZsTQ��#13`�����	:K�:�:�S��O�ѱ�Ēa��-&]um��]���U73?�dX���
R䪾�ӳ��n�=�{ϙ_x��O��_\��}�G����g���ww��6�gS������wEb�٘�R��'&<�Y�����P�7��گ���b!�ZҩRJ�@�Q�� X�*^߼p���k�P�ϋ�FK�I��N���oRB�D��NDI)+ԑ��*m�z�F-���k��(r��}�T����]E�Ҏ���G����U�M�V| )F�b����d�
�h�)����T�z}�A�(�L��X+F�!a|�.�Ɨz#ʥI��LzN]G@@Y*i�K^��~���NY���z��_)��Ϣ�x�f����qH=W����]|*yL8����)�I !��iO�ޭ{ܔy����^E {<��E0V8��$�U@���3=C�
m��&��>RʱO�]�C�"(���;p�0��e�R�4kQ>���n������R�����j콲ͧ��Ee<A� ��-Ô�B~�ʘ���b�u�$ՍX���?h{�`p�Zssn��~��5gV57�+�2�_��Iua��h�፭���J��wz���;�i��rm�17���~��?��_~ǃ/|�'�����m��Í�����W����n���g�s�-�_�}[y��g���2�sϼ�3x)�a�ڍZP.�o�o�g�P짽�~R���� ��o~\~=܋%�}�H��⼕�������&��ʪ��t��7:������.�蒫�p�ӗ~�1~�+�8����v����h�� �t8ͽ���c��=(BKH�����F6=�0�h���
�)VT�B��J!P��P�E±�����u��v>XQ9�̆*�=
��3933m Q�!�^)
�k�Ht�N�B�0�����"���	�鐅!���iS��!(<#$�k����3!��BJ�p�:M��(�|���:65�E���2Q�������C9�q�e�Ѕ{�;'+���q~˖�'R�F��\G�+�R�SS���<:����>ST()ȕ�Ba���׼H�d[���T����b�b� ��+�M��f|���iD�	����+�j��]���Z�gH�cU��
�x��g����5��מ�7B��2�/�����c&�� ��S���D𣐒�54��
��M���ϣ�E�����B���|�A��A!+�i�,	�i}C�Xx��&cDϠ�
�z���}��$�O�K�dq�l���ek���e���Qxw�p#�D��XeX�}~�Q���c�����g�j,m���7�k�A��3?������yKY>��dEH���'���{���������/.:^��~�u����-9���^����/����3s�듗�]�[,���><v���q^�7�2=ey)�g�q�=��S��*PvK�@@��@��`�W�2l����>�?f�y;]�������m;v\u��/�/���{��+ƿ�7ݿ|��͝a���j�K�mʭ�|z�B_h�dY�#K���!b
=��Y3rQ8Lx&�s�	��	�6u�g�z�J	V{�7��uq^��]݈����A(��#ɑ�"�� �;XH��Y�	�FB^BZ@AYB�0:S�3�G��NT-%覼	4q|
B<��R��M�L`Kݳ,s��46)�t-�p��L�Y�07L��PX��Zg΅7Gs$E$������kl��e�k�RJ��Ɲ�94o'{v�K�o򮌣b��V�2`�z;Eކ*8�#���Z&V��E�&��R/��$�����=ڿ��(%���D�2㴾D~�D�&���Nu�C)ܘ�[ݗ����W��C�X�?/#��uR?�'dm�q�\:O��O�i~X�=O����hJ��J+�0�i��`\�Ԇ"x�&���G1���
%���:�3���������\y>�Ժ��ӎm
�	P�cX�L�J%*�!�7�h8q���FF�^VB��0����(_���K���o�����0�7���~�m�i�c�������w��n��Rܴ��g�j��	�H�߿�R�4=,��	~���e<��CVo���ҹ�/�s����r��y0:��[%}��u!��ԫכ�v�9w]����{<Ƕ��]����k���9+�7��;P�P5
"n�Q$�Z�����k��[�ДNR|�i�1(�ф�*��hUv�yp�~����H56�T/���C�����#��<��Q�q�j4��ӷ�'^1�sI��@���,΂c30���f���Rn�YUh�b>�G#k^�:u����R��@�~��IxoO���y�W�r�w�'M'�X���*��J���C���M�1�!��$�HQZ�O�1%~��!�ν�S�#o��Hu:��ܒB�7�����-�,�Fl�X�ށ4�-�Zh=�N)&�	��h��s��=�֘1���0@�uͣgBσ@�\�)q���0�(�O��=EDJ�N�C�>k��J)��a�o@��`����8p^v4��
`�g�K4k�M\"y;�.Ш57�Ug�O~.�u�s�Cw�<���y߯G}����^�0���3S������	��-���y��Xk����ґ��7B8�i	��t��7�W)F���!*�t{n�������E�ι�����>����8 0�ۿ~���G�z�#�Ϙ���:�4�eC+�U6�e�;� �qdSZp�S#����{��Ì��8,xx9���7%�*S�T��ŪkQܩ�	�I>�ǃ����O��S�~���{l�\r���];��;2`!���b�9�#P�L�m?�I�C��v�eUC���?B�b�J�[�O��J��a�JP�ԋj��% �	�̦҄'#[�g&�!��"EX�$$�P8V*
�����
Y.�3u-p#�^ 	u	>ΧB[i#F��R[D�K ܓx06�w�3�.�@�F���F�HEʢ�d���R���R�� ��̓<^5���h��ֱ�VJ�:;W4�K�ҤdU���t]��/�?�=j��O�]
N\!]K�(>G
��]
�������R��YO���9Lɧ�B�y)�=trƚ�c\��y������7y28R��� =c
sr(�s���)�3�H���;!��Ӆ,�F��1.~��W��^k���m�E����00z!�|0aE�A+��k������Џy ��r�W����y�z���Ow�A�%������J�Z��q�ud�jM5BW�^)2s4s]]]wS����s){Y�����
BC�V6��a7'<�mn�>|�%O��e�]���g����=p��?��7_qtmu�Jwѕ�w��իu��7JAi{�D�V��<��NY��Yn�<�>4+�,)><��ak�5���m�v����^}�����@g����˿�k�����|� K�̄��o��
����rX|�	)�&��<��I�f	fgYV��I�)�4���V¼N�lҘQV'�	��2����Z��Q")���V+^ENU6����N����BB��ص�*�R*KU
C��_�ܐ�zv���A�,*��|�ƛf��{����K�">�y�͹(Bƹ΍��97� z���F��� � �)�OU`4�Z�:N�Sҡ<*�}rn�P
P^^�cW��EYvJ�/��> K������>����ܔ�p�xo4.͙� }�X֕�N��)���R�|jo
2�w�y��[�a�9/�ay��|*.�kBiꘆ�87�K�Ge[�@{Z�$D�F�iW >���a�|�9Ż%��w�H^�_�r���0=�,��ϳ��▎��&��0f��Q0�zw��+՞�Bڳ��s���z|��O}j��C���G��c����n��Cx��Ri����U���>�\
=ʫI}v�����߷B{��&O��>|�td�/�ν��\����M`1x_G&O�F2�J1!aqq!p�jU˨��W��B���x)!jՑ~�v�Zh5�m��.�r�������m
�d�M�:�q�9���V��7���k���A�Ľm�;p�9�=��㥭]�;w�ٿ1.��|���N��q%*zSo�Q�1��4+��oV)� wJ%�C��	~���e<�X�X\��K��Ǻ��䕒=C�vH_��5B�V�A��כ���_��W<΃۾=�4���hPPTF����ɊN�u��t�uђ/M�_5�c�#b�p�Є2e�sHhbYO���
`� KH�Pi!6�	��.�+�	��@�䒧�`@��X�#aAEG`Ρ�������kQVRr
O h���T�e���8D�TI~Wl]��+���|��w  �|�+P'�J�fs�]T�C�3�O�.���𜛤��K��L=C\���(4����"q�*�Y��S��엾�%s�3�|F�$���|��wo�� P�賣���"W<݆Y�(8ZSo���AZZM
�u�馛l����z+ݛ ܿ
�qX��� �+��rS�_��d-ه"�������~���o�w)��:
�{B7m���=��AתENs˽ѫ�~]�}�uӮx%���|�;�5��i_\^����>��E��ƟtsVy)6��9����~�/���o����#��Ъ ����Z�敹g�3�4�0Ԍ��������{߳�1�ꑤ��H�|W�Q�����	w�g�W���b��8���&��;햍`��Zn�z�}g�>��R��[�"�A��Ѩ ̅�/EY�Oj���T�=}#���T�YQ�R��Z��$NO�%�A8&�r��b��]im������.V�z`?���/���Xn��^�=Pʚ�s.���x�JgHi3f2R�4�V�C��x|����8eop���:�z��ܷ:�l^)�b��!Ip~M�þ�zt]�jfY�[[Y_����|��9<=Y�Z���R�����SI~A،�̳<Q����8Reiq�R�)��l$5S���7�r��@�R7!�=4�K��>�����-����@0�����Bò۽{o�te!p�.��PYZ	9?] XS����@9p�.���(2��Q1����C9s]J�qXs<����|�y�>�̭����r��P.��8�`@#�暎��4�t7�����-x{����P;}����|�~FX���s����Z�s�#�����W�ba��
�9>����K735]�_^��C���"OI��qLR"kZx�h��W��Y��|��9e��b��(9�I�]֐k(�����/�3���J�s�.�&�$B�sX��H����+�H>S��n� �����Tknֿ�Zk6ο���7�ގ�0��-`���,��R{�g��ΑWG��܍7��������J��f�����կ�o�tc�� =�«H��c#�s��5���[�t���7�+G�����Kk�`rM `@M}���e	qo\�����#��^���y���7k8���η���M�-[#���m��	pu���l)d-,l��s�/rM/;�b��r�Hr^��W��p�uk�/�����zӵ����ۣ�T�֙��=��l��2����<5��{{j����w�q�R�%s�J͵G>��9��1�Oa%����3vO��/�zeT��4���Ay��d�&�J�yhnH1�N�[[�J�N��}[�2����{|k�աUX��),g��Ҙ̢0F+�dcD0�f��R�˲Hʚ(�,1aS��lya�gΈ�F��n�JRc�>JY��P)Ek$�Z@Ϧn]��s~��~@i��d�]���|��;(**B�^-j�'N�Z�
%J�f��+�o|��� ��V�e�w87^�E7b��,���(s�F!�Y�G��5�y�}�s"�Q��G�������M�
�(!��}<H������/��2�0�L(Y�(_�
K���>T�Nu4 ;X�( 8 �2�}���5�\���qs������a��=��L�%��u�g�d͑�OF�l��<�(���e���}�֐{ ȰfxA�;���W���O]���aI�k�#�݃?���hB����мz���(�p˞�P��}
xHq~�{�j�x���}����f ���~�y�l��{_����_��)x���gxF �a_��b?��J7�7����=�'�s/8�?��=��d��s�� ��h����y ����N���^ok�� ��N�Q�8tȮǾ���Y���cz����2��!��
��X_�{#����n���Ϧ{Ƴ��v����X�����eU7y��Y7^.�����,n���O4�����b� <�ah�f�B1��3*�g�0���M�x���ug\�%ø1U�����I	�R��/�7:�R��p}/�^�7�S�4�Y��\���A?p�b}�!L��h����UO�Bu�,x�֨���~�;��U��Ӓݣ�q��(�j����f\s}գl�k��zk#�hw��?��;�}���+x��Od��V}qq��=��f�ӁU�"j�|�7�G��W�bk��.�_�ܗ��Y�y�?
�@Z�8Y cb�C�����jVx�xh[X�k��nكn\�tn@���3�F!�z�x8k-w�����~�3��^���������Z�����K @�����H�"3���\]^q;��p'�w���]��81����B�>R�Ĵ���@�荍�W�[�y.�����M�Ry����mBU���g	�no4�%��\�e���?�CS�㮨Z�٤H� 6Y�'�(�L En{�Q�R��\$�j�]���e�]�����9W�nq?^��י��_��)T�3p���s�����2��,p= �BJJoM��"�*L�����pa�_��Wٜj=  �Ї��{��K�d{��k���~�;�i��Z.V?�������g>ckD���$!~�-�5��<^x�E�3:����F!1�0�~����*!��؆[����P�<o�^���{�_��6�_�{-<�3)�0 �>Uw��ԧܟ�ٟZ��y�m�63/�fD.���e=>��O۞cM=����n�?�[��6ST��V��O|�������7��t�dz��Aw����יGĈ�x���bf�	���#�>k^��W���	s���u�<�~��a8(��{�6��e/�y�䩥-ޘ+?���/�������k��s�vר���m�Z�F��h}��񾔭���܌���v5��ft�_s3�Snui�֩9�p/ۦu7;�tc�ns��*^v�}��iWo4]��dW�۱&��X������ڶ��p�O�q���W�s�U{�c����edtnٱ�M�<e-[cƛ�qW��^��mB��ǤyTX�Պ��7<�����e8��˥���y^j�BV����o�N��xJu/(@�3Ն1Mwp�+�*��j����n������t�ů}���kl��[�__^9�?D�Ss3Y�+��`d�(�l����{U�/��ʊg,W�P`��e� �#�O�?���w�Ŕ�R6����a�oD3����*�qb6��+%��D��	�48��c
��Hp���w��MuJd��Y�"��ϔ�)�r���bF	��q��:MS���s�Ĝ}^��[��X*�%�'
�� 1�,��:J�uu^^�� 줕^��xE�6Q&�28t��i"�权q1N��"5�$e���TaV���v�(S7�O���
��>�@��$�H��+�9��(|֐У��N��^��;iUX�o6�{�N�7 X�x/�>�`&������n����}?4�/� }�r0?* :��}���	���/��Mi+dƚ�Y��/��B���X$���c f��9�};Z�G�ՊRؓ�+�Yi�ϔ\�uyn�����r�d<�������6v�I��YU�����C<Xx|��X5^$��s<� +��]sd�w����9X���7����lϻ��<��Uk1V��=��
�U���O2����TJ�}I���mD���z�j])y���mw1���5������zí��d�:�H
����:<���'����5���e��!�ǎ~�����O���q<����_�/���wϞ�S���[K�������������W�8���ƙ׍c�o�xꂗN'/�K��U|5ģi�X���1֤�,��EH�>EA$��+Y��������>���������z��g>.(zy��֍����a��V�b�-o���t��f��E*4��6]2�p8*B��lRT.���c�&�6vz>Q�'g��Ri�|�x<$A<+�R)M:(��&�jZ;E�L�*��Xxa&�j�hLi\��!PQ~�F��J�Vd�l�4qxB�H9z8JV:���Y�����;�'�+�&rb��4�@�Y9��*�X�(je�ȞH���Ѻ��YY�"�c�k��ݤth�T���#Ҕdͧ�I�<�)و��4u^����o*�&��PJq�� rR�
/*����"(�y8�=�"��g?�Y��ҵ7����ޱӽ�5��T�k�k6��o�%V��WI��k��;�(�#@�� H1Eo�5ee������R�ٳ�U�~�{���}�jw�]�8�/�A.�3���Qd�Ԥ0���=4ʰ (���/V�v�EA�I���Yf?�̛��׆���z�����X?疖��{_�J�f�; J����Yܺ�n�<g�0�7x��y�]�ʋ��)�AD�d��� k��-��w��2{��4֍^K�m�T�i�P�nl��g:������(� ɤ��E�㺽P�y����dl��Ȑ���U��*�dd�C&����u7��70+���?z�]w]�����&�?�q��Ƕ?��O�:ba��îm[]Ńz3\�\wx$��" �@�ǋ�����'tȈ�/v��9�C��ް��x��<8���ּ��x S�7�5����&�֧�F�S�?�����/�w������C��W4���S���Ξ�;h�?���q�!����4������SU��=��9���l%�H��=Z(C	�j��,�����N@�d��p��jy?~XB�C����|��O5.M���H�rw+K!=԰M�qA�9Y��D�7@5`�)Aȥ�f�knr1,��E�4w)�T�-�Ъ�<�H1�5�{�wB[�P&E��B+)Jc�
3��iq-yRR�@�ư	�FP����őHm���tt������ f�#�����C�qX[<X�|P��/�z`�+�k�%(kʹ��&1.8���'��>`��o��^�p�.4���AX�}L���?K��,��R�	^
��������\�~~T}��ǎO����<s�V�%��c�k���tT����kfn�G�:���p�bj8�+�*�$M�-xK�b�_�E���K�K8T\�Jjt�'cU�5������3��r�N�k�&�Ț1F��,[0P���y���j߾sl�!���m����e�ժuN<�.�I�4�-۟��c���؃�y\��(Veu�J0�s�����TK� ��X�J���9��^�����<窫n��?Ï�Z&ʘ����:{m��S�qt��LH�����
96
� �x�ٓ�Z�R-���8���?�1%3�Vv�[{��@y���C>��a�w���A���ƹ�)�u�����˾���~�c������X�����G?p���?�Fo��6?3W�tzVĥ�m�c��ڜD���y+���+/�!�bjܝJ,�m]R]p�Zv�0fE��e=�T�ݔ�4������C#��aw��as�o߶���PGo5�JR�����P ո�ׁC���
p���/-�-@P��_E�TWD�A�HS '/��jH���O	����	T����
N� G����[��trZ��I�8=��i�>�� ��

Wi����G~X���@�s��R4(���F�!�@ "*�hҽ�ꪫ�;��c/ 0^��׻��Ŧ�t} �E9~�c���/��/����^�"<�"g�&�7G�*�c3f��c�F
��pm�E؏=ϼA�%����_��m����l�o���bn��q�ف|�\�����o%�	�%�,���u�=�U�^z�*!���> �=  #`���1<���� }ы^d\�?��)�]9��J�-rO��g�B����L��������;|�=�-a��pZ�s���%bO GN;}��?�����F�$��l�T%�&��c���hf��@�e�����}Z��7��2
�*gj�wSd��*�-�<K+8u�q)�|���n��o_y��]�8����������VW��:=U)�	v��������5���=ec����>�2fޢ��!O���/',�YY|@Kt�ս���������#�n��f�V陭�G�^��i�1_>r����v��w��u�W^y��^~��(�s��������r�y����4ooz	��
Z1�:�Z��eZ�ѕ�B�n�K��@X��i��X�R�i�!��*�"�R�V
��ŷ��'��T�V-���@�N�I�})�aR�_��R�&a�̕<Q�|G@"��)��&e��K����F��� ����O�~��U8B�G�4��2�j�=*5�yD���Ұ��;<��^�\j;7��W�$���Q�}����c���^uM|���Ki���P�(�(,`�8 �GP\�a�,��3B���V��B(���f� �������h�yW�XZoR���C����ǀkw�O����A��<+��|��iF��Rjž="X�� ��q�ݿ ]�b5�gYUj�Gos(���&�E�	����z�jj��\  .\��D���I�� <��=��x.Ժ@E� ]\�!o$���$q� H̬����咷J�r��$]�?����<X�xƥ�3tؓ�/�?w���ɕ��Z��P�s��y)���GU��ꦲ�V�U��Wۃ����
�y��Qih�W���������#}���1����������_�Z[v�~Z�{˼[;~�5 Wؼ�n��ԁ�-� ����yx~�Py/n��,xYkv�q6.�#�eJѫ�G�Ͳ��m�m��ž��o���[ݨYw����z{d`g0� 4�v{�K�{˷{y��G������W����eُ����G���Ϟ}��~ge8|��m[���CЌ:/9�=e/$��Q���������5�S�wŬ<�ƺ���NbsE�QT�.��*w�@�~�IV�*���#�PϺ�Y����� �
%_�57�8xQ�)M%�P��y��1�!"��߰*ճH�D^)9���«ơ�S��z�d��@PZu~�SϜ�T�l��u􋐌pa%�ёv�N��⟠`S�Q�1�xNn��)䤹IV*/��~N��+Ú�� ���*k�N��1n,x >��c�G�dSƅ��#���z���!�X��~�(z���f)껢bW"�4�ICH�k��6+����G�~B��ͼ��#���~��D�g>�w啟t�<���{�A���<��:y��h�r:��C�r̔���-C�_S@��{�K^b�ŭ[C���a�A臰.< ���7��<M���F.5Q�Y��Pkļ0�\@�e�dq~���(�a������jx ������L�x�m�: ���`.�-�/��w��nnf�䙗����N��B�����T��,�ɼ��M��e�X�Ђ%Yv��=��V[����B?�A �m��BX~�z�ɶYU���3��k�:�K'n�=��e���9��k�p�������_�}����x`}��޿����~Cgm��]��ʹg�u眶��}�����sC!([��J *��f���W��E��i����cn�����+@P#s�P�y�j�����[��0r[�g��k�Wݠ�q�rf�uͩ������ܣ,>����C�W�ی��򉻿��+����y��w�~�����3�[�y^��_�q��_�R	��@�
�����dՔ��z�/(Z<�^��q�,oS��^��HI�R0�˿h�{E[�J�Ä��p)x���#��0l[���(�����{Ƥ��)e���Y��L��B�LPu[�_	��ϫᜮ-��8fi��w2(�R�KV�2'84�W��S��ƌ��b��b�-e&i�:Ұ����IA��&�^��=��ƙ6���yD�rDɠ8+�=��� �@�����M�CU�O���V���Ⱥ�3��^�7���^Sgh<z��Sr�H�JSg/�=j��EYڋ� e�q(���-T5�tYzz/�H �5-���
sV�f����������̠t�|�9E���e�g�7$$�z�	�?R�F��ӌ�������]��mҍ�}� �v��s /s�6|%���׋�@`��y�X�5"+�24�z�^`ua���\����o 򍗿�H�J-��=����^�x<2�h`��դ ��%<(TV��al��t��v5/��g�>FCŕ��x4�g����J�B�Aƴ�3V�h����jx��Xf�z�믮�Cߦ,�l�_�{��o﮷f�VW>�u�]��wx�.�����o|�ի��؏~j�ܢ��A�B��V�8����3��|��C9��m�2K�"|d��R������������/��C��v9xʰ�r�� ���mx��n��3v�֠g$�3vm���8z��n�b~27�f�덣��O���;���wv�w���ꏮ����k/|����UW�q��������I�����Y��,���٦�9�~�M{t�<R�S�����^<D���Q�����U�UPu�~n��x^�%}?�q�f�U
N$V�R��ļ��6n�+ԃ	������&&�8<��N�v�游ղ6�1�l�����U�J���W~+m�������R%!�!�HW$�����%u��x�vӷo2�0�iT�E��/��E���()�#n�B6
W�R�q����sѢ�^N�0N������R�M܏�O �����`���ZK(d�ZZX����K�y�x�~P$��	ՠ�XkB4�L�<5YdEs����r��+��/6�l?��^��Ľ�]��č7���;�.�����=��3cZg�qi���Rһ�3�`a�g��d�$K�2B����e�Ga��
��-���C���^	��s}�y�ȣ�F%����-��\b=rn�񦸗2#�2P$����[���}�;��BSV,�2�_���sB#���Dn�ڄUX�����tg�gc�}��LTj !�a%��.K�mi�S��k�ؔ�����OR�	��xo�,�]���	կ�7����Yx��ҤA��]k�����qGhK���pMEi����3%rv�䊙������� 8<���]o��ˑ�R�����B����U��u���q��nwid[��f22��Z꬯�u�;�^���ͻ���� �X��H�����lT�;���k+o=���?���������z��O=r���|z��?����_m���^vx�#�\��.8s�;c�V��lX0�(�G���ǒ��N/���Qo~��R���|�)x�I=�.E�*gé�d�[��4�����5�"Bݿ��~��G���	��z3;m���jk��9���G_sC}���_���x�+��8��_x�l��ߵ�޺`��ы����j%��W��R��y�6��ڟ�>=*}���^8�
��K����o��� ��h ���LB \���ع*Yi�%n��Q��ؓ�
K�0���PhE�V�A��-%Թ�i�<(I�sy[8�v�c�IA;�x�������_h?�������|yG���T���a/�pZ*�qJ��\(��@�R�
���U@�����PQIsƩZ )Kq�B/�Hf ��3��
�
�uU��{��U�eq]�&��0Di y�P�X��S�_�<�T�jH8��f�) r��'U�K!�3�U���P��9�">��۾QRjͫ��ZḎڏ�B(�^�,��dL�7���g��}Ӊ��5XG��o����JR��%�����=�S h��l��\��X=[���xg �?YO�݂?�R̕}��(Vվi=��áb���EP
h!|��  `bm�Q�N�����j)���#���<R���j��]��������V�;��~b�q@�«����7a&@���(>������UnL�[a�)a����]�|�	��L#�S�i�7nT7�x¼Sx�J1��M�� Z0(��y	�?�j޸�+Sf֕j�m�����'K`-�,��Z��c���V�ֶ�{�]?z`�m�ܷ�+��wnx�K_t �o��� 9t���[n��o{���wɑ��<{�<z�����ӹ�=yq�]x�^�zã]om�&otR���F�{�5�ߛx�R�c���������?�qj������`S[�P2v�%�� `���/nkí<�n�kn��/lN����p���ҋg}��+h��n�y��q>���Zy��^y�@} ��@�Z9����m�*5ps�� Z��pY��`��AU�:���f�W�f�YO&3�t;�5�7�������F�>�c�`�<	�y���c��d2na���%x�dav�m۲h��W�8+�ٲ�n�QL�����h�bw�
}2yS]��!�2 ]�>1��F9m�'t�]��6Pd|���'�c�S�4
o���	�_����^��Oy�1+~Ϟ]V�WcT��J�2�s���@�S���̓3��e����Gp�i�
O)��:l�s��]�� 	,Se��P�^�?�zA9iN rX��3J��f���D ��TPi�Cֈ��}���E�=5���'F^#݇�)��R������W}�zh��n#�·P(p�E�A�����p�x�X�k>�yw��!k/��B_��s�A5�S�ؖ��pw�v�{�������Ȫ̝��i߲9/�k�+�n�0����ر�=�)��E��l��;�s=P<�-y���۾�sӍ�WQ��z�A|	���;̧U���͐��^�z�X�L�{��(aG��C�4����9~}i�X욮�ci��cDݯ%�R��:r�<�iOq�����q{�3/�?O�<��i�=�������ױu�Wȼq8(3~���w�۳s��[鬸G��;o��yj~�Y�vg�~�yLe�G�Ƞ�=?�Y�͓��B9G/��@�īJ�+�0������uuJ�xu�}AoP����E����Ckm�=i�a媣L?��/�M����l�OO���۷�M���<�������_�У��կ|�����J�T�sP]_]ݾ���w4ﭺ�i���L)˛�z�|��=�y_��߹������׶�S��i5"d��\�����N��W^d�r��~�y�I<3S�wɥ-E��Q�[�#���yW�e�6�#k޲��懥z��jθ�ꔛo��t����M�ix `qsW*�Ju�+��̿G�i�%�lle���(W<(�/��X��!ȼ@˨�H�r+HW�����4P�"�0�<�IS�s,�%�E��Mj������+΂KQ9��	�o0�bա�jk\ҜOdPYA�/兗���=�qt2 hT�2���T������5n(2 
DY�X|d&����V,\��D|E�a%C�[��C9 4�}�ޞ�{�� �-D�T��/�	��C2�E�8Q0�uk�  ��D,y����DM|>���0�����6(c>�{(p�] D�F,�x	wz����p�{���V�<��N3�x��`��S2h N�"T^���>����D�ͅ��!�2U�35�dM���k�A��Bu��x�����3Ľa|��e�x�c٧ �������|�C��1wd�Hq_�g��a�'������6�k���}��ސm�Kx��D;ֈN�6|��~.ٻ��4�W�9ٻ�zγ��Cx�Y��Y82��Ik
^��ܪ'������q�����tm=�"Ҏy"�y�{�@���y�����ݾ�3�)(۞�� �Z#��`�Z?�;�a?�C��}��.��%�j���B.�b�\r�P��/=dӊ��e�^��p������`��Gn��H� FH�U<<���y U�U,���2�gwja�z���u�a�y��� t��A�:=JW�ꥅ��L�њ�,��|�P߯��R-�����Z�Z��ԫ��p\�iԳ/C���?�'��v�v�Kn��G\ك��W:�<$x�>w�l�`p:+�W6�d�9lJ�X�?/?��b���V�G�r7.ǆv���
�r�����i-��a�?�s�nvk�b���y7�Q�b���zm�Ŭ{����o�j��ь+֪���7�+��9�Q9d��P��V�ys�Ն�}yk�p eR�,�ɺH�.�Yx8iF�#��g����7-�0�B��]���p4���5'����#9�(������!#��0CAXI��$��>O��X��Ii��E�˱0�2��.<�ߐ����e���УE�V�c9$@Q�Pqi�������)��tU#�����F����B�r��Y.T�=���5�-l�ȕ�[��]Vt�6p�M5Z�8B�����7�������/�0UG�J�g���ɑ�E�X�Z�Ca)�o93a%�e�������+��h�\�Oa
֜��^�_(����V!6ۓ��6���E�_������{��ۮ��w������Oߒ ���ĎFP�E.�q}�+˲ʲ����
K���^��R^	h)�<
iBbM���$�����{���g�9֞{�D�U9�����w�o��k�9�s��������z��Gk�óR����~�W^�Wޭi���գ���,*α��[��1H��|K=[�  )�d�_�?��ʚ�������+_�27������	K�z�%j�!\Y]r�|�52~��g��>_�E;�v�eEq� ^==����c��$�f ���9��̹9}M��s�\��v����8����yl̝/c	�Φ�BV�+'������x�zx�\�{t�7�	�GM2������4M�}A簆ËZ}f�*�w�.^a<���0o����ƛ�Hwvv��˴�~Z�#���$
w��6!�<�ʺɸpkk����Z��7�Y��<K�:���^�Km�,�y�j�J�n�u y��e�U�=�Ք�5W\ꮹ�Rw������㏺��W�gHm���T5�\���#��%e%�;�_��?���=�ˋER��|�$�"�J���M<d����-��3j�>�%�I�%��i/al[nq���d���`���(���������fb'�V}lQFʋ�.½7����벎��KUx�@R����B,݃�YQ�2�b�X>î=��n2� E6�6�g��F��2+x�3!4P�h�1���od�Rn��!�Z'����zXB�9�o��8lWhY=�9�~��ik�K�����<��ܼbX�l����q>K��2F\�o,�&O��C{�4��M]{�n䂟�X����YYV��C��p��h,�,�|�vY6�H@}K�@�SQ��|Ƹ��ZPF�6}�A10hd߸(��1{�16pe�ڀ$��� r1YE��j<Ov��7�H��Z1~x���U���{γ��sZ�@3�xv��:�0�x�z���-�B%f�ʭ�0 #
@9��}D_ixM �˹-�ȸ����W>�^��f1b65��>��7�;|�Ơ�W���R���jY��sVԓ�2��G�ژ�ڼ��0q~ƣ�ؑ��|��Ң�h[76��F�@㵁���x/Iӝ��(�D��υ!��X_(�[i��>�ESE��N��v\�idm?��E���?�ȋzH��	�0se:6k��5�T$.�g��X�;#P�;P�ɹ�p��v��;���6���:�K'`�J$^d5�H~��� ���x(+�����>w� ߃�rѧOo����u��3�$؛j�<;s��ϧ�}=z�cf�5��*��,x�`��Oe@�ՠ�&�l�k��_��t�5A�mR1��D�S^ڮ�4���b+�Dә9;Y�UMq`�#�՟9�e$�N�x8p}\�ī	���#ӄ�"������8
�I� S��qV,�Cք+�J�E�A��G1K���XK���p���2V"p�?�.�V�/<�h�Mʳ���BQ�37���a��m�7@+�g$A[�Y�@"��y���,j��-����iJ���Am�!2~��B���>/�i�>��d��q6�D��B)���5�V״إ��k��ɚ�ȳ��Z����,�\��b�KS���(���}ˡz�eQ�4"/F���KA6���y�s4ҥ	�qĞ�!���of��3��?㛌'yIU��!�Y��/%�G�I�!�z��]��|���8,���=����w݀N���X��ψ�K�>����U��abw�7�*��<K���4���>R�n�5}Μ�>�=��n��
-��>�i�ɽ���xWem� ��9]��I��1��%z\_=�y%d䥥�N�0���g N ��1�llo����5�����i�I�	��ߠx!�c�{ ���hZ�3�� �iB�|���qi�֚�t��
�e�Bkɑ6)X��&hO����|o�ק��[�q�,`d9�����v��M�Fo�mu��hqA�M�6��%��E*÷�@�J���|�ǽ�M�v�M��p�2&��-���0��r5}N�{r|8δ;���g�Fn��CTj���'�qN��f�Pat4T�⦦�*Z�Cm�A�PU�wv{.i F4py�/��+겫�Y�Gߒ�:���
.s ��\C��%��,9���s&� ��Zݵ���s�� <�!��i�lN���0���a3	@M>
d�ԗ���p2����'�_��j" ��T�b���]�l�
���ƣLCF�� d2u�uJ����?��Mw�,\f�L��R��+f�-�X�1VѮg�S1�TJ�*�]�획c��˱ ��`�T��פ�,�ERޟ`���JԄ&Lc����x7��[W��8PQ3c��O�b�$�@d�h,4�N�k͘YJ���Ga����i����\�%0pjP3~¢o#K�5�KZ�Yo���%h�5eF��k�5^�����U�{��	��i��'�tq�s0��j�'c�A��)�B� {V�F������W�����\m2-ʘ���i	"�j��N����}���v;{R@gD	۹�c�r����0aH-���\(=b�Y3��Xs^��-k��@�طt�d�Rk�/,��F��`��dsO�@2�E�vZz��y����-�.�Up4Y�Q9v�i5�X��]4���{��+�M��Y�-9��D���իC�5�E;w��Y垻 E<tkwG�$�j��­�sY^q�ZK�/���&]x}���r���������H�;棐ٔ�U9���͖
�%��%���6ݩ�r{�w�����[;�Z��Un]ǬO�(N��4q��z�[��^�*�ڝ�<�yy�YR4Ӫ���%����뀛��5�$jLj��W�\��s_3zF��� ����Q	
��/~���r�P�/Ff0r�r~�tQ�ʢU���MՓGQ-F��'���%I%�L{w`�׃*�E�������JM�\�V\w!qSYPe�k�I[�t7��YA�i(.�Vv�	٥������+�VTu8!s ��1ji�h<��UiU�F�^.*e8* *���kŨ�����,f�]Yl��zi�lW��,6o�aKk��ȶ;5^��F|u��r�30��g��*���0JjiF�@+��3ڏ����Ԃ�Aݕq9�;��֪f?���2��=q���ζ^C���`+�A3��33\�q0l9�e���K_�4Z��Xb߈�:͂���dN��~�W16�b�0�d���`�!�.��J�$=�&��I.@Jƙ*,K���=�߷_��@�>�J0��qq �/�~�=y�J�h�{/]�~�3��`��#��	�A_s���
�q�Ӳ3na��-���
�P��������{mEYL����a�,���a�~����<��ղ0��;���������|�!�Y���� �Zګ�v���{�V����:5l[M��h�eͿ�mU�t�����z=�s?�PUƸ'�[�Ӣ�e�D�������2"w�--Sc�dM�o���Cx(�\����1 �h���Nn��x�^�i{[��e�%P��d�Ț��4��Ɋ܋<��E/�����y~��3���&^;��x�W.�N��^&�]sW�;
�2����5Yۗ��ݒu^���m�<I�$�]�0����� 0M�l�Jw���8��A��b������dc�1��V��	��?���� [x(ۣ��3��"&�����T}�c_}4���إ�N(�(�\������E��]�lgz�g�0J.S��؋`�C^�SFF����!�J��;4\��I]"�a�5�T
��,�|v(;�lX(�15I�*$>��t�$��3|��&�ʽ���qw�iך���e��{e�sq&�yS08I0�,���s�$��'E�8�yw컦[�.�]��:m4�P�5gxA�O�"0�w����q�+�&��D�QDn�ovh�ݴ��yc�E�̛O�_F��1#c�,'/�[+�B����x���i�!����x����خ�üJV:��L2w��ra�:<��m0���e���n�j��yf !n�x0�e� 0?zC���2ݱe_�خ���z���R�Pǂ��J݇�$�T��1�S�D_O��1��ƚݧ�6�F�
1�!���0���zK湋�'���c}e2�w6�m�ٜ��ڭ���ܳe:y��t^�ܰ����o1=Odli�e2U��T'�'���!J��f~M�W��}D=Ŵ��/�co`_Ƙrk�	Ԕ��ڨzQ�T��<��@g�g���
��&�iH����<�lr[�ޚ �<�r�ΰ���]YC�[>L���jD��\"㔶j�U9��0{���d����sU�R$�PG	��(�0&c|2����@�Ti�s���%E�\r(GO�GWg���8g�˨�\� )�Tg��g��5�lRh`-�B\w��Q�A�Ti� ����� �A��d%O�$}���ᯛF�UH$Fwj�
�L�԰�󟣉�� %O��'�Z�!�:���ƭ��n�:-��n^=+�JP�l�<�A2c����3��^%����� ���cB�.Va�M�2�`�e���T�׈]֤t�B���7��1��}/�ӰŸܱ��Y�c>m7.����Lf�e׳6��Ǽf b��ec1�����Ռ����b�ӬY�'�I��Sz|9�@��R7�Eٽ�7�v���K���b��N���	����ػ�0b1�3o��XZX\.�.�gB�����}X�9,�� �	�1o�>�sqv���փ����@�^�<�>ƴ��
�=����0��w��M�vm�ִ�B~6>���{��c�B�6~���U����@�~
<_�	/�J�'�r��w�)g�kø!l��+�ը�Y{��������z_�<��t*�i��@��a��6ʃ�Q�$�ƻʃ�́[���	��-��3�����xfl�*�����
0a֨n�<�����{w�Xט�kh��8Q �����+w���\���Jo@L׹�PF�4���6�]��%Q>f���h]a�vO��/�J����k�T���WhV�G��S��H�0m�.0y�ЇfY?H��y]��LZ9�Cc��� -�9�����;�7�O�:D��� 	�x�۔�R�We�yc��K���C'6�vi'?S�d���gP�nl�����;&��Z��<�t�ni�B���{|�<�Zim���l2�xX�n�r�
1���;�`�3�[;c1��s��Z�9�{ڌ��Y-,�{�}���߭�iJ��mT��U���x�m>6>�+��?�TY?F�O����?ph�;֧6��,�d��<�����c��<�k��lJ�o�� f#Z�<
�2�v�͒(��8���'j��5(�ixU�eyR��ƍ��J�qk���R�r	i��!{Vq�tgF޵�l��{{���<NM���vX���j��a����Z]����1g)w�U��ywi����E:VRB���d���?�i=g�f洍S�Ӏ,�7��C<���r�&Ғ;ca�8��3���,z��i����i�����z$�'�j�A<ʢ��k�iE_�Ui�m����?{ ��b v&�9f���约�EԱ[M5�c��fᥑ~[�LF��Rx{�:/�ҩ�<�9����+�𨜿��!Y`��~��,x�/��Cd��*�1Ɖ��&Auv�5Up��~( �D&�D�@d��%"������o�
?�i%,�N�T�r�q�+A3�҂�k��D��y��U�O�/�)yLzPxR�4{�VՂ`R���6�⍳��xG2o8��iƠ`���%�дid���`�p��қ<��+�s��*�4Ůg;~S�<�(U���lޖ$pĞ��1)1f1�/7�7�;w�b�ݳ?��/>>�U�6y�e�%��X0�e��8�]���5^��D�H?��T���Ynq_�aF76j��}�f�\3z<?Hú�a�f�Phf�VF�57�]��??�d��%�<���j�g���,&Y�[�=<������ S� M�F���g�X�*�H�v���Rњ��Y�����J�4�敩�3u��?��y@��O����~�2a���y([��K86� 8�V���T9�B�ծSzQ'��Tb��p;��1���Ebc7h��Zg��܇v��aV��tv~���.���ʺ�7�S��>���<����s-�-m��j](u��h��J�u�g%�����q㚷%�T�������0x�XK�ޏ�Zy�:�G��)�V���ˢ��2ҾGJ2�y��t����F�EE��T��\uxj(��ެ>^���`�W�G�4�"oT�m�$�4�	Lz�Nv_�BC6:ü���YIg@���AT52���� �a�K�k6��('U2s\Н�󇄶4��܌e3W���\l�$fa#�5)��`#�"ܺ�~OAPl�c��K6�Y��z��aA�#҅�q*8(��x
���-�E���uq&��P�X�N0#9�1���x�����W�V�;^��}f�cAL���ϲF��4���}�mK���24��6;����̃:;ϼ�&>��x̘!�vZX������-C�E��E Ȟ�y�,�V��I�쫢~j�g=��$ h�eKY�*��!�
YV�㺞SEXC�gCV���r�1eF�L5�N�%o��XU"I��ߤ�=U���K�a=r峨�l~Z�h���qs3�5��p�=��0�ۏ��+��T�q`������xMB������,��ƧJEhX:��2Sh�MA�+�g�4�k1��{��^_;�To��ʽ��C�j"����
^\^p;톮�:�C��h�O�$�sI(�X`�OeT�%����([�eb�ʧhs%���H�ޫC��rk��y���#�6��K�F<�~�ͩ�&��Ś�YS5PO��'�1�+�Ѱ�">V�/�u���aw�J���Z)��r�T�P����r�)7���xRCJ��0R�ȗ��zz
�Y��������v������-b����ʦ)�#��*gQ[lh���Ju�S����l�!��9�4
�@(���X�f�h�^]( ~��2��xW^�Sُ���'6���ތ_���VD�"~��k^�8����c>�{�^�r�� ,�P�xMas�<)��u���E�%�8�������X�T�ߣ}���|Ĺ���e�S�y�|�0K�>�R�ѓ>�,��!��R��.���=������s��l
����AY�X��eX��B����κŮ>E�cW�y�f��a'9��u[�3��ơ�v���������U�i?��ȘQ�M�x3d�x��ES�O��P��>A�{���Xڲ��bO ��:����e�9Cv�q�������,�k��P��kRl�0�K�J�Jby�N�1W񙏴-$��3�I��i:?�Wcs4��z���-~V6�u�@�4���Y�|���U�] �z,������ֆ0OB]�
�@�Uor:� �
�(�2��J-�*���؃#���dc��� 2�^�I1�xn���TD�xW��~M$<�����kϢ���e#.X��V��ғ�8g�K���d"`s��Q�SE�q*n��_%�Y(��Q>V�C�@�qV(Z�Ҁ��돴�\ɶ��>�}ܖ�V���_F�:�)��qa�k0�j�83E�C%�B' B	��1UտWe���4#�8eQ�g���,x��[�l�2A�<�U�����\x(Z��r3����yal��v�!�iT�x�ٰ�)�Ƌ�1�Ů5g�M�q4��a�QbcR-�����Cg<���Ƒ�67�Ӯ5��{�]8�{��۽��g܆xq�#/q�|���7�c1����Zؑ��	0�9��3�10c��H����K���K^��C���T�7SV��� �J���".Bv o\������WL������|+ ��q���e��116�a�,�A�:�  ��z]ԡBOFA
� �ǋr(��b2����Gm%�c�(����fx)?�*0Bp���c����N=}g��Vٞ��9����0Pnm]�{FY�f�F�'/�ڜ�sk:�s�`3ϧ�hV���(�Z��Bۜ�9P�T��F2CH��=��Պ��VI�B۷w�\���@� �Ǉ�p&t�������D6md�T�z�ԋ�����~��j�Rڦ�X�����K��V���њ�?iF.��@�vWo�!4��4����pw��^Zy���D<*��l�&�R)[z��f�W��`�C#c��Peԕ�M��K�Qw4�
���s,��ˀW�w�E��@q(�!�R	��q�9p�TUh:�w/zZ9��)�
��r�ja��N���=���6]w�r�����}+S����i_i�Y�FÙ0H�(y#v؁;�DzG��r��=�4CkF�$�.�j�^�]�g3���*������Ƙ(��K�V&eOɏ�b.�]��U�gb��h����O�/������;��!���ߩ�	;U�9Oqna��ٿc��WL5����� �?���ݦ�j$Ӳ e�3d,�8�F3��R !�9j��S2���u_#���k�a΁,?��h�s2P2������}�#Q�߫���=튧i;(�������J����#��}��9k��>u\��x� >�ZO�3��$�%�<����ou�}�{��i�{ p���h�a��yG��z2}BNǷ=s�(��|���c��9ډ���v	0��LA\k�B+����^k���yg�ֲL�����㢛.ۀ�������&!΂b�LH)�I �kۛAT@O�t������O�&�� ����ڪ[ۿO7n Z���p��KV����IG�R,
�̠��$t�:����z=3�&)i[�)�gy�o��*��@���<��p_X�i�>�"��b��A~2{�zen�A7	����"�P��>ivZZO�������S��z`4A���R(�4����)l�\�� %h�0(ԫ2�ˤ��bГ��8I4L��]��1$�/͜)�\���э �W�*�E
]����!P��Lw��65\��1`�a�>v	Pd)��K#P��&�7�D^�ߛ1j��bj�JP`ל͖�e��ٸwX�ԅ<���}B.�up��{J�ue8�=>�Y>3�ٰ��x̟#v�H!6�r�A��O��~7�o�޿����y>n�O��پg�}�k���Ӱ��C��g�CivX�0$p	̓b�`#�X1�n�Xd��,�x����>��o����� &��d^�X��2���?x������Y@�e��W�6�+�������'���M1�]ɷ�� )@�U8��hcgwO����J'P������4t��<"��d|���1��G<~�Z��d��ߞ!}h�(�1�n��v�~�1�������֩��qxL�2M
g��"d.za�<�+
�#%�cCZz]4︢z?&�Dp�=��e3U�0-��V<C.�Un]���#oW��W�v��4P���9�����j=0�05�rM@@'WP㳖Xsi���d���F����Q>�5���t^��G�l
?�y�&���FT%�U�ֹ�y��wdQa�6�П�4i�K�+��E*M����WM�jD��?���E�c\�Ŀ����� ��ʋ	� 9�X$. �4)ɮh�(z�=���]��*g��3��s<b�������B�,�Z��+-������J�� �`��>�|$�� 1�/6�1�?��H���8�an�XK$�l���ZH(& ��dP��H�Y�y���8�����ߋ���bz�I�w[�+ǅ#sg?O|����.�����>?W��3�=x��_��׫� �E?x��+P��t������W��7��M�`���w��e7�2�{�so��|�r�]w��~����/�'�ʧ=M ��Z����X�>V��^X���3�~�{����I{�.�{T� !��^��2�s��2�{�����s�Q�V�W���3pm�B:��5���D=@���������^��{�s+K��!4t���߿$�?v��/|��_���{ы^�u�3^�8lL?��}�M7�� {n���p��^xF<>u�*�	���Y
	�1 t��E�!}�ax�bS|�~|�&�x�S��s.�f]� \�^~�p^U�>`&��ϩ��wB�@�n��Ue�,����@�^��!e�?�=�E���u���3�"�^8r2�b�vM�.\�<$��^W@n#��5#���m�N��U��U�����^��|,���\sIڦJ��f��gI���w�����/�A�Vk��B��f��c���u�+��2��I)���]�ww"��L�7�1�VdPg�L�K��Db��d��(]�Y�/4YW<�<�z] �nⳌRkW0����>c�����FR� (u��R��~�G�)ƒ�. �"0�+n63��R���͙rSJ5��la��
̟'�wD�uF�s�g<`����{������S�D�5gHñ�����̽̑bc/�ٞ��`��2ߗ./����o����1�������bޏ�����_�jw�W�a4�����8iH���7������W��U��j����|~)�Q��|`�~�W��R@@�>��O�[o��=��Ԁ&P老�"�pQ �A#�ε<�^(�0�]w����O��}��P���n(@y�em]��{n|��.��$�r@��O ��?�q��^19�S���k^�E1	�� �|���:�ߞ��,��� ��c���^h�c=��XX�\ H�x��~)��ɟ�s��zL�[�6|d���q֝�c�5��⸱ɪ��g�{mh�8�������y��O�m�CR��)Y���(�QaP�Q���t����ވd���e<c;rՃ�*/�u�{6�Tӻ;����n�^�Q5��S�p��Iڨ�4ԥ%`dǬ��^�ߺ����2�B����"�U�Oj��s�p$h���1�<�M�U��j���,`�*�{�����
��dc�x�EX��b#����j7
V�W��E��fT�p�6L��c����虝C��5�t�VBe� |T�ř�*�)��Itb�H��	�N�?��l:)-.lY0�u�E��s%95xn4����J�ZB#,���3���4v���\(Oj�y/�.*c��4e�~�)��7�׌�F�e�@�v{X��c/��צa*K=����ĂZ֞��3�����c�]8�����W��q�Y�yt켹�5(Sug�I1Ҋ�����}�����F�$C�'3��-aE 97#Ii Ś�7���*dc任{�v��j���!w�ב���Z�'�y^x`���o�uF��L��D�z��d���B~u��>'\w����哟rǎ>����%5r���=��8u���=���O����<ǽ��nRYx
5j�y@-$���r��D���J���O�O�Y6���0d5*�w�ĞA����
��CGZE:�da4�|G��E�~��(�ѐ���{��df���sx&8���d����׎x^���#vo�_�1"�rY���Í����;٤n֮;����x�Ǿ�
�_RMF��M�B��ȝ�������V���Mp_�=���|H��>-;@5t�����R�%���&�����L�E6[u��P�7&�6��/�2	k0 �BI�#�ef�$��</Ọ;&��(m��Py~*��^�*�zNj�a"1��þے�ٓ��������U�z`�kʄ^��-J��Ҙ)!"u�ƪYb��puwww\��נ�4.���1O���V*^���uPr%q�H��$zid���Y�}p�Ѯ�&�b��a�D�m�6��x��-�^O?�������;�X�+Ֆ`��-0
:[X�M=�a��(�a�sX;m7e�h�욦Qb����o�ڿ7�l�l�ň��}���b϶�����Į���(w�Q��S��`񵾝�)��<֎��!.#8+
��C����5�7#��]s�5�Moz�{��@��}�r>��m ڊ� �\s��nymս��/մWۑ/�!��9��g����z���g�׽�u����R�D��	^���˿P��Qu�-���i�z   5�>����s��\�����@!$���s�w�����n���1�`żW���'� KY'���͒��<H�Ry��r�[��*��yիu��hM��_3n��N���c�6���~���aǼǥ�alٺb��KѨz�.��l/�T� +O4��V��U"��[�֔M�I��ɼ�!�F��^ץٔ���R��(�a��q[�;��A%i�U����[�
�y�{�� �K}�5���S$ �3&�.�Eη#�c���GGZ$rѵ�b���ļ��$�v[��yOB*� �e�-I0��tv�|�,x�G�d4B]�P��'�ڣ�KSB�B];��ۘ�ݶ�:,؍��,�]k��\r�;p�.�� r�.p���a�l�bs�-�\C��BS���p�dCvu�Ԍ{�3�n�6U�I�f�B
U��!�F���m��8��l�@�$�n�U�0��i�2�����$/�������$��1��2����q�dXTR����xR�8� ��?9l�4C�јa���Ğ3�qfQ`�q����ܸ����gI��c/����k�YIz&�)�W�о���8ջ*���ϵS�ϔ{s�˧\� �@屼X�,;�{}Q��g��N��4�;��}���pL�wSo$�k���}��_�� `�y�k_��ɗ\r�����z6���t{�׿��_��p?�s?���6���j��_�����g?���RN�p��c�{o|���*A��R��B<1N���o���$��[���@��q�7�q��ͺ�����q��?ߝw�;��t�z�(�x�;ߩ�
F�L��q�{�KՄ����~��'@�tp�>��T�&���˼��Z0�tw���u[��.����s��#%XQ�3��a=����q�a�O8��ƜE�:��C�5h�-����_�Þ&i�U� �PyD �m���E��t�E�#�GC���e�գ��J�����4���u���ve쑉:"����F���ߍ�՗�����;���!���e�����.��G���GO��ٕq�&`�_�L�R�Ld\q��������z4�ր���4[I��A=U�v��"M�E�N�N|��,x,/���d0��yO��ԩh��rWrv2�`7�=%xZd���]\;$�Ţ[>����-�uJ��`����N�8��9Ȩ�I4j4j�%A֋�v]�w]TV�ʲ ��Ŷk����Ξ�l"����6Ż /��5��4`����T�IO�M�'�0���� �v�,�I��̼ވ�ʪ���T��:��Vw!ukO�4u��#I��e�L���%�z-�R5������V�5��(�ƺR-�8]9(�� FY�$s�%��(�E����O��ĸ�dc��;�NS�'���`R"9��갑v���� �fk_��/�!di(4�j�~k��</󇍙�;c@�l����q�ξK�s��ʶ  �x4C�T�P���ɾ��XH�jEa�	`�����#����|����Şy:s#������:�O��TÍWUAeŇX1����ޮ[�kr�n�����ye�Օղ���>�9w��>m3�</��1���(S�)� ���?�s����O��+��^�8��.�7��=k������p��<��[l�c��u9 #������ag<o���|��l���ᗳ��r3�t�����<��ԛ�g�*1W�(]_2�����q��<��ն

���F����!� M@�F꺲����u�<����]%�V�\���Vd,5VW\uq���	��t�4�c��R�s5��V��e^�.��dw�m=�� �G܆�������]!��Z��Z��YU�l2� ��H����+k�
�Q@�vUӢR��F#wO��/�f��V&��5<SQ�ܲ술�d��ͺ�uto��� ��nT��"%����.[�g��֮;v�����Iw<�:��s<���l���ڍ���::q��N�{�,r�.����ڭ�K�I�y��-��ڤ5�(�U�{!;V!����RR�r��x����O�z�v	u��ך ����BV{uP���RkSeO�*Ppr\L�t��n���m�+����\�Y��R�;_#J�dgM����w����pN:Տ��"gz2Fn�vF����BB��lD�QཐA5̽��J��Zݗ�5;B#K�m�xb]����Y�H�V����eѶІ�؎��j�1✚�J�{l2��:F�43T�U�W9#�z{��ճ��V��5Z��&�B�)� w���#��L�'��P�|��q̃�_1%A<�(J>��lY,�*�zEf��]Pe]�~��֝�n~ˋ����f�FC��Ba�������r�1��>��׺�����P�B4�<+�L���ej��V����m!D���qDx�pe ��v�?�����%/�~���_v'��q�	{���ZS��xX�a�;�r�������GtW\�4wޅh*����>���5�(�z��׹�����N	��g����N��2���CF�\��yߗ��d=�Ё��1�a��
Ukfa�+�]L���0eHZbx2���V����3Uf(�MA6*�9�99�SL7d�Qf�9��r�4ܗ��Z�6l8�WU��'B��Z������C�ײ��|�5oe̵-��o
x���D�K7`��P֐dW��(��[̗���u�XN��u�j�K?��w�5W�Oe-��u�Zp}��^����'66��J��A!}��4�٢<�#�$ϸ�ʡ��i��uǘ��I(��-yn�NY�7��nT���GK� �
����c�+�f�aH*Dc������I|���e���Z-Se]v����C�4�Z5��j�͚k�4y�� �%!mm�S����֙��vw�wbo������g_���_pt��Z��y���L��v��C+�����>x龜��x�魭#����W��}n ���d!h��$ b����T�"�z
tlM�4��-T��i��`��0�οȦn�f#�������`��ܕZIt>��r0I!3��
�����.�����:"m]����׌>;ʅ�U=�6�:�Z�Ꝑ���P�	Wif�"/CJ*����6�A�Ҏ�N��kY\�9��W8�f!�L� G�	�c<f0������uH�0�a��*Uά�gj��l���,�PG�O���"n�8��4���ݚ��� #5�'U>C�$s����k��tQ�1�{���a��oַVE\�H��	^
��{�W�np�w��P &����3k��ݎ���+�b ��w�����A9�^�*�xX6
`ڴ?��^��=2v����_��_�o|�^w��i�5����Iu����{����GC4x�~��Z�;i����>����������t@�%���A��.-�=�����/pi)�\[�g�3d,���6�qds��q���-=:�71�+�$mc���S:�4�6��l���ř��k{^�m���6�y ��g�V�~4?y�m�>�R*��7���E|Ʈ[��m��ǖ�U�n����t�+.���x�ve-9��qwL@��NO�O:ɒ�#��S��xg����9&�Q�_�g�ß���E^غ���+W�[_X^_����L�����+ H�#i�pw�z� ���:B��H]r�l~rH�M6�Ў�O�}�,x��Z�٭�A�:��±���N��{B�V�Kkuɵp��ܑ�}rkOs�{��;�Q�����[�w��y����˞q��x��,����w���������s�M�}�U��?vc�`v�问�U�qf#čd�%��R�.��ZI����W���4�����$���<u
xh�K+�	M�l��JCEQ1Øk�:,,R-|��		I:k��|:-����ծ������:�2UԼ�<��%��`%�b�ͣ{�|,�YȔ���*⤀�yM����'���7�7v�&�v��b����g ���Bo)����yc̐X:zLn�33*,!�� ��� {��Z-1��v��)��z�&㙂���'�@h��3�h\�8S %����zk��L�OI)fg�ǆ����l���&�9K�~qok]��,���:8(��Pψ�!�s���.��b�.����C�iW_�@CU ?��gE��3���3^t��Ƣ�b �4h4��Z��x�d�@��}\¬e��o�Q�e���Q?������i�����'c��I'���R�/��2%�� 5�}�dcЪu�N^?c�E{�
r#<��[�i����	����=�n��u����#���Z�}/�ܬ��|8��b���%$���g�f��4�?5}���¢������+j�ٚ��U�B���C�]���ںk��j��r�����
ڠ4�,�{I2�)��������}����d^�<����,�'�Qsgs��>t�[�ۋ�{�k�=Z��yW]u��k�+<�l��'rYO�],lJ��xɪ�� Z·�-]0V���x���7�/O�#x\�|�8d�Sٽ���E������w�.��%+K���-w��	�ma��6�z����g?�������_�����������_��=�\w�����w�-�����M��{?�rzg_:�TN�1�A�&��
M�S� wk�gUƤRO1,��&��Z�H�߽W��.#����v�Չ8:a�(/D��xc���S�����ׅ.uKo8�MnG�U��Y���+���c��"���H�Y0�#~�h0�Ⱥ`'����t1�8��/z���	�����em�����bpfZ��G������s�*2.p'������>��"��}c�VBV�7ܠ�҈��M� �b������%z�� �w?��O��|��
��>!3^VU�a<	��C���F�5c�!��1�ĸR�͘ZE�y�g�!#��y8�!}o���W���Rŕ߁]�j�:~B���\�w�>���0f8,h���xO�3ǃ1EX���ȏ�����X�-�Yv��q��~P�	��A���x� ��xP���c�XY4�ҹ9�>G����@�9��]�ʹoC�} ��/ߦ�����O<P�o�3B���0֘#c^��c�w�\�*w,�f<&���<��	�g�<�{��[{��J�ѳ+���a�B���5�f��MI�ㆂ6L0#���!s(�h��Ī4;gr"kq�n�D��Ҏ�㻝����܃2���>�m�߮>�\]��K�����>��o���]���������O��>�>��Gkw|����C/W+��:r��/\^Zڷ���{7�&G�a��Մΰu������%�֛*46,�l���ﬠԓ�8g�˸�+2yz��C-�T�K&/��c��!��oY8t���W� w�#;o1�#
q�+��ng�����g��������������w҆$��L�}�{߭����~�ck�<���Z�Б��T���9��K!M^��P3��{c����s��Al����t����p��j����E7���,?Ա�)	�-
��^f3^�nǔ`��Y��K���~5�֫J�$���XU �JF鰙����C10��yؙRW���S���?x�8,��b�U@���<-Zu9Z�c�KL6�#.��O�!>�19���=#Gڂm�1��C��;�#��7�Y��e���� 	h���ރ��<fv}H�����1�b�����?- q4K�E\�@ZY-<,����>�8b�㌎����>�#64
b1�iZ�`��� �m�Z�g% ���l�Fe��%{h{��I�1�pLzt�:!D�?�ԛ� 8 ZGI�χ0�@YHUd7{���óŋv饗j�ϔ��iAyu�GX��?�s$���I��)@�`##4H��Z��EX�g�s5PKQK�}��K�'
,��OƋvr}��ܷ	P���������0�cE1ml�{=����"<^�|��޳��u�~����YX\�y�u���&$��&���9�Л��\#�W��N��Z�M�ʹlB��M�{�K�n��<@�)���p'(�0�g����n���.��7}�so���{��_�����,��r_�?���c�����}#���K_�����$�o�vջ��e�A諪w2�\&����r��Q߄9��j���'�q΂�S�(쒑��0J+0��x6ڮ%��u�<Wݷ�`���n�"��K]P�#G��Z���\w���-�%>d��n���:����}��q%}iҪ���bLڐ��ZԋPRLeho$ڲ��9�\��:!s�̋Z����1s�_�L��Ē2da9��d��ŉ��.��d�[S�k�=��8�~I2���q�!��ɮ��`�Y$`v���
�3��*�Aѹ�� v��{�k�\�o�Ѯ�B4�n�E����F�=�H��2��G�kC��0*�5xs� �]����`�� mg���7#kO����a�ɋ6�5�YZ�%#��D�Lܭ�L�"���7�Z�^�Oo���~��X�;�`��;�˾4$I2��7�dcψϦAbU��[p��A��P�Ū���m�6���0���<{G`���?x�����5d�p�$	Y9��� 	@,�o��x�~�~��R A�'�Y6(�Q�����dv >�vb��Ϳm�.ƵU�N����X|���n��uoT� �%F�t�q� ��DY7�a0��"ʖ����ya�` ͇ӹ���������<?^
�L���X4����*����fN��>�%ҧ�+�X\�mg����ɒ�A�X� ��l8+bC����d���e�<5�S��o�F�Gw{���+���y��_�һ���w�}A�w�����/}�˟�����{���^\;o�2�/-����~�&<cl�S����]��<C��$ՆY0�"�>Q��pX�$���� 8��Be�,��}�.]]sM~�-��<�<O��j�Գ|��G/��ʿ}ŏ��#7���\�ᆷ����w�r�����G��d��Z��&�D&��⇉w���S��,��D�j%��P��ͅz�P]d։��Y6���+�ӉS.�p<��f�Ĝ3���t��)�?� ��
0�����n�E�C � /�B�W�eqd��'����\]p�!�ր�b�ܹfX�;�nH9�xƵϒAw�u��tx�=��Ƌ�֛���ϊP�@Ó8	ma���0	x.i؝���#�N0�7�A��v�F��<xTh?�
�g��>�>�]c�0��"v��'l�h�f[��i�M7I�"t��糝6�c4/��RM�-�)��{N�Yy	Ό,k�7����Pzab7��U��l+~쐩6���(�����/��Ғ�mm5�,��s��d�۽�]UG�{�x��������N?������s�:|�c�r�(1Y|��
�XrW��$D�0����P�x�������R����Y[�JY���W.������O��
�徢�ɹǘ 0ܽ�/P��8�1n�+�>��%�l���a��jW�?���x,��S1��/��a�Y�����BN
T��ӹ����L�[O�'�Ϧ���̷��/��Pڨ�=�'��'z�' �h�N�'��~ֳ����^�U.����w������[���[?��#w;v����Ç��,Yo/�=��l�*�}
Z�����w�B�d*2��:<���9^���l2�qZ�i���"(M�^��&�p�n��]����)�����p��V��\X�}��������Z�m�[���;����g6�=s��{�y�+�|�f���L�AT�^Ơ���L����Ρ i���ʵ:�� 1f���]��C�0�נ�-L撬i����=�vccKk���g��/o�i],�xkF���TA�kw��~��^I��>p����_�E��A�:���'u�w����^���f˘��pӷ� 4�|�CV8z�a5fbυU��s`���߮;U��1P"�|��~��4��@��]��gÎ�g~�g�۟�q�׉2dl��������ޙ�T�6�y�~��!�p�I��� l��ø9&;g͇�l,�?m�Y�?<D����(��a��8KF�Y�G����
�^�Ş�y�4�w�����u�����?������,����7i&O�V<5�
���0y~����,�J%��?Fǿ��.���?�KS�h/?$r� �A����I[�&����Ƃ`X�\�~�G���0�,T������R�	Mq�7���^����iˌ�b�(�<1��|��=��u9+�%
]���Cy�C��zWP�0dL9�|�r�mt̐V��� X&����)�R�����P@B��z������+��~���S�A���QQ��9�^��7��?]ֈ�JS�q�e[W�o������W�q��k��f�K/JR�S�=��Bî؏Du�r]0�/�<��C�"I7��)��'��<�����0���z���-�ǲ3��%PS���ʎ�t��nE�s��0[ڿ��U�\��׽�{�W��q���>��W����<��q����q���2�j?U�O��Tv)ބQ�;䊪��� ��ca jc�ef�%����VOs��hT����O��(E�̵�!&���e
��eT)�iI ����0`Y�|�j���WB���(�ȵ�A3s[��@����'�s>��AL�4ǱKf���j�T���=/�8lla��w�]k|3�9��0� (�m�����rM�
4����9�cP�wBc�}�V�r	&�!����3D��5d�,����j�887�c���q/�ޓ�ml�s��+c�2@k�2�;0o��f�Y=fr�"��%<��>��1`�*�Ƀ�)0:���u�No�x4�]��e�9x7|�(�G������S0�y�?�`~H5
�q^��1N6@&�5��4$��Cx1y ��؇�������!�������##[�{�m�O���$�!�R2>�D�MA��@'�'��O�/������C��K<ӐMg�m�Y��9Qxv�4�o8�g����T�R	��*n^;�c:^�SQJ���K�T���v����]�{{;.[Z��g�=Z������h<Ұ}�]w=6�o%k���D�1U�( ft���ݕFs������������=�v������������͛9q��{O���%'_x��9~�7�U�eA��D#Ӷ�ŨM�������I��xy"K�,�n7�Ŧ �����J�g�3WB�@�0�J����  �h���N�__�����W���x�+Iޑ��/��k��J�����iQ�V�JQ�t���tiD����h���dvw�F�2UlU5UY�l!TC,�̣�]���ĕ�}�(嵘�(L]³qpm4�2}���em�T�IQ!=1l��I�4v�,�J2%���>���c��*��8��r��
�R�)���5/+��(�x��_�߇D�
ζ�����( D�OH	�a#�e���;h�;`�Iq8����*�Ԡ�r8,�m�f��0�>k�� ����E�x�"��q�(k�)T�=�� !$�ǉq�'��K%ِ6M��Q(�R~yp? ]��4N�}�3`ָ0o}��{�Zx ����{p��q�g8��aϒ�
h�r���U��g+�5�D�����a�l�ڌA����\ "���	� 6����)�� W�#�y�� ���m�2�̭2�i�׌ss�T�6�b����>�}%p
3����gc��w�"��S@4�wQ���c�~�@;�C��������ݩ��2G��3/�����st�Mec]#���j����(�Xs����9&S��x����?q��.�~���׷��e��ĉ{���c�;��2v�$㥠i2Vs�K�d���a���.�P��I|���e��R�k�a`V{�
lB2r��g2$D3������nS���ɭ�~�u����p��q݁g���z�ӧNt�7�kJ�#/_AK����/'i��:J��ߪ����Xt�\�]��.�4��U\�@�?(�Fҩ�T�9`�>|��?������qclad!4]�E\��TU�����?_�a��7��LȄ`�E2��B�][Yu����������G�."��+C?��
G�qg�������H�1_Ď�Un
��� <�����
^pߛA���J��q�젹o��Xʷy+L:�j�`08#,��0�o/{���@k+ 
��TU��a�%��4��<����;���iZ� }I����ތh��0詘��B4�ϘU����!Ə���u� +?���h�4�'3	8����z��ަ�Dv��O|��'~�'���x���?��?����#�O���o}�z�,��4m�7 @N��ȵ�7����1�2qn<(d'�72�H��93n���:dC�����[_]+���Yx��B�������3�I���a��|�D�	păd��4��b�13X(�~%[
dk������{{3k�<��n1͔`n@i�|n��ƞy��3�>�`}}E���~��6N�6%b���[��:���%�<x�	ѓ,�����U�E4��p��"���1h�U�������o<�ؿ���+��н_���p�G7�W:�Zk��d�'�bWl"u�&t�R�ۜ��lt��g�>�y/�,xѣ�f(عW�����D��])Š�⯌3��������������l����?2��(]��n M� 	�w���W'�#��'�G����$/	�zd��"[W�2>ԁ��D�	_M@��M���T�^>���M����b�E�E��#�2�w5�"���!��dp���Ґ�Li�Y��c�;��Fh��1,���.�)�d@�/��$����4���h�z&�ȗ)�6ZM�iÓ`��������01a�W
<+�%X��!���ei;`<|����{fԍ�b���}��F7�Ҥ����'u�}`�����A�i�`p>����DmŜ��+eG�1R�<� ����ä�@A���{����������U�h$���2���@xcL�bh�f�����[n���"C yFx��_���o
��ׁl�z.���
 �cƳE�_ǝ�����q�K���9��N�x~�E� �*��x�_v��:ghϟ��{܍7ޮ^����2ks ���r�C�75���h/���JCv�yOƁ�lc�2�L<ш��<<:|^=�Q��<������,���m~�u���#���:���<1��V��J���@6U��a��m��j���WK`�UB��/uA�q��/��Z�5�\[@xw0t�� �&I���C�\��ǜ{���O��i��<|���~teiu[֋�ւ/ ����I��N����g��'5p�8��K����k�{�Nz��
J���mHE�:Ʋ�H���5w�������}�#����&i�Z���?^�"(��8���+�������xc���P�F"s�Z��B���p�QMy �|�`�c16��q�K�e;rɰ(U�)� ލ���B	YI&΍Q%�����JjE]A��9����Ű��ᮘ\��(���G5{�x:k�+
^ 9��iF �=/�e�,�$�/��d����q�n�����3e��X�.6��o��c��v�*���gC��Eˆ��'���50:� >f�-�fz<�� ��p����G��럫�M�)We<p]��� |#n�}�YF�GvĤ��;se,u��랣�$pV,����y�n+d}�H�VjC�ѹ�r1�W^��1r�=y��zH���-˿!6�y�
�4<�E�z6�*�%f�PZ����<�!M�H���Ow�yg�Y��a<�\ъ��g볤:�����Ϟ�rQ膃�\]uŕ�B�����s��W�8�]�{��O�K.QO��##��x�w�^��`��@�i	�f�	0D_��la��0������?��>S�P9,U���]Tc_�>�<���<wB�F�Gsj�y�S��xZ���6W�M=�Q�5�v��:�$�8��_#��x�Á���'��˷m�\Z�d[ �zsAK���H��xF)�d6[0-���Oj�=�i�"�9�1�
����U~���ԐA��#�8��Y�E��s7r��ۅ{�;�����R�-������
7Nr-�u
��릃�X���ɞM4�j5�8Ԇ]�{��W�q��Z�m;� �tZ�$+�Z!IR�D}H���cKu�[YY�E�3���S�z�����B�L��P�-@����oO�4����X���7����f��*�&WƉ���-O���B�(��W^�z,V,�˵@�˳@���1�8���1��	`Ð���+ڃ��	>a< �w�{ ;��;x8f8�O�\�NBR���m�����u{��7/������8������r9`�,�� `��L�M��]��E>�]�)�n�Ҵ�E�EԌ.��Q�������;d� �g2�8��w��]���7���3b��%U���_��_����s0v8��^�:='c���u}K *��G�G΅W�~�tܚ�	���W~�W�b:$��@�>T36/�zJ��{x!�D���B�$ =�%�lP���3<� �����e$~�_�٘t(�07����c&�z���L��S�u��3� �G/�x�h��.�R�"��qش��MX�nai�%M��I�]�Q6@5U�U�_��EE��r4t�u��9&�:O�������q]��%/yIv�����o�d��I��ǬBe�Tۧ+�`V��(ey�JB1�<_}R{_�m��NQ>IRA���+�VЊ��9W03U��o�,��';�I}kwsI;����}��'$���B����h��#�<"̦�OyK\����)ƈBoQx�Ⲵ���L�튂3����4��2�����3D�hGU��8 ��4t���g�>�?�����C6��vd1a��# o�a�,�.7H������;<#*��]I�>��2:�� �1h�0�ϧ��|4)-�c�/Hh�\#���M�G�
Ƌ�)��k`�y�f3f��������RCgu}x�6^�?L� �E#C�%D�_�4
 ^h�ܟ��=
b��ٺ�'-y�2k�Dܿe�h��M9���0�?�r�3�2���끃՘��e�~6��3�8��_�Qzd��ˮ
Z_Z_����F*���@2���a�4�{&수������&|c�6�/�ǻ�GA�\�7�7ug�L����s��V�v���P�`0�T�X��[�mc��w�M�*2~h��<������?�c�d����b��}H�a޶��Ɯ��C��Fj5��Mڼ����>#�ڳ���5��:˫�=F~��ϘgPuOh��蘆ߊ���y<5�!�c}��#ߑuH��*�o����>L�����O��8�u�*�F�ZY=]]j���!�Y�������+*��m�0�j��1͔4������޲���I������:�i�"@�2%��y�Cd��ė�������@�}xm9��\���|�#_��[�g�da�m�:�*��E��FHA�<{Q����%��H�̵����Xy(9�3���.���u�%���h��Á�e(�j�f��:�cRMҙvg0��d�uT�WB:�ת@dW3z-&[���'�nms��D�v���q%��	/�Qr�ռ��<�j�\���`�y�>��(�0�1�My�˴c+�g�ֈȶ����w��8��t1��]���w����=}C��q,��}���k��tm��d���V�D�)����8��/ ����ڷ��!R�{�<�٪ӱ!��1���S����p�ѵ�a���1c�[G� c�e�J��M��D�h�Up�o��CCt�#��J�Sr�x8���\�:�l���g�kC�W�?a$<��,8D�'�ǋs�ɀPK���-ϝ1D���l�L�Z�g �6^,mXf����%ߥ��<����K��g\�t=/^�Ǹ���<`��x���L� ���Ɩ�C��A� #�����VeN�ṽ@µ��g��BPܧ��<��xv�q�k��D�`�H�0�s���.3c��̂�~��v��z�Y�e��b��B����1�����HR���D@̘�e]��=qJI���T+�"�M�C���S�G�ׯ-�z_M�<i7ꚝJ�S%T�gs��Y�+��#�v�Y]�]�'r�ʁ�Jy���ॱ���Ɠj���뱳ƈ��}�ERy�Xa0�������.-�cikc�����8��{>��Սc_��j7R@TQ��d&9����U��:Y��/b��ߙ�9'+|� �i 3��h~0�FZ��Af��<�7�\oԓW_	�d!5�HM����h{o�dN��R�J����r���f�g�\x�ť���ճ@C�������!ƅ����.����?��35?(�ٟ�Y�4(	Yv:,�V萅tyy�}���@_�%U�N�4iL�3�L�~���^'T�n����݌�h]h*7�y�l%�bXѲ��Mv�[bT�{z�k^�a���T�_�J��Zİ�ꕯTn�i���`X	�!����r� �q�<�@g8������=}1���C@'J_�t�ܗo�=/�08pPTG�  ^�䚴�vs߃r�#&1+W$��R�@�0�Ҕ���D`�ɸ9�0���B7���}�j��W��ՠ�b@���oEQ��i5�7�A��K�T���1F� ��\��wD?-������P��g���}/�>%��s��0�E7�PC= d�*�`��)BS�#�!��ɂ�+����%�?x9��U��$�"��,����7�����~��uǝ�j5�f¯x� ���k��������	�<s/�xZi��w��m�� ��[�Ӑ5E����\�>��s�$ܦ�@�Q�t��c�w{$��t���6|�������ܯUM�㑯�FJ��n�����-4��zM�=�hxhTK*���sK�n(�2��@:�+�K>��3��F3��x��Gj��������z��#./��*� ��%s^گ�R$d�T��5�Lˑ�N���$Y�@P��O��/�+����7M�M��.��� �I5y�����kŰ�I��7��ǎ>����][?����N<���Y8+���������W��+�V�%O����uiaOCH����%	d+���=̛P��D6���{�OFn7 0�����F�HKH�3ԉ{���v�Eh��,^�|ȁK���=�iP���e��cx����2(�[���#0��&�������p�"�f5K�ga�)K�5��XD�tF��b"rF*�`W�=�L�>	�"�
@!1x"�?K���-�������{����M0��i� V8��D�Ȳ���N8����s����[Ƶ����B=�;��x2�E������ޛ@�vVu��Zk�{������CB ��T�*a�x���H�
E
��v�|�'ч�W8�"�Q�;��X�N�(�����������w��Z5�����{.D^nv�=gｚo}��9��'�G����bpM�MXH_�9��ZV
6��f Ɣ��~�t�H��fzIq1C�f�"� �I��O~Z�������}�����`.���;��
p@d�c�]? �~VDu�ȳ�+��H�U�uZ��T�G��<��h���˸(̗�<��E��?��x�J6q9�4���b
s�"t���"��O�VTN1.�QH�8V!hj�V6��8q�~m(W�oy��ҽ<"0
jB��H�FePmݔ'q!;V���3/ߝ0'�q�����K�Y�tfκcb�MG˷\�G(R�Q����䫞��j-��:�|�������gv辍۝'Z<q��5�J�w4��Ƥ+����$�q�RW	�r��{ʯITs.�xy<n���(g�)R��<����冧��v��$lʧ�L><��,�sq3v;?���n��g�>��,���1���'�>����Y�ػ{O2XZu1�2��m�8ɃV�+Z�VC�%K�a	�
J8�j� >ƖӔ�Fû�fA��ʄ�����?�h� �rܕ�{���\�b��z:�t��TE��<�4��/�FpV���������<��fy{+]f.�g^D�-��)U°�.�~&�V-ec%�&`e��2_Ō����(�c|���]�3�c�Y�i��(�]�Q w*�e���q�4ܿ��ch�m�-ۇ�5��)�H�p����E޸�gT���,W����fi��I�@�8
,��9Ow�{�~��ACǢD;ؘ���� ��3�O����C�B�k��wM>O��+�F�*m�9�B_��t<I�о@��5�aNs���b��sa�r�x�h� b$kO��CD��Ώ�IH��J3�.-���]׈�����4
� alHS��jHuN��R��5-	cl�d{nyF�|�/� ΄ƈq`���d�,��y�Yں^|+���Q�$��,�d�&]��αFH�C��_(���]K��`��t�qqI٧�(rMg����-6d��r��^4J]���zӍ�dy<޽r�Ŀ���_����}r�o[������{���v�:�o��,�ne4p�AO�Њ�|������D�K�)X1Q���=���j�^$x��eyT��rʑ����(��ܮn ȹ-MM>3\�!V-�9~�{�r����xD����D�����������߿��Z쯮D�5�a�	�X^U#���\G.�Ud���u�|?W��A5V�9���6��P��bJ�������>J��f��Q��E"��[�0�8��wޭ��/�:����e�P?�5'Ҁ �&�bD
:!m9o�r��Hx��h0�� "ʼ3�=`�(������(y7�F�"����Z�?�A0� ��8�]�x�-k�%�9,RDB�������bF�f\���tœ�{6�f���#j@�ur���8r�f���J ��gs��Ӷ2���l(�^�@�{|^�&�0je���«_��|�����)��!Z �a��i%΃�Fd�9F$ �g��Qo��t�1^ �믿^��6$Y��fC�:�t���$]�7�o"qV�C��^���3��s'�/�={����b�F���������+]+����:R9����>����΍��r	4 �s'U8�z�\�|��n`��-��2ci)"��X�Y��l��ȯ�xLE��M �0V������Dxy6�s}��
<�8����
0��*�( DM�ʺ��<'�W��� �NB��ح��r�3���=w�����˙|[*����w�c7�����ʕsqV��K�2�}��^���Q���8�*5�6e�i�$�אxog-xqn���A�X-�(�$��A��Q�Md�F}R&2��.�d�k�݆L�����kW��ɣ������f�����_���۞�җ��#0����;�ѱ��nG�u�\�� ��uy@�/}�; �,Bd��'�Ntb�Q��!�@�%F��X<�j>������0�*�x���i�\^2�y��0�&�
��*!u�"�!����T���!r�,x}�����!�`!(nhm��	��6 ��>5���l�,�j�1.&aϿ1�,b��EM�e�r��� �Q⺏����3�C@g"H�������8�Y�0?IO`�4X��d�#�:�
�D�;��3�@pN�����7�G�Ԑ����5a� 9��t%T�eEa6+�f3�����!�Ӱ��\pn�@��	�oR\�6TH-��!J�,�$D;,2m&,RE�B{7ɳAH��t���Mor>�pѳ*&�1a��#N�"���r����v��k���fc>-D�N�d�����Ę~��I�)�xOOz�e:_HA�U�1P*���:�2�9읈���z8H�/~�5��U�G��4Z��"Z�<�D�Hi�I�@H�'��:�C���V��ׇ�v&�b�l�3�6Y��ɲy�)�j�6z}-#������h���Řo�7t�0�}Z�;*�^^��2�\�؊J�	̕��F�����봚N���˰�Tĩ!���N3�8���=q��?�.�|����җ��(j���^����w�=��r�^۱�Q�I�g;��!v�v79���ƾ�A�]�<b4��|�,��{og1x!\��2�e�W�^&�M��z��ƒ,
�m7ۨ�=s3�Dw�Ũd����gڮ?�t���ʞy��;�{��_x�O��cj Zt���~���S���?�A|�g,δZ;����׻�$�FԿ�:v Fx\q���w -�F2M��đ�f$�dC��%ՊM%�*��%�@��r��^全,Ɩ����{7��z��$'��Y�m���N<E��V��	�����Vm�m50�(�j�#�D{��|�(5ϵA����UT�Ȏ|�E��$�9G�d�c�-�o���� ?�N�t^  �ۀ��hY�c�q�1�E��f������.�(
�`o�=;���	a  ��IDAT�aBc�CH��*0
$K��X?���zeE�JH�I�V��:a���N�Kd����i�@���u@:��zoi9�\�͜�riƂ�iZ�ȃ�3�'����'V�P���Z��y�3@�Exx��Ei���C�l-T@�>`����7�w�y#�5r|����D18� ��~��yrD87����(����mB�cd��}���� ks���s��9���2�d��{Dix��0r���4���q� l�g����cّ:�1�Ƣ��~K~-ὁ����r����'Ni��8�������v�ܭ�#]x��w^E֏�o!`�F(��Y Z_u�O_�u�N�C��p�Z����qő�~�'?����|�;���?��ߒZ;<�C_���}���u�ѽ`v�|�ܝ��b�3���V�D�n_�ի�k�3�ի؉j]�>(VO����m�|���j�B:��D� �����r�
7#�_Zv�z��gd��Y�u��v�����]�s��z�s�Ա��Щ�{|�w��}���\x�ɗ����RIL8����^{�����/;�C�|����t�[�(���\���ا;�7������xf�x�^5PR�|?�4��9�I�К�3���7r϶5:���ig`o��.�o�(Y���z�i���D#����ϩ�a�����x���Mٔ��P a���bt��%��Aׂ�B�\�U�i��iUV���GTpL�$�#Y���#�&y!�B���J����~#c����%/y�~׌���l��b�h2W���v�t�P�����tI]���Aa���sd�UR>K�J��c���y�{ޣi��4<@�c"����ܮ%@���u�O��҉\pG�I�[ڍ�s�_���7#�,5�ߩ��P�w���{F��8|���U�~H�yD��~>�8�Ǌ�I�ۿ�[����ZR�87�њ�����V�?�'�`��Ør�w�=�p�T�����KD""M�xrmY�
}��N�w�X��|�#���u�^t��/��w���T� 9H��1���������_-���c�C� ������t��1����̖	��.D�,�Ĝ�rtR]6~ j�N�7�}c�oG�����!�c������rΧ>�;�jC)���ǓB�e\	N\�J�5���.�}�
$U:ϼ^���`��ݾkvZn��G�/0a��s��(G�Z<37��������;�tۻ~�Mo���q�=�X�8�����>��n���_��ꮞx�L#ju�^��1�vv�b;����䪣�5�,�3_UK�I�]4hL�=�)k�(�7�#Q���/��v�`���QJ�C��k'�XI]�}5ˍ�\&�8�jsV�W�Zf"�|��< ��(�G�������X=g���������>�����_<�o�=XM����HV�K����/|���9v��˧^t��¾������\S�X��;��c"�#墪k
eYЮ��@�����*����t�SϜ���"���`ц�W��)�`��>mY�����)p�*�#��E΢',�D5�7���P=<P�=�M<p�MDcH��{����WƔg�dR/�(̦���������cd�Ę j�w�[��[��9VJ������p�h�G��a����B�T�f��^z���Ac���OՐKDU 5`0��:O����pn�=�:���G��5���Q�e��,��>�g�w�y3b���ml��0�;�Up�e���`ـY�q:��A��i��/�" �"pd�KH׌�>�!/�xD΀JƙJ,���.����#>��Đ[Go�o'��6��ƿ�ClD�������B��@cJr�F���������}SK?N�bN2��� �Q�[��f-��|�˹m�FB�ueҙǏ+�`��LZ�D��CD��s<#��h���\iL������\%@��$�,3z�籯�售ͯ)��k���
��N�4�d�����H|_3mO2C*���Q��g>��{:���	$5O�2�w�,��������i�*�P�jT݆ؔ#�r��n�^�6����x���������3;���^�=/������z5����+��_����[��k}��Wl�z��[���q-ԫ���>�����]�H�̓zC�*ܭl��5�b���~~�R�c��3>n�j��~�x��qk��1Ӛq�]&�̭�8%�{��3�hV�ޅn9��j����[__v��,�A�j�%�9���~�����q��7Ӟyhvn�d-�����9��DY~��d�k���xF&�Y�S�E���{C-嫨��x�*��ܨ4�� (�^"�z
<�����KkNSPDKxP�rxd]��Q��Z~ؓ� ����yR6[<���=��Xߖ�M���!Ҳ��<GɃ,�|���Y���N|��cK����r��yӌx��c[yA�-��r�?�0W�+8�P\u���nr�3���,���B�O e՘�����HHUY��z��o����X�4d��!_�n)5��g?�pJ��엱 %e �tR��"b$����_,��ۘq.�ct_ F�u�b��k ڼ�90�7���Bi�G�w[��q���D6���1�0M
�@�2�5!5���f� �p`���5 !�c� �*{/c�(� 	���`��m�\M5�󇂱�gf�����'aUTZ=DI���C����P��7_್�p�V}ed{�/�к{�^מ����y�3�m_�'�w�yX���rF�VnO���  yv��):d��4�@ޣ�#���L�2�%P�V���&@k���������7�{+	����cG�Bm�1���N(����e>��y�x�$朎7�&���<Kk.��\簪*�D�5�*Ñ�7�FV���9���ӻ,�#������f�ө7�x����>|�<q�>v�w��o�����p�h���d\������>��?:���_~��G=�}�Nzf#�<y�|gn���fv��/8�upV��@րj>qIN�=��@"��zͭ!�������c��~���|�<��l7�C���=iB
B~6+ן�D��x��*�L�7W����!�ţNŃJ���t�d/�Vsa<N�������q-���d�ѨԫuA9	��Ѩ���2��Z7/@�� ^m��n�t�,Q�By4 �*�h��j�e��8+!5�u��G�1z0����n8��D��C,3�i���l�H��t^��.���ʥ�>�A^.��ϲH�>�ԁq.XX�m^B���1�Ѯɼ�2g�r6�p���ʔ�S���t�_ݧ?� ��Հ�4/���A�Ú��>�7S�5#oi�`�!5Cl^#�BY�6��� �+�P`�P��o���3 þ1XpPHX�ў�ު�Y��*����^�6iJ�����!����c�h!�IeB�(p\�V���5�������Z����5A fs�1R�gR��u��g"5D�%��9H�t���-�E����̘��2o�����[��m��l�:��|��g�yo�Y�R͸ �n��&T�(�Ih��번����t�_��k�"{���o�Y#��x$U���V�NDN��L����V^��Մ���g��߆a��MA���:�k$W~߽c�;FK�4sx�N8��n��Ty�Y�a�%N`�������g�	�p��⬎ƣ�!ؿg��$�����C���o[���l.�k�a�VMF��������n���p�/��g��]�L�V4�Γ���ݻ\����W�\�
����Z��"�ѵ"S�9W<K��~XaWZ����ՅEWX��M���C�*}'Nа�X��`}׼�J}�-�C&j3V����Smĕ'���,���ϫ�H��x8�#R4S��l��=Ѫ�̍iJ(���Kv�]]q��tcd�S�X��R�^)y�<p���?q�kB��Qx��~wE�;Ε7Sh:L���FP���)W��WC]bN���+J�!����1O���ɖJ�jH<4u�s��y�[/������y�x��'&Ѵ���jI�@=O�H��l���
)3-�8���j��P)1/� a�M?1,�,z��.�\�8�oi��w�1�'F�tߵ�1���aR�f�Øf	)���v�:F�ƨ���i�!���MX;ǵY��εL�.�h�A�E^�V���0Fde�"��U:��)7R;D�����:�3��"�DڌT��"}��w�b��W~�W܁�����<O��s% 58)����eߌ��^�2w��.�y/fuyE<�G�;����3F�17��2��=4��?��S$���Q]o\S�l��'��u/��ROD� 2DŴG���@I� ��x�F�P�����gQ7�CJL�3O��r���� *�3|���������d�^�o�I�v﷋�<V��v��3��LCCU+ŷ}L9k��׊󱼺\�VAH�=_��y�FxO�MsW�u�Z/�fuk����%7[�!�G�H�F�w �  r�%��;	�K�]3�hc4�w'�������`�YQg�rB�5+�j%�H�T�A�'�O��Ο�qW�?�]y�~�Ƒ���w��e.5�-�܏���?��ؽ�2�]<�y��.J�َ���<7�<�L`����ȃS2S�Ǯ���74B���=�Q�����:�I�V�53A����㡦�wh����R��X>+u���Z2�,<�O��8z}��Pd��#�R�\C�QN�
�)��YV��w��Ҫ�#�,`�B�Z����8T{X踦����;�����쳶�nQ���६�b�[��{�X���ٛ�ҚWm^�EUl��4}��80�H����DY�Z=�2��������
��ă[�C@n�u`��[�H磤ǐ2({�.�q�sE�x�R	^��ͨOK�ӂKa�������������dVǡ�dꁗ�B�.�e�R�v˂ue�2?��r�7&�>R�D	l<0�ƝJ�� r �1���m�Dǔ +F�*g��ɱJ7uQ\��L�FzF�u��$�` 8	��O��j�u)X��a�rΤ���R�R�\�q��+�We���L���扞PiF��h���d?��g���{�gy&H[�>���"Z�H�c?��"E��n�OSa��6·�f��TX���A �ߍ��BrnZ8�83&�hND^_P�[V��� ,���uK�Bԥ�3\��:s>�C:kި\1�#*�^�Mz2��uUDo�C��!�gq�͢n>��)��Dl�`cQ.7�h��f]ΰ��'����d�ù|Ԓ��i����rW8W ��Sν+�eM�P�ޓ�>S.�x�W��ءa>���P+U��I�ޮX�	����Ź�L�i%��5Yp`S�61�r�r?�`d8ؐ�7��CA��%K�������]��3q�*��)h}0@��>�]:��FM*)}���o9`q y0zK�˃���L�qU#.Dlh�XQu�T[xVF����i�0�3�6	�˃�����h��-��}{lA��i��ȪƋ�Z)P&�m�(��;=M�#0>�<��"�S�܍�jQ�"X�]3�Ƈ��b�"�oh���w���o6H#5M&�xN�<� �LtϮQ��-� y��/e/��>�uڢ�6̠�y�\%e ���ʣm�0<T�Hk%��H��#v~��SN��q2���~���j̀@Y��\Q���o������m����0��L�����0���"���/��B4��?�3�X�o�k��~��	p ���ɟ��x��(��`X�J9W�/����D]"0���9P֎
.���go���E�n�y��Ƚ��*�"4 �|�򖷨Q��s����#
g`�˴q�G1/n ���}L5�=D@v���ԅ�����7x=�(�[ ���  @ �q�����WxV\+�Ft��-EA�9���RO[A�m�Dس`sҪ��q�m��F}w��\UKk �bܳp4mӰ�*���I�MsYSƔ$O�pS�d�k�&�ׇ�ج���ٶ�%�r?]��jw�����[��]�QS�� vcq�j��5�ٜ�鸝3mw�¬�t�nw�ܢ�e���8�N<�6����u7[m���CBT^��:��z�J[1�!eX���3�Nc%q��ê{og1x	�Xe������:�	f���h+��� @$F_S+����A�hǜ�����LƤ��-������g>4�i�Џ"0*�õ����������'2�׫�ߣ�A�"t>4I84V�% ��R�=�<���L�m,�e�5����J z��I��TQVU��A�]O�X��p��{e�q3\���~����t��V�R����i;w�8hV��J ����a�|����4ed��x��P�t⁜��-%q��f(�Л��f�[�@��{�T�㕰ٸZ�i�|�h�;�z:6~�1��-*��u"on�#�?d����2���.G���]*WvoLO�H����(� Fo ����F���3o}�[5}cD��T��V)E��D������r���9`$���gT�X�aT#�'���b���{����������L�r��K��PJ��}z�&Xg�9��_]uo~��ڵ�bk�O /@��s7QB� �1{��߭�$u8�\���k_�Z��Xe�瘀;o*�H+� t7�pCQ9�c,�7�-�MSca_�1<RM���FV�3����vme �5�Ƕ�㥪���P
FDHk�.���;o�B��p@���
�YS�}w�����Eq�TOĽ�HϻQ��rU~����5��l���3snP����q���i>����Fbc��*2O��V(���U�6w��Z�w;��l�ݞ���ԵU�v�?��'�\U��Z�͉-B�#�}��y�y�t=m���(Nb�,�����g�}�f�Y}qy>ɝrv1X�\��������*f)�+���j�G�u{���k��j�0��.�I9�n
�h	"o���PO��b�.��>e����Šv�@�.��ɼ!C7k�Az�_���i`lR$�3��p_�f�P�Q'lI�5���)�9��#�j8v�ݏE^�)�U��Phs��t��x���v��L�jA�t�4j^�U4�� P�@\�PI�"7�fy�TQ�w�Pl�i�a���"�����g�*��hJ-�����Y����)QtJ�����S��t�u���@w&�7���VQ�<����q/;=7�*Q� �7���R�s)i ��R��Ke S��[�.�{`���EL[�g�}ή�^�m"2c4�B�o6?�?�������	ʴ����E�6��;�T0�>���|�/N
��QX tH�#�&�������4B������k6��/p3�9��9�W���̻��z����Kt,l���NA-���B�e��d.�}[K��/�H9=53�� � bL� bUiǎ׆��N�5[i��� H ��[^Z.^����0�5&���V S.B�\����d��&T�(�i��9�T�\��}��X1/>��;�{]g������c��_I��(�p"}�y�Qs��}�;������;-7�w�k��f�"�"��;;�N��v�ד��`�lT�,��ά��E7CĜc��V���GO�ѩUW��23u�sq�k�ڏp^����;+z&�FaY%HЅ�4)�mI�(�v#���v��������ܘ �acEjA�k���ĉ�qU��3���ˣ�K7�LV�h����4e��&^h$����6]�zI�lr���d�,���7�6�akWj��x������t�r�|��\�3�ľ�"��*�����i�u�Q�-�\WeM�%Ed]]TՈg����W��,x8a5�M=��6#�DY]����_����p��F����"	�.��j�J0��]�s �R ����i�QhkOȷb\�<lf�)V�{�RF��d4,�Yf-��
Q6�n�s-�Ě���#�Z��M#R!}��e�[I��<*!�eck�����������X�C��e�b����m����1�j�5��*'�"i떌�&���tFLD����X0���~臔4j߅�a�F��;�"��w0ؤu���0�7�G{
ՙ�g���pe0�D!(MV�R�k����ܢ3:��ʇ?�a7��rm�+��c�sLRc�\H߰q?��Ba�v �y�`E� �`DfR:D� J�������
%�Db �2G97t��^k�I$��q^6W\����e�OD}H;�=�m��Y܎��X��"�������6w�V�&@�ȓL����;~r�}���܊ V*���g*~�wf;�3�P���Q[���<��ȸ�(U���s7I�b�-�Y�?r��4�rjmō���*)��ٳS於/ߝ��ݾ�Y�@�R�gD�N���y 0��� d���ڑG�dy�G�)$�Q�2ߢKx�w���
1�<D�X����Bd5��5C>�ȿm#���^��(�TjQ1���IU�S1��0�ś�	6���TPp���f�:��mȄ�2J�d2�=�C���ɟ�Z&#h�芒�F�[u����}0����k�Ȥ$���Y@  ��)�XS0y�ۜk��[uPMlE�k�(�m�S�u���;c�8��9L�>�$���&�)g���5x�jRP��!��曌�
�V�x��̫ؔ��(����42)��I`0�+�EĀF��%��5��7]�u�|����*���vպ����!����iwfܤ�+��;x�rLb݌�U\�����(�2�5�0��9��±�ހ�ai��p�z],]��r�o���Z/ w�ia������[����L".G��ബ��fƨ0����>����*���O�S�y�;����W^��x% �����%?�b������  #�=$���Oox���AZb�P�z̟o�Q�����]��,@�ԚT=o�������G�?����?V�p���8����i��կV�9���7�?}�;���cc�=a���RD/���=�5M,��'?�)Um����D)��~M���3?�3
Ҭ�B��K����; ���?�"u|�o|���1�����k���Ƣ�?�ID����v ��!A>�\��U0}b����v����
 �ү'W��x.j8
(��<&�H���U_��x�x��[�+h��ّ�6}��;�,���}q w�dcI�.����p^\1	�T��D��\�l�fc�2��X,��>��5���k��	0��9Z�U�>0S���PUZ�]�dåT(�9��ٮ��,ܼ؞,�Qa���V7�P�݊s=�L�[���i�t���u�R��p�L����~�xog/x9 H�Ȝ$�#�O��(~���9�_��g�Jt����"P7��[(�Ʃ�L��|�ȹ5�<D��B�c^"��Tr/K_ɽA��̑�\�+���ȗ)�q���j +Q��9+��(N�.�e��}��G��p�dR�ƾ-��9Q�Ck�'5�w����Hm��l��<ao낣���Հ�8��g/�:L����H�f�[���d,=��
0 $��wň�r���-��.R�R���u�vӪ$����j�Ewm]e�=�F
��m ��S��UN[��#�ݚi0���x�ǎ)9�S��TQ���eFB�x�ʭ�s��k��-����^���=w����3gz��m1 Z��ߖz�}� {����Ƶ����0�4�{� �R�rK��> �h�h�O8&�@��� H�z�����+�����Fp��_MC�
Q�S����"���H�0OLL�QY
���t=yv�9 �tR�x���R��⸀���A%���/,�@����#cK��j"㼔ӗF�&�H�z-��y���|��/z7x1��x�y����iR���u^|���v����9��Q
�?�	�T��,7�O���`�\����;W���ޒ;�HK�bMS�D�U�^�� Pj�Q���k	�!Ғ��"�ZMb����!/��L�DU���F�jU�ɺ�"�������|uZ |��|Di�e�棁�z}7�%g2Hs��&ǫ��I:�I$:B�جl�ݢ���V"��.���a|��{��xX��|�	����e�6��'��i�k���4�r�K���k��ƅ �v�4G2yF�9.���T���P�5���D���}4��?���<t�%���T�a�}4E+^&P%!MCTD'[�$0�F`��B������d�3㠮�a��<4�Փƪ��@��B5��h7v]�2(3��-i���>�M��}��ք��i��rU
��m߂�G���軂�IR�a�z�������b���i�z�j�XM�$�B�U��Ȃ�4<���`<R���@lV%��p΄�1���k�[@i�����ƅcFĆ�F�[A�uǎ�,M�W���؃;+sgl����pؿ�߾C�S���9N���Z����5�q�P�ܱ��ڹK�]D�P:5�4H�DL�������2����������3�|��9����E��D���蠼�G~�]!�hbl\��'^�zO�DR�/��/~A���hi��nn��}���5�i:����-w��#��?�a��|ҷ0�|[�D�Ǥ=�����:#���pX����z�T��l���p�� \�9�1׈� Jx�����z9���yp6qCs��e�T��#�m.YJh�ʲ@ʧx�m��m,���S#��z��^�s��kȿUY���V-NR#�2�p�e���4�4U�>��#U��������,���3-A[�&��l�%�C���H�Qo<іiO��ʺ�;�ϪFE��\
���D���nA5 ��^5R{�ľ]�H�3��>�'�R	zV�ʴ�;� �`�wO��/�..�K�J�x���XJ�E6ն�r�Mh+Rp��O�F �E4�B�hLS&Q�F�i��K7O�3��(��Ȝ!���	�����E�s2iwK�ȾҊ7��z����|��|#�/�7�E���߇�Ws��+FX�� -���uٓ�d�[\�XF�J5��r$Ƥ�F^l3�]<o_�K�hX�)����9r-R,��܇��,�ƩI����ViԐŝ.�v�s�`p,�y�ϵ\�\�ce�S�M���9	 ��A�p@�`��Z9uJ�|:kc L�c%T9pl��¬wM3"i	h~��<��\.�[9�_���λ�3��X��H�	Q�q�PC$e��f"Vf@M���<"&����s� 3���O|�
���3������65Ҍ�`�*4�=Qӝ1�2��
 Ώ���\|����f���&#ks��,�6�#ງ�i+��p!k_@�FAN�+�����~��~N#S
��_���S�f��H�>I��o����>UZ�@�4�L��^QrMď�}��1�f�c���DKǜe�ӷ��#���4%}')�����ܜҴ5`J���h"N$�����]������zEY���A�E_�@{���y�ppzY��9�y��sM��.CAh4�/r�� 18ic��^��JL��:C�Rw�VC�� �^�&�Q��4���T6��<"�ARG�\�:O)
#�m�TD�[l�}�lg-x��&���I5W�M%���Q�	Q�����1q f�������pe��H��&�S'��Đ��� %0��L�D�/a�E�׽kX���5�FF2:��8�UP��� �:�ȫ����4"D��>N�'��F]�J�T�_;R�k?�!M74xl&�n-�?��F\����M��r:ѷl'!����bN������y��A�����b�bM�EE�	s]g� *WrX�iy���a�3ǎU����.���1���ɐ���e�H�s�8@���F �A$��K�+�����5�_�������B�㣹k��<:���s%,�����X��҄����ԓ�{�i9������n^@X������g�U�D�@�{���T[�~�s�N��1g<��"�& ��a���$�sg�8?-R�fi�c�^1�*RFky�IO�\Sy�Whh�SC��"�x��4m����ڻ��m�s���s x��{�rx�FY�}PB}B@@��*�a��3��x�a��ʁ[���X������,`�s��bs/p�0t���=_+*�L�N�l2�z]ޫ�vn}��Y�{�i��f��8k碇)�F�i���uR��H�2w5hm��}ԝqD@N@�zw�+�����ѵJ!� '1�T+���Mkc$6�j��p���E��jytx�����ި���5}o��,5�B��Q�J$�22�_|F��#cY����U�,�܋�*����E���θj�Vf���=����&7;&�1&5�^
�<#Q�4��I�TY8���p��I}j0��q>�K��\%����<�XAM�5�8F[�4T�w����r4��0� &�OI	h�)�m4��:5>m���ܧ��TZ�eB�L���#���KY0ǣt�(�A6y'���FNʯ�����qa�zdepT�[���q`0���
)�Fh�HZp�½�� �>4x��3ƣJ],u��b,l��7�8S�A��_rٓ
��m,�p%�z��1��"$o��^; �/׊Q ���F��0�J�	#h�\	��8^,BU&�NK�ݶ��oV
���ޙ"d���c�����v������m���|��	����TA11�����1�h����YQ�� �g\�g�U�;�(s��3~���<3^V�nD�cA� ��z��>g�D���1���D�GD�����b\�'s��NzӢw\/@���
@3R7/@�P�9�PbQ�z��n�M��<�9c�2y�p�;���˪��4Ud��-�hۭۥ��4�̠��+�<�[<7�M���ޑ��զ��&>��s^sv��M�㐎�s�On����t�mG��(8]�z�e��W5�`�_5��50i:��P�I�!r�k�8�QP@�@:��ܚ$��\{���z۠��+5߸T��|<ь�:�De8�4�j\8!B�[�4iD��yy�n*�D�|>0+�کHZ(A���01}"���ǣ�
�ڢV�~�8q�W�/��Hs�^�-Q:�O�e?�ė�"��SF�~&�\�F]b�2N����sCr����]��f]�*#y�F��f�@��2��������S����]���14Q�t�=�ࠕ�O�z�I��[�3+�p��+ ^�C?�.C�A�z�Ta3�ý_���h��ň�ʺ�"�k��ZZ-�y��	=6�JZIw�%����:�ϐ0�9/~���)ȕ�+�v����*���1�S�/ɽ�6�J���"�;�3���7z߹�/���KeM�Q�=ʌ���� [ ��&�`����Ɠ�n���p�=mPJwj���r����_�e�'�1r$�CpPi$Gd��c� ���H"e�_~����i=6���p�lW_u�;_@�i�X�#�'�Fz�;��>�яjE���O���y�_��&��v!�ii'q����=[UaN�;S�̾ O�=��+_�JM�Y�(��2^�|1(VB��k����)�1��J�\�8B���q \��/������>��� �⋦�</ �2���9�ͣ06�V�m?w��>o�OړjkZm9�n��h�b��+9�^�it�!��`e�}4ZpO�8)@f�� RY����	�$�؎_;00@p ��z�İ�V=��UX������7ҍ5(���!(��z"ބ]��'�X��[�͉�5�b{���qr�^_~�c�y�	K�����mg��)��#�`��s>���a��� T0�H	��A� �_�����n�7���� d؟���e�f	�$u�3�G�S=��*@�`��E�ķ�`�='f�x�)�W�qx���g�XI�h��(ӭιV>pن�"�"�jz���f�\Lm}o�*���TF��x��>=�7�ֽ�}�HG��C$�7ݤ�9}�K����bA����<m��k\�N���þ{���-���V'��ٵ�CuB0�֜������f�iM��E�eA�s����3WNOHe�4��U�$�������kIo�3},���"c[����M�B�N3N�s
�'�H��$������`�憀6"/|�u\ 8�(���"uG4�΋��4��� �Ҫ�0�T�#4�Ɓ����,2��n�M�y��u�
l�b�c�}"D-��@.�U��T ��ȋ)�D 8�a:p�Mm���yqaQ^;��D�|ܞ��ֻ��tJ�Z�o>ϸ2�\#�"�� B �D I�����Fi�BgV#b�W��X��8�����50̲M� ���;}��{��*�{�Z�N�"�l�4�)藹��q1�]���z	Tź���-�p����� '���8�}ѵ92�9."0rũM*����^=�=�1�,�|լ|~<��"u�ll~^4��cQnKb|c�[���W�'΄1E�*w��2.=�T�����ģ8�d�3!˳|;��K&w���_gU`�{)�M}N���p<qc�n�W�L 0�}Z���&v�����Z���>XT#%mE���g�7�+��}�2��BXQE�2����QE�g�2������)#=��ph 4l-��4�Z�c�x�UWI'%N�tA`�����.���l}u�TƟ'��ٸ(*]���ӆ��41I|O�A6.z
M�r��pUB�^��R�Ӈ�Ta�ස���>�y]\Yx���g��eA-�@��)�� �y��5�1YxM��4R c������.�l�C/}���;_#8_f��e�XgfMuԺ�F!-`�j�H�F���v>�1�3�&T�ƿ��Bl��i�I�v;������D�������pY&�E҈�p�P�%u����������	�@�}~�S�*�y1�ր0��x�{�s����w����[��:�c��c~�ο�����B�߯|��n��N���JSD�B�� ��z����� ,'��˷ݪz>�D_���Z?g�>�S~+�O=`ՈP��ÃlRCp�8>@��q1'Kh&V�,�]!�dϗq~\p,�d��fd����^����t��o��/���ԙ)?og*{�Fw7+3O�4�mU����5]O�tS7{�R��3S d�J�jݵM�]���/�\*�����ƭ����'��ʲ�I��! ����o�m��2�����1t�ʆ[�[( �ΛtR-����;Q�%����aժ�Q��C�/��7 ��XWj>���Ė6�v�7�'�*@��!?@J6�q'��M���q��-�>�{�wO�sO��/lY�z������Q��)浪�|<t�Q_������T���(@XNv�j.���PA���sm��!�0�U�%t:�G̼�A`P�_�����^|J��JK�j�y ���3�h�vR����Fݾ>�u4h�q�V��K��8�y)ێ_ɫџ�ao�'��[X�@����JQ-d�|����ҽ���Ս�kǂ��w�_zٓ
��2�B����'r���+��B?m67��u}]�9W����%�M����c��B�r�k�E��s=.+�����X���Ԅ��HeӮ��.�	���ǧ���o��[��S�崢�`kX�<P�>��w�v{兑F���(3+���-�j��ǵj�Ɖ�� ( F�8��M�n�yֳ�������*�f}ևPCڅ�L��g����>�W ���l��O��5��A ��'_�6J/�jD����J+��>����W�ʽ�u�S`I4�&����������Ā+��|�;�Y˳�(Y�U�\R��#*� �T=�F��+D]ʕO�k��1�0&5��0n��Q۽��_�����>M�� #��˻=�Zu4�F�sf+&Ϸ�e��'IR|SD�m��+��,�9�41��"6�� � �&]� �}�>=�hעrZ��P`���cq,'򅸖x��Y�t�q��I<t���F2�+����qLj>J��4s�I�I�M�4�x��'Q"+g�/�E8��=L-�N-r��FO<wR��\A��N�H98�s0�:d!�נܻ�Q.�b���;s�����n�k./��<���D�0ʄ�_	�ہ��*we�s��:��\#��I�ل��m�Hnu}�w]"�7�"�S1��K����j����Q�U����y��A���n\.%e�z��7�I��]\�L2"�I��l�&�?�L�-@M^"����¸x*�G4+� ��֯ܪDG��Jf�͛f_� XH�Q!<nƏ}X�cSC�b���.��+�N�����)�)M#�� E�AX,��(@��������ٽ۽�~�]z�Ů% �ģ���Z 0\�L�)��gB�)9��R�f�kO���c?/ĸ�[h<��cL�ў3H���) $�!����(E����v��l8�7Pc�b�=l�;w�'_�\[����];wh�� ��~ c��2t�
 �9�} d UuY��B*�~^ 4f � `C
�.z�!�8k+�.:�*��H,�<�f[��3H�}��H���b�p��8D���1�hH�����U��5O{�{�s_�)�ʬuߑ����;M��ļ��I�s�8@���jo5����A��MYE3β�"cl%�&Q�9s�D��b�5=��E�Ъ�ʠ��F�w��Tc98�L姁K��3a�g3Bk��{yP��j�E�����|CN�d��+>����o���e��)�	h�]3nh�J������X�/� ���E��O[��|o � -�պ:�Z�4ǎ2z�[�;���psXW;�1E�y�R�T�� �M˫��+�;Q��S2RU����)�+Wb��yBF]��b��u��6;��P���/ ���
0q�����nYP/�|���a{Ur�Ji���q%�u��t��`{y��bi<�U^�ܳ�ӌ��Te��%ͩ8O�UB1�0fy�i:�SQq��FT���HY磢��x�s#)W���q�4�K٣.<�-�.�q\��~�x�R������?��B�H�u�ޙWo��.��c�wyr��-��W����>EXH��F���N�/���l|�x踠�P���c�\��_��W
ȸF�t0T}몋w��+�ʣ��(�z�!���)��3@����?��j��F�VILd�s����l1.W��Wi��nnee�,��Y�T�����}�����Ɨ��r�d~���=c�[�A3����^= �'��^��ۘ�]ރ��9 ��>plʱ9�s����1�� k��߈V�~����tJ��~��;f��7�q  �4P,H��� �AZ�@�E�,��),{f�\��*R]D`��nȰ�3lNJ��(�#��1�cd�gӽ�����}Z�D��c�*�9�_�3�p�K�n�3�і���G���A|y>�#u[�me ����49S�6���#�h4�D:^֯-�X�4T i�̆b#�k�I A%8V��ۗ5\�i%�5M'i�R�'*��y�n��� ���&Zժ"���P[���|��Gz��6|Y���N��Omq��5�Bu��5t]"O7� -V�T;C�E�Z��&`R���D�7�k���R�׆l2��3�D.)�T�����]��Z�2Zڑ��xϺ�gIH���R�2�T�Yy-��[����]��r�H�e��ZmW��ޙs��;�7]��Ċv���
�ٵ�Z��������N# �L�h�7�4�D�G�y4���i�竊�2"-����"�o�aR�����w!��ڮ�� 6Tw�f'-e����a�󄹩��iZ�<����Q�e���]{�0���!�_�fff5��j�`�:��]���`����z4��_,䍠gA��~=��/L<�H�(aY�����i��k������k�N]L�l�x�xDX�,D�0�j��]9 ����ʱ�6��8e�)?���y�f�����Y[��o���vm�EvN�o�;v=zm�D��kH�P����[�"dq�)�c\L�v,^3cfcX%m��?��Zy�oV`b$]S6&�hd|�l��[� J�
0�S~�ou��:K��e��h.F��K�-�Bt���\�^_��3;���\���3��lMg�b|��Ї���>�o��o����q$�}gu�e��~�� �Q�q�kA���L�]�-��H��P�4Zc0� E@��?��?���e�+��8o�����p���eu�(m�0[G&A}{ӽw��x��֞lӜ.ϣ��R�hZ P���F�Ǟ;~�uPZ�L\��� �J5�3tJ�o7!�)�'��Vd]UBp� ���ح�z��t�c�O��6�VHs7j��7�{�Ԛ.F?�J
I�S&�'�x�:�d*�߈}��A5V�Z�2�~�9�}��N� ��Fn$�]5�B�TK�5�y�a����4��^����Oi;Uk�}�"�'+�>��A{s��_�e[�	�D��*��)�D�O��v����4;`f��v}�p�cwjC7�x���h�d�Ϲƌx����I#��O'ݐ�'�|�E�k��G�A�`U�k�����x/����W����i�Jo]� ��ԓ��Mv���>*s,�%�尫�U�)�zX�}���<���!F<~�|�8|��ͫ� ρ�������?���,�E�P�� �ch�X�����æ9��p����kcD���=����<1px�,vp0L�~��F=B�
Z.���׿��z\#pv��֊���r��y�ge�v�6#Kھ����3l�	�S�(�1��-2���M� .��qeH�`h�R4�}���!��p�O�?���g?�|"++k2o�
H�� �h7�{�� �*���ؘP6m	8�i�X4iye9���j-, Z�.ǧ����8e~`RDwn��N���i%Kq���q,"Ǿ�k�s����ދ���t,{��Q��s�1H��%"�V)*�%M1I��Iw���}�<O�0���#G�}ǿ�Q�F�V�*3�m7綂�������K�	t��f�i)p[Ƕ�m�,�S�^e<C7����"
|��<4\���m�JC�������-n�=h�e��ytֲ�S����R6M�|<pI*�)7q�;1`^�߼�8�xF��G��(�����ʪ[�躶�W=h"�u��d=�u@��}}����ז;=W/|�(�VZټ�'j��Y^�qʪ#�4�Mc��Ń�Ě�\�I-kr�'�DAJ�C9�v�p�TR�ƌ�n�������F���HG�`�؜N�㥕����Y�I%i$�f��FcYه���G�+9.�-�j��aB�����h3�,�,sR?I���6..���V�9ފ�h�߳l�Gb��##�ıieUWiH���o��b��Q��UI��G�wYt![�l�W�+n��֗w��߻ɽ�]�"���1U-/� �I�X%
�0��+��)�EI��o=��o�B�w~�v50G����,����ߧ�O·n�\� �v"�q����6�*[Y�=�
l9ed�b��F u��ag �����nme�Q��|*�(�{��^�v��\1�vK��U��� ��w�|��s����s����~I�z DU������p J��H�ā3b�G�3 ���g1�L��܃� ��C�4b6s��;������ހ �\��'�J,���}@��d���Z*;u>�/an�Ӥ�������Q�D��ޠ�{[(��z���I-�r��o)���3~V�d��ϛp#�"���Y�u��2v~�JB�����U�<�ΏӀ����{���i��4p��6�5��u��L�w���;z�@����&�������,�4Q����s�qN�ni��F��_�ym���K�(QT��7d��k�<ߝ:"*Oevε�˿]��ҚO���$a�8���|�=ׯ�sT���yT2��
�BT]�>)��P��8��W3�gGsMh��UO4�_~n�#�;:'���J?�CK;�Q-}?�3/:��N�*�/����'���]�Qq�xp�N�5�ge�͸9Q�^W>���u+CA���h��?9����A�+I�ÕJ}=�d���ڬ ۽�$��^�\�i5�%�Je�͛4����)�1��n8�|?��X���K�@!Φ$.���wN����U�k ����q)�RV%UP�N
��Py$G���9۶�C`;[$�ME�p'������t~��D��˞�$��k�Q�����.�H[���j����I��_���a �E�R�x0t-�ް�S�p��t�˄KqɅ�c�i�X�݆�2�9ΣH�à����haH1�IX�x�rd�,VWN��#BZD�c��K�Z��*q��Nn���/oe��"V�N�(z���}��W��a �6���r��}�����<�1�}"^�y�{��Z'f���?��J�%����YƗ�Cuqd��
Rw�F��Ϛ���S�~�{��G�/p>x������������>߽�5�v���չY���� #V�PP���ݣcC� ���Q��<���Q@���/�m^��w@�M7�$��Fq ��������"�� �Y����F�l���EpH��S�?Ƃ1���1�����tn�3���Czu�)ּ�"lqS��q�fpbY�3EL,m�f��,g�9�ґ�;}}��$�ɦu	���Rū���N�{�nC)���Ltv��v�s��Ɍ8M�7Z�Pi"kw�=\��wJ2%=C�eH�Fָz�᪲޴�\N5`�^uk�YYr����a� �t��-�g����Ѿ���y��Qs�n�?qҍW��`uE#�u�#�4!��5l2=�3��x!�yR'7M�)m"��*v���Z��F*FK��5Α�O]�Ԙn��֚��h�-�dX�Fϵ������k#�H���cG���hc��Om�ݽџ|hva���{����_�oU'��/���S����,�\���C�\���`3I�5�h�l�7���=.]���|id���X���	�6�&�.�Q�]���*��5��(0�E'SA,�����FRsi�e�P�����]5	��{���Р+���EM�}6[x��9&���j%����y;]��j�#��f��my��h�$.現�U��.w���s��@5 Yois���Z���U%.D6 ,,.�˨H���<�x��bt0��!X��]�t�����bL��7��-������iDUR6�6�x�D�Hm��o�+D��{����:1e��t�7ȿ�&p~�L�ff=gF�aR)�K�����r�gk��tn���V>Ay��5�j� ���;�g>�Y�,F�"$x�J~ yN���Ðy+!���q�ܿn��}U�QD�F��e�Nϥ��Zs/|��UdR�C<�/��8;w�];v��R����?z�5d�]x�����}���y
P�~�C�7~�7���=�^�����
������M27�9c.Pv���!7K���9�=����0U����k��:��}���.q_��+~��w�T��`N��.�s�ǹ ���P ��|�-�b-��}��n�������YA��ʫ\��T^�S�Q�}�$żP�*�C�9EU�-�4��U[ED<8L�E^t� ����DK'��{k͆?�A�S�$��r]�cn�-�8��}��w�^w]ɱ�*���1��w�KT$J�e-�]c��ݕ��[3��u&7�ڲ��3��ę���Fn�:��
�����9�ڽ���r�r�'O.��Ʃ�ȝ0�6O�?ٗ��J�'�N5��,,4��5sΎݭ�L�V�D�欛�&�Çܲ��EqZ�J)��C3����3%sroHkk�g�v,������e��`E��{og-x�ϮFT�Ԃ�2��h��A��?��P�tY��NK'],`Rcq��e=���\�.�����s���\v�ާ>���.v�$�#���?���㝟����_y�ȣ����;.�����lw�����[~>�e��J�fM+�������{3��IL�9��(���^B:t`M�)��(H4�R0�Y��I��ĠhY�񷢼�l���m;�\�3�
��r��t�3m`���喇Xl_��W�k��LO:Vf������A/%+��^�0�"+|	o0����$(�*9����F���P��tZ.9/ǀ�?���x�*�/��ɓQ@�C��/|�f8@JB��N0�'3׋��	�:�6�e�-���Lw� Cy�O����z+��[ٔ�M��L����7�[YZ�t���G���\��x��ts5��R�`>3�.xTD�0ހCƄ
���_�4�O��$N�F`j͖�K?qL�.M`�u����Keۑ��,zO�k�f����[7�ƃ7B(���6��%���Dk�����̹ �!�� E|�4�Y�+K2��ι��5�E��f3pΆEU)%���$D9���,�(X�p����V�5�n�,)�&b��-��R��0E����U����N�uOJR�����^)���Л�Q� ���\wmU��*k^-s�ȗ%#w�g�|�����|VL�kɚ��=�љ�F[ ]GSK�F��
�J�+�sʑLf��P��!��}8����ٱ��pR���Z�p��p�\g��l�vT;���dmy��[|����G.kD���ܳ���u�k� �ڠ�r�c�@5R��J�c߿��ׄs�%>O�V�ʤ
j���8��{y��������"��7��'�����OB|+T�4�kɳ��5+���ྠ�%1��17f��c'V����e�����_����߭����D�����^�{�;���/�M�W˄yZR�[}x����"r%�� K*�r�Z�y'��R�_gA�qL�4�L\{&����2�JuS.�0�>om���o7o[yQ�plꜵ�Wi�̎ㅪ�|��x9��0�v���m�޹K��.�<���������K�6au|3`���5��0�2�g���^��+u&����� �B��&��t�㒜�!���
�ɂFx�HdAe�ea5�3����F�����,2c����{�1�d���RH۽�/.l&*�6�f���M7�K.��}�\�+�6�d�Z)4E�ה�����Z<�i��4��{��)gK� /�R"H
����o��{䑇ܞ��T�`�!����zr� �E�{�ڝ�{�^��.�'ܗ��y=�@a:Dl��VP�&2���O��@aQ?�3: �o�QS��"}ddnxS�c�+hϼ�-o�q1��m�[5���x1O��DC��0/-���Fr~/�{B���4�Eqt^�8��8�Mw�q�;z���

hW�{S�%����;�q�-y�S*ƩQ�8Dg6w��ʡ�kEV� X
uJl�VH��+󫬙�u�/�ڳ�����u�s
�� �VS��r��gժ�ԫp��<t�a�~�QW��:�5iD4��& ���Þ[�o��)��% I�#���θ5B�-��y؝��1���W�ki=�u��k�����sΝ{����W<] ����{�u_�����8t���Gx�����3Gn��a>������_��ǎ���#��¸�zM���b�E�����rX%b� :��0�d��dԬN�W*����g�J}ю~6&��*^��6���c�5��ga8.�ѡ���՞�����,��򫮺�O��s�����?�S����w������?p�����yO�u�����cn��S����C:�5��mPs�Bo���osР�F��I��m҃���Z�)A�!�2y�/(�Ip�L}?���Be�Û�2e�]�@�XQ�n��έ|����Aa����wi:��j�����J�{��/�D�VR>������T
c��x�M�����������`8M-��Q��]=�> �B�l�zŧ�X$�LE:1��9�jXd�����ܬ{�^�����u�"��Γ�vC7p������z�J�M�m����#(��6�E�	�|�͈�FP�J*��QM���:��{��`�k�~?���d�؟i�,.��21��I T�y�(o�2����w8!��u�F���P��V�k9�\k�՛�
�cp���Z	>���d�M�'��3��{��}/I�}a1��  �Y��`�6�Q��Cc���3����=6��n6`��0�6����$Ui�R���s������FFfUa��J��I�2##^�x������wg������8pm��	5� ���:C���n��c?�w�;3��Y��?���3��}8?��\'��O��Oܭ@,��@>���N�[�6���o�k�9 A�{�>��9������s4/�x� �W���F�N&�&�,�|�
7Ș3�K����o��̃�Q�h;�q�O���)x���TXN5��^&�}���B�x��;�6ՋM����*x�o.��Ť���V_�IM>��o7[Z�f,Q�3��Ĕ+H�,	����>1/}(��ý~R�����ۓTK�n=��{ι��{�y�o�����"������+���Gn㹏���7|ǁ�?q`����SO�v޶K�Z�-���-as�[T��JӰ�c����t��EJ>�&���9/Oŭ;1������Ũ�B�'|ފ;J���dB��tՕ3.�<'����wnѵHg�b����:������.����O��¼�����?��6ݻsǛNX��ר&�h�f�e���V��D����ƥ-�z3��g!�Z�$���$�b#1NY��Q����r=jT��:�=?���yq� �D/-k{ҝ�x�1inԐ�rb�����: ��$��.i�v>�`,���v7�z���j����oԵ�0���-̀��Ly���w�o@���2�6oݒi^h�D�10�k�f��Ӗa��&�JɤxR���ϔ`��y�OR-y76�8Vm����t����1.��<d*q�(����B��6c`��sY)�w�������&��7;�y�ll�
O)��2LJc�f�:�n<PH�������4���s@Y5Nh��G*5 ��
h�~ah�0~9����g��8,NJ.�SN?M=`g�}��b��<�B7�'���;}O�x��bsY�Ǿ��֭[���u[�{l} 1��(����9,���� �dC ?6��s1��C�#��·���a6y� b�0簺\�9�#�MR�_ZвT+�Ii�Yg���;�^�wFp���i��2�{���T��'2 �T�A6^�[���l�����d�{�la��� �r��Z�,��-�=�w�֒�4�2�Vz]�6׺C2�N�-����j�s���T�^ ���&��FM^W��N\Hܢ|��\t{����NX��{xoR��/������}�w���>�.������7
4�⭿������;v�fuO8e�����0O1Ӗ,�z��Tu^��Ι���d��
^�^��8���(�9xy*n���A���2K�,!y�Z��BhD�j�+MN	��]2I>.�~Y�ɓ,���jf�K_���������K~�����,�?�����G��9s�	�a�<!Y���r]+Mw��/f^��n1������y�b�&��S�'&�b=�T�|H�e�40�CC���ܾG'�c�����"{Z�=&=ȉ�S�u�����!�:�r��	�V���M�����$�C��a�m�����(M�4��i���I0)��ʆ�{��u[���a
���H{b(8>+d8�A����E��+���^�w��X�k�OFS5�L�낁�O�0@>�����t������)�n�* ��wߣ4� /�+^��z�����?�q5��w��^� �뮽V��@�  Y9��w~WA��3}��\?�ˁ��$xP�]�n�)0���-�Z1��{��|��m��\#�����A'��E����_�tl,����b�)�k�c� B.�*����c�\���4�D�����Ա��!5�Ț�,����q86��9�\�[3��?mC���i'����N�þ�,��U+n��	���̧�UC�q��I�Jp�pP���s�ވ�v�|V���ld��l &��|vb�=y�<QON�U(呂	��2PQ��k]�f�[����ۻ�5�7K�6K+iQ�-v[nV�OS�Q�ދ���a]^�v���v<�,v�����c�ɩ��쵯��i����c�����g�?����ۮ����w�;�̉�O8)(3��/�rI�gH�TߧS�|�<���=�
^��)�ӏ��4ݎ[����Y��Kl=�$-FE��-E1v��q��4�l6<���%׎��k6=�i���\x�3����HL�$W<��g���?�����_���9G�5誢b1�h�WW/=��B>�d���$�s���o.�L]6�\5::9�9��G�|z�^����v�5�4긱��L�s9ϯH�-0Q�w���L$�e�[���K���N��Y�ɂ��0굎�4o�վ)�H�&��tƩ��f�W��3��T�2�L��x��ܩ2!N�Qu)a��Ih@:�=��]��ɑ(�r��Xݝ,�Z���>1�p p�Cd�{�j��&L/Dk��o�d�ݷM��ǁ���g!Y���B[xK�K�����[�/^
*2��& p�=�u����g�_SVfl<��ʛ����!��a �\��d<���)�k��D����_��9BPs�M��Q��=�^�:LQ�}�3A�Tu�������}:��^�	z0���f�������0R�X���K Bg�qX �]F�,2��LLNj������<���G��TLg�r�{2M��E^ ���;�{��鯳]`�<�޴es6	��)00��-J��sH���k��Nj��4
n,�ms� ��H�b|0���	fA1�֛K�������0FZs�̛ݒ�/6[nz��5��9�+&�j���"��n��It2o4f&\R��D�����p[�r/��[�S|dlj�/��՟�����]A�	,����#�.���w���v/.]0'���+qGk8+�J�\s���Jh�h1��,�li��[�s��T�����*5C	<
�F]M�k	xa2�OL��L8%1�2h�/͹y�"�^sq7^l�O]���o�z��OJZY\��w�;�����K�������k� �N�N>�t�D�������<�5�ȥ���<(�6��� S�x��?y�]����&���[����M :W%��gf1I��F>�ɒ��ȋxB4��$�>�KE��*���x<H��G `��YL(�(Y���Ʋp>.3&l���� ��v6cD�޼?ZH/�Z��pg�%�w5���M=�BVxo'�o���[-(�%+]�\a��c�%��?��� ��y�=3>\��uZ��@e�2��� �׼�5�Z�a��"����!T�Bi��8R�'^�?39���r��R�۶��@���Cj�'&��z���ȵ�MԄ��l9AI��෤�	1Af��"�i.�J�Gx'�!���i��o��>S8�X���������3��/��|�p*�Md`�4���)?���s{^h��E)��W��em�Hd��D�܀�az�\���S���#S� �C�FV�9�X\{���@}t�:��o����\���)��� ��̤�}vi��E��]�Rׅs#������B�9%d6^l��a9�<�IX������g<��v�G>�x�oT�}�������5���'>�{��}N^��"٨�]�W%1B��ӥɶ^H�yE�QäT*���������?l�-x�=��K�~R,�|�{�U���/
@�ٸ�uf�\ ���Y�$��%+���*G���ލ[7]y�/�<�2��|��ң�l����n��W��.���_��{��؇ P��u�"%�T����"��v�-K�cT�(==ƴT���H�{�5��V���4����`��.nXPo�{�C2�A��V���lr�0����e!<k��'��G������I��z,t't���ڒM萠�81}`�u��D�����QU�L}5�3N�w��Ej{z���o0T���Z�j�/#۽c����5['U�I2�F����"��k[���!�"W\3�
#���2MV�o�ەx���9��  �'�s���җ�Du��P��>=6�:�>�Oij�O1��/����/��K��z���߾\S�O;��~�<�m-��ֈA?�Qs��\��w�K�K��.��կ�v�d��o~�mݺY�]K�C  ��0�'U@&��N=U��0�dD}��_V� �{��/�T�u8^���+_�p  ������/����ߪ'���5�l�T&c����ѝ����D�u�ƍ��0�_}���M�Btw��#Γ������s����`}�ḻp"�B��c��<,�ɏ-mO
V��A��ƛmp
�]a�c������<�*>Jn9�p��@�ʘ^M�lA�:�n���c<��+V�>󮌵>�?�{��&�~x�����"�j���7�|��ϻ�E�>Y��w����w�������=qp���Ur��ȋe��;K2Gtq�K5u�9����]-���9���SskͮK
��[,�����ĥ��!`BZ�z�[�h����
����D�KWK�Wk宀��kW����K.i?�m���?�o��[����W'W&%���؅�ģf�����(:_a��_U�6LS�'a1�P�)D�yB^2�ҕ�)Z�	@�T��X�����~�Q%ލ�\2���~���%��'��U�7�g�2��8�1�O�(m��j�����ϭ�[>�*kW�M�>ֆ��QK 0r�r�0qYY{�A��Q=g6�$�:1��پy�x��C��G�ɱ@���O�u��{�����Ï*��$WM� ��s�a �+V����y��?���<�F�;��>�B�F.`bՒ1�x6�n��Uҷ]����:��>5]v�8�Yn��9�i�r���k��0,���e��B�0e��|2tLSE_��{1�� �i��
��.������j�����ǃD��ӄ��} ���E�k�7�x��mAB_�ٸ%�}������_�*�y�F�1�x�\sY��Sd��x����{5����I���c(N����[��G���
@��F��ԣ�6�m0 A�}�o�2(c�+*�YM�ZC��K�q����Nz�/�-h���Պ�KJ�����b�,\�v�]i��\�v��o�/����?��dm�>�9�m�����~�<6�b��t%I�V���po(�8ų֒b9��⽵������)��ΈU�J��y�p��צ��H&�E����ݒ	�Oh���\13��̆5�-K�&�[��*.�j�Ȅ]�blb���E�E ��y�V�$��x��8e��;��R˔�wIfXGc�V��a�
	!�C���Q?zߚ^����I9/A��H��E����=3i�Aw�q`,_����'�&�ߐ�>�sK�����0p�@$������4��u��w:ƙ�Ƀ
�a�A7����g�le ,�d��W��s�[��q�<Ii��_�M����Kxi�86�[ߘ���8�u�o�w!eZi���9Q­sY��n^`oBx�w~q!*3.M#LH�4^�J٧�s-Ⱥ��w #s�4�<�7��!����m��d��C�ZJ��Ӵh+���]���	}��{�,<��n��#�����zm,-6J��閗Z�̗��-'fYCdT�8H�&��_��������l�*��^�����V�p��^���\���9ɸV�f��� ���B��oy��s��×zn#���|�Ca�ѱ3:V��~$x	�x��5/ҡ�Y��������x���:]�nM��L�H'�������.{!�A��������jN��q��SB��V��'i�Q���{��L�q�)'�
�������pÝ������/��_�%�B��heN��6c�(��t��--K���+����<U7�"�I6y�I��'&]�Zs���.��Ā�Z2i45uwb��Ȝ2�q���[W7Z�m+UJ�Zc���
`�C=d[������U;5܁'#<��E�HCS�7����V��g��S�fS�8.i�)]�+���I9/�����a��p��h�Mpv�(��F�|mK�4/�@,-��[h*	�j6���_�����6�f.n�.GhN� �3���AV�(�'����h.���"���ަ����U��P�n�a�0�x+X,��g�A*�gA(�}�X5^���}&��wƭ�dد~���� ��>��!�8�A��7��{���MM�d� a��I-�^΍A�K������;��k�M���� �o�Z�Y�X-'�����;91�e��^�A������!�)F4��'�T��߱�����A��Hy��ަ�K������H����4��絯}��!���yQ�����Zb�i���Uף;QoDE	���򌇕�&&���'3?~�㣇�F��`��P]�Щ��O0���K�nAu�u
��5�9
�V��������@�N �Gv������ɕ���K.�ʹ���^��Ρݔ��U�� �r9	��������g�?�_��������Qt�%����c\�2BM���4�S�SWW~��Q����Y[�?=U�(�A�	e d����BF�#��`����WߤnF���>�?�6jK�M��.��0L��Zҗ����%�bAAK���=X����y�-��x@�J��B�Y�� �r�K��y�$9Rl�Ν*�J���(�҇a�kd�#/�T�|q?{�,�'�l�~e�&$Yʥz1��������Ϣ�{K2��`�2����V��8�}����.�>��R�0�ɇ�Lg#�f�l��Hw��~������$ޗQ���!/ f}a���x!��O���
�����cާ�.�LI�p/̻$O���q� �b��7V��>"���YJ�O��g��3��[os��N��%� L�&QZ��6�@+����/���Rq:U|ӛޤޣ<��X�zIu'e�f�e��P�E��C�Pfli@0�z򀧐�+2�8�����]�r�x�;�s��;)9=�;�6P�J4Rd�?�h�r���K���gݭ?�E���XX^�@6ǳcy��ӝA�8$6�K2�L�fZ�3:�6�q�o�S�/��:Y��t)�
�~z\�;x3�ՑL���ЉF͍�A��7�](׸q�[+ h��c�-�����6�(f:�IC짟
bo���Rc|���^��sO�656�����v;��7�j/Z��>������t��:O��/�n7 eDA�b��=5�Q���b��̓�O+qȿ�T*���-Zd��n[ԏ��~��e��d��A甇;��e���"�\L]V�˸4����<T�^�Diztʿ����5�c��J�z8�cբ�����ť�y�I�X�{:�8il��)Cq�p��mމQm���|��RT�;v�vl;�'���}r�]����@�����CĖ)���C��9�g����G������h������;���Y�G��Y�h���a��#�N(��c]K%�1�V���z#>����-�� ��So��j�r�ZN9e�ۼq����IZ5���Yu�#V��rg��P�$^!Ҵ5�&駩��zz�� �5xC�s}vݍT�E���J���θ��G^
@	/�eYV�:;i��,@.әQ�j�+��u����*g�Ρ�W��ɉIW�<�_|���=��CE��hce�����9TAY����s�x��V�woJ^sjtL�Ҏ3 6.p|��˅X�r���;6Ř'�"M9Q����������-r�`G�y�@��j2�V�5��)�=i�#�lu�N�좋��̯����i�ʮ�cP*�K�ʿ_ݠ�W��mGq`z�����|wz^i=ǡ��/�Td��
zg<��q^�(.����<1&'���>&^�]�Z0��f_V_=3mw��|>~��w.n��œJؕ-�]X�����b�:2�
=�d��p�D��U�ʈ��h+�
u����L�R��!ה��OXy#g���w8E�S��\�ÒQi���	(��ML�� �,1����ގaF6?�YF�M��r���}n����'�*P1����v,���˧lg��.D�b��D��Э��>�� -��Q��-Ԕ?g�4�� ��/^�;�%ƹ &�*��~%���BH�x���H�ᴺ7�ðS��ңW_�=�g�^�|�/�h"�®yG��`�{%��`t�d�z��nl��^tɋ�s�}�������ݏ�[�6l��^�/rk�mp=����7*�Y!�_Z�Uȹ. D�SO;MI����{�5�V��<������ ��M?�U�q`4�J�?����{|d4�/��x�
)���x�;A���+�>v�س�'gQ��Hvh�\�l�Ɩ)!�&<;��9�l�AIV�%@f���_�p��Q��Ђ�7�q� @��Qy���p����ʏa;^����F!}R_2L�7O�r`��44�h���^!P�6D
fʕ�,
����a��L -7^�����̍������pЋ�K���;Z�egzA������4=x�BЯT�QR+ի���.P;sb#������M-@��>��<' ~���~6!��g;n�Km���R���Jx�zon�%L&�Ε�����,�di��m���6�Ԙ[\~���>zB�����YO�v��W��w=����M��0H��㞦���� �PR-I�!�%>s�4�b�Ӑ1��J���Ӊn�PS�Ҍ��Z<p�2���DiX�Mɸ��~�j���عd��7$H�|=�m{>#�V�F�4��O'�K�۹��	\b�i�$im?��ϼ0�H��s��3�U2 `�a���נɷ}��u��~h����m��4f��\(��'�
��E�
i�V.��fh�gdY��-����Ѹ�+܅^�@f^V�;v<�`�,��.�/�j�����xm��좀�	�n��� ����}8+��sNw���R��,K�W�[�"u���R���z����<I! �~d���W/-.*0����u��9�l�]v�|Խ����td�� L(Vy�嗫��_���_�'��U�(+VN�M����q�)��U�2M�;��e��NǺ��\s�5�ȋ:��nW���_�7!s�7�8�!.�xn����-�vK��z}�[�r��ޥmn�����p�cat�-���F�!�yͰg���칷�*�^AUs��z�HC�)�M�R*|.we~�r\���T\*�k�֡�!G*O"�����Ւ��#]D��� �h��⸶�8�����=�
�ԅ�\c������ͥ���`B�WY��Ir���"�ݒ�S+������%T5�X��ʽ��l���v܂�Ņ@�J��SvA��jŪ���UKV�kW	@����q7+���b\l,+���f����Gz�glߓ$W�F`��hխ�|m��}'5ʕ)u����L����Ң��K]*���J�ۀJ������T�ͯ�Y�0� w ����D��BX,p�A��8u�B�3/�q+ڤ |a���T�ML�+�,�&(M6^�˧+"Q�ɤ�Y=����X)��e���Z9#�쾵/k.��qr1�P�G��A�n|&q �=.k��� ]��c�
���Z1U�RO��~Z�2�y .�l�3�0Ò/�i�n��>[f�Q�ON�#C(�P
��ԇGW��/�ʓi��-���1��9ֿ�x9����8� �3�C��B'�\�~}���J��Y�ct�΍熪� �5t����۸a���@�����CbP�n���.c�S�=1}ժUm6��zp�^�0���+�>�ig��.����]7Zv��§5���!�r�V�qke��.<���&|a�N�><��������=�n��Fw��7*��k2���Y%Ǚ��t7��~���[��DC���T�F?����#;t<*��ʕ38�3/�UT�B�
����}Z�	��b�Es�C�������po0����16��Uuʏ�6�^�J=\��b�2u�9� ���bO$���( �{���h��;]ȁꙋ}-2�}��g,��H��:.$�&-�Ȍ�,c���4�xN�c�׋\ F���iwH��p�fD�X��]�1�굪�t�]�Z,@nj�<2W��^��l���g=z��o�)��'q{���;���E�v�����b/ve��z$��A%�}A+~{e�ꘌ�FRqa��'��g���v���/��	��@�5[.hu]%�j�q��z��17)7ue�y��5.�TVb[��f����k���W^�i9���f}�����W?w���ܥ�Ri�-+�w�-���� ���Q��ȝ�[���"A���������y%2��/1���!.��ǟc%
{f~~��f�+*�����2q����2q��{���s�w���{����c4-����t�m�{.�hj����؊.���T�fĐ�g����<v�殷Ta��|�E��i(��`�Ǳ�N���A�ڱ,�h�vy}����ݧ�������h����ckɆ!|t�9i~$���]I�pcd��L���޽{���?���Iٹ�a5���� w�9N9�T�����W+�&\<$�?����s�Mٵ�1������k�ɧns�F��FI�M���e/S�qםw	��s�7��6՜� �2�,��ۥz*w�~�,~&��_�R�J��_��z�JŊ���[���� �q��S�$�=Dx�����G?�����n�4ӊa|���_��%��e5�V����?�4�d�Y q?L�:IA8�Z����W.���9!�;n�]�`�j�m޸�+��Y>a�pĸб��aK۲g7;���r4��qI	V�ԹG�O�C!�@�L��̄�Ek�� ��8�̓|�x<�z��Bbr8e���RQ�]�U�[x\��L_�a1HKs��{��/��O��%���I����߼����ӵpՌ<�����=�)1^��H��b��'���J�ж�~|&�q��ॼw&
E���tu�$W�h&�hwZr�ۮX!�Tq�Zn�1����ʉ��'�����X/V������׼���~�6}��/|�+�x����n�R=u\�HHĨY��Y��.�pP�$͜q��b�)�*��ĵ�B��lE���V4G��F�6������Iء�:l�e���7o�GW��a�z�bm����xOGI�Ї��n�@5 ����d �켣:,BD`@T�H��^$��î���T�$GF���������>��a灙�;ڷ�ώ�.����Wʣ�ɹ4�Y����纨�G�P �D��J��'m����4���;nw����ݷ���T-�{�����Fb��V�+0z�+~�m޴U�> ��}�������������^��ԓݯ��Wܳ��%\:=_pq���w.�������{�}�{Q���"1���w��>�9�|�;ݚ5�ܵ�^�>��) ��ki؄�Z�r�bo����C�q��u]�Ύj�HY1N�ϔ��|�8��> � %DsL@�eRU�^ä���Yɉ<7�2y�^+W}�{��k�u7\��&��tq�T����i&��+GY��Wan��g��U>���$��S��y1m3r�M@p�l#t^�\=���l[�xfj��_KE�_���sf
	^tP��RwL&�z�-`?���:ه�S7�V�>������[�v>�dp_���'x��/�G�_�b�^�&t�b���)V_�&ch�J{�n�X�'Mڒt��v����Sw+
a5LL_�t�>�=Ae��k��KE�g��R�m������b����ч��YV-{����o�����?K{��җ�?x�����k�Fѣf˫�"#_��)�i����bR��'�}:bAs�TҐ	ފ�O#.�����V����xr����·IF9+�i���z��Q�-��\����*�����M��ߙrk�+a�&[��l&�o)�y��M�y�vkS4�
ZE����4�� �	���f��h��4K$����y�j�_P�:�]���<��׶<�!�1�����,Lf�B�ct�c�;�	. Ƌӵ�L�gM�vgH۩I����ك�9�Xo��������%����y��Գ��~5���;xHE��<�,w�֓�JyG��|Up*��|�:��<�=p�Cٸ��d{��Wk��c YCdP���Z<��V�f%,��{G_���RS��U;������Z5f�k5/�GEiH��Q9�Bm���^]�?Wx~��h%� ���뙄���R</�! T+��ϓyX܀d��E�H>�hF\~̸l��=7'Y;�s�yIԓ��F�/��;��J���z��I9 ҇�$�aA^�-���a
IW�=���,2���@�욀�j��xa��2��R��p���v����^�݇j��OIk���v�-�����O�~��/s�ֺ�ɕa���(�RL��?�e+�E���ɜ��OI�[bZA��<U7��*�ߋ
�d�jF�̘L(�ͮ[���wՉ1|�
F�N��ÇMSMTLM�rj��l��~����]hn��w��?��?��O��h:���={����w�������ck��VǕy�eR(��Z�])TU���LX�A@i}��Y=i�%Ӗ5�����u_%���xݔ�d��D�+m��$�Y�c�m�b�v�^7����<�&�4Ί��n�|��"6�7�b������L�L���Dm)��J��R>Kˮ��[_�o�� �!��|�C>���b�c���ͼbQ:�{�� ��ӈ�>�{����N������Qp;J���6ƌo�[�a��A�nݪ��V�4H��ӆJ�k��pbY���2t >����=����"�t�W��N<YۂQ�@?��N-��H�Pt�Z����q(FlBñ����L�p���K�xuB�۹瞯 hI���+펿G �����o�׫�#��Vw�~O�����p^�/��xx6h�$C= c۶���  ��q�u�v�b�+_�J�p���Qx@4��7u� �b��$p^���p��$!(�s�'�܉[�j�) �r�����[=�i˪���0�+��6�|<#����ET��n��@~��a'nt��y9���y�\��R���Kx�J%��B�\��ā��+S���nn~Q��dH�b|=9f%�=4�����S�1���/tڤ^��ډ>x��Ʒ�����+>�;���G~�@������7���X=1^�����]&�ߗ6F2�:���ݲ���ˉ���� W�Ov�Sn;����<<]A����2Hܘ��F�$�L2Hk+�e �\�����n��$�^&�9��}�$X��v����/Z�?������b�%�\�c��?�+�����6>x��/���c[Hb�G햫������CA���L�Ӫ�տ����grd��}�K�`(i�n�V��
�ɑU[G5>FC�]f̎q]����n�̻���4�.�e$؄�_=��F�w��b�^3����V���9> �b��6���&R�=���b4��h����&P�!c�ù� #+k���[W�����2`a^�ibg�t7@��-�f�l�͵`�9����k4�k��p��gKv8����V�|�s�����W˴EtE���*���/}��d��ur/��� �h�iu�O~�S��}B%�	���|x8����;x�
�'�W����D�Zs�~�y�m�X�s+W�Ұ.�� �F��v�xĽ�=�q�6m�{����5��7<��dX^LV��)����o~��ꫯu'��U�Ư��k}�R��x��>��[�g�ş��|��o���/��߭m���/t�&� 20l����O��l���bW���EG���η��n��v|�^9���R�-���t�}�/m�6} J���\���18/�*[�ɮh1�=�E-a��`%Dw�ﳟH�n/�5�hfr�M
�e0���~>(6"�L���
�I�ѓ��ˋ�:3�j2�"�*K���^_����������=���W��W�^������O�}�}��^�����Ԓhl���(�=}�J9W�E�K�(�%]kF:N��-ż�E9e1�Y�ǵi�����
eE�0Aه�`��2��eP7�]]��v��ؙFõeP�]�wͨ��;�{0�b����N[�=�������wl�����߽�m�z�8#Y�����k\�Q�wb��}S���w�y��헅��y+'&N��T1��e�>�޻29C�����.@��-Ƒ���
o��!�JĽ�f�ެ�U��Ѣ_��eŜ'�z`��i�y/J~�,�z�C��$�$˄��=�
ͽΖW�5����yg3v�"1xZ�a%i�zZ����k����R+��3�y�#sļ5&Ff��Ӿ��� ��d��r7�����3��%�L/��D�@k�4���������00c�S��k�-��Ä61�GF�O�0�W���V�Ǹ�Ǻ���4�Be���< \������g��f
� X����
�/���!���ഔw21>��0��nϺ�f;#���������h�0�gh'�P��b�hK�Ĭi��+i�0`S+V����>����98{��6� @�OE��{���ׯ�{vB��\< ܗx@z�Z'�?BWpM��]x��m;��޽Ǒ���pH�i��p�Yg��@m�����]� �_�ʜӼ���	�ط?�(�K�۸e������u��Y�NI�)hn����[Cx�5�nԫb�Ϗ��@� ��J�-z�y����I#`ih'���	ê8�Nk�nW�V�x�{nb^�)��(���_��w!�������<Y��e��d,U����`S�%�	�2<��R�n������'����o\��o���?��?t�3_��e�]��*��q������y��������'+aa�����9�<5�?�����3Y.U��|ZȔ�X�%�Q��Tb�T
JOw�w����SQ(��2����y��M���鲬�x�QQ,�knfl�p191斖���U���<#U�N޽o�[�?��y���M�c8_��{A��LˉO�6�'D��I�8^_���~?�T�7��T���� ���� � �z��.Jq�� %R��ɺa��ôrt~�?Q�&-��rT�1b�F��ƃ�m���g���C]�yi�=�ܣ.n\�Ȗ���~E�4@�P�_���<�����s�Yp& p���������A&���K ��0cb�
6[ǀ��u@���������j���/�w�q|�-�I��r˸�\���tR�˲��&��߲%�ֲ������`����B��E/zQ�u͏�M�z�F7�/o��lV���v���w�>A���� ���+b�.�D�����{�L!�1Y6\+���ɷ��]��'�o+W�V����n��5r/OQ J��א���oe�i-���L�)@ 3>5������2� '�x�+4D��݌7��8' ò� -|��d;�3�8�1�= 4�9��|ul�q�o�j8�A?2���=O�;��  ��W�|��F��,�!k�O��z1�EMU?|ࠊ�����tN)�d������j�%�uˆ2ss�@m:�~�i��<&���m l� �i�D�9�ǂ�]�]y��r�p��R���W �)�u��֢̻�̓en��Q�t����M�bcZ�*��\s��ɋR�J��韸���K�˓2^�����N[}�@��{݈���k��������y��������X=^�lo�S�>��f�e��K���� ��* 7Ѕ�¶�g�ji��'�~�ŘdsY�Fǵm�I�����X+%h| ��v}1�<�	�)���u\/��ܼ���+e�#|t�E��%����{���+��S����-5�dX���~$�� ���2.Ⱦ<N�X-  ���g]C������
��Ґ�X� R�e���ݧUM5���0L�+�(�%^��d��*���G��B5fh,~�����jaa��2L�s���Ǳ�ɟo|l2�`(�ë́N��UW]�n��&�V�2�ḼTˀ�yH̍L�M�U3������u�.M�P>m�����0N��p���?�����5�I;���7����3\���0����ap9�bcUY�J�1N>�l�X��~ \����X�o�R�SOe�y��V
m���1�ȡp�yvv^��1 ���?_������?,��_%�v40cF�ƏmJ6F�E���b��������⋴c��H�1�'lޢ�ܼ\�c'���7��u������.�w����ʯ)����v��s�������[��V�CЎ���ۏ\���N����s�2 c��S+����!��
���\�s�{�o4^�ϟ����X�\�7>;�s~�3��1�1w�#�7��m l��?�c�3.)l��v�J,X]$�`��/��=��B�Z׭���j�*��8��@@얛nv7K��E�ʽI��;b��l�ydta�e�
G��#��""_߈y�x_��o�0[�#5��b%��3��Ǹ� ��1���� ])O���=U�ȜIձE~�6�]���.Z몟��x��}bG��a������"���N������2�����j�ШUV�|���}��	������n�V�~��޶Պu���[Z�~������{��!���b�uz�Zܴr�V;uݚ�Y'lq'�����E������QwE�m��a�TFD=K\ϼJ2�9�h�M������p;��K��'j<rC#-�z��P�Q�dɗ�o-,�@ne�ᦕ�P�A:��T�G����xPj��6S)��dR�$�	!��,�aT��bG�yyJ��6!W 7_�u5�Ԉ��!"��x��D�:mJ&s)��NoT�{��I�@Z��o�.��ǈ������M��OB�y#d�-�\,FO� ���w6nm��L�֢M�Ÿ"^Q���3���a40F�zyXxMXQڄj^����|��P# ����mUa�@�s?���8�)�bP0��}���g�~�<�� \��&[<Bp0(�,�!׭i�r|&�7��I�Q�c����ԧ>����/��+ǥ�B�< ΃C9���'B���#��p��M�q`�P�T��-|7%��,�&�����S>^ ȱ�=�"��s����O	 �{�'�ɳ�u����P��~%\��� �ʲu8�Gw����K��K7�s�7lX���9��pz8 ��|!H����%ZXh�X�L��4S�8�YUm+pɱ�lI��b��sawt\��;C��_ +o�w%���6�3>6�&�<���(���\�?_�5w����5�5�
ijf�U>�I8+�eˇoF	�A0(fz4/^�$0��s�.�tN�e9����k����a2(���v�}B�#��h��U�n
P,�s�9?���}��W��a��CYaٍK_TuYp�Z]�/�=ץ���Ű-c�ĥ��R�y�c?p����~u�P�{r���ˮ��4iE�V����i4&��rq�x=8c���'��N0]k-��C�ݡ]���ؐ����s��_�O�S�Q?2�NP
��
U�4ߎk�"��}�q�]V����&6��b-�HY�$�Rqɡ3֨*	�X�KRp�b
QW��J�;H�� ��)�fYF5�Y#Sj�{)ȻZ�,�ƣ�_Y����^QIg���ՠ!%OKũvd>��bqil7Y��;�l�)�E9�!`�8ێB:VPh�����Xxj���܁t�1��k�?��?�����7�9sͳ�S5o��o���(�;��P@���%�\���M�`�A��jf��z��t߻�;r+ۺ*���6 ц��������&�*�\݌%��_�����O��pF`���ƪ��5 *��`�6s�\��������`��i���P`$	��ż?x�0�xe~�7~C��g՜	� �'�O_���@>lgc�h[��ze�@yf�
%�"ϯ�.b|[���w
�d� 4��g��F=H�b!(���]����'5'�B'h��\�ʕ�;��s�B��H?�s�����g��2=5�+Skm�&+䞻��j��V��Ҽ��L��d���4�Ę�k��^�K$t�O�g��S���;@�Й)>G1޹�7�|���'x<���)��b�̫�jf^�gm< ��Ȣ9Ή�	c��L�K����l�G�6"�ϱ�\3}��<p|�iq?���Qoh�W�����"gs�� d�M�ϓ}Gy,:�%~Ag��|����L#F��k��|@��vy�&��zE)��%�i�r1��;(�z� �y/f���rx/�\?�Riu�D�����e<�Zt���,~�����Z�7
��no�/�'��P�g�.�nA@d!�,�Β��w���xƖM���\]�{n��9xصι:�R��*`:Էa�@��DQ#�w���Tَ[��=|8Dۗ�/ҁ��+�0��/	H����v�-���rũqטh����jUA�Ų�<�����Ey�Z�Vf}P ���+�d�(�Z!J9�4#2iP�-�H��5l�v ��S�Q���Ta�u`��$����B����OR#也��0��pZ�(9�6�ܐ;�w�������W/�L����uo�+C�
�ɩ�ac�dǸ`T��	��{<	oy�[0�c迼�n1]���)7�<pA L���)'��a�Gv>����ئ���1 @������HI���Yg�����p{ n_�����S���q À�Ƅ~Q���d�_�����B_�ɂ��ɪ�Z��s|��֢������,,�3v��bFC���M7��OS�����;�S�s�#Nozӛ4M�&��j����usMٸK�:Zx�Џ� GY�m'�� �w~�?e��1����E%9R]�.��ey����W�ݞ��2.aIư�0�����*xa�\������X]����0������oh ���k�+�x�: q�Ws�WN�`�Y~�b�SO�����א����ڥ/}�f�X�ҵ;^��g����l"�����q���&��\��Rj /�L���7�m�� Z�d8#)?���;�T�#ƙ�#3ʣ��e�%�����H�UEV��~ۍWKnf�J��][��s>�8���t�"��+�)���bOmܨ:!�$-I�K	�I��NN�G�!��|�~�!i�a���	#�ɏ+㵒����x�y�<�gV�Ʀ�)�׹Mbg�� ?��#�.�=D�
����R��-^�Ac���Ћ�`�'�f�Sm;n�Kkݺ�xOA#��E(���)zNsC.Jd &*VEl��Rˑ��zcL��������<��Q�i(�_��D{"���A�6tS�k{]�wY��r�����t)cW�}
^5�!&&� 6�gbC��t\H|�T������M,j����M �7lل�d`\]�ǘ���+��xH�0IeEw���������MX���	<+a�N� 򒗼Dɉ&v���IVy�~�I:��$̄�!%�¹{�zӒ�- x0,F����Ť���"&{�:!O	V٬�� �~i�Y$\�tsdJ�2�/�e�Q৤�4Vx�0����qd8����}��a�1��Lf(�$Z��Q�S�+e;/��<��ؠMxh+����\��@��糰F�����>��ә/V�Ʉ_V�� ���}b��2~���c��
��њ���\����vz:8�(�!�]�5R������@X��e��=Y@����o����������?�B�i�[�j�z��{��	��<�7�I��@�I����`&��--�T[-^9��ȓ�	�]s�պ__�Z��S �˦ ��l��-�Ƈ���3�Y��q�E��G�ޕ�EP>|遵�a�#�s���(�ϼ2̍�[�ݑ�f���>��n˅��nj݌ ��-�v峦��.y%EB_��gy$�aQ�r���$Xt�)_�����5W���G�S��S�������q�, �)�6����i�E�m�@�U��	�~j�m�MibI(������0̺�ZU��q��UJ��0��0]�2���³�y���i�~��;�c�i����MYƑ" �QQ_F�"i?1�*��Pm�	�����r��/�]���
��

W/G���ad@�Q7�ܨd�Ġu)�0�1��P� lu\�xv(P��j��i�UU�R��<�%QIg)�Z�1������҉
߱�Q�l_�#J���g�����b��l^�n�Y4�}�>��b�_)y��@wo	���W��f�;��i^���G�>����x�_�����e@��3�%�#�q�H����j�|�{��*&����x�H�֔r��	�ª�0ƙ�䬽���/�Ƚ������]³bZ!fHi}��4��m�MC� �%�|�.������k˃�<��e��N�?��7�2󚨧I�1�A�n��/ƈ�L���G�#����B؉1����w<泳��[����iXZ^P#x���O!�ifn����B?��w ^�˸��5By��x�g������E�~q�8�/޸S�$�c������{g� a���s*Z���}D�����@�!p����F~�ڰz���Cl��P槉�Iw�3��V�]�a'��9_�Pd5�|�h��я�D�8/�]���$���7�����ێ�c�� ��h#]dƂS'Wθ~���îw!J�V��D�ow6ϙ8^�rJ"�|	d�9��NB�HP�Q0+�$�E�ZY���e�@�'fM"���Zn���BQ]l@	%d9�Jy6WNLjv,���	ם�ws2�,8�:�wM�������U��UQ* �!P� �CZL3T��_���<%��={�~��W�q�J��y�Gq��S�HI��7*��ц�۔O�m��츨#�I0*�y��ĕ'W�(�O��@��Mמ�Wbo����cڮ�a�
b't1�F�a -CKc\�4�z�Q�#�i0(�A`3�=�`.�GLF��˷�]�����s�Ցm&�f���T��\�I����h��613����Ӳ�8^&\��!�ہ���w��k��R.#�Қ�-��*T�b�y{�h n����o2�I
*����aη��Ѐ�	#����)ӟa3В���B�}���z���N2�U�VY���I�W^��j����sS���V�Gs�n?�pT�g��p��I�2�0�vnSf�YX��~�^�O�df�+ �R�����{�fa��|������3��{x�{�I���_��_i��Wa�i�TS����׿�G��׽�Wݡ��z�����}��?��. D��T���}�?��)�Ae���������z=W^�5��+���������h���>�V����V�q/|�%��m�j����_븢����k�n�c�W����vQڀ�e_�d�!E�\����ڕ�ٵ�	w��k�b�k֮���3� D�|�;L�!I*��dهGf���qe���̻�LH�%hz}�@I�y���҂��;�&��oe�]��g�6>�f���'�;�/5e���bs��"��0��g���$��j1�4cS�;��ڑ�vJ�|F��t�ظ��>J��9��B�)��0h��Q�/ɳ��n���[B/i~�U�~�I�'TZ/W+�0O
-���+E*{0��9��M��3������-
����Ձ� 58��AJ'�AyuW<"�5-C�]h7��bGK�C�£xi-,�2eә�仞 7��JM1�������MkR����3�x-:_����!/������"P`�f���U&�0J�H?R��Q��5l���������V���G>I*�&�G�h0�c�mk:)����e!EW��J��ti3^V�!�E�,��~s���8��J�RWIǠ0�c0Lj�s��+�|�rՌw1�p$T9VVp�V��ۿGy#k�yPA����
_h0���saX0���y�l5i��������o�Nȡ#�Ee)�0�.�2�	��7��`�8+V�}�<6,m� k^�utU|4�b�f�~MLO�� �`�1�l�Dl��=`����|�=b� �f$i�O}[ F�7�  �3��1ޱ�!��YCx���0�P�����rǨ�tH9Dz���^T>	m���p^��nݺ5z~���w%x?�����K�0<g�!�x`�]x�E�ިj�B�l�+�(�D_q�~��:��+�7/���3�j?�y�qB����m趝|����.�X�X��t��{��/�6lޤ� ��q�F���D�0-�x�yb��r�7w��<�Ƌz��Y׼���4(��]ה�����O�y��$?^����;m�inz�
-	A�+<4���r}�q-��A�1A���f��4.����̻�Bɵ��i/�^+�9#�C<��֋S� �fLlATBA]�(BP2͓v]��}B�������.Zh+/v��՚z��n���d���J�I��	�v��6��~�|o�-xA���{S�xe=�?�AQ��n��;�����]����"\�k�5W��CDn�~/�T;�=5�T���*n�N�J]�]d����>�r�bT�`¥�^�b�5�Rڕ���X���V����ɸ(LFV?LBe��� �ste�^Z������H�y��Q������BВ�>L��<Ԛq;]���R��ރ{�[E�.�I��(-Ԇ�UnE��k⿢<�x�4[�O��fpܢ�>���}�osc�2E�|�L��bb�!x����YR�u_I������\ ��SFsi�5�>3M6
t*y2������.��z:��S�+~��b9?�������P�=.wB
�>�\�t \���'0��< ��hݷo���7�o|�zm>�yn���˩B0���s1tg�q�{������q?�]_q�g,��s7�t�ۻg�۰~��hK�j� -֖�����qb�:���r] .8-��8�e"�j�J�x]���Q��J���|v�O��D�LQ�F �A���n��6F�^�] ����L5V|� t�{Q��)���-�5����?��}�}T�p�m�����iX+@��������O�Ç�I�W����z$<s��!jjX�d�l�r�{��ߠ$�V�����6ʹ�+���I=�C=�CۿYuf%+fծѻ!y���)O�{��c���ܼ��ٟ`	�9��T�Ҋ���
m�(����6��l�S%b���es�������tR��H�I��sO�y�z{���n�|�ס\�Y���.8�r����y��zQ��3��?_Zq��pmT�e.سp�m^!ߏ7�;�|���7�W�bC���[��I7��̽E.�8������-�������q�r��{ˮT[)ꂚk���Zʳ��@Z�:��B���&�֪*`���$��z���k�����V�lTE|�	�=B|A�E�z���FO��W�7�BP�t&'���0�����`���<�#BZ��I�rH>��28ˮ�����K���؎�(�$�!��k~U�������J�)�}Oo���ޓ�=���%��W���f�u��D�V-+I�k�a��}��r~�cnW��p玆���	�ӶB�F��̇��9]�O4�tg^���W��tjB����Ou՗���µ~�)�ʊ���N� �|xG�xX��$<�>&󖬌��xK��b���\������W+�5�V�u��!5�bp���'�@6���L��9���2φyC,����F�5�>ag8B��-t�Z12��n�:�,���X�o�ZQ�)coʲ�;�~cz2��<8�k�m��F�6��: /\��>4�/��G@~���.<W����Gٟ�����,����ۦ��4u�8�W #�Y1C�$�7{o\1�(r�p�U9@<2�=��SN>MyM_��?*�� ?m�}���[��7\�!"�9D�W����_���+�7Y-+�9��u�{�z$�mDV�0i��hȚ�ޖW��U
6zi��@��U� ��l{"s�����
�!V�����j�oٴ٫��|?q}?��b|�~���� I[x2Bw0(�'yg�i#�&�¯����6
�Q>T��K�~�C�U��w�-��m�@�xS��l0����E�K�<7��d���u�:;-Y�tfK�-�BE)H˯0]��0R0�y����L]:�jUY�F�.��e��8G��`���E�O�K�j�ӣ6QAK��]�E�\�Lc��	�ڠW�>35N5\t�kʙ,�A���gr�w&�ŧ)�������-(�'�^MAb�oVT.��+~��z��wEO����K?����C5����@�Bfy_�;z�B��+���97�.
C�T�?�o�"��;�)�?�
�гq�1�_��-3D�@��zU��6ر�o3|� �YRTQ�#�6ƒ�)e�U�`(sC�bw(��,�E5�8@�Q����,��!K�mP(TӚ2=���-�$i�1�D�*J
Դ��_#�E��MT���N�$�k@�����t�L����Lɖ߮IW�lkEQhţ��a��sa�O� �
�\/��� F��#�h���������c�R�T�g�TM�^[+��9c��6,̖�@���k��/����h;��[9��(��\7FU��� ��)(�Y �dDmx#�SV���!�$�c�-덶b��[49�)�"4n
�hY&��; '� ��K�X�e�[�>���ᜦ8��kg� 2����7
��D��۷�/���z���:C�˙�T�hhī9G���w�sVv/Ѫ����ۖM���'�P����{���aSO�\�U`�\�zj�F��ީ'�QO﫥2ɯӿ�#S��T.��y�Cg�DI>���d�&�,��",?Ǚr2�V��{�"x{ifY�f���k��hG��W�2�E������ҨC<�xb��l$�֑W;�8mi{K�;.�|}:�xy�2_Ʌ*Wf�" (Di�Ğ�XL�
J"����=f��D��]D�"��`Ay��b�~�n�5xd��ʂ�zT��42�ц�Yq�I_�0�J؉�p��W
���Q���2({*��c����8"@�`����0�^}�v�(o�S��#�qLڙ�l����v�3�_��'#��~��v�0�^���&��t���5�j�eɄ)�"Koi�����Z����!�����b�B��̳NWoK�������4,��l�,�Ba���;�$΋�U���^%*�b1x�_~�N��(�ˊo )�\?�1c�_�׉�������p+~�Y��mxm�W��4�����1��K���UW}/����-��{h��ƭ�<���(Gatˇ�>Y��� ����:�m�=��\�@4R��L?r,�7!(~G?cd��k:;�������(�~�06�����@�h�� ��R�.�?�8��C�j�g��y��1��aqO����� ���ce' 5V�����|KI����c�V���e�4j���b*R�6 pjbR�ୡ����yv 0�?�n-�����yic	o��M�<�t<FV����#���~>��Kn���l<�!S�MǦ��嫰۸5��& ���YM(4n�յ/� uI��砤�U�*j�Q�zg�'_�)P*�y����+!�!����Q�DXiR�����OR�*��#�}~ ʇ���8���$]Lz��mBVE�������f�/�/�ٳZ��_���9/O�A�B�|*��Lx�G����L2x�S�O-ż4���{�.I���f������궤��[�{��f���~R��A>�r�߉3Ñ����b͸�d���B"A�><�"f ��H'Gٱ�`��i��V�MW�H(���ږ��������o^��J#�ܛ�����>Y���:=K�K�-7��]���y���z�$3z�H��=I3���>�4�n���;$N�\H�ƭ_����VY�RӇ��O|���"�f�Z�E�D���ȱAl��<-F��<f�Fóf�
/t�qC*B�h;�p��d@N��Rjg���$n7�R�o��4�c�-��o~��A���{e��7-��q�=X����1Qk�j3����s�V}`@��������=m����0�U�漌'kw��� -���'Փs�9g��"�S�
�@�s��@7�\�q���a?��%�@kz7�{0�5�I���G����]z�*X��w�[��@��A�,3��}��$�	�B�/�+���Ϲ��В�p3����jw��w�M�7(�^ŏ~��
t~�e/�~� ���Z��8Gv΋ԥ�_��B�y��{���\CۼR!{>2@S8z��y�����JRY���@�'�{u�'i����BW�\ܠ�
�<:>�(�)ܖD���ePx�,&�ʼEW��]Q���������D9V_m�WAN����5�$TW���4S�痒E''V�;����u�J� rm������v\��0���?~��1��&�bZ. J&i�Q����o�i�-Bfӡ�Y?����L
�4�^CU�q.G�6�E�W-)4�D�l˼*��y���$%�\*a�}j���?��`�3���l%1I��0?�x�0;���f�_�=�M9�f�7m�2�$d����Z3V>`4����j�tz���<(�I��[�z�d[�<-���y ���*���|�U6�g������غe�8�nMU�v���^���bYQ���8SMÊ�Aw䢋��N�Z"��;������r'mۦ�$;J���r� ߗC)���`l�b�a 	�B6�Ō�e��o�=/Hh�C���n~~Q�[�v�z>4�;5x#�k�ΏwЇn
�(�"v xxU4*3��R�֤��#���:���y�miU'��p��<9ݼ�P��DMTŨ2�Ҩ`�*��'�B��ц���/����m�k���x�-��(����T5ܚ�;gޜ�|�����Z���wN�|6Q��vEV�<����o��Z��[���F\@3�6�<���h)7�m��Re���v%��1¼ž-r�:G���d��׊�`�Ea*/�{X՞�}�_ $�7���BG����t�C��������o�[t�O�Et_^5�
����w~[���CH[
��}�:���ϒF?�i�u�
ץI l�#l-�2
�g��(.�뱔s ^�KT-�s� ��_�0�E]ؼF#�G.b�;*.��&�Y�5���G�$|��
w�_�D����u��d�.!��d&��Kg�4Qp���h̀�$�ʰ�kA�F+�AO~B�\����ǻ�E^��۠("D6PJ,�Eλ�boAt#r���G� (R��ޗ���Z8�"\V�H%��t�G�6
h���O��0c�r�v���X���	�����!�%,��;6|�kzʎ��Z�� dZI�{�'��d�Ad�P�CAx�4W�R��N�f�?lHӎx?(�������uT_��WHZ�𡣼�kɣT]�G�a] ������s�d-����ñ�0pd����Pd��5~�F�F>0?��x �Xڳ�7g$*=P[�a�����K��D�,l.����kF
�0H��0u��W���@��?��?�F{��0��$��O~�2�d�Ǿ���3���Cj�IFڶ1�1~�ED���t ` �=kk`z6�'������ڀ�i��m
 p06 #�����7�)�G��c�!Ղ���V�)�f���] ���m�a(�{ls
���~FҲ��ag��[n~�21�`$�n+B
9�@�p� �C @��k��y~�P���{�0ޗ����R��*<��O����}U�S *�#�sco)N��Q4rC���q�\��s�R[����Z`���O����y�Q�`��*%W"�����VXGd]�#�BB��d[#}�2U�"�K���\ R�!��zM��	�U"�L/N/��
8b�:½X�'Y��e}�>�ӵ7�4B,|em�<��-tjs�#�X��{=�����Q4̳h��ψ �:r�`�Ng�4�!ݟ�*�čr�\Å�3¥lmJJ	e��W��QJ-N��E.|W��_���"+��jj��
��ɑ+�v�#���,'s�^�.�v�����[ɧ���n�(�BM���ױpX����Ǽ(�@��8,�UW� �5W	x,���@^�%�|7��g|��w
�ځ��B���oG��@&^�Y�-(!�?\���]�i����)r�j��ix�W��Z�l��k�_0�0�0f0�07�4�h"�E�R4H�@)��ǅ�؀cC$?����h���.�{a$lr��-�b�.�7m�'w�z׻�sa�3�w�k�8�~�{�%H�g�jA�" RA������4*�PNB��{����sA+	T��8�B�"W �s B?�#o ��>�7#"z��S��6}�{�+�׃9
Æs@�A�����.���|` �Zoy��ro <-���!�� �-;/�MŎ7���[��D�PI����a\$����q֐҃R6�GK�Y�ӢhRV<��UG��\�Nk#��\��E'�hE_�S��:�o^����8@�,*��4:TH� ��#*s�ui�8r�ɑ6�e=��`��T=�#�Op���Q80�S&�H�|!�&d��9�g���q!��r@{�Y��$��Yq�+Ҝv��F��-�(ʆ���-��.�-�+E�O�so�5x��a V��#�����LL? �o�i�2YtR)1��]|GH�Zq��x�"��<vlZ��*X
�b"n�"4.�B�j*���MY8L��c�"�J�W�B����E��Q�]z�qIj3�:$X������JL˂�!�ʪ�X�U��:�x:0��t
�9��=�6SoE"(x�}4��F<�zU�$i�й�5B���~���@�s�N[��/�	.'��צ��V�d�#��])'M�gM��J�,�1���f�����p�߫�c9O\?� %��b`� ��_�u�uY����X x�0v�c��(�+�)����#���+OH4fqa�GB����'&9�)�P���H�ρ��u ����(��E�`ȵjlZ>#^�3����q]F���^Gt?h�X�Z��� h�8�O�c���8"�`!������AY�)6�>C��>�#�{[���$�gDu����+��6�`l������5�D�(��u�-��?|�>�����X�@?�h�-TiT��k��k�V�g�O?�� ]3����& xkk[˫���9!�&�F�\mw�ɴ�FL��đq�ɢ�y
�k��I����cZI�ޑ���dƃ��Q�~�Ӛ.�:�MD]PI���@�����O�Xv�>�&.jx�+І�7��b\ t��w$B����G��"�>w��;�=B/"�)!G?<������p��f �S(��F�1<!)�H�&.�1�f#��Ι9�a�ԁ�"I+e�ųt����<��ˑ���<|+Y����Dk�eb����82�nA>,����"���|"�4r��}��X��B3	*<��s��TS꥔^p�hx�nT�h���#\,|��i�.����W���di! 
��a`Q=��!i��:���c�.��M�ʹ�
��	x�Xl���lӓ#��g�R���Dt�̾}��P@���"C�R�z;�E�[',VE�� <x��ģl<}��U`��0h /��pP�gp�0��#z�s��,�)���������1sF�`����a0�:Y�a�t�*��yx��t��s��{�y��F�)4D/0�F@E�`���|��j��<+��Yd�D�p��n�V�WQ���ļ��ɝ��ꪌ�C��=��p.k�%�`Q6����r\���zB�ЈkH��؇���	��<6n�5��³a�� |2�\4�P�蚥�p:�V�1fl���}��tq v͉�t�(�9��U�þ�V�敵U�z�3�{�ϱ=aj����2��b���lw�O��m~�:51M���֌�FJȝ�"mR���v�5�)�:U�ifj�fi�9+a�N�G��Hz�� �R�.�ph���U�B���V�B0t��ީ���;jm�=v�:�����4ab$�~�+5�B�B��������jC��Z��ET/Ś�"� ��|c�X��=Qo�Y�]���W��n�Q$����n��D�9�)�������@�?����dPъ��9�HFki��(�<�<�l\�T�L�6W�8�8*?o�B��$5�!�b�<p��o�9.n�i�r38%�x���R8]���+�L�!S}^�AB��a�O�_}�3A������뮥�J�C,+i\�l�E��{�@�bjzI�:x-���IJg���`�=��;��'����.��KK��HEQ��[E�I,r܃��BUuWHZ�3��u,��7�
 #Qnm��6B�����Ea{DT�X�l�n��7�c�F�M��Z �����5�oe�!W`7 ��2|�RC���f�J�s���� 2���4�� t�F�f�z��_-�/ l�7�*++�����úk���1���@��Pd@��Rn H�� ���C����o���!J%ݕ��"�Rp�'����EV�@�k��k2_��{�c`\pm(�����*� �T+��������D���ϻ��P�) ����]��G�����2B1��!w���c�	U�I�
���x�yի�����G?��r�|��8.sݸ/�|�FJ�y��3�0Ҳ
G��.�k[�B`:Ω�1`c@�&�BE�|I��#?GZ�-��ե�ϣ|$������b��P�8!���JR�>�!��T�N�`R-L�3���D@Ŀ��k����N!B���{��X�&�!r�W��B5|�'W����#TQ1�L^��
J�Զ�w��"v�3މ��6z�n|�����ǲa\����"$�QSC�{�C��C>�:7K���Ęq�]d>�����3�X�$u!G���*�K���&#�4�?bP̳}�!�z��y�>�X�Zw���,v<�Z�Qo<�9xx��c��֟�����Q�R�N�데6�Eu�{�`���m��+)q�DK+����k��>�P�o3�b�]*����.�F T�����s�;��ޅ,���`L���-�0�VU��40���㼑�@��E���5�a||Ǉa�y���׌���PYtضȏ���	57�-����F��s\@��ٰyb� ��c���j3���3��҇��+   �����]�A\gp"��G��}"�p��*芈!�;�7�"�D�c���H�ac������9֪(�/���7����i�(�]��i� �@k�EҬQ����m�s��d�C��C*����j��	W"��a�!}��h��'�'�<��"��N8Boa� �$��VQ0G�}��4N�	�6�J2p�G������|�����_+˶��ک��mk�q��3[�j��Q�L
�ɘ׊�P:i�
�� Ge�|ӴZHqH����n�:�vu�l� +	��t0qL�n�73R�d��~M����SE��Dc��j��P�AJc�FUTA�ʙ�U���]ᵪ_�]3^R��DߍM�5繴�3u�2�����j��"�/�(4�%l��?�^v���H%N�6՞���]l�2�b�3(�(��(*�x3�@fJ&��4�[de��(,;�D���)���.4Z�����Qn���f.B��VN>�Fs���E8������#>�a��kU`���Ч�U�T#�TB� C����/`����Y�q�V���a��MLOG�eiiQ�UTVlmm(�F4+3�R່܀C�ϘA�!�Y�À�,[�W�f����{�c<$�շ(�.�	��ma�'E���� TS�DF/u ���t��X����=�ߓ�$���\��r��Gp�x�ɩ��0޸� c�	#�NG�渉�%�̸4j�Oڳ`�r���b�0��0�]D�L?c(τ��@�'|��Z�]|���1��d����g8��֦[�6�j�!�@��ݳg��׆ߦ�j�&�ۢr���Y�MSB
�zs�����rh�B�"4��೨D���c��9�>���[Wl̍�
*"�b�>K���{�f[�BI��-��&Bi�U�:�]�"�J#����#*�,��z~�y��$j�<��4�-�t����!�nD��H�ؑ���[�3�ԛ�Z�n�f�C�р*�Y�xLT��1��kR�_G��FmJ�)�����Zg�uq�F��D�D{��C�w��d}�*��?U	B�.�v���
�~}�X�cƸ�9���rǆ��rcU-Q�B%��D+�B��Ǖ��27��5�#�"���Y��FV���<�n���(�HK�xc������$tz+���5�kQ��S���o�T��F`�C�(���0��N���ʎı�^�dUJ{���[d.� �0�?��7��y�
���[�G�E$�M�R���8x��Y������Ũ�H+*p�EH5\Rϛ������>�/�T�ԫ2�B���j<�\Xi3���|��:�'<X�u��^��y;`!�4E{>� ��::w�7�~`4����u�����{8/D���R8��w�j� ���TXH�y+O�C�'@�/���~^V��0Fb\]o!#"[�?�Aj*U�1q;;��ǰ"�ŵ���{��"1�T��8Wp����x�=4r4�P�-� %� +"E��
N@6*��	��_�;�`�x����_�I]WY��{q�?��?.`s�Y$���&h,���N�Xˠ���o}����=tܕs���z��G��x�ǅݵϓ��`�n������qE�z"���Պ/��v��J��2��׽��p=���?��x@�ׇ~@ ��ñ��]&�B����5�;t��z���˴q����bc�@���J���*M��Y���i�6?�Pp6,�y������\��������ꁑ��g��Kʶ�ޘ�y�{�ۼXu���B-�7���Q������c��Ԇ�l1H����9��3I��#/��g�xy�n�0bF��^iׅM�Ic^��:�:4Q�J��GIQ1YI=fn��G���Z��;`�BsIEQF4�`Ӈ���sB."�o$چ=�}B����H�Chu�A��n	K!����oה�D�%|O����q@��9<˗��%�@��o�����"V�`�]#�Bj0H�Ѵ��AZ���S��E/�M�*�V$�o)�ۤR����Ǥ� +�:���ph%�`�Z�r�}���B
FǕ�v�?.�EZ	�v�M(�t���a@x�g�/�f���k���~aM�Ut)��'�r@*-���� ���A�4���g������h�����C��d�}r�$�2`'"{.�q�����k�3.��-�oϖH��w�_���������d�9��q�"%�s?�sr hb�hU�XՒhu^ �ő����t͵W�>��OW�=8z䄀lp�q�f�Z;64�q���ƍ�A�E���;��]ҲN8,��D	S�j�xl)��Ct��'}�M�;� ����pun��&1<~�
��?�s�o��������6I!s�̡��3@m�Ưn���9r���Ϻ�/5��O �1�͢T�E��t��Z�g=���>E�f��Q}F:xW�D�>�e�Mԫ���Ђ;i�raM���6:=Z�5������7��#67Mս�4��Hi:>�%�O��յ�b��`XT3���thi)�7�M-4�Z�G�U���x��J���.�h*9t!�,�h�t=u{�L8�(�]�Y�]��i�?z�5����P��~E�X��U�f[R���h)�z/���v\�Iҹ�!p�_���E��p�DJ�U&x�}�|'F��Os�cdQ�/W2�6w���t����:d$�-F�����=�蔚dU]�R/Ns4̂�s#��]��o&Qoi�(R�#:|�مY�/��
�cON��m	����ģ3އyUY���f{0n t�����籽�)!|�k8L�(�roM��<RD+���Z��O��|��
�67}`�) 0��<%�lA*0>�OȂ� �*0�J��aH���_�'?�I1H-�"k�GM*��Qq�W^y\r�f�LQ��6�Bǖ*B�� �HM���*�`��A<���|E�7+<(0�j�w��0�ftL��A3}�0h���k�����fH���D��"-v>؇�4 |p϶���{��"g8�%�m8pG�z��ǉ�t�bks]	�Q�W��x8_��  ��m0O���� �ai2 h�������nv{��'�E/�Mz
A��妛����f��:Z�)L��222���O���]��(�����X��A��NsF�)�x./80���tsF@����_x����$�W$c���b�L�3�Ęʈ��upc.ᜳ��L���:g�1o�S�k�Ղ�.߃M��v������� �9_K-�>RGk�DV�V��������'�T�"�Q�"5�nF�-Z0 ��y}!���m�b�z����:w�.����V���=hu����o6���F�ڍGER#�����=��������Z��=5�����4X�9)]�;���l�U}�j��.�[�l	`��#L��"/�ԭ��"��O��ƱFH�g�>�0�kd�K;�&.�� afZ*�%r����D�U�5�ʡ��HU6�y098�P��bu�bx!m�<s�m���Q)\ۛ��+�#"0����d����"#O�3#��"��'1{k���@��xbmI�/��F*#Ҋ*��ba���{�F�=�``Q�poꈗ��baL��u�^�W���wi���Y�J��O����?@����bdlq��n�����vѮ=q�^�}H��̲gS�Нw�I_���̹Ӣ��u쩢'��l�
0�Q6����o�����o�߳���!�x� t�����2�˟�	z�K_J��;���&/��l�y���'�{����~�#�䩧$aiT�|�`��Aoy�[���%�a @�'����xx�x 04�  ��,{t�ky�_E�>������9g%������u�|�-��׾�^xۋy.ht�fl��������k���2ړ�Ն����X��� �VV�mcU��i�~/����8Pl�r���  ��oQ �7��uz����a����~S�7� ` @�c�������TU_�+<'��
f �,]��ǔ�\ǃ�����U���A���߽���k��ȡâ��������?��ph�]8O��t�����|?,�8��b\;��������q�0w r�����\��8�^ܨzѹ嵺����A�Ǹp~����?�=Kx�>�5 6.���]�f��J�����I�ò�p]��BhZS⑦9�z��n��Т��Ky�"��%1�2M���W{f�|vz}:�r^�b*� ��"BA�Q��o(g����߯��Fk�f�[�� �Y�S�w�����D�(�[���5<���������|��<���~�"�w;�$�,���Fo�R$�C|w/.,>��w��lX��ޠ���;s~����k7{����+^p��S��m3`�YڋN}>fc5IE���d,�,F���Z���T�D�F�Q��(�����3u�$I^T��[��8v�X�>I������%,���#�Mp@�FZ�B�li*�Z]�;���!��|P���Y�@Eę�\�B�Z"-�+�.4�"[T~'[�fg�@�Q��k2v!R]HU'r!�3��>MA�8���~A�����\�*���aQӮ�"-�G|шd|��.e�_��/�/��/H4 ��a�1I��`���\��uA�����e����:����+�:N{U=Vy0u*�gP���O}J*R������"��^Կ��7�j+�5�| .�h��8g��a��?(��|\7JM���ΰT�Y�7��4��}{$�
ȢN��60�ڴN���jᘸ��NCZ���F4	�TĀ?��E|�Y�d2d�k���ɼ.��c�y��)��y��I�ى�Q@�VVI�r��`�0�7@
"Z�����6�kHGt�$�c�9`�R.���>�1��5��>�Q��5�%���O'�=�A�A��
ݟ<� ��o��Ο_��&�>@;��O��O�=Ǳ?�{�/@����~G�?��%C`������;қ #y��yI�����y�����c���y0�J�r0x�P".78�!p�r�:����ΞjIb�GJ��"�S���؍'��"�j���d�����hOF��CfYG�s�s�)Un�Q�VO#.��\E�e/~��m{�Eh?�f�<��V�T
g��
0��V�OmDǧT�u&���;i۽.��ޠ��Vڝb���Z��F<�����{�욛o��m�<���`��������L(vZ���0}����<y����o�����y�U�-��q�R�
;�h���65T���٠Hd ��J+|���_=˷���̣4.P#1�+�LH�eSx���0�E@�:d��뇚!������-!-b".��hgi^(R�H��Uy��GPoM�&�ep�@#�e(���*|V��:t'5�ŧho�ܵy  �I�Ah�G�i�$K�u	$����9������-8�U6aØ�79Mt�� ���Rf���xQ23�/e�-\mH�X%j��K��A��� s �|�;����Fq��>r�1^̦Ń�w�{��g�t�M7JI��~����F��B_+9,UF��!~���#}ee�x��E/z�7�T���)�K���� :��"Xu�H#������r��^ù���|`����/�f��K�ǻk��Ѷ�Dq��Eqp�Bb@Q�/��0��]�	)]���Wr2Ȱ��˟1r�U�`�֬��ꊫ��W_E�Y{<�R�g"�}� �u\�i��a�1N&(����7��I�ay0�������(w'�>B�N�V�V��?�W�q��'|�.Dю=,s��2����R��׌��&I?���$�#V��b�y����*_��X��fsNR� I+���r��������h"�Y��� ݳ�C������-���IS7�C�33B�Fu��)Yq�p/b���$"U�W��X��Q�`O�#� �2H��qp�0�� ˂h_(_��
ʐ]��� 6��c�v;4d���0G��,uy�Y�w�;9O��P�Z��ᠷ�<^i���u/|��pÍ'����v��ݱG�6��������k�����p�7=�0=;���2�5>ɫBG(2W�"�������K�r��¨�8г|�l�&Ɲo��<��H�(���+5���x�L\�kd�ʑ�ɳ�=l��}Gb2үc�體3�3��V@�I���	@~��C���ʇqJS;4^�ijB�SV�
�X�<��*Z�|�HyVZl<	;�	�Y��B�
.4%$uD���pkBi���-�k��$��Ɉ���-l/��>-�	� \X�(�#$�!b
���Zh@���ZP����SHC�6<z(��h`�������� )�&�K/�ċ^�b�G������]Uۂc�H�
�-؏oq]G����d��6�0� -���R��J��:6��Y�c!�i3�1�,��P O����u��J�O�,J}4��$� Bg����v�cb��eJ��4R|�0r��a��H���5�`)QO�R�����yOb��ȼ8����Xn��`��} ;D��)q�r5Ƭ�`�ʹ-beϝm�^�w��}GT�����%�s�D�c�c ���`�,³���x��y�� �B6RC/����]t=��\'�{��d'�l͟���uki!�ҭ��Y�Bĵ� �ˈ�YMl���?�3\j�ŸU���}��H�����k�?����5T���#+��A���!0WMD�ܢv!PB�h_B��)u�p/�fi�1E����A��܍\�mvd��@�%�nP�c�繶�ݢ��-Z��bm�s6�t����ٹ��~�m/����[O��5w�~�ݿEO������������7EO<�$�����i,Uj�(浢�;���H>SV{�+��Q���Tt0�q�xy&oQ� o#m9��5��ڸ'�#A�VD_П�!��AEd���.�h˟��w���@z�=��n_�
{4��OF�?�]�R6�c�"���Tx5�d7~A�.���E��c$�uQ"]$��L
�+�K�� �P�Ἂ�Hte	u( �9]�X�d5�I�/}�w�C��V���a�	i*x-�*�x���ixحv�{�FLŏ����l�810���00zM�t�mwzrO���IA��O%ڳ�P����Y���6��1�����Y��Q ��Ѣ���������"������y"��JX�c)%��)��X�Ζ*�g@���C"Q8�
������R��5�����cC����*�#�i#�:	����#�����0^�P*@)>g:'�|�'W~�h���� D�@�F���5�|���&Dp��~��������׽�u *�eO5f��J�P)ầ>et͵W��G������������?.@i4B���~,=,�WV��=��/t��1�_�������XP�� ]H!� �3?�3����a��s7@	 !!p�=����*u;}IUV��4���	�{Q 8���ؔ���C��Zr�>JK|B�#¶�Xdٯ�n��[a	�w��Ԕ'*�Ɖ��( �*� �2�"D�$�?��#6t
����+���G�Z���y^g���R����&k%ۂ.���^���7��Us��SU�dS�<��9v
6F�b+N���/��C����~��~p�?�ޟ�?us��Νw���ї�.<�����7��fgO4�#��J2�T��y*�D9�l�ej3���.��G���/q����\{rҀA�5w� ��Op1�U�  ���>r��,jUbJ-������p����0x��[B�N�Z���V!�vY�4	��%��dv���RY�ʠ-N��
�� ����H�uL;C���i��+ȷ�(s� �Is[��H��LpT2�����a⥶0��`a� V7<��ғ�Ɔ��1���Փ����� �m�b'��	��@g�`k��%Gn��(�HL]�e+��<""�{�C�f`�<SƆ��{����	�����ؘZD���$��9=�y-D	`\,Z�o�>�#_^l�nhW��0��FH��b�_Xjo F��iTO��j�
��D�.^\�#G�R�>�P�f��5�3P)+b`���k��)-|)4,�i��Ѯ�`c$_�����0�/~��A�M8"F�����RV�BaLq�F�U�~L����\�����Θ�nz������S$�5��X�=���o���+N�&��g��zM'<1 D� ^l��;h٠�Չ��`�B��O�5{��n�;�`ck�}V��b[�KѸ�_��:���͏8O9[$����س�#��X��c=�V��	�*�s�wz"6�o�������7�ڬ�ܭt(����<m�Bc�ҬCƈ�˸��A�~�;3�LMS���.��:��
��/��^�5�V�i��~��?�B���o�c��qW�S��<���]3�o9���:pZo�A��Yk�)��d�|�4/��E�-��9��3yd���"W���a��Io#*;㏦Z�)��;������ ���ɿ���2a��g�XK���W��G�f���	>�J^��*������1:4 N
�|xK��(�Jɲ=�C�l�ʌ���0�BH�lT����G>�=��Tg��H�_*�	�uC���Z�¤��Wj��;��p���`q��"�����H����G��yL�kՠF7�);&��JzM�Îo ���G�"G �EۢEr�]��q?l��L�w؁ٴ?���{��=��o��P��m�,̏�T�.��Lj M�I �՜�q�C����=lط7����y���͡<z c�y bi����l��V�h��O��^���M�H�i��D	a�����
Ƽ��-_� @70��B� �o�Da �P*�q8�	ʹ&Hg�KA ࠫ��Ç������|�'�@c��)(�D�� Y��A��k8o�'c����!�g�=�^��P=?�H=���
��x}k�%����E��VBJ
Ƕ9g�1I�1�{�^��Y���R��m4�yT�W��5�Z6�Þ�㲄~|�����bY�e��y���(�ژc ϼ,wP����L��J��0@�kp{ئv���f��з�?���� �S��pj Rt�tm�9��Ya�r�L��  �pIDAT�X^v;Y���k���?�����_?L�#�;�yG�O?�_�o��`�'~���W���U��^��\w�U�p�i mm.r�n#�,�.k�g�BB���N1�|�a 
I��!���g�',&��DQB��M^X�@�ȽW�!��WZ�m�G�:�,u����� >�SG�x��fj"B�	,�a�AN�^@�ّrEX�!Z�H���E1�[��p��`J�Q��cCf��2WOХ2�B�����a��$pN�ôG��7�h�g^S��ԓ&%��cF�Ϋ(�(��g�ٙlQ l>d��D��է��e)[Xճ/�@��m�/��@��m�d����Bp���"L6��q;�y;f��J�,.��~�{�6Mō|�	{��I�c���l��42>� ��K�� 5lk�HT��T�;g����h߾%:{���}��o���_0�(R/�QXfC��j���P`�Ŏ  ��WW7�\+�ܓu@���O��O%:�4$H�F>�������<`�0H-�#e�1��_��_�.H�!�"uf�1� ���_�w��k^�j!���S0(9E������뮗�#����y$�: �8O<߽�^�����g�Z�R�����7�I�9�F��0>�b���k�). ;�w � �p-+���p-��i)9�y�1�җ�$�g@���a�����,9,�}4���b�Y	#�<O�<���k��hdC�� m.��y�������om�՟�_�T�U�����Z���X��
���U���.�=�zeE��6/4���|�ݯy�k�'M�gy�}w�ǿ��>~�}O<u��k�޷$����V��^����
7IE%q�H�>=˷���`�<�d�<�.݅�|����l��MY�Q8�SW�[�������Y�~��'vc���>��0/>{y�����Ce�]�E�?�K�E��26�S��� ����n�Bj	 ���*�K�ߑn{�%W	/�t/�������h��QF,��R6�\T��D�\b7O?^��'�ЈK��e�R�.F���JM��" fP��)�(0���:D�D�'	(��kڮ�Ul�?H��1�ٺ���6;ǖkFg� ��s4FL��]�g�_��L˄~�����k�a���t]���1#����mBV��9��Rx�i��<Y�,�8�}j6g��^Mo|�ظ>�?�������J�<�Ǭ����z�5���&y �Ǐ��=�&����u骼�  �l��L[��~�V-�� �k)Bl�&Dc`̱�}"(3���r'Q!��w�A���m�}@�����h&~pQ~�_�M�
-��_�6�= 
G�8B��v��!'���%�f�@|z���ꅲ� =��-�h�N8q�Zm�5�X 9 h�a�#\7�6f m =�'�=����� �#����Zkkl-ɰ:�K2������"(>}�Ӑ�a)_ZZ�L9�X�����Nr�?��Z�ҢS6��ϯ�K�;�X;zO�'���H��p�*��UiT�@��G��b���T���+ƣ�_wӗ���j��/��l��%�<w�޻������˷�<��t�X���F�`K�H��b�7X��ِ�U\߬~KӜz^}Na���e|�01Ӻ����-��]Bks4�b��9����U����=�O�s�� ?ߤ)�&�Ԙ�������[o���]z�{�C)/?�����<L_��7�K��[�:}�*����B�|�H�x�u�[�~홞��i��CYA���.���DM��;�ч2�#B�),,�ND�,��K�&K=`3/ڼ�0�o��L���m��FA&�G�7�l2�/�������d�ʢf��(�����ܒpL�}{m*#S�8 �cGQ��0�d}�,��#�1�^���4��+v>V}V	�d�ݶЋE�~�����t��k�}֫�&e?#�[�jM�Q���°ZWwQ5u\K?a��c��Z=9Gi�p>� �pa�2Q��c#� �o�B #��A� D^q \%#0��r�7"?��?-i"i�歛�����쿖#rqL�h
PH�@��G$߱(��P\?")8�� m�������wH�ɸZ x]Z?��z��~L�c�1 0��8~�^��V  	�V��F�l����7D�p��q^-��h���|~z��ӽ?��,x��lHj=Ҙy9_MZAx ��3�����*spT�%��'��b*p��qv��!M���������ƴ���B����_9t���Qt��%�����������{z�i���f�k�����oSTQc\g�N�:��8rQ������/q�G��	��$0 �A�e(^t���S�_��t�sB����@:Hǯ��n{���1^h�[m:��L�{(߷�:�ɧ�Q��a��#��@4+���_G?t� �y���K_�"�ŧ?M��NS�to_����J}H�3��W��( ���:���	p)%m<VH����l??��2/�+�-����"ء���1�b�aP�"�5�����A/'���1q��|�7��b������ �o��nD���T�F$����A�}�7�ש���&@�e/�����1 %�.�����$?G�I�}�g�K��ݸ(IZ�^���u)Lk�: �}��1²�cck�Ʈ�n~��B�d��ϕW_I���u3�F}�����o�%��D�҆C�
�m � v:]Ii��1*�0�������ʫ뮿�/�=Iǩ�+�ƿ�n�R1?�8.�&�����T���J�7�66�Q� �"!ʀ}-,�ɵ;v�����tIO�q"����ͮ��F��k䜻��QV�6 �|±k����a�gp��g�}Sl6rmiUБ�����Q]5�6~ ���k�&� {�{|]��^���C��F-r��I>����OZ���*b�Ȍ��Qs��Ң���8<�W�(�>"]�RTr-d�4pB"�	��%Q��*��]B�;�������S�FU�����IR�jL�~�e����=ސ���{���Ao��Y�U�a>�#�b�_��j�E�� 8�w k�Z���g�v���4�&����cQ���Nj�K�v�C�s	�j���~�F�4a���,����[o��_�B��%/�*{4��/P끓���A��tjs�Μ:M-���<A�r�t/� ���z��륌��)Z9w�VN��GﻏΰGU����LRe�a$ތ�kU�%y_<��xY�x�N�	� ��:U�'��#����<�Q^�T�F��O6�K#^u.�~<���W����v�0Z3镙a�H�,�Ad���ƭ��&��,xz���,���M~?��?!8�<���,�n�2�O�q�ƣVa�G�ŵc0�M��	�*�UHaߠ���E��E�����cmQ�F�h]����y��v�f�K%�Rp��l�q��d�ԏS��[������	K��Ǣ�#Jz�L��>�_V(��Y����:����������N�ҬDR
/&�nU�lɾgf��9 �F��J�d���bC*���Ee�p��9��3�f�*���:�[�J����ZM#F 2��ӱ��h�0/��Qy��'^=�����$/��{$F?������س�)8{""�R��d7�<�]�^��Z(M4!:5C�t��g�x�4d�]]�Hq����zWS��S7҄V�A R��������y�l+��Zg���|�w|O�.�����@Z�� �|__q���6-wےF��[F~. �BR�`N�Bz�o�5x����"����DxNo�2m{���������7|#��75MW�t3��������2�{�E�i�����:��iz��ǔ��r�N�w/]8w^��g��(�7h~�MgO����ЭϿ������������t߷�A#~ N~�[���:͂�;��h^f��i��Һ �\84�C�$7ކ<T�j��=ȉ6T,��K���.az!TX���EG�g�[�l3�O��G����!E4ƱQc*��}�c\m2~I�.O]*�1��2�0IH��9%B�M��<߲;�8ȳ����@�qH����;a���Ovq6����k FŮc3	-�c\��:J@C��qr������v�=)WF�):��$bBs�j+U�������e�rr�9�M�*�I�U�m���q��a� l�踎��m��8iL&�֨���!�9D�a���/��֜�N�xF���@UXr^aϾ�ʹk�*{acѱ{kה�*�`�(���J�n�tڮ�.�J"\�DQP����f���"Ρ��Ԙ��;j����g�y���s>K��ǶQ��d;^��G�2bZ��ǟO;�O���j��#����n��S�Q��A�H�"2/뮦�P�<r��P��`��gr�����3�������.�O��h�g�3����@�={���?�k�K��5
�����9�oz�� �g�vY��"�Z��/�Y,�9�E`��;�<�QF��iZdr�k_M/���Scq�N1@���W��!:un�?u��;r�Z(K�а�әS�iue��
-.�!H�[=����ڻ�����5FҤqf~���3���.5F�M+�:� ^�s�R(��y���UwDU5�Cp^r�7��M����醂b��yL����	�U�3�F%�"4nr>~�/�(�S	���J��;�0�`�����	����m��h�-s��UIƥ��	S	Nh�q���؉ZcC�l�Pdcc��=/��f
�Ǽ�p�&?^GX�f��hFy>��$�D�s��^>��`�+�1t��A���V)���zQ\��۱mlD��)8�{���6#k��aң��^l����K�X��}���@��Z�MCG�5��������}�3���	��,���-�e##�� |�1&����6�R��L�G��ٳf��vm^�쀁�pMP�3�9��$����D;��	�vNQA*a�L�F!����	�[��ߥ����NS����k��\�i�p�*uHK������1 P��A8�v�+�v�Wq4���+����Rڨ�����lԥ�rU�3���x�QY��y4�[��ϕJ?���j�J�'z�QwW�OX��9?�m����9:z��4{����Z<�Q��]w�=���3����V��FK��tJ���u�4���Bx�;��{9�=����/,����7]GW>H��>Ai-�? ��|��[]�F�X�G��7�����fUOC$��߉��nF.T*�OD>/Q>,�A�;3����d�^������p)���b<xI0^�� �4��F9�X\*�3�wQ�c�M��D��"]`)�J��FL&�8�g�)�8)���T�-���yI�/���h�)0��H�)��k$�����r[��	y:!���l�C`��Bp�������D-w(��X����щ�g�	D�@|���!i���J�<��1��pPG�U�ZYW�Ȅ�TƁ�����s��cʻ6&7�Q�zQ�m)��d�"N�̄��2])H $$ h =,�T7Ny��	|�(<�]r�?�őK�đA4 @Oދ������I��rH�g#�l�8�4a=3B��s`��y�5/��g��3���;|>�K-,~?��@��zPg%М��H�@�P�=]�ـ�t�E�5W��q���ݨ�.�YA@E�H�蘸����vyͬG<g*Q<���jk�Q����rKy�ʩ�g����z�GTp]RN/)��s�V�fuc>q	����s��g�O��P�yh,�X�:QF�X���T��]����y�x9e�s4Lkt����o�M_������	�(Ua�l�mR��M3�T��u�vD��mF��:���?~�=y�}��o�M�?���%��5��+^�:������cw�E��D<h�J��4{l$�p2	eƅv���l,BR\U/�_VS��!Б+i�4缴�*K	�w���|��'�:���+,u��/"�N�H���EJ�� �Z�'��fB}�݌o��sz��>B �Bl?
JQ�#�����œ^���w�w�M��� ���X�*�x����0�d`G��p�� �3C��!i@[D;��n� ��X놂|T��F��-���>� ��<�:�p�0"�.��-z.ip%���V>�M��rTL"�x-�p�0�VE$:K :�4	��<��;�ʱ�GY	�ɾ��C6����:�+H����ȑ5����Tӊ��\@�E�l~X���,ZЂP����0��p|@-OK��^
%�J5��`��ZN�z�Y�t��U��h+��;2�r�Չ*�&!j�5cekZ������v���͙��IC�)�ߏ$�22�J�޸�i"�;XG$�Ґw��;E�\�:x1lJ��3��=[�k7��o��>�-�n������O^�nm�k�S�X_��{NЀ����f�K�y�gE\ $��噼1�7\T����x�@�e��e��=^T��fic0���=�<q%�����B�=�(=��c�|~��:��x��[�2�Qb�ga�6.�Ш���+���� @w"�OӠۣ'�_�G�?I��/��{��sg�_�띴wv����&~��t����ą�T�MӔ����� ���(S�X�%y��z"�4-�JE��`�B/��V$E��w����2�h9�e[��t4zD�U��3�W�mn����O�hE��F��6�|�`J��@&"
v�̌����B;��L��x�&�_Sk$�:'C��o�6���L���8�"Z���A\��s'�f��l���a�,���Xګ$�](F��n\���*{*�,�}!#*����Z/��_�c��r-�Eʧ�x=��a�Mȵ�8�� w����L#?s �چ@�gF�����t��62UR��k�XDP):��Bx����9���msL*Gp�n�*�Ҹ�b�y��6�Us���ް㯫^)����O���5�/�(]פ�V&�=FlkiMf	
�؋�\=�t���BjU������i	�^S #b��^�rNG4Y���*|��(wϚ�:FZ�0)��
i��'V �]I�P��+���4�NQ�3�[{�G^/��g�"�V|@>� 	Ϭ�L�NNq*S�>��8��쨍�1��Z�	�{E�R/�n��
.?ܕ�.����޶܋��_翧��MO-Q/�h�٠-vdk���je���|�����/|���^��a;��{�9���[���L���/G��g���R�
[Q���޼�'EM�m^\������ �e^F��)���+5��l�$F7�A-�?���=�t�8�N�����O��~�Qm�0�ToJ�a�P�'IsjZ<�����?C�<Hh�^��/.#�37/����y�4�?s�O�^�����\%���}Kt�M7�����n����ō5J���(�GrMҐQ*�H�1x:/������M�x�H�������3Hx[DԘΘ]:�ǈ|x[����`�A�y2<��?�O/?���n�_?�r!��~O^_�������L��'�1L?�{���e�:$�F�����M���t��dt-`!��6Z��q�;��e�Ǝ����ԧ1�2��\O1�a�*���F���ߜv��4�q>��i>
[/h�
�^K�u�c:��y����%u	?�����*�%>
�g11�b|��E1�G.-�R�����ڎ ��υ��ν|�9^ߎ�N�.;�|��i����ƣ��9�G�BS�Q��V�+j��bLb�,e��<��e�yIsR�3�L����g�N$�8���U0�����e �������7�8M�	����^��o}����O^��=��H}�k������o\;{��դ��[D�.m\�@��&�W�R���\
UӇ�6 ř�$Z}�o�5xɊ�R5�c����P����,E�s��O�4��6����q��������4��: R/����g$ڂ���*u��t�Ӣ��>O�.{oR��i9d� !�K��-�w�U��FJ7�z3�Z���]�P��*-�+�u��yi�8����4*��=r��4V"�'��.SA<�[��t4�L$�sre��pL��,�\�����
��Q�H�����܇TB�|}tD�{;I��5Y�GW�IPT�а��c|!-	��xR�R��<��<&���>����������@El�U��䀢�Մ#$Z�]̹�F��4�g%&%bpa�~'�uٿ'����m�yC��!���P���SQ�H����D�TtQ�M�&I&��z�q���}t���b�/.E��'�k�!�����TE�K��G�t���Nm��p��o1���}ֲ\�PQ�Q�*Ax��\�%���~. F�ť�r�fdJ�w�'��$G�����&G�VC�8(�y�%'�Yw������E-u��J���� ��my1�������Fzv�P0��Z�^՛9;�H�	ee$�>{Ƒj/Z#jҌV�e%i)��L���V�n`�}����;E�<'f�gD�lx���ti���������ǯ����i������/|��տ������o�y�����L3n j��Q�E	�u����Y�'����B*$O�a��u	=���`�s��(�;`oiz���Ͽ΅bn��R�OO<�$=��z����M,�0�dh�1��TA�|-����m^先'�(-Ւ��������,-P<?KG�:A�^�����6�$����I��"���z���[Wm�������x��B�DZr]�GV߹0��ZP"?��-6,�bP�c�Y�����'�����x:��'�\�_�������t�N���N���">�A;=�0zQ^O��n���K�h��%Qq@��|�P��I����`n\���EU�s�1�|!/�����oe�p<E!�zV��T;f8������LF��8�J�����9��N��X�w�������$�ʤ�\4��R06 d���u����Z=/'/��r���y���G�E߬���ޟ��zR��x	��%�(��.�4�G�����s�y�F�44��X��Gi,c���B��t�F�t�N�3�l:S��v �3Xq/)�.�ىdGs*�/��Y�$�O�������ʈjH��ͩF��б�g������S��o�����/��D�������׏}�K_|S}�x��&�����N���%ed��JZx@�=	��t�x�bt�=yy�oC<s���〸��d�5g�$��E):3xYk�評5z쉧�̹�TkLI�D ���>}Z���х��A_J<��W]��:î,K#5��S5���^o�j��xm��E:xp/���uM7hv��{� �//S��Qg�"I�,x���z�q��� 	g�CT���鴈�E�<Uׯa��)_�i�F���Rt�:R�.vQS�-�Gh`K��w)��ax~;�	����0\j�
OB��Tڤ<��8�>]=v�Ÿ��?��D�{��g�|�>���t4RO�.#4Bq5��H��(9Ft>�����)�뒴-� �ߪ��S�*ˢ{ҫ�y�f3W�,���+�rΨΒ�FL@��heM!MT�ۙj2!�(⍒��%z�v?�=�T���PPQF�Q�<��S��,.D�ҩVYd�{!p�c9�r��=%�����&��F<�Y��M7&�9>��R�ݵ�'�
'{��~h���笋�`~���Q2^������n��y>���Ԑ���En\$G֏���	����w	�u�H������G�G�HംcO�*���nsu�Z�@�#�̔�Jf=��;��BU>��v���Z���u���ހNo�Q�ˢ&/�y�?���������{�'��_��'��)$ ����_�����O���7�Ug�A�N�Y��N���I�*��lA��h! ܟ�㋉X����Kӈ���e^�"��"#�!?	�S���R�z<!��Y�j6�Ties��<s��/�1�9�Hk+)�e���Jg�_�8�G����}�(�z0�S���\A��X�ͫ�W�'B�.*xHP�0�պ�j��ff�hzq��-QRK���ㅓ�~.C戒����",� �E���p"�������{�9Q1�V�ޫD�c�]1Ch���-PYx��{-0Pr3h�|���8��v�_���xrq,N%�ƺL{�L�L�s_j�4�����C�^��u������\����jD*�G�	��y������ıg���Ű���L�����Y�?���v�B����똼�>��+�i��(�"��K{�c����}�l��ѱ����n��X��$ �P�w�{�� Q�ǃ-4ݒp��y�������bQQ�u���Ҳ������ꝝ �_W����7�X��4�bUE�j�p/��<P��9	�;��T�ԙ\H"�ȹQ����:ݟ$�����yM޻�W�Ak�E=v��:Uu���9��X�@ܮ���9��o�Cx?�m�y��I5+�Ơ�_{�W���mml�o����;��ַ��i#�����w������<��[�*����-!�ܷ�L�R��w�H M�1�)!�bB���\HJ��ų��e^�fEx��(�)���8�/�J�%����-�O�ՍM)���d@O V�&>�~\�<ĵ���',��v�7�{�,�.�����������S47Ӥ��^�F��|��.-J��Z2'Q����Z�ģ_o$T�Jwm��8ƿ��y����N酄Mm���}���#�n!�	I�F�c���9�_�yB�4�t�L���0p<L�$\8�ߎ�I�p���z���Kɛ��zhT^X���S�G9^����h�O�.r"��0�G��P���sAԋv��":��L=�t��<��L=`v �c�8U�-D�'*�9�C��a�<0>���X4��D'X&�^�� �Q����f�lb��բ�:Q1����
���ȥ1��y�93c�(2�\��槌N1�b����=фN�M1�>�f��ae��C�(s�'UF��t
��ta�pK6���M� �&UnNk$<Ws&�����%�,5�<}�0׵�R�jRU�<�<������8xV&��5���ȪI��9i7����l�h\��X �q�D�E�KK�O�����!顩#ff�I3ق(K�>�AN�|E��D�E�\��{�H%��4���}͡]����3���NQ�8W�ى�sgo���/��핿������o_�oFw�7n,��zw���l���/_������/�=���zzpc*Yb;q͞%Z�T)�ڢ���DըP"�k
���q���i=���лߍG-�5��兦˓��ࣨ5�L�쾽t����+�Ɠ{e}C"����pLv �=����!xE�m�$��#);ͤDS-�By�����NZ,iU:F�;=z��'ܚj�&Y��!๹ڬ��0�����$�.e���G���eÏ�U�Fdȅ��i �#-�g����#^%�wd�)a���P�zMy8*���U0�ڤ��� آ����bz!Q4��Pb�Cc�( �#�,�^�r<�Ԅ������ h!d�F,���1B��ݶ0r����a<��B���|�א2�E���@%
@M�ZZ��z�;�'�a�YpLm�II�����Iɗ���n�2b~����o�H�J4��ǳ(�a@�-�H/B�H�oP�{j=v�Zw'����Dq	�ȝS(�G�Bo^��n�6�����H��&�o�)� ,��xk�'n���3���
xe~��7)��pUEc����\Т���85�~Z(�1@�=u���t�{o�f��߿�&�T2D�I$��5�oTi���Kc'�/�ȴ9�	*��*=�u�|f�kO�U�Y���,KQ���b0U�y���Ug�Ӭ�i�k�V֧}�9je���dc�A�`�߻���^�������k��o�{��?����G�]qxછ����������g�v˃'��h�}����R���S|�>��^~�M����Ƚߥ��WaۄqD�H���'�
��7S-���⠒V��K=��"�ة��H%5Ro�҈'_�Ǡ�٠#�`�]}m��~�>�j�f��4��a�A8�����)�`������^a-\����#��E�+0a�C��� ؅�b�����"�{�u�>�扵v�u[]ZZ�C�ssT�mI�(����"�j���1�K�G���gp(�����hi��/~�?�� �..�pBOx� <��	��q�D�@�Z�����Î��b�X4Ea�e֔@�a ACAtʖt�7��q�Ů�D�f���En<%�7H� )���#����	�/��;� �,��L}�/Ls�`�W���8ԄA�k4Y��Ѳh�o�Ph��s2��q͝!�� H���@�d�L�@v����842���w�-$�q��H���;M��w�%wO �Xc����ED�ˉ�U+54P��6�l�-L�h*#�
�*ӑ*K�Q�
��S����Y�u�F�@�~��d�`I(�.ET�C�@dg�ư���؎���B
�{�WT�%�}N�q`D��d�e�<#cM8�H��M�*q�A������}Q���v 1�b���q]x߈ �w7;������E3ub{%�� '@8�qK�RY��Q����q����:�Q*Tg���>���5�+kH-��1�������-ȶ>Rkb��p�l�y����8��:8�n��*ٸ���F�{��M2;��D|1F5׭���V�z3}��lN�(��v<�uDB�i��-����!u��������K���C4�V�%�97�J���������ݭ��/�=��|���tcR�|�f[ۇ7VW�ڃ}i���Փ��t-���Q:6�@�y}�B��ɋ�T��ډg��h�9�sIJ�yͫ� ^��E����HNӳ���K���Cv����X̠�����%H+�.Ov[ډ�����+�H��*|��ǟ��"`�:�bdA��jr��Z_���$�$�x�A&���c ����+j�]���Lc��g���yr����*�����4��]�&r��fr��r/���uz衇�hI� D�T�䱐(�,�R�ܥsJ�
����\KwI�@<Z�4 6H��8�ѩ�������._�lL���eU��(�*f�SSr�R�2R�Vt��~�K�\�ra1Ƃ��+�W�6RT�Pe��}Tk��x�
��b��2�nV�R�TK�	�	��RO�"�|3w���TI�ky�
��b��"a�2GԆ:�� �p��
8���R)��
�L~��
|�p(box��HB��ڬ\����{.K�]Yz�E�qE���(TA4h8ͱn�F3� ���9�0�hd[Ӭ����ACP�:�
�\pk��qs��,��WD�?g˵�*,��-���������U��"?�)��:���jp.����u�:s���߮������JЏ+%����k�#�^]�-����u��^8C����h��;}��� V�UܲS�RFu�<^K�x��5�x>��}-��D)�C�Aкd%��T��g��N�� '���.�H4���M\�V�ɜX�Se���}�t�R�H���r�gO�����N��L�p���H]\P��*�;���ڧM�Nf��s�l}�WϾ���N�\�й�g[��4U&��*/���S^� Q�R���c�y�};�Ҳ;���ޜM/�Ϧ�7�|ra����r���;K|�-h�m-F�U�{������q_���Y�_o��r��:{ry�����g�����/�G�i��NW�xw$~���6����k�Ӓ-���ِ�t�������,���bc�eh�ހL�	��E۳��ؿ_��	/_�w�p-�m�'O�l2�{vU��>*�?n��2�"��˙8�R���H�P���fړ9+��=T�hz`̜LG:D��&�,K8Ù �f�9T��T�/q�8�Xu��ش2�v�v�n�6~��G�XQ�O-�����f���>��?�?�ߌ,��x��K9!�k��ƫ	�Y냜;N���i��4Qb��+��Ib[#?1�B�/��6�dKGa�̍M������GiJ�t6����{:���,��qO���38�zy?9��p���=9�6���BY5k�ei�&t��:6�j���������3����Z�^^|P�׭���}t���[��G,�{��0�����~O��>�>��3�N�OjMd;P�*g�lٻ�(�*)�M8�i'l�Z_S6VP(%�6t�BN��� ;��D��]���s�=� �Ϡ���<�$����C�H�"8I�P���j�'m��8V�Hme�'0��ZU	GR���Zw���Z��e��7�/����cp��=��}��N�֑W�C=[@���G-Fڍ�(�A�w������� VCaz��&����@"������a�*��yÇ�>����g�� ���Gr��������<��:�D6&���+����'"�=�;���U������%:�*W���k?l|0�
��3ئ�s��c��Sj���
�)`c��1�qRNɃLn�`���{c��~���oC^��ɨ���}�$�X����C��^�q
~m�_]N�m�.������D!_���E������� ���OCi����2��uh�+�tg�U���	��L%��k�5m7|��"��}�_�������gY�0��gDѳ�y���zs܅��7*?n,z�]�?�x���s ��2����+9��ÝǨ�����pT�.#hQ=A���A��]+�[�S�a�$;�A0m;l�ل���mK= l��L�'e�����"���B4� "��{�!����)&�Ll�A�k[m��Vۍ���?do�싶��(�>��"�\.���9AK��h7Is&��:DB-ޗ��k����&㇚�jB*�|�O��W�����J%���^�k� �u,����3�����Y�yF�b��҂���\ee=7Z;d��aо����s����E�=��T	"k+bP�ފچ/E��w��{kk��#�6�
~���h�!4��,��m������L�5P�Ԍ��qtEp�T����N,ɉ|0a0p�b����=��3Ẓ��كW�Si��߼M'n����w8'�h�_����SC�K鎗k��0Xs?T q0I@N<��X���r�\/{6E)PH=~�.RB@5�cR��q`������,��^�ZO�z�ޞ�
�p+d�2}ֿ�����`K��G��E�SK&ռ�*X]���>���$�>�*�����l�>̣|	�S�y��1� +�ZjG;��(08M��u�����8�x�~]^IIzQ	#�����EQ�jP�O�*AJA����+2E���֓r:/v>�����?���.�+�y�</!�$������+U�:���ע��E����;Usɥ���-�>BL@�㹏��K`��_�+8�Yn��ŋ�p���p9�
c׃�Bs6�w����r�g�ص�veuPk���,��Ю��b>:������}��ḽ�f����wac~kDbb�6>;��[#��*NX�"b¼b�l^��~��ӯom��{d4��-Yƹ���?���߆������pss��{4=�!�����Wn�ز�)�o��v�C/�C^��2�f�d���ڈS	�#/�pv6��Ō�ojN6�vC����X�t��1}V��!��6�0O���K�ǲ�*fg�YX�����{�Xr�b�o�$R���a���b��t
�]a��KrVp#��+UaH�]�g���}dB�1��o�vT�,H�*�f$�f�sd�i�Y��z��&8�����Oh-�,Z��$b	 ό��̌=�8fY8��
Z�#�C�eg)׮����4%,q#XUյ�h�Κ����N�E��q���^)�wϜ"�d�;�{�CAƥ�哫��[�77T �(�|X��9�������y%gӋ���AN������f_ǅ� +���+��V�\�
�����4�sI�^�XUI_��u�^x�)xQ5�
LҔ_z�	nze��	�&��E�q ��E!�3L������י9֖��w�~�LFQ�b����~�H�S�o~7M��<�B�_G�T��c�s
v\�E6�X�L�~U������sK2��ݻ7�^;]W
f�6�ş�F_G�D�]߃%�;	;r_CWj2�'W�|H�/UI�(0���ώ�$��o*T�u�k3k�j������&��d���_v��QnB�֒�m>���7�8}~[ʾ��Ws�ρ����T��Ա!,�?e#C��m�@��@;Q�NfB�$kv����D�lZB��Cyo�ɳ����>s6��O-y]_?��Y��|֋�ʅ�Jʚ��]��_}?�w?������w�Co���2,��a��E8�yz��gd_�{^Y�Ƅk�e�S�b\�u����p:�Y([���w���^���D͇#�+d�백Ás�,,��07�����:<l}�y0�q��b��ȴ��L��C?d���81$�e�vP*�?����9Ӟz���~���bx���z/s�/�x���fbYR��#38�ܝ��N�^�.��Rq�����j
��<ʢGr0�񮮟(�8�Y���?�8���{��u��݇�x �a��t|2��Y��Ld4 .S�=��#jԶF�^��Cm�Sz��_�8Ȍ�BS(s,��bb6��1W�;�9n�gS��z�Tx ż���@���4�ڋ�i��Y�WOV��?�&J���#9֮JО�G�~���9ƶJ��(���|uijd<�v���}_?_5�T0�C�go�&�*m.<����~w��z�^Y�+��x(����*��;�ժ��K�����Ojh���I�R�Uv7�x��d�?E��E�a��ӿ�1��k	���k���B��:kw��A�����̉�ӳ�T:�ň)�=��qF��[�p���p]��J����۷o���T���ϲ�	���΄`N{���v!9ᙍ�6�,�X,��Ж�:� ?��	ä�L@�,�Uǫ�5��?�S7`�Zvi��7���,������D%���:�'�3l�����ZT.�Ru���n�M�%l�c�4i�����ٍBL�\�s\���զ#���Qą9t��y�L6�=:�>�3UL�����r�+
�� A0J�	���S���q�[2�;V"�[��#R	w��w�'�.,�Gmw'^�FAF#1H�Ւ���R��i��Xb�>Z�}1��&л��G�h���n��w���)�{�U�������������������Csokswv旆�V#�;�v_;DL9q���J+ɭ���f�i)�^��0/���a���U��E�!,�dvfi�8l�R����*��<��_�K۸���:��̟\���(���	$�e�_\:.��n�%�v�mt����U�Ѵ ���٫|�m��އ�U�L�	�T������$���t�z���k��՞��;\���W_}F�����pn����L�Ҳ��]�`��BO��X�"h�Ra��VG�x����*=t^����e�e�vP`�Df�hE%@)�2w�%���D��B}Ҽ����A�xZxeTæ�O��  0enN��.�)��:k"�{�B��� M�d4̩��؍� ���;1�3ϲ۰��@֜����+#�����~��2n��E��Se��R����I-�ur̋�C(���_j!�@���]UwN��/��ql����n޵6��
e�I-�eQ�I���?tՍ8$ ��"7P���'|V(�9%���Mm%ր�r��PNm>��2�!����>�}�Ń4*�Ӊ��x_9ǳ����'Jzo�h��|g�֤?��*b`����6$��jӚ�u��L災G��k|����'U��y���,������[wo�eJ�cg����f*6$+������)7�E�����-<PL�c"�a��4��t{[��(d�(0I��lb�Tvg��.��kx�������}`G^��O��W���:����u���L\�����������(���h�i�NT[�����1/T�>χ�p1=�^~�`*o�
�>a��U۩�#��H̨hYB��3{o���jm�d��ϡ%}��0>�
S[���W�΃�M��[yK����Zb=2�������&4o���vo�ff�Ϩz��ŵ��"�=�e���zH:[!t,�4d^���&;�%x�3~�}�qV��9�p`��.�p�&��lsJ����/�~��	/^���߇w��ǐ)���-�6LGaa�}n�E��˜��� dr���C NH��W3VW��K����;� �Qj@��
�[/��&��p414��c�B����dhx��h��2�<�.�a�RV��
��?����@P!e��?�(���?
���� ��Kb}�x�d(`l<*C���Y�_[fu�u�>�������ϗ
R:�CLy��"�/>=�r7ʟ
RM���� x�>I�'�Q�U�W�DAr�i4c�J�`j�3�sj;d����`3�n{eT�S���ꠀ�J���L����S��dq�'�m���_����70��:c��(�����l�l1U>zqr���3���]"�J'F�4>^�YtƩB��a�F�a���ޞ��uB6rmk���q����4��Z_Yp/���9��ޞ�����cc|z'M��{>� �J�2�D�� f��M{p�iF���m%��Ͷ��Џ�*Z=<�
\��ce�J�*�h��2�g[9��?���}�̟#|r�	��+�^��v�嫫��ڮ�����a29SJ[t��k��`�:���j\�v�q_��~#��p��\�j�σ�e->����Z/Tգr�σ���Gz{8t�A+��ݻwz�C��ˋ�l�OH�>�*;+�N�y�M'��]@��WĠ%r(9M�M��\Hv��Ǟ��qF�(�0[@�,N�e*�<��iwv	�={�g@�L�����������o���?�c���������IL�'f���'*��1Q8�h��d�����C��^����tj�S=mr�Ƒ�QZSH����(K�[{sKVw�%	� g�{�f7���f7�?���-@5�@w������_���7a\��yob>�m9���U(�e��v��E#���eG��'�Ť����B���/�/U^ʼ-�}X?�ä8���Y�}�,,�7����O�����Ë��a�]ڿ�R��u�*��~��yz�D�.�W�E���e;�P7Szv< ���"�Q����mT���kZ�8���,;���Y�^2�=�d0z��0�0�`&v��^R��k�:8v|�D"��t���-�f��x�(Ͱ��=�?~��"r��e;����E��_���3�ͩ7�L�xR�^p�wT��[x�Yg3b=U^�V�y�F���f���(b��2�u�8E@_�|�d\}�;ke��X��y�=We�U��m0v	��ە���5��6�h��0Cv��`��91hK��CWQ![�9U�(��� 3 ��j��X�o;=�Өry(�\̞��z�kW�vBCsG�o�>1l(���2��I�M'�,���GU�Y������F`'=���5�8��J��ob�WG�x@(m/W^��3s�����jg׶�&���̲U�zY߶�lhΨ��qne�����03������]�֝�L-	�tt~��0���:�_�:��6�>� ��1�	akAv�$�9�����7A���7�+��`����긿��Ԏ �{o_� �'�U��s=�R N�v$ޣ�0��~nl/Y�b�Z�
�X��F&`�Ǳ�Y���>�u�cUe@A(����JA���9�h�$	A���'Ǚ�HekW["7$s?4v�B��/W`� Y�,L�T�m��£"��R^y�X>���JZS�D�u����g�h�0�h��ބ�r/�,���5{Ű��9�#�öZ����_}�\��w�^�[�fޘ]��7_�:��_�J ���C��~�ӟ�|��p}}%��z6���B3�q�ʹ\��e����+Q̙�Z�jШ�e+k_��т�v�z��ls��0���3��?�OB�oBN���fggʒ��l���",w_;^���l�	��(�/va��������k���ꨒO�Y��ߦ���&��1AD�%��^������l�o��n��6��~��om�2�|m�j��/�sA� �~�̎��h��l<G�m�|��*<�?d��?}n�d)�ѫE�4=��Sߨd�F�ƌ����yvq>as�b��m1ت}��eԱ�|�i���??���0�����?�{"���P�}�?a/���j|Z�f�z�<L,���,�e3��,|����������V�a��woo�?���9hx̞>1�37w7a�[w����8�eS�W�V�4�I�Hl'�����+qKx�+U7
�������8�4)�Z8�*Ne�b����Cŕ&���G!����'Q�we���Aۧ�iODO�##�%\L�DH8T���&2�������2ӔY����!�E�2MW�
��j�7Є�;��E؃Q?�*ڰ����i��0�UȄ����ֱ0�\�����s�z8�x��~��4ҝ�Y+	!r��d�5�ϓu�]s�l�Z�-�*5��Д��^�=��= ��0�,��֞E7>ކ(�P���:�eN\X�_N�*�
������K��){���v�ؘ��iZ@U����
��N��(�`v�	�1��8F��4t�$!o�Ū�O��)���;U<kIi����+N���Y Kj��͛W���n)��T��c=��U�����:M��O(���.�r�ήH�:�۰^����g��Z���:����h�^�p��������2|������^�eD���ga �>/;��ܮ�	#�z�*Q�#�M��a�����>����[�3�����K�������ԗ^�Fk�3Y�ڏZ�2�C Ȑ��s��K�F[��oL@x��b���M���Q��:ַk��a'�Ii�ٽ4���8v/860�	#H�X�&�Ѥ�'Ag-��C����[���\Y��8�)D�w�E8nv�r��GQ�6�a�
�����C���Vv���"4���h�ͪ,��M�k��k���qd*&=bP�^�b8,� �,��H[�go|v>����|����ӧ""z��R����ZY(���tҦ��Ȱ;A�%*Ɏl��ZvY�����ե�����&2�c;�^z�d���r�'�k�/?
��x��\�jK�'��"+�BԒ[�ZB�r��fl}�G:k�uG�4f���&]C�%�29�ʉ� �)Mz�jH?;���7U,p�M�N�?�9�{�C5CN�0���јf�I��J��#VG%@��a,���PT�����A�Q���Gf��D�BJ��!��&rt����eTUV%Ɂ�MTr���� �++O�+jɀ�����^�:81^���*-���t݌�
8I�<v9����a�(��u��0,�/��H�_�U�L����0Ъ��Ӿ��D����*'=ۣ�+aVZ����Y�{I����X`��@�qkGc���}~a�LG�خ���#�ҳ����m8踊R�(�%��x4X�,ό��(~���O���j�A��IU�ģ�F�S`�pG�h�;v���\ �T<x�Z��w�4- {�L��u�-�,^�Cp2;�B�9��:�:��X��D�6m^���Xt�t~�v,�W�qn���G̹�4��ԫ���T��",W�ў�!��=M��JP@�t1:_��'�����I�[p����ʧÉ����}X�--�p.TաB��S�6(����Z�m����|�>�D�֚*fɺ�To��C
�"ѣ�i����Y�M}2p̊���>j�����Go�����(XzELVZ^Z�k*��^4����ʑ������w��.�$/�c�o���^x�Y]�M�Q��{�yV�

��J�/��Y��׳�y8���D����U�G���P��T�����u�y)��`�qԎ� ���,�ɯ$)�#��ڡ)�g1���O�G]�_��g�Ҳ��b޿	���U�f��<ކ�^�Du�8#�]~l�H�� E�k�.��ׯ��G?��f(�����_��`��y���O�0�&|+¤����#��N糙0	d�8S�xDJ72�����d	(�G``�L�K'B-1�b�Cp��"	)�ȼ\w$�=���>OI��2��%��c�_�`R �1XZ��]x�@�{�O�EY�p�id����iD52Le�'��?iy�ŝ`����Q6�| uAI�d�3>(Л�/)�`�9^|R��X�]�I�S���+���Ϣ�W��4�02�c�yz]u-��~Y�ݏ�6�KË"�>�;P;ikN����	�R��*��?'0w�T��q�>�@�	� ;?i,% u
8�%k���'���*��Kڹ��:�b�pL��;N��8��u,��c�9��x_���(9����Yw�፲`$$I�"p��5�V�;���o))�n�I)%�-[��z��^U���7Q(8p������Τ]5m���k��q��H��H8�E����&>��٢B�`2�U��RA�
�J{clA�Ă� �n��_c_����;��o��&\������@��M6L��zF`�,� x����Y�C_����Q�W���Wfυ��".X�K����qT<�W�� G�
%I�}�2�8��a���)��� �/p@�ȡ��[7�Ԕ�"��{���������'&�DEUx,Z�}}k����N9�=X:.z��K�CF�W�n�jS����am���u6����g:���F��N�$_%�{�F��yc� �~N�������ZF���-M+�W��g�G_~���?�>��忄w/^��a.��P�?��b�[?�, ���7�����b�@R����O>y.�
 '��Z!et��Yn�b
�[�%��C�<���0�&�P'ݛ��ĳѣoNe�p�W�nrF
NDk߈�<�+�i���H��`1&ú�*PHIʖ�D�cn��">N��Zh�Lw�ι����J��ذ�?�L�c�ڂ�P�z_2�]̸ K�A>�q�EO����(���Wjs�Qn�G���{Y}�'$�lF:p�$�bY��������[+M{�ry& ��M�����HS(Q�fb�}v�d���>����^֡�����4���ux��&8��ݺ��qj� �'��/xy,a �E�3r$�ss���n���_ir�!(�.����V�Hj'�H�qF��$�;k�/=�#���q˫ce��C��D�����������@�s��'�C9�,����WP�y���8OK��;��9�Zc�2������vN�ǖӉ"@U�C�dH��"h�b���q�m$D�����E�OЃM�,�	?�-�cWQc�tc�h ��T��0<7��矇O`v���b;?��O˫�ps�wo���w�8z�t\�9E(~���W�	S�T/�x���$�s���=�:��mvacvb��jr�u�*x�i_1���%P���%��}`���2	$U���̫�T^�x[;��O�1QKC���o��ƾ� ��m��ۚ��?���]}k���oF��6[#:D�J�l��,��Yа��{�o�������]x1_�W+�HHնR���s�@(����hl�ق��)2!��N،�>��6�M_aE��V}��������o~^���!��`���b@Dޔi�I�t92��i�l�ڣ��a�al�
���^S
pü�揺�O��}���>�~�J����e�|v�>������}��]W�W�ۜ&NY�;��!�*��ll� aJ��z�k�}��_�{ P��ȝ�Z�)�f��y���]3��tݭc.`<V)���몑���0z-&^��WFd�����@����H��	�l6���r�d̉M�̛gA(QK3F}sΫ���/����*!v�d��֍�㥆��H	8:\M7�p|b������R��r�1�E��1FɟO�jOm9H�>�ҤzX�*n3M�h����Sʨी�5p��4�2��K�5$6�Dd�^8Q���{����Wp�j��8�cڜ$x/oIf���)�NY��i��j���]��H:��SO)�����EDw��'�S�h��'�� Ġ3�:��6;�!s���FF���"pOg'�����=I��n�|�*T�J�@z��^�;�"w�W&��u�?� �7踃�1b�'��0>�UŎ�� Jx��$�8d�I��fĻ��9o1Z����	Ƅ���}�G���
�}}J�;�E�Ñ�u�/v.��fW���ǿ?�������o�ݫ�a��}cS�L N�pYýY�����k�D3xqsvZ{_'��]��k�Ϙ��3.mOf��,��UTu���i�� Qm��S1�P�"�N��x���'c���<�lW��IE;8H����<�A���Ĥ"��(�c�Bh�y�?�1H��F��C؆�˰�����ј�B��^����ކ����p�~�:̘��w��J��yv�`0|8�L����m�H�� �V��M��χr�hj4i�E �C=>��A���E��雰g�i���O��,�'@B�����Fi~�woR��o���e��Jyx��$'�U�y��z�4nǳs�$ݲ�����8,ß^�-�s��Dmh��VY-�:<r�1�Mt�D�rc�����̇��2��z��j�i:�ȻL� 	�	�a�;AF���@���Kً��H��ô���c[7]ࡖC�dF)K���d��>W�df�Ӑ�`0�t8�M�*�w[ׁY[ ���N��`5ЎJ�ú9�[�6Ķe�D�~�#��ڞc�����k5�J�@&��	<�A�Y$g��I8��o���h'm ���	%�G��h_��"�I�Mu�JAO��I�b�ȼ*�h�{g
��TN�TAr� ����{M/.���'ƨ@%�'�5炃��i�89��J��T9K�Ci���
r���<D�v�ޥVf��(�	�L�DŅ�HAAq�$$�:��Y��.�q��y��K�Zc�aW�LU�$(J#`C�t��sӁ|C�~6@�υ�9K�?�T��zjQUQb�-U�$T)��P��un������`���
��K�j�3������M�e�F��؆�1�*��}��M�#��V�ITӊRӚ������Cf�
�~�Q�z2�������o^���Cxj�♭�U��� \Y��ʄ���/���A�,8xħQ:����wLxQ����T�=�q+>Zy�R�;n�3-�H�dVb�.���Zw�W����"%���AU�6K#녰�`�"u<ʞQe+4�X�������/�'��;w�|d�9S9fnW�,�CߜT��q>������I�7��bq�2��W_�gϮ������6O�,r�?pʿL��dQn����I h����}����wpb��]��*4;� ���7oÜ#g��T��pI{ae�#}Wp9�K�f�aR[�U\�@�����2D<8�F�e7� PF�5��O�=���9���2m�IT�l��T�b�LG2B��m�
�h�������3xA+O�𪔴-hz��I���DKe�0`�~ vL�2)&�y�C����q�b�c���J�>���T%�Ip�3;����V�^��,����}������ENgsbhm#?OA�*�
�\v��	���a/\��p�N<v�ζy�	�TP�����`0V�3��x,�U�A\���<*c=����Э���K[���1�M�<��7�f0��ɡV�����F��(*�~�ͫ����p�쩂��͛7ae�G��I-��d�ɱw e�}�)XH�ޔ٧)��t� ����#�@1s9��4:�m/�n|]@W;���`�J�Z��7
��P"���)��ħD�7	m�Jp�,��y��*1�&�d�q�7�%]&*g�/�_�����v���'��6�s��y�����#e�[s߇��9�O�}�sjI�ڃ�x��W��Y�N��L����NIA����������Y���+��*|��Kp���O_k=�����o�mx��}��W�	����+��������pm{�ʮ�
��Ƃ��1��x����/VL�9V�iv�$9OQ�*�Z�����r6/�&�]5��8r5)�?��e�B�@�A ���2�E+�����]�UU�ƃi&�A	�g�ˡk5��jog�p�^/��~�/����$� 3ٳj���N��ʂ����;MQV��Ռ�_}�y(//�7L*0/�>��y8��NF���ك�F6[m�6����A
�iV1
˭g�q��j��%M-k͛���/oއ��w!�`bd��A�:��Î(�T�]6��s�ݦ偱�cx�`�i0,�pm��h�n�jC����2�Cd�]o̠��hʣ��� �N�h�4��C��O�Ko8�AҰ�g�е0.�(7gj;�ܼ$�D&�FI������gw�cf䌃K�3�E���(x�J��c�M���벱`�z���ǉ�(m���p2F�P',��DyPBF��.xq��HB����"Ǫ��N�&4�#����a����}���X�KK�����z�����:���T9������64A@L7���VH��c��?�v,����zT[ gmA?B�I`��>N4�S;�8-��.>������~��������g������_[]fy��R��Z'��|4q�FG�^�+F�~7z:08��&UԦ�k_:;t#g�ɩ�����&r���M����a�d�e�WW�~���F^����^l�[�撐�*����v��Q#餌�@���񫍔uW��{&8��G���(��q���y79��z>�L�Z���U[=,\�p!T��[0.�H�H0���� ��7{�y"�.0\@Eg2+�g��qo^�p���W�἟�����ś�C�Z��ْ� eZ�n}r�p�C�Y =�����u�~|������@��#P��!wԙ��k��L�b��*Vu�&����L8K����G	ς�k�k�`X����;��X�}!�-̦ �q�>RT� Y�D#�q����$@l6���?���Ȳ�]�_��?�W�4y{���!�:�Aٯ���!�,������7���*������������p��0`�M���0d���Y�QY�䄗	[������K�P�і1g=���'a:i��v���3ۄ}{���w�~wf\ v� ��'c[��R)��L:��QB�$�(�a~w�]L�>"�Y[t����z#⻡9�:	�s��g�8�� ��N.�ѵ�%����`�λ�ircC��Q��8p�����k��fÓ`#�;��IIJ�]ٵ6��@�2��1�"�:%1�r
^�Qڞ�tras�`ױG/_oyef�n�/|�8j��nl`.^m_�x\R� Nc$Ǩ̾u�I ��fdD�b�#�'���ˉ�"VD�-!�*|�@Ձ�qS�����m=�-"�wF%0�z����$8�1`�}㕂�T�{���X�H[p���Wгx)*���p����S
�ȸc;��@��B��ulͤ �+G�!%���~����g��8B��\��۷�J�T�b�­"�a���S�q������J�*s=w0�3���$`X��b	}�RR�����=,��1�U�	�1Z=]��@��i>�g�m�v�^�
��@N�j�r�A����!�#��bFEFj���ْ��Hv����~�b�s�8�v�ĬC3��C���?��b�4TeQi]`b�<���B�L p��(��9l���"uw�{�.Q�QԚ6?�]�A��}e����>�{�
���e&���@����x0�V`"&�]�]������������6�]M휴��p>���د��/:�B�YҘ��O����@�lʂ�A���F�?^�$ȕ�i�
HR[���u� ���.��UE�
�ج-��Hl��o��Cc�st.���:����5{������Ql!���W�,�r���q9_��_��?�Wo����Ç���l�R>j�x{g��2�������>	���_/�~�e�J�/�B��Ձ��
�S�v���j2^��v�FS�?���`�k3��N��#�f�_���I�%c��ɩ�>1�dSjӨܟ�\ s�#��f�Y_|.LS��ی�����az~F�@��T3Hui?��%���}���f,��5���A�1�}�%UH�_D�@4�ΥB�U��̥���,��?׎�u#�S/fR2΅3��]��gD���&"r'�Jx�����<�F�D�]���5F�62�p��%`�V졍��p���>x{}��Բ3��s�G~W�3��{#uKi��<�*/u�i0XpX3�n�2��u裍�dq2ײ�(����T�qr��"MB��o�5��x&\L]A��V�1C�YC����P�E!��*N��@���{soW���d�H�b ���N�X�RsH �X���wF�,<@�=��w��D]��+Y��L�'�w6�$�>l�s���j8�8iVxfb/�g},��%?�8w�b��/�4Y�Fݝ��)��v�-ߖJ 2!�p�=P/>�A�W��9�(4�Ci<8(f<l��߷�L\q���b?�4-�.�0�s��N|~�iƬÞ�q�渗H׭��uв��{������x�S{���[.8XGUt{�eL�9#a��J��@Q�dbA��Q;��� �L��HE����y&ĩ�&KD{��Y��Vx�QP�"��$tp`|�+����L�L���l���>�4첃��2|~�4|��:L6Uؽ����ʮ	R@[[�Ɍ�c\-�z�<|U�R��D�2�KT�h�r�hs#�?��%���x�h���Z�(ꨔDT����B�6�8�K�, ���6�W>�����?s�#�u���AK�:�Qs�X��d���׷6x������DޥS+2�1\
��ѳ������PQ��_���'��|/�z��2��9�BeȌ@9w{��LY�Jz�]��>��5��@�q)����M���ڬ�����E�c�e���m15C�3���49�H�x�ޮ+s4
Zh1�)@f>�'�]X`��_e�xeY���p�P������cA�2�mfYv���)bԓS&c�d�m}�NR����m"�H�HR�������h�7�U��N���c���C����ٱNi�	��aW�B����1a���,r �NdE�����4���3�T{0 �g��v" ��&:���(VbZ�i��d	h1:z����7�_�+�僰+,#��x�0O��FiڞÎ�#�b�.��e zK���P������5�����Z\
j�Sk����Õ��C�֪hĳqҹ��6����̟^?Q�㥝�����Wsl�>�ʬ�F�e�\�r�Ѳu�p?�Ȱ�Ё%��� ��v���Jѳ�@r�ʠ��=�2~�ڲ��D�"Ek����n�H��@(�L�Xu�c��FH�Z����)dՉ��w��f#��_���7>y���A��dx��`�J�Ҳi^D>�B��:T�zTWϥ(X�M��4@p��˴����g�f�]E��3׎�0�O�@:�{mص���+#�C}����r�7�c���ܠ�q���J��E9�;b`���Y`���?p]�X��e�\p���/�4b32�<��l<Մ��v�m�q�6�T�[����
&�Hv�>�||�qa��/ӧ���܂��%��+x�eo�V���7�/����M��������&h���̂���R�����(��Gg�,�W� �R�Um#֫u 4kȽ"X[��v�"�=�b��+<q:���@�*��t��6�EN*�"9�@ڼgvg��n{�;���/�p�ك��*�0�9��r��=��V[���`����-�'33V��ӏ�����g*�=,V�=�[����/%o����ߘa��ŕ2x�
451v���7�ݯ��7��A��;@vH�{��:��~wz�3�0F�)/(!*ww��z9G��e����Vv�`٨A��=2v=�|b�J���8H5��
�
�FS�-�}#C�]O�L��u;�/�,V�ۍ%(�,ؚ8G�9���.����w��*�BCZ�,�I\��3YD�gnup��ϯ�{�d�&R���%���KO`7z�HlC�7��*\��#j�8�(6��g�,p�P nr/���r|�Og�R�#P�F��x���[�� �x9�^qp�mS($�*�DeZ/�%�^P�s�"x�e�w\/d�ƀmQ?�F����b��K� �7�nWo8's���[�D��2X��Q�L�{F�+���RX ��Pq��Sa�|1�R�7?�?z�����
����<D)�u�$E����>h_��*}"@#�bj�J�����g��G�;���jW�'Ȃz�G��R~��������jE�r"��?��{p�-q�|��Jk�%����7�.�on�܄z�nX�h4���;����l�đY���W���Ug������q��Y'���ٗ��Q��\�'���w�	�a�ͼR1&�9F���`��w�l]Z�惮����Y�"�d�p$呛	̕=oΗƇ	����4�����jCm�k�m�FSWނf�q�T9|�y�6����I@�U��tF�>�sx���W�w*�ך�:��ZT}KΞՁ}�ǳ�ep6���sb��f�����β�8fO�a<�M�\�p�ifs<�8jX��)��*���N�V$Y�b`�-mk$"�|Ĩ�
J[�$���a�+_"�"lL?2,��Lef�M:����[}����4��̨<�2�[!e���l�� ޒI"���}�'�|bA��Y^��+�D���ǟ���@0O�gacƋ>& ���=��ؐ�M?�̨olS����m~ۜ��2ܼy'��~.-�}B�	��_d�J�]�i�0v�5@�TL
�=�F�������&�� h�㦜��=��o��uj����ۛ�!�DƵ���U蠋-8x�GB��9�Y=A��� O N�1�1қ�*DϞ�ՌXNF��̓��)3e������u�%�SՈ��9�1�7e+�r`Z���E`h��+��CP����_E�+��#}辀�Qk�v��BS(����sAU�$j�#�	��Nw&��6{����'��֥t����F�ђqe�iS� =�04�W!>��L�8��Mu����"F�xծy�]�!���p}T.�6 c.��RJ��V�2gw�����b��=.c�lNVɈ�F����X�JYv��,���d�nv�*�N�1*^=�GS��UW2."��t+v��D�������1K�l�3`J�L��so#琞�}�)>�2�6ȁD�Zb���x�V�G[���:X7
��=��L֥VI���h��r��}�M�'wd���$ ��9[�
7�#�2��%+�k�qV��[d��#ey���' +��V�2�n���u�*�A�����:j��_�݆�Yi[����4/�I�Ӆ�B��I��%��ͨ�Lk�kײ���[�zz�G����tQ���2�9w������l7���f¨ �����Qq&��g�gZӮ[mÛ�;WC�ގ���^nv���<?�۫]��w��-�ep��|�6��'.;c��yLQ|p{/��W�f|��S	8����
�}�_��,u�H�Ļg�5�P;?�I�?Wx���:�u��r��~�`k%R��rn���b[N�k4�w���^��PQ_n���9A��e.�۬K�P��Gl؃o�=m�9
��K3�_]��z���*����>��a8;��w�-ؙ?܄��W�(#�b�����;q��r�da�1WY���Dˈv�Zb/ur5F��X�D=�À<�YoT6��{���wc��z�q9tU#*�X��ai;4O:���D F�3�ʕNI.����1G�΅���G��<�
�X!�3g��#�?m���H��*=H���h����RN�T-i�A�XC�ϐ���_�\�)c��>�C�ES�I��d��6�/�tFV��{�4�u$�J�p�^j])s��tl���q�p8��!l (�)S؃�1/ �{qʈ�<8���2q��aJ&���C�����`�5mO�X����;�Y�@q@|T���8�G���tv�T͂��֥9Z'�Ҥ��yb�n���X�{�ȳn[�&�
�G��\_������;m��qb���snN"5ISŪE�Dk[����:P�̒��=��@
�
���L8�W�n���Ǌ�k�u#\I�fDM��c��qӤ/���4�߸��pCg�%�u��\m'�97�ZF�����W�Q��|���k�~�4FK�EKO<H�3��"��>M�����ғݠ�"Ҵǖiy�f[1UW��?���ZU
�_�wbiVCT@����&�E�՗ps��6��l��#�u�4aOh,��*$�dV����4���h8���j���[Ȅ�0N���WkN#pF�����l�\2 �7�Ӱ�7����| p��Z��i��EC�`(��ғ6[G��_����F_��9���AĠ�!i�NCOq�&*�;v���!p�R0���5�q鳩��N��x��D�l��02���@ޭ���H�)��`?48�٨
��׷6x�U�Oe��P�{�Il�� �k��!ƣh$sV�=�9�������
L�a�p'C��6��
}X��_���2�d�}�_�����í"����e>S�DW�a�j���ڎ�0�U��0���籸F��"��/���	�rYX� �������U���\�_��s�4W�ޏ���~����A��AS��]�"1a��`�pZ�"QR+yt̅șx%�h�gI�@>X �k�^E"53�}�r�~]����01��D|��
��J~ץj���a�T&�j)êz�JhGx�'�j"�W�����R�J%�V{�}���x4�t�s���>�s�o����'U1��H�T�	9 ;�NF�o�z69�A���N��̠��c������^���<w��	�S�s�L�Xr�ڟ��>����}�k��˕pE�x�<�q���ց`6��;	�(�#���뛄��Q	����.��[և�����"�� p4�t���[=O�@g�����R�CǑ�\��js�F�ܶ������E��s���	b����#i �/�Ǣ�ƻ��.z
��l�&��/��D�^��s���"���kY�Go�����7Y�&>Q:lw�\�m�T��7�LU���rˁ�o�<�t+�E�Wދ \AO�w��q}2�f;��	t#Ac��}̚6#|H����12C�6'�ai߻���`�݃M�m�]>� b(�^���qLM��؂l�lt./fbD�07��?��,\�z|�������a~�.	��J�§"P��kغ��E ]�ֲ�&mRr�
�v��C������h�\��;w�w%�J�r��D�Wr<������.�ۓh�Ե
����齩�Rq:;s_�]7��~}k�����zM^
��@>�$}P�b�'d���_�!���_��]D�C>����<E��v��/�׫77�Vk-ױ9;e�T,(��(x67�pa�����lɦ(��΄�M����l�����?p.���Q��uK�Bu�>��|>zra�?��xvq..D?��G���*Ƈ떨dD�s 0~���l�7�{q�(c�`5Yd��I�h�>5�"'H��"��,Vtxp����s��[H���Ft���,��0��`�6c����t`����:�VZe>�A_m֚�J%l%k"���RH�P����������4i�H�q���g�!X`�~�]�Q�ǥ81��>��O�8pNr����W���M
��8m�L�ly��4-��# B�]:3��&��̷o��s�?�L#�E�����-4U jϋ��P]������ {=��������X�}���?DV�{c��`�9i2%��,��p��k���@Q ;���"��ђx���ޓ l<�tNpҾD&���	nS"�$aE~b�E�uM��o�Z;b������Z	bV�I�����\�)H^���jɝ�1	�&%sޏϻ������"�G&��z?��`J?���)�+�>���$ð��U�$\H�H�o�ud�&2J*��H�8�8׺��,;�*O^�e���L�������g��'LǨ�ޛ��T�9�=�;����'I���l{-�2{�۷�ĳY$�8�g�b�>��^�O5����'W"ţ���$��Ƞ��y��W�T���w�
���ې�Wa���^	��G�q.&�޷/o�l>�����l�^��$������5�L�WG�Fe���,k��Z`.g"ED+�<��s]5:�*L9�=�>ڞ�{?��
���A#���@���w��-^���jGoD��\̆�t��>k�&�90��f�[i�lCeY��b2�&�9�8ڡ�A�H��K'������>��z��m��~&[s4K=�	�`"�ت��5�M��d���!��9�B���2�P�6b
$9Ш�ʊT/�;��/C�ٳ��2�J�%"*{\���{�ɀj$x�C:Z����PA�UF���$v�m�ƌ.D�+�tA�J��^����d��BĶ�yu�=�6M��IL���u�>98�7�:-�;%��ᮢHY�4�b)��PHz+ ;���$��\0	�xGb.��]�gϖ�i끁��s|�u�p6�R1-�R��=���y����R�`��D�������ŏ\��_��H?�CU�I��r�-�G�ɇʟ��#x����.���{�?휇��Gly�p�#踓.�e�(����C�*t�±�1������n�M����K��2��l��uG"W�>!�a�7��W�B~��a�T�v$�� lf�M��};p�4�&!ɬ�RzA�1P�ECg>�ҙ+��k�Q� ��'�L�L�^���l�~�"~��};��5m���-�=�~��W�z�!�1* x��Z�R��1�E�Nc�w� �/!gr��5��'�n=_�*��;IP��-Jٶ.<���8\M���a�`+x?F�	*.ϼ���W7�,�'��cr fj{9��:�E�-�uQ-c�.����S�w��i�Җ��.T5�c����i���:�Ց��f�֑ ��mmہ! ;��"`���ed{��y1�ߝ����o�۷��̮���<3��C�(9�wc�.��r!T:�I�$�!���0p��J�5ad��Ŋ�OAH/\��!�f�`�4Nk�i��	���K�2v�S���_T�iGo��}}{��m��D&2�:�T`��[��Raݷ�Dxď�U����<����=Ԧ�	eC��
C<g�_� O�ϵ8�j8*�.F�'m#SB���1�"۟��f@��F\� Ft�k,�(�xD�mN���a%F ��?�4�߿�L?١�[f`n'i(��#y��ќ��b�C'j�DkZL&P�d�x틝�.�V#����T��/���Z`�zw�L��(�ҒA� �w���\t�"�AKB����8(��&Y��Yv8��HBk��$)/�oc�g&n=e�$H�Ϟ�~�T+�:q� �T�ȶi\�y�]�U�`	�O���G�� �"\kdH���l��c����Μ���>�#�,R_1U%�ib*&"#�jm��`�0�M������#��i|��+caU�����
����ւ��ٳ�ULs�)kE�����]{bӂQ�R'i�9h:��r{�-��c��HYzFp��mcu���ȕ�5Gg�๒('`���0�wӃT�&��>#�Z�T`�:��g��ѩ#�Z���7�ڋ󰟭i��`��b6(= ��a��ٜ����vc"'�AmN}�[&Ȁ�8k*���iܺ�8~���J�'�E�I,R�h�{۝g�v�LP�^RۈV�0$��Z���Dg��\_g^I?C5e��s�ބ3d0f
�w�ȶ+}'[{K~T��硱q����<�}b���xh�9��u]j}0ξ�Ib�3��0N/��Kf���0c�o{fL���8v�E%����X��a�ò3��5m�^,�l� ���1���ĝ�:C7��g:Ǖ���>�l�}<9� �c���ً%G��z�^t��$S��gH8ܓ	l,	I�$! ����1ޟ~M�?��ij�2�0�u9�<��	����Qy�Bbz��L*��s�z������]'����[��:���<K���Ti@^}�8��1������Y��6��Q ;���!��;��
�j�u"\�mʭ�,��,�X��ˠŃ���)���nD�"�?yc��d�8C�M2�ҳ9�'*!L�e2��������;��р?�
};쌅�0�M�����.��<���v\�n�w7�r&T��˫�NX���4�������:?W�Y�*ە���Z��փ�î�C�VPdZ�}��mN���4��h�Pc�]�.bN�H���5�!���D���^�#��_��1�v}dzL�`�Bya<Șɔ��ٵ����\��ޗ2��p�0.TPD��������.Hr)<N�7��T�`h���1~�G��|n�4]�[�K���33zggo&��c��΂e۵�DNh7��	��}\�	�ί.;�z�r�_m�D���֢>;���]����%��H>��N�٢�b+nV��T(�g�����lyl�j�gN�5����!=ʞ'�}���v���a�?�Z�$�Hu�`��[��� �Ǥ2~u޵.	���\�� ǃ����	t�K����x�"x4�v
��U1i!���qPp��&{w�:="��y����چ�����p%�\��cs�B!j� ��fіY-V �]3��%��G�^l�7Ջ���i�5�	��t}�7�X�}�U��I�j���̱:L]�0͇}=�6WxTet�K��}ZqA0�ۨzFE�
L�$��x�Ir8��9��e�8��������[��o�25�����SxófO�TB�zM�/�?�R�E�ŽdU�5}��KƯ�F�A$:������JqSG��*��WH�Ҧb���|nh��@��	#��j��u�l\g��[KS*��7j%�r^���C'�/&.	\��Ȏ�Z�����AA|��x��;��V/u+U��`��'�3�í�唹|����q��}y�\�p��2	��!��n�����z{���}��NKm�U㊌L�=S���3�9F40
�1�L$��������љC{�ZY��ھ�q\6n%�8�P�yXB�� �)r$0
Q�G��<��s�U��uEl���an��ˇe�o��#�m�H�&fNs�G��=7��֚���~cf}o��arc�΃�]�%���?U6�"H���(�OH����@�3�J�݃@��(JU���A�[@�r������~���E�wr2��n#�B�]��7�aMy��:-����b�O�y��Mk��:��>pk�
��� p�h�8�#^�7�t��G>��=	�)�b�
�K��:�(3��
Gf_[�/5��-�/X�Lm����!<��t-	�ɢuD���2s#���;����޴���P��[�5��xЈ9���!#��zq��2p�.�6��R����Z�`>"nI�e�������de9��C$
��$���*M�񬪾�%:~0eu��j�P�����3�q�J<l�~� ����[g�y�c@.�ρ4��:	���P]��d�5��@w��a�We� G̍%H$4p{;���sa[�Ϯ�"�M�Ԋ�:?9h��BI5c��M���h"\K⬻W�O�C ��G��]5p|/�L���+�r̅k81��A�I��U�F�����5���0Q���~�\uA4ρ	-����/�a�T�W��#��M{`e��K�#�@^F�	`�a���Y�W�yѮ�t ���T5)b��py��X)�*�x�k���Β^�G�¶x����3�eAA\ĵ�xB�~�]��:>'V1�.U�1�M�.���e���n���8�D���2]5�b-N���A�U;�U^����\�<��ew�S�i"��:�ۡ!GN�ڤ�ȉ��� �J�C2<�ھ���)d��=D�1(ޣ�U,s�*�YGݡ�h���6l���DL��8e�����
ky��шK��5⑑F��M�4V+˲x˂ �Iwh���
��Wz=���Q�f\����� �1�Ʊ�#�������t@�bR��svH2KFf+&F �"C����@\�ԗ���&��� F���<:S�9
�Y׍�I�-
�����}��s,T�W����$����j-6Ue��/��z�GgI��gP�bD�pt��E>.Z�� ؃ ˲=���p8k��T��0iD<�3�����#�6&��
�#�Q�>���U�8t.��{�-Яy$=�=O�(5A6�@U+ ����H7N[� Q�,d�C�D��<M�`��,��?C�.�4�����[��p�Q۬��y�O%��6
�M��Ζ�F1�܃a�!kf�"`���(�Bɝ�~P�0+*�2�s#�CPs�a��r���>�;8��Wb�Ȏs��T3 ����F�Y��[J���M��7K�6�h���Ld��S�S�Fge���
#�,%b�F|�X7�(���Ȍ��k?�d|~.[�4w���9�N�v
�w��ΔF��/�\;��u|��ZN���>	�L��I��������Fx6��o����zY:p�����b��`=pM��*�P0�]X@F%nj��.�U��"�<�:A]hD2��Pkevr�^x۫�ek��M�?�m�ad�@������SU���9�>�XD�T���ek=u!�"�J-ʁ̛{P�^��;��D����&��[�f��ӡ��t�o�X�Z��~����������W�ە�7�����Y����T�h����G���r���&�I��Qx�yţj02�g/J��f�lT�^�c�BrT��$�%�]�(� �#J0����"J?k�/#k��zt��ܣl��c@�M�h,�J�e�{T9ާ0ʦ��	���SD	��'��D�@��h�hH9>�er�PG	��g��I�۞}_���V��.��向����au)w_O�<���g�3�la4=�R��mPu������Z��g
e�o:�Ca��L d4��|�v�j��<N@d��-Ɓ A�X�W�O����.\/d^ +s���B�d�o��M�C��/Nc�Se��� �����0ս,�4*bH���W��F��ZU>�IG���86n� �RIJ#���!j'�q�8��%9�p�&��F?ׯ|b���&k�)�6>s�c`$"�Gsp�kMc��ٹ�0A,<7�H��z������6��D0��0
n�C`�4��w�P[��/��M@�01��U^i��ʥ&����pl"n�΃�W9_�牕^'��k4�H�^�y�6��6pkW륂�	�T#��jgӨ����iQ���̻����vh�sT������
�Wd����Z�1D�����/Y�,ˮ:�m����"�E�Y����j�a��_�O`VU?�`L���	_�L$d`�dT)��h^��m�9����"�dL�ȼG��2��_��4��k%FF�Ћ�T��*�p��X���.�W� �濘Q}a���\��H�coy�,A��ѰI#��=F3;=�
�B�2.�~�2�+Otmn;�N��`)h��SP5�q����'U�7�������BR�0��C��Vh�D�Έ�{5�
SS�Zs������p�d���<�G vzv�j1���{�?t��| �%�~�� 6bo��{����=�xisv�bŎ�?#-|��v3��I�U���NQC��`���;��,	'v���c�PkT6WDA����Z�K�@���N��&c� �C+f�"¢{��d��`����d�h5���-��(�b�@�C�,TV��(��S,Z���=Q�FA�id�
���N����C��:`�eMƤm���G�$�	؅�W���LT_�����d1̨������N
������,8��� 4s�~�I�FM3���a�D�d@>(XDP���0�Xڍ�@Җ�&w ��C��k��ز��E�n@��T
I��Q��2%��`��N�So��*@>C�Z�z��9�?(�* �L���=}0�b0ŕi�'���3V�l�j:Cך�d�
ˑ��K��=�ݵu[I!�2vV���=�S��d�RQ�n�5�TS��
cc���=b��T�!9����jr�־%y���Q�<i�$�C<�4�0�DHE�,G�h��9M�Ep0wZ��)�&UPtr&�����:�A�Dy�0,G-���;Mu lb�V�Ӿ��D�3"��	33 ܤ$��ԩb�2�FwAH43lќ��E��+���A/�F�{X�3�r�^��gdW�ÕvԔ
,��GmI���}a�!AY��F��m������f�)D��je�s���r��+d
tp�	uT�[���Ȯ�D~��g�%x#(Q�k�p�@�:v��pB�b��6q�� 5%�G  ������<!���da��#��&���b��	��A#*f�oS,:�N��c."��c��%dO��]���'�����N)T�"/��޲,Iġ����v���KhVH(x��f0-`�����]7pX�hS�\��O�d��3�T�́�lTn�S��@j�����F�]��4<���O�3��HtҤ�	|k$ωNݫ �2l;��ds�| �I���癬v�D���p³��\� ������6�4���&'�L@����}9t��aB�F�C��0��G��E�evZ��I��cN1�5L�0��-��w�x����l!\���*@�
�!+Nz�C�7���S�]H,�EQ�T�j���	:!Z�2��� ��}���1�Hk2�C��
D���X0�FQ��bU���V�j������b�)��V]�@gp���P,C�A����!+��VY���*,��Q2Fs��)��ϙ��k��p�c�2��E$#s<��0E����1��fvq8���s-S��F6���kAhA���F5kJ%<!���)��	�#'*-(Y���B��D�rD����K�(�M	�B�9�I�We�Ț-�<�����,�l��X���ia*���;S;n�(Pj���R�Zё��pQ���&M�1WO�Y8����?��쑒@�ZT ��xH�)mE�i8^A�v�h�l@���
]��w��V�9�7�H��=4z���5s��a���8�U�ĩ�"C�v�j���)%6S�p*0G:���T߅1��3�]d'"j���'mUF�šP�N���Q	'��pG��Z�T!���=����Q��r�z��i5���`FM����8�(	��#��ir
��q��0�5:괂�G�����j������#dO2An�FUIwa���<K��wv��O�6ڷ���ާQH���Kɞ*I�P!�ǣ�DdBETt�ܰ^��$�R���h�@��Ъx5�����c�ԑ�!��V�9Z�T�|.�^����z�437��g�B��wddN<ظc�a5�8G`�� �Kx�P��J<�Sf�m�L2�4=k5�siߤ*F$,#�9>to���i (���[<��#b=�Z��Lo��a�5h�J��S���]d߀�-�2n��S5��0`,�=j�^�@f�fRcΑ;I�D�-����C½� ؕ¶�L��YD7zF�A-Ҧ0y�15�~�N�{j�gG;2��BU�ӱ5�U�Ga�T���%lx���0���%���&��Ć
K�hdR�g��E5R���Y�c2��,`�y��7���1X��y[��3���7��5c�#饅W�(�)�XKV���5Q��"��� j�pfFb��
e�:1��i���K��� O��F��L���i(���C��(�i��r���[(�o��SeVi �Xy>�sJ�An'$��n�4��}cʭ�4��NOќ��0�`h���3*�!�~X����;�Z��g���,�hc�ۘx8���0wx�Q�S�h�S�b�l/�Nt	������-J4���G΋%F7�^3��������h�/��IA��A��i9Hԁ)��(�OpŌ���O����D%�9C�=��Zm��&�Pu�8��i	�r�t�T ]�6f�߉�D���W�/��Lu�u�00���	�L���y��~$��֠X�;����֏������a�y�ĖF�'S��d:���CE�w@H.�:�ed]D��]�#F8�9���xo����q#�v�
Wx�$Z��I/����ܛ�+"�0��OZ<�M�b@O<�=�	[�Z;C+ Lm��8���.(Ӕxg-�H4N�D3�3IM!8���z��k!fNr�2-�� �i(���S�ª�Ū<D�Yh�	{[0U>����Aò(f��˝�lн����L�G��P�O�|q���b
�f�d԰�!�Y%*oKA7{;,� �QtT����Q,2��+G�o��u�� u����܉�ga�v�����6�9q͜�H�ҌZX��W�#R;+�b�jYr�m��B��-p�Ѷ�3�x��ax!�}�x�,���u9c�9
���) �IY�Iy�R���^��ű�n���{`�!�����r�H���>b�،Me����4�\S4wߩ燵�,R���Bma���D�O1��� ���w<<(R���=i�(<��˘'�t����d_��$�[��cf�;�� ;�Y�~�	E�w�k�``�9
���Nͬ$�w�R0*[��D��Z��H�"�ZD��I�RK4����|q��*s�:��v�h�
j��\�e��.�����'�|l:ٷ�o�1mS����	��a�3����F/"ʹKl�Ҭ
*8c�Z-8�a �gL6jf�<�"l�d�uC��E�{7�#�Q�&a�2�J�XSDDe��C�h.��r���5*Q�ut� 2��5�{�.�ɯ��m�(�H����'B�.
�q��%�0����<�6�뭬�H	�͈Ļ�(�[��e)ה��'g��F���H�V' R�� 00�J7�6-�L�3����0:s�����+#�(�/��=���'c��34Sǵ���j�$��6�)�v��|gGq��X�_��D�����QeŚS�&�ȳ�{ Gʺ&[.B����y}��'t*:9$llx�kE�- S�v�P�f
|��&Gň��Π��uy�P��l�$��#�'f�O;���A�=�o��ᄴۧ��^=d<c'�$��˅���C���pI��	�2��¦�����L&��gN����<���x�%��)70�������
u"�����il��-�H����lh��^�ptx�*��Cp���r�z繝����K���44]\^��]�n���x8��""(
�}��Ѥ-��o.2���"�NzB�F�N��A������ {tu�.'{k�ycn�LU�3��bn�͝`gL�^1j��i":����9L��Q�A�gC�v�/��s���\yRJ!��|Ƙ@��y�m)����Jq�i$x�<&�i�z�N��OT��.��� F�uіg�#��4����L[0BdY��O��O�ٹkg�ڋLݔ�%��E\�ÎH��<�xD�x|v{g����#�|�9u� wV*.P,�Nj��l��j<~������qov�DC��KmVӣ�K������
?��umHH��I���?2������0_��ڼF�W���lM���FƤ�ɘ���W�����m�߈��ʖ�����#U�GQ4{���Lй�u���}45��`t�o�ZP���n/_&2Q��䇌NǍ)��}Y��P����k�9�ȡ�{g�"�����"�N�DYACs[�,��6~Ce��m���K���W���=1������M4�^� �'���1�i�y,D�]CI04�符�'F�5�;����	@�9���A��,Y�ݯ)�uS���%�5Rt�:�w5c!�
%��ږ8C��:;'���O�x4nZ����Ţ���G��2T~v�&��V�cN�J��^a�e�5�9�~dή.͹L i�o2�}�����٠��TA�ͳ�%(��Z6��'���ϟ��2��(G@��DQM��g�RRhxx�
'��[�
��\���n�do��3�V:�v��:�ő$k�hQi4�?��̅�3;�o�ɝM��1CU��<�����<42�,t#( g�?xA!��_���Ͳ�m�|���=#L��M  �d^Z����9<=C����C��JF_����ڀ�A�;�����͕�I���ro�oߨ睿c��CV��K�qj؊���J���`�IV�y�Q����I�{Z�n�믿��ty}m�W���79�ʹ������(>�N[���֩
Բ	TPE!�s�\�smL���T�����R��\�HZ�s(}�c �@��3���25�F���5oݷ�Ntv)@��ĽC��L��px��#/�� c �[o�T00[^�:��]cC���@���Zqp �4���uc������}�駟2:��g����+K3�.0z�C7�L9�43:�s�3�@��c����L���8��8Ph��3�j��pQZ�����E�d5-�����G�]����`�����U۱8
N�������r���Y��τ=��[ej�Ȇ��-S��R�>+*E�u%ۥ1�d]�-Ӎ^����xm"Ct��?@!�?���A��ye��9��:�dv�|R�"�M��qb�GA�(�}|�b�}�5�-�Td�s1�0���77oO@�L���**�d��F��czI�w+{�������ݙ��� �z�}�����G1C7��?�:"]N_�̅ds�քE5�aj^�s�v2�X)�V?���-Wz��V�k��F�Ǥ�f����3S^]'I&Q޺zS��/̋-Č����������_�l�7�Ӌ��;�lk�eS�J�ean.b�a8�eq՘��cs��h��N�$5��+i٠8����,���1��3�,��y���������{�].�F7���N(����!H73tz�b��&+�l`���A���N̵!wv�N�T|�1��ιo�6��&i�����s���u(�R��"���O_<7��h���i�ޜ��h?}P09�dg'fa8�^8��󹕑�g����I*��e�d���ǽ(�3�i(�����G������5�����˅Ό(�[�ym+�3�p�{�/��}��&��Ix���g����ݙG��+�;�\s�~�ܬe^���ɳ��b� `Z�sʇ�"cF�-,cae��	���t_��`x�s�k]�}�"�Ȳ���r1����E�'�ms%f�eާ�QL�cO��z�5���1'�K�� y"�.o������Gb�8�چY�m�&*���@aÐ;�2r�ܑ"�=�D���T�(��AT���c��\�_<5��*/fP���@�:���.��Uz��l���$`NϷ4ư�i�9@�E�ye�	E�rod�n���=�|��_H��~��O>6��%ѓ��,ɵ�˕Y]�1�B�1/���S Edw��Ù����>}�TU��T|�}�{'P���� �g3����D��Ĕ���Ȗ.�ŏ��:�Լ��Ks!���x������8�>�ي�!�d>�׈p� ����`��>�`�Z��E��~��파��id����3"I4m��v�wf��Gfsuͺ*D~�y�P8�n,Հ|�=sރ��:Ǵ�\��T�sG#�;03&��A���X��7G�\F���0�}�ټN0.g>8�҈��.�
d���Ρh��\U�y]�����zyo������_�ÿ��b��g�C���i��v
Oc���zU��B}�B���l�c]�kd�|�A�o괺ئ��J"��"l�~��yF%1
�E��g�3O�U�:�'"�//AϊR��bT��Y�ع�����<@`�b�"H�D��Gz�ιT�UhJ��	_W�e�#�$B2��@�Lb7�܉$���.��� �m��đ���|����5^�,,�o��yu��gv_����+�HC��a�OQ�"14�x���3c]X-�e#ޏ�U%.�ʎH!���u���q��@_����J���æ������5�n����>�N aW�׋�y
���*�@T6��{�	�USYQxb�V���.)^�c]�$�m�VFJ!`+�ىX�d�_�?�#B5�"�Xy�t#
<���)L���[Ղ	JFs�ٺJ�%k����KHo���"
7�C*�߽FD�j�N9�������,�/�`]��E��hF��L'��Ltr�8�4wAT�{X�9�ԅB�j�?h9*��#��+ӯ
7ʅ�X�pވ�yf���`��#Y��y�P���΄��6��\�f/�<�u��#x6h��Oĉ���x<dޚ�y����R^�~��"F�;@)���۵�O��s�7U<��C�w'����9�I2�Z%6+�\3Ğ@�QS�-����������uS4U�����1^��Qx�
\k���9,2�CS��g߭��m/�
w~��G($٘Ë��4�������/�l�(�1<����D��q7���b/ǳ/7�ٗq�\��m�4�F�~5��+mڣ<�D\[ޫ%�%�͈�[W����4y�[iBq!�����ZN���p�9��c=�׏CU�Al�1���$����y^b
u2?N�<䱽�[�31�|j��ضc�C��G�ytiK�)��qP(�zUr���- � �8~��/�M���f��rMUX@E���Ű�Y��}�Z�Nq�XV�8��b����'9�2�WgG�ƭS���A���4���9��"3S\�J���E�SW��a���Y�эP�P�6�o�+��ÿ]���c��������W0W��/�ǯ�G������c��k?:����b]>�s�lY�٠��8����)�.s]O�lQ�[����8_�����Љ�S�b���`�#�áM;s�FI|P(YH�a�"	,q&N�ė@_Bt( ;c�x
�"�X�%�M�Cs�l'8֊z���j� n�b��=�C+��;�c/���w���ڱ�k�h�d��㞼�Bθ��ç��I�_�<�BŋDde�0v,e�R�Ll^o�~ 0G:�l���x����m�S9m�Um�$?��aa<A!�H�J��{�NKxQ�1MV�Y��y�)�G��{����FT��n�����[{w�jY���˰Yo����l�Z�*�\�{<����;C6 ʪ�0�)��f+N�\~�q�#D����{��&'�#�����c0��W��77�Ư�Z��ۡ�b�d;�A.�̋���eN�,k^Kt�R��V�ɶQ�oVU�֫�Ⱦ���?apY�}7����OS,]��X��Ȗ�Iny'{y���6V��J�=�=�8��Sa���d�č�ݓ��Dp �e/L��Q6 �HL([YD�/|�������}Y�U�W!C��e�M��#��������*���mW��(sts+���?E��4��/G�ɋ>i3��l�C��<�F���|�l�R�-��`}{pm���b�O�=��2��Y�b�N]r�=��rv����b܀��ь�l�)��7���ށI#O���]�L@�V&kG�(Q���Ţ��M"`�$��,�H�8�A����_/�芻����c���eG�]}���g�"�@�
��eovb�tN�V<$�&ș�	$w��&�v?tź,<0]@Us#�����'>���ĐN�x�r@���`�� ���}M]8{f'���b��Q�������F��SY��AdD͓�c�]��vj1���4�Ţ<���!&'�!S/�k��m���*��W�n%{�8v�'�����ںj�.+K��*,B9l�]����w�s�j'+/.��_����z��R^�La�̪�7�����t9��5�"k]�V��]���|�ZɆߊUޠ�Z�:�ч%��\�����S�ߤ�.�"�b<OQ���D�2�����x]x^�(���g'~I���cUw�����O�b��w��?�qo~ �6^�����Fx#����ٿ�����Owӱ
�{d��Jvc-"ȥ�g��x!��}ph�l�T�翪���mVӐ����(w9bq� :P\M�^S��A���*D���������e�����Nk'v�(CQ���~qQ�J<թzhia�O4z��=�z�ТZ�0��B%�[Sz��A�=	]��m��+��S KZ�'���䚍y��<U]G���	�GwB;ȿw�U�&�Y��g�`�J<�^�r���S5�3>��;ɍ���V���kV�]�A%J��4��b<���ӽ��^@�j�z�d�r[�6ދ��WV\?eR�܊�]���]�^�h�$c��w�c)�#f,R_�	'u zU�5ӥ����ʧ�z�0�Mc�)���؍{1$�6��.N��f-��Z16䧵�p�ks�yI,�J��o���и��y�ߊ���x��qhl1:z�v�X��Y���U��s�A������QG!��0 u��+q�z��E��<^>7`?9�ފ��q���o1���2c�&w�"�)~�㞯��싃���KƔ_⅗�i�]������C�����)�{���F?���o��m�4�:�t�����;�~�+�/唤���:n��+(qC�%�2��k�*��w���N���X�AL����4�u�����o�K/��lo����E?ڕ��;��%/��`�U��"�n'�J1L�g���|]�ym��K��+�|�R�!<���?�������|�7��C��)��(��=X��?[�o��X�2��|�~]�y�:s�:�ks�����g�-��n���KJ�=K��������ޣȇ�8��|��~����l�y���~j~�k���ϫ�J��[����N^���/�����F��ƾm'�tbĞ��Aw��\��ܦ�Yz�F%��7��k��¦]wn�x'����Mj͓�x�:N�T4/�~��zu�����L�|������3�Aܭ���3��$�!�}����z��7I��%���y�?�����im���X�7�w{�?,���,T�jo�~��[�[(i�G�RY�b-r~%���"J"�|�b�8�jX�/�vUZ�)&]�a��c)�q'�TE&"�= ����b��JS�x`D��Œ���W�{�V���[��_�G������~�#.��^/��7���D��_�����,+)�_��u�?��D���._䗿����r�_��������fĿ��!m�e�0ƻ����x�;{�A���7�`��;�����o�o�_�5��?���:;]�O�{u�>�k�ݎ����^%�x�������ya������?~e�/#�����]�2~�c���x��;{x������xY�2���e,c߯�/�X�2���e,���e,c�X�2ޫ�/�X�2���e,���e,c�X�2ޫ�/�X�2���e,���e,c�X�2ޫ�/�X�2���e,���e,c�X�2ޫ�/�X�2���e,���e,c�X�2ޫ�/�X�2���e,�� +�����    IEND�B`�PK
     ��Z��_2�I  �I  /   images/5f4f8fc5-f884-4b46-b794-7d87214b037b.png�PNG

   IHDR   d   O   �`�   	pHYs  �  ��+  IfIDATx�Ž��u-����:wO�9g� ��(���"%K�D?Q��l�ߒ�,�K�����DZɲ�h1I�9�ȉ�3�0��=ӹ+�}n5����̷���i8����[������{;���+��8��%$�Y�z�9
{������i�<�4�����ۋc38p4�6��ۥ��[��Q���S���j�Ϸ�{%�u~7�;§�-iԦ��:��� ��?�{��#/����k1��v�;�	V}�n�|�IƋ���4u؉$��$R�M�V��+ch��u�zGu2���!��y�4���w"�?�w��h"�,�5w�6�CD��hjiGi"�x,��ON ��0&����)�s硚G����W�?4�قiE��s�m]��㭥���|ٞr���cz��Y���n�=�͋�����w�Co賣c���������2����~�Z����9G	����3b��y>'�q��w�0-+�놡Y�e�Dߚ�L������o�������'�6Z��4����L���]��ܬ�h������j���� _�����l-jE=-�k�V�c���멶�S��Z��{A*�2��jb��� ���1�/����J69V<Mx%��!	$㉄ܟ�i����U���>{s�q��5���Z��gg�⭾�s�x�JS�g[{�{�Է|)�8��8;���G1�
t/\-F�P�8�ß»��89"�8촁XG?��ezV͍i�u�Dz��?������t�'� �Lq{h���{��	|z��a���8���^�V�]���(��L��
_�t�fi��xY�vnG��0Wݎ��v��F��0���o=@e�z̻l#�y��]v���;����M���!55�HCq~q��g����kEN�K��E1?���qE�H�Y	����c�{���3�4�C��}��� �ݮi����G12��d Ǟ@2��F�ty6b�t��W101�����ih��W,v����ۨ��am!Xi>�� �����"��QI�Y�q� T���uiD�W�?3a6��X��i�N�DĂ�|1���@�Ћh���hP��+#92�9�>�4�0x�0�r	��f�3ǟ3S�����8��?��d,V+hH7"vzM=���?ǡ�_���qD�CG�*��c��W0���^4�!o{	3eؑڅE�fŰ���ij���sA�Ĕ6s�,�F��;��SC|��,6���8vx��]���ڙ��"g�x�$�Ύ`�i����lǃ��^Ƣ=\x~�\ۖ��Q1Z1�.�`t8P�|���8Q��A$ڪ�Q��ˇ��u7ނ`lz� -���}۰�P�Ɂa̎�A�y�r�X��A��?�������$N¼��1%�[�D�RFj�"<11�AF{���`]i�p���0��%�a�߀��v��5�[?z7�������7���o �;B猂��
|���,ᴵ~ac�)L��f�E�� �Y��b��Q� sc���Y����ܹ-pb�K"�#"�m2U����aj���^!��x�y��Y����W� ���a�z=�+���<�$z��o���%�~����eK�f�*��	�y�1̜8��(^A�������=����'pEW;!����)B���𮫮E&�F�RD�{߃{rH�Ms��ǟ|�XK�݄eWm¹��J9�e�tǳ�pnNl��x�j%�EN',n�!㠯7��b5����a��;��ʨ�6��G��U�=��u6m�ͷ\g�ADh��_���o�Q
n�l%��Ӱ�x��	��v\���hlk�]sK8�Cw\F���+fa�5[���x��8w����],X�˶\���4���a�(l��2q�ַ���Gkg+6m�'���>�"t�o�#PV]40�645�1����oiFe�4�^F�o"�46o��\�k֭�S���\���c�K��h��B:��\A�JE�d�턲V��nxfsV-C�lU�QuP��E�G(� �H��-�Ld��;�����Т��/�~I5���ѽt!��*�߂A�`�<�x�4)���2\�XUѓ"��i\�O��M�:'�pV�#�X��-8����l�����Y�7
��l��4��&>y�^�����䩣Ȓ �1�T�N�c�p;�s���������2zV53�Β����>���w3�s�'�ʵ�<�JI9L$j��.&B[��TS6p�'O�aҥ'Z���c����蚷��è� _C����]�`�����L���$��������_t��Y�R�d��f�'`�y�� K��j5d����qx��/�CR����Б��X�%<İ�ҫp*����"r�1�2��cNiC܈��Zb���h(�1�D�1�M��C��N�_M�Q��@�V�3|�Y�K/��g΢%��μ��V`���/�?zQ�jF���l.D��YD*3*R��\�ӎ�����,���ڎLt��}
#G��H�T�H5�����fӇO���tÔ�ݐI����6��{�a~i"�.�)AH�ҕ���&�hm��\��$đ����KA]x.�j�����4�8!L9���J�g"Fj=4t���hf�%�8*dS����3
h�DGav�Qn�J�=}d�0I���<K���ys1~����Aj�:9rEx4��+�DgW/��s���	�}v����W*�����h��Ѻa�DH��!���DgF}�`�3���D��:���@S�&�y
6��/��w�޶p��|�PCOn�	��h}�����1E_�V�PD��Z�	���~0R���\U1m���K|F��a���Ř�䎜|m�(R�کSHRd��lR�X̄�0�r��FQa*���*ɗ��я�,C�Ճh?{v��P	[�>�;{0�z�Ze�j�XB��)k�q���"��VT4��v�
�Z���΅$*������~��2B�8E�z���^�I���Qd���|�b�'3� +P�#^�mlC���8Za>֔��J���(69EWKw����h�k&x��V"�D�X�O��R1�?!�p仺2�N��J^"$f��hm����]>7���n"K�DH�C#	��j�,�um���X~�ep*��tfc+�Rt�5v&C�xK���0���N`eO���EP���̅dt=t�Y���J�%+Prc~Re͋H�>��6�N�4��t���������4����"u1'�/ZBS�:�I��e�k�iX	&��(�I�[�uÑ�Ř<gg
4��aFr����S�9�H�B�,L����	�W�L���|��zU�����uI�y���Nx��-��G��2	����y�t1�X���H��F��z�0jg*�]����r6��gƚ�p��Y�:���byO700��߅C�����GY]��-�8AXn��
ĺ���xI�" K����1�m�YOp���X|�%�j3��1�S�.#�%Uܹ�e�-6]��>J�3��M��kє���ҁ¾"�'���)�9&�,/LC0�Q*��m��]F�@O�!�'��K3�!�bz�nԘp�.h"������"vp/F_���0�!�HH��#11�s��Q�!E��nz�Uj�d�N:")n&�x�Ă�4�Jk�܌��P串-�h�����3�>�_<�n��zl���b:�V6���Rf�p������M�И��v�P�\y�D���l�S4�C+�yX��������FaNw3�{T�v����<��A�W#��ד�)9�W�dR�7!���jjb>!�edƲ�k4���D�)���c?���
3�Oj�l�\��l���$�e�u���| #D��c���x�	,X��?�KV����("�G᢫�	m�=82����{;��><��ǰ-݄��1�)�.Z���4�cg`��O=��{�Ҙ�r.5`q5�hE1[�*Ē�$�dVϟ?�m輯�ײsf׾kW�t�sK<�br�e�:�Ru�`�&�1|�$V��GҤ��YaGF�(���*.�*^|U��|)�ǈ��" ��t*j��\	JF��>c��E�j��s#�x���a�L����Taj@ى������}��fJhan+d��q܏�������c���~����0MB7���L��/}�`%Ȥ%{�^��l�k$�#i���8�FSG{+�ZF�iZZ��/� E&�j�צ(�LΎ̟e��[�z�o6���?s��z��F�+�Z2��"��A+2٧�ˌ�	r�\�b"M�*�gz��p�MU4�N��W�Ph�z�j/��ȟ��*N��Q�2R|N�.��H�Da�Vܰm�J��G(Ni0�b�����]���~�B���r�j�s��Y=�p5��F��	gdT:Q;��AX�Y�66,��g_މ��q\s��sct.NJ2�BŇE������"��e��\jÄ�/�� -j��� �ݕb1�l�br�����k���N���4#"J�!HD���hE�<�d������݂���(�j���.�F��),��bmW���x�����~�Ԅ�f�Yu��{A?Q�A�J=�` �V@<�FoM����^OO&9�կcٮX�v#��7[��̮���71c�07�c����ћ�y1$JE���$��
���,�q���p{k-������jhV���lBǒ��d$:�s".L��YFu�b:�ʣ�f୾~�A,R��@L3bے#<�<�+Z���?��_Z�Ƿ]�.a}�)�A�PD#�G
�1B�4���-m��]��
H�.7��!�����v��k��B��	AXS���BY��&ٙ������@�wа������;�"^��J��s�#L���s����ѡ��hdnz4�Jk��}XHX�;AC����p�wQ�$I��qŇ>�iGkH��Qk�i�)z!��PbA��[�������a^�T�=M[̎�p�$I\G��5���AWjt%�~P��{���a7��Bf��P����)(�p�!�eN;��J�ikM�TLeF�L��v��O�p]r�h@�1$�#��P�HJ"B�i����,^�C(#�gD6͙��'pff�#b��6��A-G�]0	'|�_���A��
a)�hɃԞ���ڮ=���Zs'�D���oP�X��pl6�
�!���Q��4���G����^��]ާQ"$Ӻ�ӽ��<���E�,�[��3���6��8=ӯ%l-XR�:'7��F2��	��^���4�|�7����)x_%x�rh2�*���KM�tٕ�3Wy�E|���r�(F��D40�ښN��.a������2��^_�h*wdQ�^Ņ]�MU��U12�Lۘk.?K-#���9G�tDW��QƱ�"$������i���E#�C��C�jB�9FU^����(�(��t�r���i�����.��[q=Zɡ9?�~*�
3ӬqR������L�2�8-b���(OK�+.D@`r��iFO�T�_�kUOVm&u�%RDr}�(���f59ռ������D��H�͏jhi�AcC��E�	\M,�*�H����6_�Y�L�,��A�!�Z*��Q+��T��Liv`>��4�L�s�ԣ���zKtl܄�{_�A��(���I�^�^�Fj�X�6t�A.�t�Ql��1��#�SI�#����`�K�q��\�I��Ec���L��I����]P;�ee�J�L�RUP$�a�Mȓ�$<��O~�u�;Y��	Pɝ��%6�"5�	E��"�%�)�����L�I��k��ϯ�!4��|�����u\�-7���|[q�_'o����)��砷�	���V�c:�j���3�������&ч�D��`�T��5�{���9��S�o���@��k#���;���z8�&o�JHzmz���F��	�T��+�Қn/\a���Bh���u��$�/�)YE�h(�!j�Wy��K��W�d)N�
�T��z�YĥF�<��k�q=\}TUB�D�U���)�A#K~��c�\���y����6t,�s�:>��9��F��6��ɜ1�߸�ڻג�̧������ὥ=��Z��8��R�MF1N���ѓ��)��
��7fǞ�OO6e��I(��7vP�H%�=<�&�뉎�B�(e���D�!7+0ζK����a�J��&+�d3���d���\O���L��`L�DH��Bkt1�)�UݩG'�+Q�Ȫ#!FWK�a�GږĪ�.p�)a*�Sm���m1��'G���7�1Q��]����w��.��/c��_R�9�<�3��p�N����Q2%b«����s�ڇj�����	���I��Q��KG�y&?��	V����4��# D�L���$"�'���\bq<��z�&m?B�eq�bK�+�Ւ�L��wP�|�5)�V�-;��M�������GT�Y}-�9J�
Ī��d����e�4q2���P��u�P�w.Y����D��+�������o�N���V��s�;��� "��1;R��ژAGֻ�G����^|��W#��d9c\���5G1!�S��*�U-E��J1,#�������5��Em�Z��'�|�}��EP� �`n���� �ɘIp�nD@��GͰ&ĉ���W��Η�5ɢi�g���fG-��a9F�L
��f�5�2PFTĈ�Ts�����Y��j2�D�"]O�Z9�����g�b�����jL���I��9�J٘ڷmx�5��m��8eD�w�JuUS����h�6�W��k7wƥt �:_`1�T֮�:ܪ�cT�h~F��yL�s6Jp��P�-"?���9��z4n�]�a������������|}}-�U�bP��.������!����a���i�Dt
|Ս*�!k8Z}A�&�L����^R|fe���t)�Je[Z��յ����-[�bjj/��k|��&����i�z���$Fڶ�7��=�P�v�:��~]Έ_��Tǥ����2C�����]��NA%4VU9�uv�g!2��}���~����dF�t�����0����Ӆz�/G��M(ɊaFF�I�FEQ���{*_��&Pj�WQ��%q+�
'_��IyZ���q��69�٤�J�ٟ��x}�!KT�D'�I)�',�g~��h
X8s)H��Y��\��\��D0s>-$��q�87�C�L�]E�褨i��=y��|�l� l������&a���,Wu+�vv§ʕ��X	
�(j��K<W�Q�f������Y�5��=�,v�ځ��v��]�VK�_��/������?�<�ŋa������x��044��˗�ƛnR��`?ڨ3���w��� ��yʆ���:<p �W,GgW�ZN��¿�(WȚ(��B�5$�Fq���c��`��U����q޷a�<?����@'wE֤�{=�F"{��1������l�	�x���^^�8�I�y��82�f�7!ޥL�ңk����)����̈�D��g����f
��}�Z�詆4�����Fq��	�����4�g>_��y�p�ڵ�3&'d��Y�����p��1���˰	;�}�3�я��?�>�k|���'��O��=�����MMM�3g.}I�Q���a�LnS�1��N�.���[y�E:S��#Q)�1�����ꃜ�M�[���M{����2C�":CkJa�5�q�|!�E��:5y�71��"�n� ;�qLkaE%�Q�j��!BY��g�fa�t�<<���0�0G��N�5m�l�`�.2�b[7AoH�ˊ��O���شi���o������-,+��E1�����o�v+z��q��q,\�?��O�m�-���UFx\�,V�P�U,���3����jt6�A��P,
�.���P�MQ?�H��B��>澃t�)F|�рc��}5;r/_W=y�I%3�Qn�r0S=mxa��o�=��/nY�}�1��;+�':�m��BUlܰ`8u�(!�p�ǿ@ln/fK$��pl������yc ƌ�4Y�D"s�C�)�?�Ӱi3��U.�p�;%*���?�y��׿�k��� �I��6*�UE,bϐ���C����.í��B��&&'19=��.Ź�#����l>��b�ҥx��	S.�R�R��HOi� 6#�p�Z`O'< Ķ_y#>v���/�����*��ۑb>�$��C��M��\�A*�"�N�e��D�����߿��EB��xձ�G���F�0�p����6|��2��Y��������9(ϔ_���ߌ��ϢᚫQ�i�A�y|N��P>�q>��u)���>__��L&�h��;��sF+����c�%��	�+U��D�RI���3���<��S������?֯_�
���X�dn{��0���������<�����/~�g��2j��^�dϤNX����wl[�����3�}���Ld��?�#�ۅK	�N���Ǯ�.B���@�'\��X�]�O��2�ԆD��X��I?��'��ҋ��m^x���zM�3'Am7�IݩI���'���F�ɧ%=��N���D��J4���U�K��*Ά�'B�"&�e˖��%Zb�8>�g��]ct��{E��`®���m�����p"/�Q.]�6I��������ݧ I�m�6��׆�W��V��f�D�1����%��Dq��
�Ac�����g�$#ԙ[/CX,�`���P���e���	���X��-����涾��1�h�ᛚT�1�A�������'Hs�K�W���U�7�މ�w�&M-h�ֆ�*+j��`�"�R\bt�pF��Xz�5�ۮo]��SU���B1(�}�9�g�o��K%P}c>Bj��*�6�E��j��^�BH�����_�J�YV��e��Q��ӑ���i|����]��#�2��p�?����B�5]�P[͋X1�j��"�ղdU�c��1������ɚ��l���ȴZ"�j�,1q��eյh�]$7mT�6V+"�(1H])��iT
eRYK���?Y$QE�T�zŔF�"	 5Cծ�"a"�D����R�T*�R𫔩O�鍵J�tZ��5i�P�I$U^�͈�|���^���&�/��j�LM*���]�{Dý)�%3�aH�:�D�l7�O���E���Q|�~=I�0����(�RT�U<���Tp,Kl)�@_��_҅tp�G�J�����j�����ZތlK��ÿ�UWn��CT�^n<�Na�%�(JZ%��4>1��HOe�w���x�:`3���8r�(�-_�3gΠ��A}�x}��	�w�Rד tV j��)mmmسg�\}5F���������������k1;;�\.�X�^>�����ŝ�U6`���hikŕWnPM��SC{S;��|7P��6:��L��L6�Xn)2��8��˘Կ���`���hM��Z���B;mb4))B<U����P8j?`X�P�$UwzR{G;_뫟�۷o��4@o_&9Abo�.W+�$�O���0o�֬����*�+�[�(�Z�
Ӝȅ�%�--JC����h���ΝC3�R�XT�U^s�$d��<6���[oU�����hinl��YG�;����ѣ�m��VG�e�?�����ᖢv|RQfq߄#+�3�S�ǨTR!�l�����%\�ה��J8�Wq�;��x���VG��B_v�`��c�R���!JѪ�7i��)x�Ţ�&��*,f��611�"CZ豔!b�P�ɤ�Y�o:����2�����*�n��f�8����jrQ�466*�%N"J���{��^,Y�DY~�+�b#��#��Q�&���Ǳf�e�kH
d�w�څ[n�Y!����.5���(˖?U��Ј�9L�$��L���轓e4I�9�0uU4��.��I�:M��k�v�r�`n����`����+ے��J��'�U�[�4���f�x�-��at	;��w�K��jY�ju��	u29�7oV<_�W�D�@`#��թ􆼏�E�]��W]�8Y����)�]L!(��/p$Ͽ�J�8�܎�4Ѐ�W�QXvj�Y�F分LW^�^E�\*u�2�2�id�_��	���g�Q���_'l�,W�3U*k��%�.��ʂ3�WD\K�v�7Z\�Aj��ղ�̦,�M%0xj��M���-d���3�d�����_4���j��@��b�zo?yLmC�뛃��!Nl������S!��)$GHR��L�y8器gg��#�wt�6��˗@����~�3K[�h��x�@����$�IPُ��hm�E#�E��-#K�"��^J�W���
I��2U'��{j���c������:Hf�cz��;�W�4ݲkN쏃@�L�e���4�Ԩ�N�ٞ��u�x$Y���я��4'�U�CS�z��Z�$}�_$z��_3�o�Y��2�=��&d)��Td�9�K/�����=x��Մ�1�[&����ʈ#�H�h�k�Sosb�1B�$f��)�|�ޏ��;�S��,�r����+����r�J<���X������3 �1jV��QD�W^Q���{�.�ȹHs^"�-���Q�f�4r��'��yz�<�>�A�2�����,�L9)�C��l�� ��w(�#�I���1>�O7����yv��߶��|���ծG6�HU��� �/ˣ"��5�ع�	3z�<��IS�|u���B2%1��{�%.�B M�f������ ��\2��<��
ޒ�<y�D���\�=���_ێl��4:A�0_�,1� x饗��c��ƾ}{��$�K	���M9�S>�R���bN�Q+�i���jo<�ny��g�����޿w���|YBpj
4T��GH*�8�K���8�?��Ɔ�情�G�|��h���,��m��S6n��	�O*Q��prn��&)��%��
��XcS�ڎ�+W*�
�(SC5��mioU9H�� aS����bh�[$��7K��~�[�R�Zü �p��)��Z���_|i��嗭�l��儹)̙;�H��u���3�v�����2��a횵8�� ��=<�@�&W����#F�'qMߜ�>����=�|���荝M���!�$e�^�A�x�>��!VR-_J߿�w�t	�T}q#���e�,=��7j�{�5�g<��-pmWamԊ ��,�:�k�/��T��/o���h _A�<�*aQ���֭�\9��}�U,�K�	%��J��{�bk�^��~Z�C������R�v������uk��4�}�U[���-5>��뮥ଠ��O�Ğ�n�7�r���Z#t@Y�$Ἒs����,Y����et̈́����k�o���_t.Δ	D�l���%�:��\M[Q�I�4�j�d�EU&ި�Ҩf_�Ֆ��2Y��+�&)�E���2H�V�0��B�$`��@53�c
�P�
3��	e�#?�����~��%�d�8[Q0%0��ܤ�Rn��v���S���»��.E��|�I��aW��u�.eĨMK�J�2Iqi?���4I�1�{쩕�^)�,�^�OR9<�댨[��kSmJ>��L^x��9�0�Ն<g�<[�J>2E1KXV�)�1[�AxI]�F��Q��)��'�Q⫤�z�Y[�9!F��E�ɈDy;��F�W�ɓ'��8J�2�)���_UU���_Of7W*>D�Ԍ�V�̩���w��$$�\r�r�:�T��^�ɈY�R?_���^z$��LJ��q���t� �L����Fn�&X�4�yـ�_D�D:2��3E�_��hI�l�v�j>ښ~�5���^�=E��/K�J�Q+�ִ�Ύ@-V�9$ǉǗ���;�RGw�J�R�,�!Y��6@�0�F&��v?�9�sԲl�7*7&�Z���h�t�����O˖,Gq��5��S"�J��(��pfHw%Y������1���Q�9���?�#�����;Q�����:\\�qY/�'�8B#E��}oQCC��8�����6=�E`;nFZݲ�7�r�DF�4����]>7������ҧ��:�wg��S�u��V5�Kֈ7�=x��*��( e��^`��R8<��a45d�
�ɤ-M+W�Vu.�BuE��k�x�i��G>��<�"#m���a?'j�:��~Q�T��;w���O��DE����W�������3�<��У"-�ͪ������>���V�^-����P�[R}t#P{ѥ��j��:��w�?Y��l#�IM;�n��n�V��d�9S˲��R�A�tEig1�:���?_?���=�����Cr��ԤCIzn�^������X�b��'�B880H�9�+7\If�Zy���A?��1�.�����4(,Y���=$�梹��!7����9�r��C�1LZA&��O~?��ϰk�N|�P�e���U�W�`[oX�"Y�����p]��?�4�﫩N���6FTcXΧ�J$,S��sw/�w��/�;V԰׶��4o^�-2Z�f\�z������4?�b>iJ��p?��^�̜ES���^í�eSq��Cũ(�%:F��I�H2���;8!&ޫ�ؠ(���I9E
�)ޔܬ�����E�M�S�a��];�r��?�����-��5F�)j)$^w��=z�@�U��Ff��k�����cC7�|����G��կ⪫�R�G-վ��u��T���{Z��N*~�?�X[��m�vY�T�"�ܢمL�0��,S7/� )b��x�]����l�KE�9|������Ԇ�BaEKU��m�'���E���p� ��,yBnz玝`�]KO6��uS���%���j�څ���(z��^��͛U�q	�.&F��׋�݄9�:�	W��i|�S�)�;r�^~�et�Zs��Ԟ�Lc���i���-�/)H�"���Ռ���e�+lYU}�a�d����x[Kveur��b��ޔ�躦-{O?���5�фz�Z��P�8v�S��@~P�a�Yao<�r��=�1_A��T��h��	2�!�����M&��$��6-Z�m��6��Ǜ]��=$q�˄H�+���܂�]CW�K��E��/&�}��F�C�SQ%6o��F�ݻ��,������O�}�l٢z��;��WmFߜ~>g���B>�"V��+�8������+7� �;�c��ږ��9=k�gm�i`禵�a")k׮̳��.� �X{�m�D�@ᶄ��q��� <�C�1�����&:Qʐ�<�
Wk�q�=��]�;}���n�MՑ�2>}j{gWmڤ�[�T����2j�zS�jMR����n�TT��K.U�5�p�/<���F^�@8�z�M�j�F|��������N���L�@�q��wc����A������y���'�㠮G����#tȘ�c�uYGU�me$du0naLQh�҉19$�7�$Մl��˔���
�R	�T.W@��!%�̂
i2�8�������P" IgN����T=�����4'�̜�o�ziA%�Y��\q�M7)��B{wQ?M�~}Y���O~����$zd�P�eF��}]��8'���>>�����_?J�Մ�+��{�QUb��kI-���2l(��7�(��!�ɏ�]S��y��:���f���<#���LϘ4٩C�l!��2]ʩ����Ď�1���0�����OWf�F[��.d{������e]$<��U���ي4�%�u`�\�e��u٥�zMnb
Ǐ��b�!�)b�=#{����.�Hh�y�m�5�=}�V�W���_`ǎ�ɏ���OU�71Z�����J�339<��� ���7I�Y�����(xS�(�'Fp,�O �����tPN�vt��ٞ�]���� �<����jA{c�&Q�j��$�ݙ�v��������ᦥ�o���n���~m���V:�e˗C�Ť� ��d3��D��a�i2��IN�^���Z��3O�~��J�;q�v�QD�H�ee���m�7_/���Kzzz`�R+�y�&�>{�o���;j9@T�Y
��_=��������BY�����]���%�7ijv��(W�2C�P�:���)����H�����}���w9V��[�q��t�싴�Z�1U..� ^"���1�(��(�r�R���5=�ቜv�����+#���)+�J��'\��VlEZ����>� i��\��}P�2���u{w�Zf�H��{?�b��8�S͓���s���-���G@��4�y�;��уG~����&<I%��Ǟ���'�ܳ����~��{=� ���R����3(r���Ȯ]��m�\5�ɂJ�UӪ���ILt6�X��̶��w�]7_����`�K�Z>�6��R�5p"�̅�*�+���ye27���06N�(1on�LL3"����;�t&�h�(�Mav5�F�����3+_2�R:����\9!H�dX�ɡ��J$a�B9_��s��j��Y�Z�l)�V?�����T�٣���`��Uص{?޿��|�R�J�	�RI��%x�՗���㯿�78�{�����I.�kE�?�:�rl��⠙�jkk�̵�r%�g�G�ya�Fn����P�23f���l��jQ�<����6Q�&�Oh��9?����pus���fz�ɛ+	���4�v���,���s@UR%��˗h��{Vy��C�U	}�b<��ӪQJ��T�[�l�m��%)˵v�\I���"�z�i��=X�t%�Z��~O5H���~��5���	<�ȣx��g�!���?A8������Sa����K�n���L3͉�󞢈�qZʁؕW�h�ֱ��׹���eM���_�"V'^Ԛz��C���%����'0۔�q˼�������(�z8C�B�����Zuj�n��FG}�\ĝL���w'���������ߤ�!5-�"'��w��E�K���S<\Gg�^�v��S���O|�n�)dk�֫2��}��x����O�ϥ�RW.W��T\��#��\wӍo������&�.}� #a�`�ʙ�=��2Mx.�g̭���?an��S�4p�)-�Vbj��F��i�g�Y#m���L��V�rP��3��s�qӗ����(��;�TE3����!"]��w�A[k�x�\v��pz��+Jv� =�=���X�h1��%j"eeq.�y�+�e��a�����Z�����XE�5�_�vZ��� C_�j��*��5���+����!�P544�<t����!'\��6!<*J�T�`.F�Ebj�)k.�����b�)�qjV"��@14ul�{�Y�HsW �����)>>��gڵ'�*3\�MA�����I�����p9�L*��tBݘ����$�J6Ꟈ6�^
y�C%�x�S�A����z6�V�"��x��7� ����� �/R��h�2�4/̝;_��W�裏���{㍃���)���j��R(��d^��+�:o�B��"��[�/��y+B{=ݭ/[{�ZrRBra1���Xع�[*�D�K�������� �Z7������J��!.��Nu��/�+Z���0oniB����SjRW�^��m�<�N2!��çU�$��%_H���ʊ�T��,����o�=���/}�KJ��!��8p@E�H�d��3��4��T���7���)QLv���#�eW��l�c�����~���\���h�h������%p�2(O6'P�fJ-e7�<1�%^���9w�"��e�U.`��\u�q��pΧ������ ���l�7���[�l�D�=�X�4Ȧ��'�sr��7�~��/�9!O<�jb�6�t}/HwO7O`מ�ؼe˛��i��G��RW���\�l�R�	���P>���v�*���3���w(�q�]Qpv�[U������Ov~13��[S'JH�G�j�Ȑ5[H��&�wB�)F�s);+���}�+��م���z[a撸'2�H{��q��L�+G��J6����k��b	4����,�ڝ��q�Y��6��p�ۑ�<�L#�ܰ��(�)�YQck�;oW'�)�[��Z�	#˸[�\�G0���/�&>���Ů];�E����9tv� ���"L^��#�*�h��݃��3��]��c�U��航Bϟ7��W�����X�w�G�2�x��UD�Gu�k�|S���nH��jyǏw�����zܬV�3���yMm�tk�x�ůiZp��EliS�-I]�Ib�����o݆�G�p�7t���c��������!trD_���R���a��Z��|��d/JX5����y~
��+���c�ĉ��E���Q���9}��pe��s���Z��
u���.���ݽX�j�r��c�x%?0/���;��\�>~������)ND`�����@G��,]�#�Nc<�<㵤]��Ё�����.� �=��,0I�T*���s��S/a���������;�x;�nڄ�_=��h\հԹ�~Hue���+��}���V�x�o�����ڑ�6�(X�=�r�\DW$%��jC�����}����TeY��Ȉ��7�R+�"��y~-�~���q)AZ������_��)�v��=�^�����ݼ#}Oǣ����p�P�s��M�/�Tz��N�>�� 
�%��2�����Љ!DIu%
ҙ8&���՚Va�ΐQ�!�ꐰ���@��,t7CA-@k�)/uZ�{�x��k��4Bu�oub6�tHP�")�ӌ�ڙ��r�VݛU����F������ІZ���h�/��z���R��X�����9[ҩ܆)gq1�:k.���H�f���L�M5����y#���qL+�GU��"�<#g��O>)j�*��)�F#
�"1����p1�~+�>kC#���a��&�+�(�P�z}����KRU%So��
����T��R�Տ��K��◼&�V��K�gY�Z{��
�����_I��Pa%��r2���	���8R�SC�b���

�Ѥr�M�X!�EcC
s�/B�29?�Γ��Rsp��4�����ԶYX�D��'�O��43��ŜJ�cғ&8�2��),�Z�d[�*fΐ��;�h}�ENR"�L�JN�1�ɶ\+#I��j�ܤ���$���5u�� u&�'}��Z���nM-�J[x*������2�Ҙ�tJE���b�ni���ֆ�@�F�h&k�D-�ɗ>��Amo����Ũ�E�*8TmsG~��B�F��j��EF���UՙI�MD�0'��As�A���i�C���`��-m5v$if�(7�1��(�x�M�HqV�v�;�K>V����U��(�����]��곥��Э�"��A5�:�8���pʾrߡ���)��]��fԙ��&Y����I��X��*"�ʅl)n�+O˶�]���l9�9��:�՗���PF�O�ē�i�Qi��8�6�p���@�N83;B�9'qL��@�1c����"�t\�>��h�`�d})��\YVG�p�(��4�=�|N|��dɶ�W=��&�V*����ܠSmO�9�U�N�IZO�j�7<�/�u��R>�(��#��:S�<��	���ߡ�����(S��KS��ۣ&��-�]���	����%)��e��8��	�o$�%,9hIS'tK���L��ld�h�d�4��n��U�`��<3	qQL�Иm ��q��rC�]�F�#�x?��+=��ឦYB��9�I�N�U���[9)٘��C�795� �Q�!�����>uG���W������/ܣ���l)��D�A!p��b��f_Ux�Z��*�3)����TS�W�8kE��j�g(@�|옜)d@�ThJ�1���]&�6���'�i��|y��a�᱁�F��߇^3�<��R^-�ayB�&�P>/K�/�?�c��U�mLf���?)���IӐ7����)L*��t5�Qݖ�z���4�ĥ�Tu����ٔ0$Wл-Y+�=xr�#�:,��� �Pw�e[�h*`Sȑ�.!�|!��K����W/3wɶf�/�d�$�0QG9Y�|A���y&�R{��غ�\9��/�Uu�x*��`Y>�U�L�Z���ec�j_��?�+,]�M�MM��0+Ҫ(���e*֮#J���ԇɖ�K����+�����A�{o��'������ZW$��٢�łLK��,:A��ln:"�N9!�1�r��[wjUͱ+�ѐ��%ߟ,ȇ�h�l:bWm-��Z��5��*�m5�t;������d��ˮ��34���Zfd	dc0YRP�dO�L��ON�SZ���wr&��Y-����
EO7#L�ߚm6���@N����0�̻��y-���$,�}nJ��"ѦT$Ax���nŮz��H4�bnV�-�f�6��%
)�D�t���M�$�r��eE�>��J=g]sb�9n���?2!�Bw��~Az�TS����Ӗ(�|Qr,^䀘�m��ݰ�/��r@1ī�e��j�G��c��Y��c����@����̀�W9F�	�VD��B���@du81���ꦗd_.��E���G��˸�>���'���:	۝��C�y��pF�3��Ɛ�2�q�|]�za�a6���D���B��9�@�/��R����r���!^bd��p�\��O��A�*��8x??9���G}�������iw���K����1�o����s�b�e|��1����39��ҍ�:���/yа�Gs;�    IEND�B`�PK
     ��Z A���J �J /   images/36e83e0e-fd9a-4553-9782-762f273f5010.png�PNG

   IHDR  �  �   �2%K   	pHYs )� )�;d��   tEXtSoftware www.inkscape.org��<    IDATx���wtUU������@]EED`TgFѱ*�4یPT�U�23���`G�JSQ��K��$��{�{�?�`�)7�[�<��� ��s�3�51���a�&"""�*|����К?�k��B ?����	��~^@����|~(`������(�w�4�Yŀ(��<L*�"�(�Bi�ߋj��y5��|n~�59F�
t�� 1@T�WW ;Q@g�#��گ@7eu�~/֫�L
�,� k���, ��_DDD�P�.""M ��a'�� 
�����zdZ�����7 ��� �����,�Eq-�""Ҟ�=�����0���E���Cb��(//�����FII	UUUQUUEII	V����
�ʫ��U\\L��fWTTPQQqD���~~G�O4���#g��������?>>>���E�N��X,��닿�?������Ҋ�*+��P���)�-dP]��Rix
���H��]DD��z����Q�=tvփ9t�yyy���S\\LQQ�%���V\|��EE�k&wHH!!!|��!!!��~-<<���p"""�ԩ�3c� )�$�Xj�� ÙiM*�ED�E'�c�_��7�8�<//���l������#77�C���999��呗�Geeek=�C���!<<���0"##	#<<��Α����(���	k�G�Q]�'c���]�`;Յ�����P�.""�Nu!~vN�����c����V+���ddd���S���߿���233)--=�ǈ���ETT������Y��QQt���0��QyT��o��6���mTO��/H""�r*�ED�:����Q3:^�S�Q�Z�ddT����gF�����oX�-틟�111���W���{ll,�������Κ�}+���Fv�ƨ@��d ��.�b08H8�+++#--�}��.�k�򬬬?l�&`�X����C񞐐@�=��?�U��M�l��&`m�V�]DD��7���O��)u���VXXHjj*�����M#%%���4~��7�Ҫ� &&�=zЫW/zt���G���Ȯ ،�暢}=���i�����
tqTw���`0l��k�.RSSII�.�SRR����aq�Ν;.�{��EϞ=�۷���%�L��H��z`iwT���HC:'�0�ti����c�v��AJj
)))���jD\ڜ��(���OϞ=�ݫ7�<=z��b���c�_0�끟�.�""R�
t����Y�	G�z�f�l6���IJJ"iwR��II;5��;ӷo_����q}��_�~���G?��0�	��5�n��6A��H��E��ñ3���n�ޜ��æM�ؼe3;v�`���X�V��i+����޽;���甓Oa���-i?��`���9+���x�""�7՛�����~�ȍEEE�ر�M�6�s�N�l�B~~�3���+�������p�~�i����� ���k�ů�z���iaED��T����?^�`�<L���=W�����;w�i�&����m۶��o�9;�H�À8i�I8�~������ȭ���|��z��*gf�R�."�>�Fa2
�7wCyy9�v�:<]}�ƍ9=��)  �~��q�)�0𔁜v�i9rk���
���Lv�6M��H��8;�0�+�!/--��_eӦMlڼ�M�6i����o߾8�SN>����ȭ�U5�r ݩAED�թ@i|�.�/�)��7wCqq1�����Y�~=�����v�'�Ve�X�ի�b��!4���`Gnݎ�2,,Vz#'"��T���x�h௘\�hr������$Y���6PYY钠"�:��~��1d��r��׷��J�^��X�wzPi1�""���J�Z�a4syFFk׮%q]"?��%%%��)"��ϏSN9�3����!C�ׯ�#G�m��,� �Gǹ��x�""�\���0�3й��999������O�[����פ�6#,,���s��3>|8�;7�c�&_ba1��7Q�."�z����\A���F���vv��Ebb"�׬f����綈�D�^��ӟ��C�`РA��VE��������@����� .�YO~��X���BI\�ȪU����qQDi�BCC<x0C�s�!""���v`#&���>��5)ED:.�""�s
v.��R���:&%%��?��5lݺU�����Y,N>�d�Έ#8�㚻e� � [��PD��Q�."ҺN��X� ��d��ٺu+߭�������F����xF���sF2`���6�ۃ�GX� �좈""�
t�c���I��u�-�W|��+V����""-����u�(����OS�S1��v�&��H��]D��$ ��l�6��N$&&���Z����"�%i<�Q��s�!00����1Y��w�=.�("�n�@q\p&c��4rFyII	��=+�Y�ڵk���piHg���c�С�w�y��&�P�|��B���a*�ED���	��@��UTT�z�j���+֬Y��juiHW���cĈ���a������5ֵ
X��[�"��e!ED��""d�ag<�P]����n�_~a��%�\�����)"����ӟ}���֬��1xXJu�.""5T�����p5&7���u7z[�|9yyy�M("��BBB8묳u�(���W�� �c�.^v�0����R�."]�;�O�5�i���,Y��������\ץi�:w������Gӿ�ƺ����>
\PD�è@�������0��o�Svv6˖-c�Ť���6��H;ӻwo.}\p����u+��S,�|Cu�."�a�@���0	���u�Z��]��%K���w�QU��"��4��ϧ��___��Û���aY,N?�t.}�{.���#؃�k����.("�F*�E��3��j֕_
4�sю;X�l)K�.��@�+E�e���ؽ{��Ez{{CTT��ੌ^pp0g�}6�/�����w��a�
U�vN���W͎�gee�x�b/YLzz�kӉH����Nvvv������S�N.Nնt�ޝ����/&**��n���oY�K'"�*�E�����\�ֿX{4�ǟ|�ʕ+���tCDio�lق�fk�Ohh(			M�.�>���.g�ȑ�-Ш���K*�E�=�L��Vฆ:dee�����g������t"��9R��Att4111Z��.��R����55����^�^�p""N�]Dڲ>ع�P}\�4Z."��w�^rrr����M\\�;w��t88�^���Xx���""�B���5�\L������b���,�xpy@�x*++ٵk���-�/00���xBBB��������.��1Wеk׆���75��?t���*�E����i�}�a�>X�����G����ddd�������É���������s��+���Nk�����H��]D<��ع�	���***X�l.����$7�9Rqq1{��m�h�aDEE���-Էo_���*��׿6�����Xx�,D�c�@O5�)���~S����O>�Å�����t""M���dff���IK����!66V�ӏBpp0_|1�\}111u1�%<�pm:��@ObFcr/0��;v����|�rMc�WVVFZZ���-�700���������}�X,�1��W�e������X�����h���x�"�	�I��I��+**X�t).��ݻw�>���10M��r�����C���ݺu����	��?�������|�e�DDZ�
tq�H�����01??��>���?x�E���x���
���KQQQ��X,��O�X,NH�����sŘ+���+	��ɜ ٘��f��!�T���{��ΝL�_ܿ?��._|�E�7Y�t999�۷����{}||��.G��ߟ���o��fqqqu)��,<��8��tp*�Eĕzc����_ܵk���֗�H�WQQAzz:��Gw�WPP���Z�~jשO�4��N:��.v`;\�ND:*�"�
j
�k��#�i��[��|��U��OD�=:�������<����É�����c4p�@&N�Ȉ#�P�,�)�7�>��t$*�EęN��~�o����l6�-[�;�CJJ�{҉�x ��Fzz�Qi�X�ҥ]�v���cԻwo�_;����/���Կl�b�*�E�IT���3�d&0�z���je��ż��kdee�'������#==��G�}}}��.ǦK�.��v<�]vYc;�����gG�vN������ .������>���o�';;��DD<_UU���?��+BBB���'0�{pJEDD0��c7nAAAu��9�
�&��J����s0yQ�BII	,���;��""MAA���X�֣��Ν;��Tmi���p�]3�+�����׌��vq4igT��ȱ��40b^RR�G}�����.�""Yk��׮O���ih�3i��� ƌ��	�ԩSC]V`0X��h"�N�@��q"&c���<??�?���?x���"��iG���ػw/G�������ڊɚVZZJVV6����J����ҥK��q>00�K.��I'5��� ]MD�8�"���3�+�#�
���g�[�Y�p!���n�'"�>��v222�ys�N�:O@@@+%kXYY;w��n�����E||<���N}��r�W0a���^~�1� s�ݮO'"m�
tqD7�܇�u�w����,\��7��&���n�'"�1������vL/B� **���������($''7��H׮]���sʳݡ�P�4q!!!�/ہE��\Qi�
tiJLMa~#pĜĲ�2,X�[o��5�"".d�&��������q����������7o�|�qq�JKK�u�֍���V}�����2q�D���J����_���,<
d�!���*�E�!A�m��1`����/x��W�i�"96����ݻ����h�������Q۲e6�����<�}��W��ɹ���b�4�mZxx8׎�������5���<WS�������D�c�܄�L�Nq^YY�ҥKs�����s7���'..ܲ�2���HII9����g�e={��4�#r�l6rss[�y�&//����.���?�������1��I20�zK�D�c���Ժ�y@���v���˗��k��o�>7E������w��c���X��]�S�_ZZʎ; cȐ!����f͚#������֭���������Y�������Q�."�1y8�����D�y�v���X""�RYYYddd�a������!>>���������t���1�ѵ�			DGG�3ښ^�z1��)�1���?cp7����"�1�@鸺c�a���Y�)))���+�X��M�DD�hY�V����*x���@PPP�ﭬ�d۶mGlW���'�x">>>���2dӦN�o߾�/��G��]�LD�M�H������z;�<x�_z��K��苈��WNN��ﯿ���t�ܙ�������dggSPPpD��� �u�v�Z���b�p�E�����YVL^��#@�\�/"R�.�qx�a2��{����w�y��o�o��DD��l6���M�I�(///�v�J�.]Z|,�i����a�Z���uya^ZZJnn.EEETUU��퍿�?]�t!  ��Y����窫�b��׿���C�@�SD�]Q�.�1���ऺ����|�����K�v']��U<==����-���G||<aaa��̹���ؿ���#""������υ��(44�	�'4v4�N�_�!����
t���&�.��o�������""Dee%���k���:u"!!�V���d�&�����nPW�at�ܙ��X����֭��v;#G�l��G5ɥ�6����
t��);�`08�7���T����駟�MDDܩ�����t�V�1�aDEE���W+�;vV����ԣ:r����k��~:���q�W�R&�ba.P�h"�D*�E�SslZ��
y��WY�`�6��પ�8p� YYY��y���������魩������c�����Kll,�;wn�dG�b�p�0m�4����_��`�6ջ��H;�]���ɳ����UUU,Z���^~�U���������{����$$$�*����~k����i������ϛ�����_��T`���H+S�.���a�!n��_��/������ݻw�)���x:��~x4��~/'>>����Z�i����9m�S�0���=���[[�=�~�t�<����옼��i�X6�6M�H�v1&���6fee��_`ɒ%n�%""mMqq1��ɭ��;�f=wee%����7>|8W_}5/��"۶mkѳ�޽�G��~�Ygq�������)�f����KDZ�
t���_Ma~n����r��ߛ���ۭ������o������QXXx�������K\\����޽ۡ��AAA<��S�p����n�w�aΜ9���:�L�0�ڵ+111nM���c℉L�8��#⾮�Y�)t"m�
t��% ;30�8�ƫW���=Ɂ�MDDڊ�M�rrr\�qhpp0			�2]ZZʞ={��l��=�X�p!'�p��Y�V^~�e|�A���~~@@ ={�$  �E��!66���`����/�0�� �O&"GC�H�1�f��������<����."")//g���n�iyL������h����y饗�})���ͬY�x�7~aaqqqt��š��v�Ygq���еk����1�X�X"�B*�E<_v�`|�ƪ�*.\�_�/�����&""mHee%;w�l�]ۏ���111DGG�h�xnn.iii�nfgs��e�̙-ʕ���m��ƺu��'$$�=z�dC�����3a�&O�������sC4q�
t�en��Q���j6o�̼��g��$�6)##���Lw�8��Ϗ��BCC��{��A����l��� �ϟ�W\qT��v;�=���w%%%����E�n�Z}����۷/3��I'�T�R3�����"I��g�ɫ�Ⱥ������ګ,X��ekED��ؾ};eee��͝7�o�>��������(����8�cΔ��7�ȷ�~��=t��//��;;�a\x��1�����_����n�&"MP�.�Y��[kF�/�3M�e˖���O�h�Zv���7�;F�� **�������n'55����f��ի˗/��k�L�i�ꫯr�]wQTT��=�����у����;�@�N����۸���/'(��q,���mOD\B���8�ׁS�6������Gذa��b��H{�믿�}�ys������%44���d��Y9��X�dIC�����T&N���ի��k׮��ƺ�8�Z��Y�_��z�6�!��ԣ]��|�;1�?��3������<r:����=������;�C�hv38���?�E�9}��n����ٳg;��#00��={6:u�������ƛ?~<���JL����~�#�Ω@q�a����۸g�~�a�m��X""�����s�N�
߶��k���7�t��[�laܸq�����X,�����d��۷/�~�~��տ�����O%"�]�]�3����;�TVV������/a�i9������vC������|}}��������LӤ����WUU6����
��'oӧO��'�t����rfΜ�3�<��ˎ���w����9��ۛq����Q���ɫX�plὈ��"�7��@���[�n��G&%%�M�DD��8t�����l6	%$$�U����J***(//������RJJJ���l���G�����f�ԩ��y��믿fҤI8p�������x������q�z�b��0`@�KiLF��".�]�u��3���yEE���
o����N�v������J���    IDATJJ���=��=44����.��		�ΡC��馛����'$$�nݺy��t��¥�^ʴ���{�v4�����D䘩@q��kF�O�ۘ����G璑��X"""��e˖/�:�����O9����o��ӦMs�86�0����k׮��{||<��w?��~z�K�0� �H'S�.�\����;�k�\DD:���2�o��p???f͚��w�M@@�����d���Z~��g������[�nsn�a\v�e�1���޵;�?��Mq�"�����#^C���<8�A����X"""�STTDRRR�}�����SOe�����z���J�͛�#�<��ju��Ν;�����9...�9���SO�i]�h�N7�i�T���>������*++y�7x���4j.""Vyyy�ǈnܸ���0�sl޼�ɓ'�q�F�����"66���(������ŵ�^�?����/�1�<	��V�5g�wgiOzb�)pp��dIIIL�:�����ݜ=+""r4������n�e���;v��S���]�r�u�����?����y�4),,������@����X�͛7�z�jN9�"""j/y���0��w[H�vF#�"��
L^�j�v;o��6/��r�������g�����7^�}��\r�%.L�\�6m⦛nbݺu-�ϓ��{{{s�����X,u/bp+������+*�E�]v^�`|�ƌ��<4�ES�DDD:���Bv�������h�n�Jtt�S9WUU/��"��?�g�X�ҥ]�v�_��I'��Cs�[�n�/-��&4�.rLT���30y�]�`�&.��瞥��܍�DDD<׮]�(..n���#��o�>ͻ�effr�=����o��>ooobbb<b}z@@ ӦN���{�K�1����D��A9:0�����Ƽ�<f�7������J���p~~~:t������r��0��s�e�1t�P֮]Knn�C���v
������''m\ee%k֬aW�.�rF�,���0��`��@�R�.�r]0����j�}���ر�}�DDD�???*++)--m��ڵk���dȐ!.L�}��ᦛn��Ǉ�����������R\\����[g�ݻ��Kӻwoj�-��	�o�"�i�4�]�e.��u���k�^�u�&""�Bv���۷SQQ�h�0x��י<y���VJJ
S�Laɒ%-�7<<���8������1�a0v�X��>���v9\|�h"m�
t��c�qn�zz; ���g˖-n�&""�v��������Kn>��c.��"&s��>���={���>�0���"&&ooo'�k�	'��#?���L���?�ƧK��]��c�P��/���=���<iޡC�HKKk�O@@ ˖-���vM(7��l������dgg��^��Btt4]�v��˫�� 00�{g�˅^X��f���K��P�.Ҵ�1y�m())��cٲen�%""Ҿ�۷����&�t�ԉ����N;�E��'77�Gy�^x��ڢ{}||���!22�m;��5�Y3gѩS���E5G�}��P"m�
t���a�)n�۸e���~8�\"""�i��������d���(V�X��'��d��̙3�裏h����������tM���c�#s0`��L���]@��<�t *�E��&g�6��ɂx��g��ln�&""�~��Irr2M���/�d���.J�~�֭cƌ|��w-�7((���x������i^^^�r�-L�0��h���)�).%��T���bL��_5������|�c���tv��ݻwS\\�d���0�/_�g��d��fŊ�}��lڴ��������>�l��`�)�\,ry �]��7v����R۸s�N�y/���wc4���������f7beٲe�y�.J��v;�-bƌ�����^wn$�c���O��l֙�i���@�8L ��6.]�����m�lVq��Ʈ]����pHHK�.eĈ.J�9���y��7o^�k�����%..���'�k��Sn��رc�_Z��X@�H��]:��1y��m(--呹���W_�1����TTT�����.����|���9�E�<Knn.�����矧���E�v�ԉnݺ����t����y�L�6gap5�KÈx�ґ݄��wmCjj*3�AJ��+�V�����fG����������K]����߿��~��_���*��3�.]���bi��Vҽ{w�q���S��
����]Dă�@���;/c0�n�ҥK���<���ܕKDDD`�Zٽ{w��þ����3�E�<Ӗ-[���;[�����?ݺu#$$�I����Ϗ{K.���&`���eaD<�
t�hza�	p��T����O<�g�}��X"""���FRRR�E���o��&Lh�_G���s��w���Ԣ�"##���w�&rcƌa������ۼ	�ˀ4�q3�ґ�Ss���������3��n���X"""���J������fO=�S�NuQ2�e��x��7������q�>___z���ҳ�O>�d�x�	"##�6�Y���˂���ל9sܝA��`*&� ��lm޼�[n����4��Y,���)**�fk�D�/����� ��t���ˋA�q���S\\̆pd�������\L�$88�0������|�՗�|��t�ҥ�9��
�G��q3�����өs���̬�fQ\\�d"""�b����������ooo�:�,��\����=����olڴ�����+..������`����������l�2����߿m����,C�K;�]ڳޘ|>s�j�2�y��ګ��v7F��U;�^RR��l�}������OrQ:�ֵkW&O�L�Ν��������:t??��Ǣ9EUU�׬&�PC��}-�� �"�Zv�H�]ګ�0�
�Qې��Ŕ�SX�j��R���H��I/++kv�o���08�s\��Y,�8�&M�DVV[�li��4����f��)�;v�`ݺu>������.��$���R�.������d����zۭZo.""Ҏ�Axx�CE�ʕ+U���e�]�i��Ʒ�~KII�'����RRRBXX�K�L?x� K�.��N$66��9��"=X��".�]�/�<���h�"�7i�j�􊊊fww_�r%���4�E�چ~��1a�v���Бl撣�������/����.�BLB0���T�.�5i/�1y����n����|��X"""�*iii:t��>>>>|�嗌9��~�i������u�]�����ѷo_|}}]����_�=w�Sú��
\D�IT�K{���������̺ok֬qc,q��{�6{�whh(K�,a���.Jն$%%1n�8~��f����ӯ_?���^�3��y�R��W.F�ҥ�s���:�_�S�gdd0i�$�"""P��݉��l�OAA��_X�b��R�-}��e͚5�x���-//gϞ=.=g�ڵL�4������0Y�L=i�T�K[v&�P��'P����&�����X"""�N��%%%\p�<��s.Jն�����+����/����dߒ����]Z����3��ɬ_��nsd�)>\D��i���Ev�`6p����?��y���f��1����x�4INN����e��Ǐ��矧S�N.H��|��W�3����&����ЧO���^��ǇY3gq��y��Y,��H+P�.m�?&oW�6��v�}�Y�y�7�OSUUŮ]�����G��|�Mm׈�72j�(rss��B�޽]��{]'N��[n=���,L*\F��@��$�O�������f?�����X"""�*++IJJr�H7�k�����_DGG� ]۲v�Z�;�fwx�O�>.��`���<:�Q����6���߀�w�*Х���R��ᗙ���q��޽ۍ�DDD��UVV�{�nJKK��C=�?���f�_w4_|��_~9���M����������Eɪ��ۗ��z����\ �7r���P�.m�I5�y|mCrr2�O����,7���������T�֤��ӧ�>�(cƌ�0��o� �}�]&N�HUUU������ի����GEE����зoߺͿap���aDZH�x�Q�,�dOLL��P\\��X"""�eff���Ѣ{��w�͸q�\���S-\��q��5�9�a���ҵkW%��c�cذau��1�X��0"-�5g�wgi�DL ��K�.�ޙ�R^^��X"""�VDQQ��ǂeee�駟�p�BBCC9�\�S�':��0` �|�I�#�EEEX�V:u�䲙6��߬ .6��;����
�L4�.J�x��<~M����G]zƦ����?���t����ڢ��999|��'����q�'����Ĥ����:�O?����d߲�2


		qٿ��ng�ʕ` A�j�-�E��tI��w�4^�y��6��v�x�	>��#w��v����}��QQ�򓸢����曙2e
NH�6lݺ�/�����7��b�н{w��{]r�%̚9��%
&o`�@�;މ��
t�$��|��m(//g�}�X�j�c���H{f���������G5S/88�믿�iӦѣG����ݻ�ѣG�m�6��GFF����ҥg�}6s�[g��14���@O��b`DmCAAwN��͛7�1����tV�������������UW]Ō38餓��г1n�8�����ЫW/��v�'����?����tǷ�q��	�`�X۰o�>�L�¾}��KDDD:���2233���=���ࢋ.b�̙�y晭�γ��vx��͛��K��BBB���.HW�[�n<�̳����mހ�_�l�i�
tq��|>�2%%�[o���l�|�)//?\����#G�d�̙�����γ}���\�����;�?,,��ݻ�l�������g��`p>��"P�.���/��چm۶1e�

4�HDDD<��j��������i2Æ��'��.w�����رc�駟����C���	ur�j!!!<��Ӝr�)u������.	!R�
tq�A�,�j���(--uc,��Y�V������i���X,���j�ΝK��ݝ���X�V��n�{�9�g!DGG�����y��'�8��`4���ԣ]��L>:�6|��W�~p6��:�BDDD<[UU���deea��Z|���?��~;��w��F���O>��sx�{@@ ={�$  ��ɪG������6cp9���ԡ]\�⚣�o׹h�"��2&"""��i���Kff&���-�?!!��_~�.��	�<OZZW]u�����X,�����d�Ϻwƽ\~��u�+0,rz �^s��qw�8&a�.�[���o���O��+""""�b���DGG��jmшzaa!��.����������ǉi�/,,�I�&QYY�O?�����iRXXHii)!!!xyy9-�i���a>�>�zꩵ�����t�F��Un��%��?�}�Y�~�m7�i=���dff�x��SN9�E�ѻwo'%�,?���Ǐ'99١��������%KƎ��;�cFm����y�?\:<��
��俀��c>:�Q>��S7�q���222(**r����p�������[�r�-���{���.��B��`�Q{�;�g��`��T���݅ɓ���l6��>���[wfq����������C�:|,Y{��{�q�-�8<�   �޽{�����\�F�⑇�{6���]���`��T��3݃����l6fΚ�ʕ+�IDDDĵL��СC8p��5�۷o���.H�9�������Y�z�C�����ѣaaaN�5b��x�	|}}o4x�?�>X:,m'�2�nqn�Z�w�|�����$"""�r���EFFb��(++k�DD#G�tQ:�Ƅ	���f���͞�c�&yyy��IHHH���*==�;wp�y�՝�>� V8�ҡi]Z���0�]�myy9���ڵkݙJDDD�#��瓖�FUUU��{����ݻ�Vtz����q�Ƒ���P���z��Uw*z�4hO��)o4y3��P鐜���t<v��/��~��s�aaat�֭�����z��СCٸq#�Ǐw�QQ;v젤��i�֯_ϴ;�QZZ�{��=����*�
ti-v��`VmCYY��Fbb�;s����x����&w"�'\���t�ԉ��z�w�}ס�լV+�v��СCN˴a�n�r��/�c�EjN+9V��.�����\�P\\��Sng�֭��%"""�RSS���m�alܸ���֔��dƌæM��Cll���|��<�̳��h�"nT\�1��;;��-����[T�����4!**��k�i2{��F�w$�{���d	����HKK�Y�[�l�[o�����F����S(�
t96v��������s�-7�}�vw��x���G�����石t�R&�\̟?�����l�C������n�Gk����|�������h0;O:��ah��=;�`p_�EEE�r�-�رÝ�DDDDڌ���������}��i�&��Ҏ"11�1cưo߾f����ЧO�&����}���_<r��ɿ�p�S(�F���ؙS�8/..���nUq."""����G�UORRw�q�y�!C��~�z�=��f������v�*))����ӱ�S(�ל9sܝAڞ�������֮5�""""-�����ׯg���p�	.L�ق����k���`�ƍM���lᔳ�:Ć������ǧ���l��V��kA������y����L�6���""""Ұ��`"""��3a�~��'%j|||x���y�駛��^\\Lrr��6�ۺu+��~ۑ礛�f8��ni���L��������Ӧ��/��3����H�g��ضm[�S��������ݻ������������N�^���c���<��su�01�<ﴇJ��tq����a�ٸg�=*�EDDDZ���=z�h�OVV#F�`۶m�	ՆL�4�E�����d���<222��cӦM�u�]X���&�g��#�E��]1�W�j�2������n�%"""�~���5y6:@ff&�F����\r�%陙����:-�ڵk�g�=�l��&���r�M�4�L^��8����ޙ���?�9����H�OPPP�}2331b,pQ��c���,X� oo�&��ݻ�����X�f��^w$݂���=T��Ҕ�0Y xTUU1�Y�Z��ͱDDDD�'��B�>}���o�_ii)cǎe�ԩN;B����K�������qv����亣ܭ��d������M^���㴇J��c֤1�1Y
����G�|�r7�i�,�������-��v�Z֯_��ѣ�-�;��O>����&w��픔�йsg�����BƁ�9��gx��k��S*m�
tiH_LV ���x��gX�p�#����t��ބ������l��{�n>��C�F\\��z��C���o��~��F�X�Vl6aaaN˱{�n
>lxm�p9���=X�$�R_&+��چ�^{�7�|�}�DDDD: ooo������ov{^^���'((��C�:mD����_�ʪU�ػwo�}j�.		qZ�m۶���é��Z�\���@��,m��A���0Y��m�裏x����IDDD�c��l���P\\�P��.��7�|���H''krrr<x0iiiM�KHH ::کY��9�����n�F ��`i3�I����r��˗/�'�pc$���o߾܋/fРAlذ���چ��H>����o�>:��,O=�_}�Uݦ>�|�;���f�@� L� N�mX�v-��Cͮy�3��ݻӽ{w������3|�p�ϟ�t�o���������ۥ��9�H����~p6?��C��1Y4}��tZ�.ޘ|�_۰i�&��1�""""�����    IDAT	����ف���J>��SJKK9��s�<v�#�߿?UUU�������_�#�G�n��r�JN?�t�t�Rۜ �`!�5��֠wtv^����o�����<>�����Ξd���l���ZD�jk� �W(�j���jq�+��싀AV��,�nA@d�$��}�l��G2d@�Ifrg��_/_�,���R�3���ø?�C]]�7�"""""f����.��6x�`|�駈�����|������G9��������n��h4�?B�>}::Ê
c������!�E{��ɓxl�c����fLDDDD���rÕ����_cÆA_<�f��@nn�ӹIII�zu]ll,fϚ�����N�x��J>�	z�z"���<��'Nx9,""""ꌆ���z���W_u{�r_��ڊ;�_~��ӹ			HMM�XRRR0g����ػD`^�=�|��t=D|@���O��	����rXDDDD�������/Ƿ�~�Ѩ@d����w�}7֯_�tntt4222��=�~���?BHH���� l��e���RDp���(�h;���s�29'"""�c��ؒ����ݽ{7��Ţ@d��`0`�ʕ���۝έ��F^^�fs��r��!����j�ڻ���K���X�=�d@�f g_<z�7�n�:/�DDDDD� """����;v�jkk1d����Mj�w�u:�Ç��5�ͨ��ADD4��c9q���������ޥ�X���$��=x�@�7 2��g��ݘDDDD�~[uu�l�;w�K.�E]�`t�G�V�{�AYY���#;�j����
!!!0����������ҳ�� n��% Z<�@�9<������nذ~��C""""�����l�w�EQ�c�=��'O*�oR����������\�Պ�Ǐ����[by���p��ж�N�;�O��b�عs'�~�i�l6/�EDDDD�I��!,,��Ւs���������_��|� ���������u���E�e����K���l�J��,X��Oa�@g�k���y��q�;���ތ�����RYY���B�9_|�n���9�d͚5x������tnwUx�̏g"''��S�KP�y�>�|
���D�}ɼ���F�3g�)���H�HvNN����������ك�n��N�r:744YYY�j��!11s��u��^���,���g���uD|lo455a�S�����T�;�!//�?ύYGĎ;0`� �s���p��a455y4�ӧO�����f{� ���GD>�	z`�h��\��u������G�z9,""""��J���4�9o��6�mۦPD�!55[�lq����lƑ#Gd���<<������@o�>�|����س�`��7�7o�bHDDDD�mF������V�#G�Dm-��v��?��Ǐw:�f�!??ߥc�����8v�A�� "=� �:&�E�^��b{���E�y1$""""�={��Z��?v�}�Q�̃�F���3���o�~��JKKQPP����y�r�JǮ~����o�@b�;����o�>��_���j�fTDDDD�#�j5�Z-jjj$�9r��^{����������W\��kע��Uvnss3����
���=.��2��ײ!"6z��u��8F�� ���ݣ#��;0DDDD���?.���T*�Z�
��v��Q����nCQQ�ӹ!!!��ʂN��ȳ###1o�<���vt
��=� �*&��Z��
� 1j�(���{9,""""�Ef����b���o���R02�Q^^�;�۷ow:W��"++���yv�^�0g����ۻ�0��y y�A����ɹ�j�?���s""""���jѻwo� 9���C�űc���$$$��o��#�<�t��»�
����u�쮅�\����c��ߌ��y��㭷�;�����p���SvNEE��3g�(�����7o^~�e�;��
�ǏGee�G��}�vL}g�cWL{n��W0A�_D́C��e˖aٲe^������Ibb"���e�9r��r�_� �}�Y,]�z�^v�(�(,,��5lK�.Ŋ+���Y �?- ���=�^{c�����FDDDD�TFF���7]��݋!C����Q����������"..�����R�8q�#�}��7�o߾����G'űH��	"�@�����=""""�.�X,��矝^6x�`�^���Nq0;|�0��R����8��������X,\�			�.��ۋ�����2 b1ړs�Ʉ���oLΉ�����4�����hd�mذ��~;ZZZ������?���tnEE


��iee%�~�i�L&{�
"�tkaRt�k �=73�)8x�C""""�@��둕��J>Eذa��.&�2����i�&�r�-N�VUU�����$���x��W�b bX4ί0A�l���p���X�z�C""""�@�R���_���oGss�B���ш�k�b���N�VUU�t$ޙ�k���h��`�8���4i��c �<�/�����Ͽ�������mz�!!!�����w��q�޽��s�ӣ��J�Raذahnnƶm�d�677�b� 22ҭg~���8p z��a��� �wkaR�����!b=��;///��#FUU���""""�@UYY���B��n��f�Z�
!!!���<y2^x�������ֳ���p�BǊ����n-Lݎ	��K��}h��d2a츱|�������G�t�MX�z5�t'�O��'�x���355ձ"{�0 ��:���u.P���ԭ��o�BD.�½>�u&�DDDD�������C�_a�ꫯp�m��t'&L���S�:�W\\��g��ߏ�����K�}�w�}�oB�p{sժU�9k�7#""""� 
�^���Z�yزe��nޓ.㪫���`��_˟6���EDD��x�>|�����ɱw�A����E�[��"V����c�0r�H^gADDDD^Q]]�ҝ�Ć�Pd��^��ɓe��t:���׭"|!!!�?o>z��m�!�. ���(u&�)"�����&<��#.� """"�.���~饗b�ƍ���W(2�����ӦM�����l������E!44��U��0y�A�=z�X��� ^{�5&�DDDD�u111�ի��w���G\{�()a=29����.�9uuu(--u�9'N��˯�����>�	����? ڛ�����/�Q���hddd8M���g\w�u8y�B���J�E�᪫���w��)��׻���7bŊ�]�`Ûn-J�#���ʊ �C�a��10�Lތ������jjj������{FF���k�w��<���4hN�8!9G�ӡ��P���Ǫ��0g�\t�E��I�%�b��;�!b7� ����C?��q""""��R[[���|�l6�y)))������yv�؁k��Vvs.!!���n='%%�.��h�w5@�  ?��0y�����X���\E�0�&�DDDD��"##����Z-;����^{-<�Pd���+��[o�%;���n=����_��x���~������L�}�S���\�p!���;/DDDDD��ш��,�I��ӧq�72I���O��{STT���g���,Y�ı����[��G�����+����c���b�x3&""""�Nijj�ѣG�������0`�B�����J����O���������8����h0k�,��Wg�	E���n-Ln��w���Y�FCC���sLΉ������O�>�j���Μ9�����ؽ{�B�����X���{�sJKK�����b���=���F{� s$��0��	��� b�X{�k����Ή����o���8Mҫ��1x�`�ٳG���˽��+{?��lFyy���)))9�~�8�X�^�o������ƚ5k�a�/�CDDDD�>W����*�x�صk�B���w�y�tݶ��2����ꫯ�~�zǮ����S�0A��A�q��I���|�F"""""a0ЧO�t:�y555�馛�w�^�"�iiix���%ǭV+N�:�g�>��s�`�
�+=�8u
��)�{dm�~�;?�����"""""�,�Ʉ��<����΋����͛ѯ_?�"�������Duu��A@�~�dw�]կ_?̞5����q�@�ۋ�˸��4>D{r �?��䜈����N�CNN�z�켊�
<�����'����I�6E���y֡C����9veiY�\�te=��;v��'�p�#�/su'=33[�lA�=���577㢋.:��yz����h���R���{��+������n/N.��rzC���Fuu5^���s""""
x:�}��qz������QYY�Pd�/$$�'O��s��IX�V��e���¤PSS��)� n/N.a��D��Ey��PQQ�專�������j]:���O?a�С����v#F��e�]&9n6�QRR�g�9s/Lz'�#!b!�;*��de<���
  ˖-�w�}��p������gOҝUw߹s'����F�"�m*�
3f̀J%���9s�cjl۶˗/w���'=�8�b����B�K�FQQ���ZDDDD�t:�����hd�m۶=�_	mw�Wb�ر�s
=r� ���οz�u �=�8Ib�޽4�E�@�]�/Lz---^������{rrr�V�e�^�O?��BQ��)S� 99Yr�d2��ɓyVKK&�8��=D, ���e�&��I��C�a<`oΝ;�ׯ�fDDDDDD>A���h4���r7Km߾={������7��������hnnFhh�G�F?}�4.��R{W� ����tA�f���"~@�'Lyyyxt�0��^������w����رc�I�V��_|�n�A��|��wߍ+VH�k4���Z����:����Gvv���W�����Lл�"v���ɄGG>��G�z9,"""""�SSS���|�$=&&{��AFF�r�����
\|��(++���T�%''���wL�C�@ �y ��wл���
~�!�s"""""	QQQHII��SUU���&�I��|W\\�͛A$����y�Z缼<̜5ӱ�/l�������{�o �   ������+/�~HDDDD����`�Ze�V+))A}}=n��#�MYYY(--Ş={$����#&&�i�|W���àA������!�*������,q��p�� h+���Cz��"Q EǏGmm�켕+W�;�P(*���ЀK/�Ǐ��c4���#���4,�d�c�|�@�ۋ q���������erNDDDD�"AЫW/��Ǐ���J���]F�,���������yމ'����9v���xdq�ݓ~�퍝;w�^@DDDDD��V����)�t�>}O>���Q��������?d甕�����#����Ů]����Y�x��C��@_ hii�}�߇��/�EDDDD䟪��PPP ;�G�ۘL&\u�Uطo��O^������K�"44��u.����A�;�`ËhO����crNDDDD䆘�����Ι8q"Z[[��w�t:,\�!!!�s,


<R����}��cW���t���78�e˖y3""""�����
�^/9^XX��ӧ+���߿?�N�*;���^����X�d	�����!� ����A�G�ݣ��h��h2���������專����C}}=���$ǣ��q��1���(��z����'������Axx��������OC��ٻ~��+ ��^<Hq�=O��S�Y�g19'""""���p٣����x뭷�ȷ}����̔�SPP �����
1o�<ǮKLt{� ����?0 �ѣG1���NDDDDD,~��'X���GDD���QQQ
G���كk��F�����dgg��,�Z���O�>��V��a�B�A�D�B{rn�Z1���LΉ������F�Abb��x]]�Ew0p�@L�2EvN]]�G�G�Z�x��W`���]z��@p{� ��k�{cѢE8|�u���D�+��}�]455)�o{��'�^AWZZ�����u��!,^�ر�w ƹ�pb��y= �e{�ĉ�x��ތ�����(�T*$$$H��9s�f�R0"�&�Ν����9�("??f��5�>��C�<y�aq� �텃��1@$�����_�݋DDDDD
����Z����7a2��ȷEEE��O?u���f��#�������W_q\'6�z_'1A�� �7V�^�}��y1""""��V�ewы���h�"#�}W\q^z�%�9���8u���ڽ{7֯_��!� 7��pawׅ@� � P[[���555^�����(xX,8p��(�9������?�`0(��EÆ;7y����,DFF�����H,�l�cE��0 @�[	ʆgў�����erNDDDD�0�F#{/zQQ���(���-B�^�d����nmm->��cW6���h��kr b? = ���;n���iQ�L&���O�?����#//III
G��v�څ�����IxXX���A��-i*�
�f��]�p	�#]^4Hp�m��遶{��x�&�DDDDD^���dw����1y�d#����o�-;������n=�f����^��b�w�!�=�LН�z{cѢE����b8DDDDD���,[���?�����?L�0#F���S^^���*��s��1���:v��>�<�./"� eee~�p455y9,"""""*++CII�����ފ�k�*�hhh�W\�ÇK�Q�ո袋�*��ϖ}�Xy��`1/	�A�c��hO���7�`rNDDDD�#d��^�n6nܨ`D��h4��>CXX���Պ��|�j��hjj��S�9R�^��A�	��A0�������w�y3"""""r�R�гgO�9&L@Ko�:_�~�0k�,�9���(**r�9_�5�o���!`���Z4��'M���|� K�@KK&>5���^������������&���UUUP�T��������W�Byy9v��-9���Z�Vv�ݙ��#��Nh�Z�m��b���w�/l������Fii��!"""""))))��S�L�}�:����;����e�<y���]~ƩS��p�BǮ���q�����QRR�O>�ě�����0���H��L&<���*��z=rss-9GE���;^��i��?w�Sě ��-����φ� $ۛSߙ*y\������|CJJ��k�6m:�����.�J%��L&t�C���VL{o�cW
l�G�`L�ϕ	�7v�܉͛7{3"""""r�V�uZ0�BEE�B��[o��<�윺�:���u�����gϞ��@F�@L��x�h�V`�;S��*>>F�Qr�������ȿ���K���e甖������Ϙ��X�V{3���;�c���F �����8v��!""""��JKK� ��,��U����T*,\���I����.������+W:v��.-�J  h b�_mG7��N���z9,"""""���b�>}Zr<99DTT��Q���[���믇�l��c4���#�a�����\�������p)��W��Ao�g�'� ����������d�t:����RL�8Q����o~�����sPRRҥ������̏��ץ�wЁx�� yyyxx�ð�l^����������yyy�sV�Z��o�]����(�>|8>��3�y���]:��V�������̴wUB@��N/@��n�$�'� ���o19'""""�s��ላ�����㏣��Z���� �;w.���+;�������^�j�⭷�r�m��:�{��c���B    IDAT����
{���f<DDDDD�!)))�j��㥥������`D��h4��O?Ehh��������w�څM�6ut� �w�#����x� �f3�0������j����Ι3g֬Y�PD���/����yRcc#����������b9[N^��B"��� �ao���v�����H�����3f�l��`7r�H�9RvNyyy�^8q�V�X��!`8����B"xto��s���r@DDDDD�RSSe���9s�Ʊ���3f��K.��STT����N�=s�L466ڛB�I��	�= ��7�Λ�kՈ�����Z�Fjj��5k�`�n�I1X�t)�F�䜮��^]]���;v]�]
���5kZ�8 h;�q�]wv�� ����"TTTH������DVV��Q���K��������N����b�
$&&ڻ�@�� �]
�O��x�'� �����������z����F�=V�U������ߏ�c���9s�L��Gomm�G����c���[���yyy���/�)D�V###� H�ٲe�z�-�q�M���.�LvNQQL&S��]�v-�9��!�E ]�oW�n�?�=3�w����ŀ�����HIF����=��������PD��`0 77ҹsW�G��l�_}� ���H�O0%�=!�����۱s�No�CDDDDD^�������q�Ʉ|�KɃEVVfΜ);��������"O�7 =��_
�݆�>�y��^�������A���K����C����[��������?�IvNii��j.9�sl�W�"�?�����������둗���x�����ȋBBBгgO�9S�Nŷ�~�PD�i�ԩ0`��(�(((�Tὼ�<lذ��C�X �n��7�#A�� Z �X,�9K�(���D���K��l6<��#��HL/^�� 9�����ŝZ��;&����/�x��X�jJJJ�������j����bL�8Q���O�����k��Ω����'O��ڵk;:�pQ�"�����x�h+�0g�/DDDDDD�B��!55Uv����r�J�"�O��_0x�`�9��zm欙�������	�� �7�-[���r/�CDDDDD�&66��Ѳsƍ���2�"�?� `���W�Y�V��fYYٹ���%]���v�.�5�����1�|/DDDDDD�(--Z�Vr���#G��Խ��&!!s�Ε��___���
�ל3w��uw*���V�>.��+ �7�,Y���*/�CDDDDD�J�� =]�P��0{�l�"�OC�����e��l6��^ee%rss�� pe��qB�~$�k �m���~����rPDDDDD�ˊ��dwx�����?�w��
F�_���q���СC�s"##�����z���X�z����] ��#�=���~ړs X�h!�s"""""r*55z�^r���#G���fS0*�����C��HΩ��EMM�K�����O>q��wn�3A1��euu5�.]��h������O�T*dddȾG�e����{
F�.��r�����s��I�?��d�'������;���@L�o p��1o�<455y1"""""�'F�Q�9 ��_��ѣG��?M�4	����7�L.W�oll<���� \�V�>(�t��n���*,_�ܛ��JNNFHH��xSSƎˣ�2�z=>��c�T�i��ӧ].�l�2TWWwt��w/z�%�W��]���:��'"""""r� �ի��Q�͛7cƌ
F����j�5Jr�f����ܥ�����d�Ǯ\�V�>&������&����m���ۉ������N�:���R����P�߿���
F�_*++ѧOTVV^p\�V��/�Z�v�VXX>_�9"""�]� `����@�A���9�VD��9�#))	�����MMM3f��ˈ�����?/9n�Ze��s���x~�[\�V�>$pt���l�2oFCDDDDD@�U�7mڄ7�xC���ϸq㐔�$9~��i�z�{��%hhh���/w�����_
`���d����{1"""""
!!!�ѣ����w�V("�c0���K���fTUU��V}}=>��3Ǯ; p+@	z�� ��4�S/DDDDDD���Qw�ٌx��2&L� ��(9��k@[Ap�W��c=�~h�� ������/�CDDDDD�ƕ��ǎ�SO=�`T�%&&�G��oiiAmm�Kk���b�ʕ� }麟��݆�����҂O�倈����(����gϞ�sf͚��k�*���8q"4����ӧ]^k��hmm�7U��i���>Oг�?) �X����������:+11����s&L���$ddd��{����Gss�KkUVVb��� ����ʿt�� �Ʉ��z9 """""
t����j���'N�`UwO?������.�5�|��f{S&��w�s�� ���֭Ù3g��V���4�9S�LA~~�B��K.��]w��xUU,�Kk�>}_~�eG��� ���k�7A��	 !  �"/Y�倈����(XDEE!66Vr�����_�ȿ�}ol6[�6_�/���fo�������k�
��͛7������Q�III�Z��_�v-֯_�`D�cذa��̔?s�DQti���Bl߾��CğѾ��o�5A�,\��P�����(i4$''��y��\N4��J���g�q�ٌ��j��;/'�:^��'����!��y��b���ތ�������T||<BCC%���ۇ5k�(��x��!9ޙbq{��Ł::D�?��'������Y����z1"""""
f�  55Uv΋/��]�ǣ�Jot766������>Y��c�7�ۻ���_�.v��?q����;oFCDDDDDA�h4"::Zr���Ҟ|�I�T�iigvѿ���<y��C�3������_�J{c�'���yE�=d�_|�E�"�/YYY:t��xuu��=�l6�,]��5�o�
Pa�����G ��n�u��y3"""""" @HH��]�o��F���ǓO>)9&�b��\[�f͹��rH�O	z ����~���V/�CDDDDD���.�{ｧP$���oD���%�;s�ZKK�-[��5@�T��$�6<@ ������DDDDDD^�l���?GAA���A��OH�[,�N]���e�����\�/�K���֭C]]�7�!"""""����D�1�Պ>�@�h�ǈ##9ޙbq���X�~}G��GD��b�%A ���l�g^�����������d�E�={v�����=z��xcc#���\^o��%��� F��B�!AWAğ썝;w�رcތ������HRBB��Xuu5�/_�`4����3�j��xg�����c�޽"�?�}>@ ���y ��O�z1""""""y111�j���s��U0�������K�WUU�b���ާ��:63�rp
��]�x����[�n�f4DDDDDD�A@\\����͛����`D�c	�c6����.��i�&���vt��_,���~ ��7>��6�͋�9'��������+��2d���%�;s��f��_��f }��|;Aw�Z�������""""""rN��!<<\r|����|� A0v�X�����N��j�*477�]6Ho�� _N�y�����Xɱ��"lڴI�`�Ș1cd+�w�ʵ��:|��>~�/'��V@�e�DDDDDD�"::Z�*9��]Xtt4�.9^[[���V���+�|5AWA���Ʈ]�x���J���(���˗���F���ǓO>);^QQ��Z���سgOG��	��\�'�p�����jDDDDD���577c�2����.�W\q��xEEE���?�ʵ, 7t9�n�	��q�/��˱e�oFCDDDDD�%F�z�^r|޼y��g�\�X,���vy�͛7������!��%���'���X�j��ߒ+�}�v����
F�?�.{��W��w+� zt9�n�	�c �@�7q��k�Q����B�qމ~a��G��ollDSS���Z}����n�|-AWA�{c�֭�C """""�3��D�7o,�����\�~gv�O�>��۷wt�ˉ}* 7Ȱ7V�\�H������<D�{YY6lؠ`4�#==C�������juy���V:6{�Ǌ��V�~^q�s>� """""�SQQQ������?J��l6TUU���֭[Q^^��Ѷ��3|)AO0��X�j%��Q@P�T��������;u\;�:������Y�V�YsN�3�*�K	�8�;���_��Hn2��h�"��*�
�=���xss3]^��`-|�X��$�*�8�gq8"""""
4���		��1cDQT0"�1f�h�Z��������;:|�X�O`0X�������\���G��o�Q0�ѣG6Lr����S��/P,��.�A���;����=Q�pv'��3�ƿ�?^r����l�rn�8���+��8�[�z5��Q@�h4����_�z5JJJ���t�M��Ζ�l���k�vt�@��y�/$����(�X��z/�CDDDDD�}���%�,fΜ�`4�C�bq---hhhpy����:���^�� �'�bGż}�����؛�u+��([,n֬Y�z�:��5
:�Nr�3��'N���::D�Ws�v���
{c�2S��������.zII	�L��`4�#!!w�u��xg�ŝ��^�O��� �&�6�����ʊ�DDDDDbcc�V�%�_|�E�޽[������G�1QQYY��Z7nDkkkG�������� �A{�믿���DDDDDD�J�R�^�f6���0G�������ׯ��xg��744`���F��y�7���<�NDDDDD�$!!*�tJv��1<��3
F�?ƌ#9��ڊ��:��:/M�.�&�%趎����y|��������^�GϞ=e�|��X�n�B��Q�F!44Tr�����~����D�Z�8o%�p���v�Z�}NDDDDDA'!!��(bܸq��QQQ��{$�kjj\.g����_vt������[	�p g?����DDDDD�222��h$�KKK��s�)�7n��(����ry�󎹇��ˁ��;	���/8���B��ADDDDD�mZ����s�O��;v(���kd��u�{~~>:��!�wb�*o$�) ~co�[��)�����(�EEE�Vu��l�0a�V��Q��Q�FI�577�������M�G��"o$��۟k�Zy�9���Th�Z��={�`���
F��F�	�^/9ޙ]�7:~ �F۫يR>Aq���;vt� """""�@�V����";��Cqq�B����86Lr�����S���سgOG�C���L �7(�x""""""�#[ս����_����݉n��P]]��Z��W�����@��A  �L&l޼Y������4�Tҩ���˱q�F#�m7�|3���$�+++]^�o���d�7@�]tet�#[�nECC���'"""""�uz�III�s&N���=߁N�Ra�ȑ��hiiqi���z���
sW2A�@{��~�ࣉ������GRR����C�0{�l#�mcƌ�Z���L���r�KH���a�%�6�o����[�nU��DDDDDD�D�c� ���ϣ��V��|[jj*n������J����Z�6mBsssG�M�j��%�B�oj���������������ሊ��///�+���`D�m��ђc�555.���܌m۶ut���M��
 Y��ƯXЀ�����ș��� 9�����ѣ
F���N���K�w�N�ss�> .�r`��L��p��/����z$&&J��L&<���
F�t:z�!��:�
�~Q�ܦ�.�	� w��~����"""""�`����F#9�r�JlڴI��|�c�=&;��k&�	�}�]G���{�J$�p�������$"""""
j�={�������"h��W�����J���s?/w� pIW�rU�'�6�e����	�w���G���8���J��ڵ˗/W0"�%��n2��=�.�~@SSSG�w��3ݟ���-[��x;Q���Ȏ?��s�X,
E���~���I�w������!��������o��qDDDDDD�)<<�����G���9s��7���㮻������fsi��r� r�
Ή�N���3�Lؾ}{7?������(p���S�ڵI�&���Q��|�#�<"9f�Z]�}�֭0�͎]p/2yݛ��G ~q~�������:%$$111��N�´i���7]��HMM�w��{CCv����!v�1��L�{dolڼ�EDDDDD���ewѧL��r�T*��;����t^.{���&�;�;  `�ٰe˖n|Qp��tHHH�����믿�`D�iԨQ��UUU.��i�&�w�U��c�ݗ�;l��۷�����("""""�`����Z-9����D��|ONN$9��)���*�߿�����wW��w���y�F�Abb��xKK^}�U#�Mr�⚛�]��v^N{=�h���]	�� 4  �"6o��M�!"""""
N����j���3g�DAA����|z�^r�3��hq'.)ݓ��0���#Gp�ԩnyQ�R�T��C�^��l�k���`D�'&&C�H��UUUE��:%%%�����p�y=�;t�lo�8��5h�Zh�z�����"���OXۿC��Ύ��zh�Zh4٪�DD����dw��͛���|#�=r���f3���\Zg�֭�H�"��p�({c��m��""��!�T�i���t�h5�juPk�P���Q��mɵ�3���l6�,XmVج6X�VX,X�f�M��ͰY�yuA����������f���˘3g���[o�qqq�����xee%"##���m�6�=�ތp%�힊�݆�h�p������#�����V��N���}�[��B��A%S��;�T*�t:�?��wS�	fS+Z[Zajm��dr�8 )#66eeehmm�������O�O�>
G�t:��>L�>��㵵��Z��U��������H�m
�gt�q0�������#""

� @o0 2&	=z �Wz��Azvz��"61���!�'睡R����a�Gt\�Rz"-�72/��^HL�B���(�	� �.��j��/��`D�G�fs�Zp�͆~����!���ß��B�	{�_��7n���DDD>G�RA��#$4������t��]L--hnjBsS3�a�y""ň��C������j�@߾}��w���?����"""����t��C�b��MRx��yO�dg�ٰc�/ODD�}����X$���W����@lb��Ã29 ���Ș$��D�>9H��D|�$#"�����DDta��O�<Yr<�1Br�����������<���ر��������]����[�Z-"������^}r�ڻbjcet	Z����HJ鉌�l$��"*6:��ۡ������H��������
F�[��~ɿ�EQDMM��5jjj����������`�v""�wZ�Q11虑���,���cD8w��@�R!�hD\b"Ҳ2�vדa��A���:On�f�aʔ)
F�[z��_��ג㮼� ۿ?�.��h˅=?a\�hol�������漤<.)!�� 7�=J��!2&)�2����d���C���ewї,Y�cǎ)�o���{%�\=�~�}�m9�5n��s	���x{yyyP��NDD�EP���^m�"�rei�ڳ�zzV&�bc��x�&X"�`!��n�X��k�)�o>|������g�9s����j�K��b�r�֭����|��`@|�$��n;�����iu:�%&�Wv���`���;�DD��l}�KJ��    IDAT(((P0"�ѫW/8Prܕc�(�����<����t gk����2S����G�V#:6陽�ڻ"�����O���
�eg"6!���Q����$�1�ٌ7�xC�h|�'������������F�6�{���вDDD���������,�&&@��X=�fj��q����D����ND���h��9s栨�H��|��c���ܹ��5 ���y&A�����B]]�G�%""r�!$I)=����11����a��H镁�޽���DDA��E7�Lx����wddd���/�w%A����ѣG;:rbwx���7v���%����N#"�ֻRze�0�(:�	��H��Șh&�DD�̉��3g���T��|��1�����f�k�ر��!�&O���b g?�ٹ�	:y�pv�5I)=��9�G���Յ����11Lԉ�8�Eoii�;Ｃ`D���{�u����ݻ�� ���'��[�&�	���DDD�cO�{��@o�;��F��".)陽��9����N���裏\JFMFF$9���d߾}0�L�]nsw?A;�ػw/Z[[�^����UaF#�2{31' �F�kKԳ2�wԉ�A@bb��x}}=>��#�Ϊ��W�ZZZ�ݠ�O�7�+�@D%� ���4,X��ݘ������KL@HX��CQ��j��d��b��l���n��-m_�����jKJ5��U��B��@��B��B��x����֖fT�.Gsc��C!"��͆�~�I����D�V}DǏGVV��xVV"##e�x�����7k! ��{�$����UhO��#"���h����Ȁ)�f�X��܄��������--�hin��d��lv�)~g�T*h�Z�Z�CB`1�`p�wh�p������h��G��r��=�HDT*PRRr��ӧOc޼y?~�yWff&���#G�\p����i��s�N�=�@ ;��<�tnD��F������sk9""")�  *&�q�P����KD���h�oDcC��Ѐ���c��l0����ڊ������t7�h4"���P�j?�����#�hDmU5*Ϝ��DD�.>>eee�Z���71f�h�䄕�СC%tW�?x� ���qv��Fx-A:���ڵ��Q�	E|�$�d���E��V��ա���55����+M&L�U���:�'B�����(DEE!4���aA@dl£"QY^����+�DD�K�V�M�/$??˗/�}�ݧpd�5d��J����hmm����f�a�޽�����!�x��񸓠������jDD�ij�q�	���v(.1�����ՕU���A�vƻ�(�hlh@cC�JOh�i���BLl,�cc��(�����ޝ��������>DQ$u˲|������z�Gv$E��(
d���(�_�s�o���@�#A�$�ѠH�v�-�n�4�M6���z��-�,�"E��c������fDR���("r��L�Ț׼^������uuaavnc=?Q�������������o���l~��������&K�Ӻ	:���'�� � ��	�I����y��~��BU����03UQ�\Jbi1��b镕V_RK�E�_X ���
��������Ow H,ĐZZ��Y���@(B<����k��������M���q�\x��7��l���t�pX7FM.��
��4s=���T��Z;�������EDD���p�op^�5��+J��"b���⨔��ڱr�,��,�O�@�e��a��#��k�d]�eD��`af�#���6����Cɿ����U	: |�3��Mз��ѣځro��]�[k?^�r�O���h��݈�[n��T�[M�c1�;�,EQ���� �2z�a���!b���ۃ=��!������k��c�\.�A,--my��>�'�|�ӧO�|e���oj���(�˺��TUŵk����~����F5����յW�]m2���_��f+�e�����F5����)���X��d�½�AO(d�!s��>x�]���ω�����k&��j��w�1�Z�̙3���(ktŕJ�m��_�vu#A_]�n���f�� ��^\�r��0DD��y�>��f�ƞ��rss���b���U�9�� 6?���<<^/�184����K���������s�;u$�χ��.�h�Ny��w1>>�C��|e���z�D4'�k%���� ' 4�(ˍ~����l6��ω��a�$�w�C{F-��g�iܻu�>��߾���D�l��ُp��u,'[�K����AC���]""�����c���+_���W�zz���I��ܹ�|����>����8��ɮ_�εxDD��Á�{�m���T2�W���s�1���>�FUU���q��K���E��̴|-��;�����r�[zDD�xu����������"���z�r���7on�����KX� \���v""����Þ}cp{[�ʬ�*�Q\:wW>���X�e�B[[Y^Ɲ��p�7g1=9��b������^�֚�@D�S�����
������x5���
:�L��i	�� z�^\��qDDT��pC�{Z7��i��������Աu
�V>�ǃ{�q�׿��㉖%�,�oh�C��$�L�#"ڡ���\.����ַ��K�|���h����fxz?���7���?	(�˸u�V!��h7�d##���Hn�&�?:�[׮#�͚�#�R	���[��w�����s��vJ�$�*z*�·��-��u����M�oܸQ����*z�	��q�۷o�.�'""��p:1�o�@WK��ļ��%��~���i�k�]��2L�'"کp8��Cǿ�ۿ�9��=���޽{��hF�.�����NDDz�F��¡�>g���2�^���y�*
��>>w�X�����v���?0��DD"ɲ���^��������g��5<:] [�]ژ�V�F�^ ��^\�q����.�0<6j�z�b!���o�Ӌ#��d��|�Lׯ\��O?5��$a`x!�["�v����ͦy��_�j��r"�� 7n���� ��s[h4A?��ן�VB���!I����*�?�ų�03m��\d���>9��7w}��z#���8"j[6�Mw��{���?���Wd>Q����Vw@;��u4v�l$��q[""�D�$�"��k���+�>�p���t;.j-UU�dr�Z�������Ȳy���D����}�����&^��DU�����W�:��٭4�WD�^�d���v9I��?<��`дsV*<�?��_BzeŴ��s9\�r7�\E�`�`#�ߏὣ�u�D�����p 
i���p�����NT��S_���K ^Y{q�6�ۉ�h�$I�3b���D,��?:���	��Ӗc1|��y�E������`xt��ZN""���rMUՎ���M�o�>�歪b���|��� 6-p��s""V������o����w����+(�m_hg��2�޺��W��T,�rN�ǃa�NDm���K{[���G���3��c�j�p�^�m�`_��m$A_��E��;w�*u"Y�14�^�ϔ󭤖�ɹ���2�|�9��t�<M���t�V�d�NDm���O�X�P����m��<z	z�n߾]�_w�{�	����>11�L&S�W�����l6��­�fKU��Ǹ����rOsjR�Xč+W1~�.��a�v��c{�p:?�(�`n�[��7��M�;��MoiR��t:����ň�∈����(\n�-ID)����x��ך�ѩ'�|�c�Lx�cw80<���t"j+���������&^�9D��59�T�:�zt�Sk/8 ��h�Zkkwy������Z���L,~.�]��4>9��y��ew:1�w6��DDF�D"��~����\t�^�3��՜z[�&�'��IXA'"ڝ$I��Ȱ)m�3�Ӹr�RG�ё5T*ܺv��3�F��tbx�(��Q[�e�HD��͛7���wA&�xf����z�Wo�����b>��ʈ��c��>��R��΍���N���5czj
�?�l��w�˅��QHr#3z��Z����$i����;��x"נ���8��WN����B(�����(��]���ʹ����X(��O0?;k�y�j-%�|�cd���1<�G�����
�N'�������{w��5�%�ŽT*���o(8Y���KХ��޽{^��p_/�����ȤӸ|�c�,/z"-�\�/~�d"a�y�^/��������m���*��o�x5��� ����x�)��SO�.xa�����F�����X D06�K�	\���ͩ���2�}z3�ӆ�� �3%���
�~?|>������H�P�,�+� p���'QG�]O�~�zO#+�DD����C����瘝�����\>E���*�߾���g�#at�h��Y�^=���{����Wc�kЁ�������;�$�/���(Ju=u,�˅��C�p�O�����Uu����p��m���~�>ہ�h'zzz�t:5���?�J���WdC*����~w�6���M�٧����f��8""j6�C{F 8mz���s�Y��twn�4�!�$�h.�ۘ�DD;$Izu��D�Q�����Wd#֠g2D�э7������*�$ah��:O�wDܽ������n]�ՠm�d��{F s�t"����^݇�_��WL�cl��金���Aq��Fփ�,r'"����1&�����ۘ��2&>�A��v�
*�J�;�dw"�$�͆����K�.�&^�x�%��9��> �ӁXA'"�l�`�==�WUܽu��[���H2����נ(C�{�>�D"��&"ک��~��_���M�c��UЁ ���o�������:���Fd@���N<�s33��'2C2���+�kwE���94�����r���[����c��ϛxEb��2��]��]��^�O$���M^Y�,�6l(ܣ�q<�d[;u���"n߸a��8IB�����DD;���Z�X�w��]�F,�Z����L&7����'���ڏ��CDԱ����0h(��G�z<aHl�V��/���ۆ�.�l�zt"��@  �Μ�o��(4��hF���ު\�z��O�%]���ÇM_YWw���.CbOON������4;3�q���<����5""j��ά�'O����3�j�1�� �=�x!�y���%�2���^LLN4}ADDdM��~�v�������}v_Qg�NM��Ĥ!���<>�!�����u�����7L�q�Z�<�K��"������W�*�'"��00<I��|%���7o�F��b��#6� >�$a`x������l6�B!����>nݺe�Y_M. 0��Y��������Ď.����%��k�~��\7�\A�b�VTDV��*�ܸ���!@B���l�A""����|�;&]I{x��q�[�m�u%�KKK��爈��y�^����V�eܸr�bQxl"+S7�\E.���Kgk#""���nt�̯��~�������������Z��NЕ�}�����ڔ,��DO�VUܼz�tZl\�6Q*�p��5T�`�;8 ;�^#"���d������1�j���#]i���i�;t"����5�F���,%����l:�;7o
�~M�e��JD��`������E�I����Z܏���x�	:Q'p�����4+��g�X�}��?����_�_x\"�fH��[E�u�Ξ=k�Y[MN}L�sZ	� ���`���=I��?4(<n.��ݛ7��%jg�Ǒ\Z�op�,~�"�fD"H:K��u�5#���a [>�����������u����v�Y�Tp��5�XsK��TU��k�Q,�Ƶ��o3=���,��`P���ﾋh4j�5��v�-vE۲�}�=�� ���*""j	�ÁP�vZ�����P8"�b�o���u��6`�D"�f�m�V*���}�ī����Yd�w�h AWpx�ǉ�	.�'"js���bc�󘛙���$Kx2!x=�$�w�_�����,~������ַP*�L�"kRU���(3�6��nM������_����	,U,�q���1�:գ��J	��r{�7:Y�ް���Y�����Wc]O�<�x!��V��*��xzzZ�E�y$IBDtk�
ܽu�OÉꤪ*�ܼE����āqDd�p6�M��7��M�ƺjr�t��� Q&�DD��.�kU��&��ǅ�$�t�L�?�f��'����,#���ч~���q�Țjr���"�*A����t"��$�2��L���&D�Etj
�DBh̞H�ChL"�f赹������&^�5���n�no^e��������=#a��vqU����PE\L�]���;B[�%IF�_�DD�r������<�O��O�~y���3m�	z>�GB�^""2��nGO8$4��LK��@�#�l�����������HD����~򓟘x5�1c�X,�B����:t�z@�X#"j?=�H���Q�b�s��SH���(�^�b""������ӽ���DWU3���U�I�%Np'"jgv�����ܽ���҈DQUuu�B�EoW܂B5J�$�B�|?��O��ۅ�������������/-.b~nNX<"�S)�D�Bc�XE'"�ks�T*��h��XOU���^�[���[�2�X#"j+v����������GD��?@�\�����ND-��x���4������g��j�Jm��~g�
:Q{�	�Iof:�t:-,m(�J�z$v`��DdzU�Ǐ�����Wc-59vU�<��We�Q��WDDd�Á�q��J���
�GDϚ��B>�o��Ή�D�Z�P6�M��n�E�*�M�G�~PU���]����O>z�R�(,=KQ<�CB0���Q�,���G���ﾋX,f�mϬ��fggkϵg��}�`"�@�7fDDmA�e�=��r����SV����G*������������b����G&^�u�E�R��o�$�
F�~d����}t�!봒5j��]=���l��[N"I�u�9""2���Ggp巿�m��Z�r�M98�l�	:Q��i#kT.���쬰xD��d"��Ғ�x�`7dY�v�DD�Ы�߽{�ϟ7�j��&��IХ��:t"������t��ś|�شuXD����a�d��C#����!�����~`��XGU�-�A_��b�^��ke�e��g���%R�$����x�PH�Ƙ��hv�A�9?��Q(L�"k�ɵ5t�����Y�����o��#VωZH�Zt���OܿDD���}ii	?��OL�mf������ؔ�oN� ���d�NDd}��  �@���0?;'&5%�L"%p-zW�[X,"�fݝ%�2ͽR��ّT�k;���؜�W-N_X`�;��I���nq7�ѩ)Vω,��䔰X��.��va񈈚��Y���CB��f�0A6���[��(��6�'"�j^�_؍w�\�ltFH,"ڙ�X�lVL0IBW  &Q���b������0�j�f����E��b���D"�R�d¥Q�����F�(����Q�TU���a�8͝�Z�������;�x5[3��^,�T��i�
�����NDdm6��_L0UET`2@D;7��,�X�t��ֹ1&"2�^��?ly���t�&�V�������v""ktw{��Ő���""1*�
f�Qa�DΫ "jFOO��R������6�j�efx&��_�a#A�6�l��""��t	�5�dZX,"gf:
���tqOt"j)���׫y��w�5�j�ev���]B�ڏ�+�}[~���,��p��ӮZ��ć�D���f�J��'���p���!Ԟ��_�b�*��̮��ŷ��oJ�K�Y#"���@@����n�Fda"wW�4w"j5�6�t:�[�n�x5��~8�T� ��
� ��&[܉(:��    IDAT���/�&[�g�������Q�Â�m�D�bn��C��ŋM��j-����i�e-AX��[܉��i���-$�R"��pDW�T�07'$��f���i�D�Z>�O�X+t�נ�$�N ��F�޷����9WEDD�wu	ko�c���-��]ցCD�$��&^I5�
��G[�� ��t""k5�]Q*�o���,+�L���������!"j�^�~��,//�x5Z\A��{&AW�Tʤ�""�zɲ,l
s"���I�DԘ����8v��SH,"�fx�^͊��(��OL��U����<�����uO&��?= "��y|�Hu�OD��;��b��Z�f���3O�Um�f.*�
VVV6��)AWл�.ןY��'�ZU�cq!���"�ܽ:�DDf��8�"�Q;`T�ފ�t�?'"�&�_�M�b|QضMDdQs#<>��R""3XqP\+����ޛt	��w�ɤ�EDD�s8��֍.�8���bB�H���yDD��K�011a��<Պ
zM�6*�=k�����kIUW�Q�YN&�u����!"j���,˚�ϟ?o�լjE�*��6�����t�ԋ""�퉪ve2i
!���\�� )h)"+�D�J�$�Vѭ��UA�)�k$�&�DDV��z��I�9���%�uy<��+""��%��Ν3�JV���^�{W%��k�ŝ��Z�v;���X�n5D.Qq�\�b5���ޝ�ڵk�wv�b�^�	:�E���(��8����Y�Y!���ND��WA/����OL��ִ��<�XO�} �G3A'"���-$N*��}:LD�!%h���3DDͰ���8f�Co�=RM�����i��""�U�b���3�m���0A'�ֲҠ8����M�� t""+�$	.A��TJH"j�TR���n�C�|"�f�C?w�TU5�ZZ��ڪ�3t��Y���D<�U��u�l&�R�($�S�@"�f�U�1>>nڵX`H�����\��,g3i�K%!����V=ps�9ɝ�Z����f�i7s���l��l�zu�^.����M�(""�&j$Q-�Dd�~�����U֡�bz6��=oP�����d915G����ʲ�8Dd+�b~���Q�m��,��⮪jm޵�� �zNDd1NA� %�$AC}N�a�!"�z�U�o߾��I3tZ� 
���^��LЉ��C�e��b&,���'"k(
B�JH��*:�����L�E�ŋM���ο�F&�59�G�����d�DD�B��w��ϣ\.�<Y��oLЉ��l6�:;J���ު�*W��x�^��NDd�SH��u�-��6���CD�,�u�f�+�l_ib�-�DDVe���iuOD�"l�C��@"�f�C�x�)���M\��
:�U9�b֟�CQG�f�B���[CD�,�
z*��͛7�KVй���:D�����#r9!q&�D�Z.�K�s�7�����`�
��
:���4���'"k����8����VkD�rzU�>����[��.q:�e	ܤ�����C������oI��f�y"��K���_~~�l��w""˱��$y�q
�T6"�&Q�Dͼ "j�^��F199i������ŝ��b삪Y��]'�dyAKXd�t"j-��Y�.N�={���[$A�� �w�/����<���P`�N�����ND�&I��vkF�CoU�^(>�����`��uDDd��=�KE�?6D��ʂ~�e;t"j=�6w�'��*A�T*�_:d 6��DD�"6��ן�l�����յCD�z	��[��H$;�Et[U��(�a'&"����Y.q�QG�;�w"��߯����s��vnK&謠Y����2+�DM�2&�Dd�,���h7rz���"9t""+u�\*q�Q'��	:Y�^�����-�����NDdIb���N��J��y�ID���ҥK�mު�fP;+�DDV$�b���+QgS����=LDd&��P(�ҥK���XԞ�Ѳw��Y��?��
�CD�$�ލt"����˥yܨ6w���3A'"�"Q��:Qg���9Y�^ݨAq��NDD�DUЙ�u4UU�$�[܉�B�KЍ(@X$A�8""+�EU���N��DܿqHY�^��L&q��-��d�;+�DDV�
:Շ��D�i�n7�v��q#֡[��nc?Qc�*Q���9u"��CoU�^�LI��?v�DD֠���Nb�*Q�q��*<Y�^���_�Z��Z���t
�e �5u�������|�&3��+Q�q��iDd5z	���4&''���\.k32A�y�Z��_	t""k5ۍ	:Qg��(� �(^�W�߸_��WB�W,5����W4Q��ŝ��!�![܉�j$I����<.:AoU��H���ȊDU�d�	:Q'��t"����.�c�RA�Iй��Ȓ�-��!q�Ț��!j��U�DdAz��>|���)a�jՐ8�����=1�fw0A'�d�SHEп9DD"��~�U�4�V%�-YC�,�f�������g�NDV��:�?�PعXA'""M��!q't�N&�KF�CA""����E�C/�JVWf�NDdA��Q=D���ZVCD$�ޠ��ɓ';>G>��=nd��w"�6 l:��u4at&�DdQ>���u�Lзjq_o�5	���vF�zP��%$Y��%�w�R�n�$"j%Y���z5��hs�.A7��}�j�1�@��hgDU�\n��8DdMn�GH�A'"+3z?�VV�ݮ�{�� �~�7rDD�P)��
�����ԗ�Z��s�7���������#��(�^�n�}TM��d�^�j�""��QU��>�%I�����#I�$����(�����(F�C�KЍ�^��gYA'"������m'�LN���G&�DduF�Coe��[A�M�u��E!qD�Q%"ku���v"jzm�~��b��Ž���"+Ce��Ȋ�%17��'�DԾ��I��0���Hz	��{�033�tl�Vй���:ʂn�}~��8Dd->�_H�����DDF��|��읬C�L�kЉ���T�.�/�&�����%�w�\b���O�e�|�E���C�Z}=Ag���:����8�6�MH,"�Q�b�	:��֡[h�{N��
:�U*TDo�$xu�8Q��;b�PT�BA��@""��u޽{��u��]�t""K+
�qUi#"k�t�\.AU!�������u�g�6�B-�Yn�FDda�*[]�0"j?~A����R""�1j�����d +k�8H���ZD�Ct��!"k����f{;��u���/��Y��9��
zM�,H��r8ls'"�Q-��@�u�@w��8%A��̲�:����c�r9�cF&��g�&�t@����X( ���8�$�+pED�jn�.A�E=$"2�v����_6S�����-60A'"�2EQtۮ���Qk�joW��BDd��֡���lՐ�-r� �͇����r����סu���=��AСCDd��NW����p�V��JЫ*�GDd-�����F{��O"%"�u��I�s��m!"2�^Q9��޽{ųZ=���t""k)�.i����:t�6�t�����v���!"2����~�h�"����〔Ƈ���Ŋ�"*岐X�HXH"j�P8��WTU�=�#"2�$I���Fס���^�C ��/ &�DDV$�F�'�����"!!q��"E����֡��D�R�;V�*�z	�z��c�;�ՈJл��a�ۅ�""sI������l��ۉ������$._�\w��U�}uTй���z��LK��Dm�����)$V.����U<���F��-2$�-�DD�"��	[���CD���
���*�i&�D���r������;�%Z��ծv�����AA{k�Xٌ��H_��O������B��s9�?'������={�t��8�{,#�jr�%`�����nOO�a@DD��	�x��v���""s��~x}>!��uްY�ޠ�b��_��Wu�iU��^v8�%��F�
񦍈Ȋ2�4���%�GD��;�ԍCD�jN�n�[������nCUU�]o����*�ˈ��Ǫ�
:[����R��P3�=�����Ho��8J��B� $��U��I�����lF�/ɲ�����o- [$�6���∈,J�`'�ÁvL�����]v2+i���V""�Ir�ܿ�=���v�ԍJЃ�`m�y`�x����,"��",V�Р�XDd������ea��������&�?���u���������
���#GDdM�|ł���޾>��C���$I��+���� ���B�����jl��WA�$ɰmֶK��u>LDD!��.�2�YE'��P$�K{ R#�i��Qg�[����T*io�������m��&� XA'"��̊�6���aa��H��aq��+lo'���}ee�ϟ�<�WA7r�{M��ӽz6?��j��t""�*��(�Bb��~t�<u&��q8���
��T*LY������<����L�X6��<fd=���r}ɹ�՛lq'"�6���YE'����!ak���ۉ��鵹�������D[�׋�gT��B'""�ZI��6B�\�� ��Y�$I�3",�r2%,��%�7o����Ė�ZUA�J�խ�M�H$b؅���E�s�Pa�ٸ��b�����x�Ī�K�qz;u�@ ��u�UEO��`��fk�-tѵ����""CdElxt��O���1#{G��ZN.����:��fCWW�����{o���ɤnL�l��1���'k?D"C/���v.���R��r��g�,�;D��D↨����'Q'ћ���n�޼t��^��|=ߜ�od��6w""�SE�k{V숨y{��
���f���@Ddu�`P�X�X����g�oE����W۹�_A��ND�D������C��<^/"��V�Vωhq:������jz+�-r�-+�3 �{%��Y_.�E�Po��~a���q��m��T*H�!"jzm���?��J��@$�%h�^0��%""���bBX�@0�*:Q�x}>��l��:%KPEX<"�v����b1\�p����e����IU��vd�zi���DDd}+��3O�wb����bQ�����GD�����n�<��;�T�n���ꇱӛ_�&��YA'"j��"�X��;�P�Ut"3y�~�	��ZI&Q.���#"j'zU����U�E-���ճ��M����T"��x߁�b���	��'>�#"j75[�U�F��裏�_[`�N�.��NDԎ*�
Vt��4����������@w7z���w�2�ya��M �M����S�J:�Fz��;Q�k�u����a�.����K&� qEt�?t�v�N"2��#�q�sVωhד$IwO�w�y�J����IНNgm�_7A��M�k�����yd��Tr���3�WX<"zV�� �t�J6���!íՈ�t�����p��Y,,,h~�f�A��hM___m\��������/�����X�	]�>:6��%,m�e�����X��GDԮ�ks���w����f:#.###�o=���6A����2YX�P@z%���d�۱OpAD���������!���OD��$Iҭ��ۿ�&''5��ܻ&�^P��`�Ņ�U��a&�DD�&[EF0�� �ǃ�}���L���#"jwz	���"���h7,A�α��*A_�+�DD�(��	x��#G$���ݾ����s"�Z]]]���o��<fR�{	������-��B��^���Ƅ�#�������9ѳ$IB��oMiqW�I�e&�DD��� �����'4&�ncw8p��sBc�YVω�4D"���gT}hhh��`������?����kq!EQ�œd�}^X<����s��p:�TU�����%"��\.�@S�-���n~��`���]��e$Ŷ�{z0<�GhL��"c`H��+�e�y�1��:M3Ut��-�:�ȭ�J�'�t�Q�X�/�\,
�y�C���Bcu:�Á#Ǐ�����`1���C���Z�%I2�Ž&�.����V	z�� DD�FTUE"����e��p�S݉p��18�K.��(�J���h��$	���u��rA�>Q}�f��	 ���h�]m��^�DDmm%��BNl��+�����$�TC#È��cX�r��TbIhL"�N���W���F���o�h%�*���g��3UU�0;+t�5 C0���x<xN��v ��/ID��l6���Q�ҷ�b�J�e�_�q߾}�/����V��Z\m�$}��]�N!�2��<��t�+i�����$"����k��?C�e����Zƽ-ϯ��;k?�X!!"j{�1��U�.��pܐuZD�������>zE��ܜИDD��$I� �v��V�F����ٽ���M�Vщ�:��(�͊���B�w��D�lh���n� 	��&�G�ٲ�>66���C�;66V�֖	�V�� + �����O?umDD�"��jk�����V�������8t��𸅜KU��v!�ӉÇcyy�t.�>�o�����)z/���sZ	�
��� �o�t"�N������M�9v��Yqq�ڌ����' 	ކpmأ*x�#�n���ܨ��jr�[Z������z0��u�r�����6�'^zQs]Q�[
��x��^��Qȋ�.���̳���iխ���]��t"�β�J2������Sb��Dm��ѣ�l=X�呈Ņ�%""�T�A��I�7-Z���8GDDmnaf�bQx�� �?&<.���;x�C���*���hTx\""2Owww��h��>[W�l9u���ژ�(���X��70�}�KdECCػߘn���J<H#""�lё�T�!��ڋ��y""��l�D�{��Ǡ�LYI(��cG��YY�r2eHl""2OM.�0��Y��`|���ޱ�^Y��BE��O>�<z���M�j��n;u�$	�])��03+<.��&��@�����M��YA'"�L��bv:
�R\�p���F��&j!W^x�E�l6C��>��b��$����]g�;���*7��m x��\����2b�r�
���"�N'\.�^/��0��!"2P�X���G� ����$��ɓ�q�*��b�����ŉ�_�ݠ{����!����|��x!��g�t���}}}�BH\�X*�0??�X,E����ed�Y,--aff�`CCCp����ODD2+i$�q��vK��c�N�����J&��'2���Ʃ�_���4$~zy�Ē!����|�H�v��U��۵��|�СCM^ֳ��<�ܹ����g��Z��bii	w�����T&��#�I�f�ᅗ^Dw0hH|"��=�z�4\�!�םu�-:�w��?_{QU�߁l6�{��T*5�=EQ�F�����""2������A����e��q��
��Od�ߏ�Μ�۠�\�T0�dzۢ���}����K�����^*�p��}���c,//c||�I:��Nl6��x��^C����WN��2h���b~f���u��U%�W����	��Q�QA����Xg2<|����DD(�󘟎�+�6�p�$��O$Jw0�S�_6l  ���YY1,>�NU]�oo�I��
���؎��%�I$ZYY����DD��t���N I8r����w�������/�f�n�n�R�R��u��n���n��)��RO��z�/���C���m�o������DD�!�H;QZ������БÐ$�������(��:i�>� �]1�!�ԡC� �U)��
:p@~�E�m�L�L���ngjj
E��""2D|~������Q;y��d���$�Б#8x�0`�C�b>��h�K���:X�.h9 ��}������I��Ƿ�P�*�
�Ѩa�v3UU1�A!����;��é�/��rz"-6��O����C�S.�03��ۉ�:\̀�XͭuՓ�@�
0    IDAT�J���^���ic��%"��E�������������g^AW `�y�j�=�x��T�%D'&w����F��&��F�-�跕����333����h��T*�N���<�t�z�5�H�_{�.cU�eD'��rODDD�%�2<��\��{uƿ�����ž}������>�������?�����Nu�f�����S)�13�e�I�q��Q<�X���1:6�/�2t5 P3SO�EDDְ�~x���o]���f�$��S؎;V�����?�S��?�#���/7�= XX�4T""#�K%D'�P1�E�h/��
�������p��K/b�s��.�NM��7v�Y����7�,Bp�����Փ;���-���$�ݎ���e���w��/--q�
��JŢiI��+�ӯ����~��E�C�����*B����RUs���gs�������&g������U|��c#tUUJ�O�:����@�@ _�����.���:�L6�""j\�P@tr��vw`��y��	;yv����Qg�$	c����2�+CQ�>�F6m�6�DDd]U9����~��]�H�<O�؊�bC{|ִ�K_��z뭺�?1���VLOL�T,n�az����믡�'h���sx}>�����oxK; (�
f&����B�����xcS.��F&���l�#�u4:�t���_��_4cee���Q��֤�5������ӧ���A��mI����=8����}�ڎ��ډ�v��6�m�[�$�w��c��ͽ�}dd�����/bpp���R���z""ڙ�$ݴ!X������7^GO(d�9����~���i:r�l��T�eD'&9��h��
O����$�
�O�OZ砸r����d���������:t""s���<����]z�^�|�e>z�k�i�,��w� N��A�C�
<y<��Ԉ�v�cG���c5��Kc�����[Aod�9 5��~��o(ס�Oy�ڛ^^��âH���0�|���w^���P���:���Ʉ��k��,�'&M�HDD�VUAW�ooM�e\Z�qxx�:�
����rm���>���>~]�L�J��s�Ω����(����u�\8z��t��ݦ��Z��v����p����zM=wzyyu�A�w�z�H��+\�����sa�G�n��F+�Z-��H���j�qTUe�����ffL?o ؍�Μ���'�v�M??��f�a���y���� �D�љ��w���3��Jl���h�>`z��u�Cot�nQg��/~��b�ND�Z��f&��6�M�c��-ٞ�:7ҁE�A�$�ك��zc��6n��b>:���<�s""ZW�#O�o����Os~�_|q�7��+�3\�K_�RC�����G���Ų��Z48�f�c���x���`dt�۲u I�004�3�y��?��i�5T�eLONb�� ""�q�ԩ�*�5����T$�]�����p8�'h�f(�i;q����Sw�r��L&�����H�R���������r����x��oatl��z�$	���8���8r�������9<y��,�8'"�jN��z���4��;����\.9rD���%�ft�+J������i(�܉��AQ�MG�o]K������ᵷ>���Q����Պ� μ�:��<��ײkI..bzb��-d��hw8v��՝]�$���g�۵�;l=�K�0A'"js������0�q��8t�0���gq��a�8L�rlv;FFG��[o����-M̕J��å��]Y_Mn��v�1�I�+ش���S:[A�/|��x<u���r(�`�#i��Vۄs�#f���~�>��qt-�<^/=o|�8h��'�BO&&[�<����GMn|@�Sr���l;~�X]/˲�~�v��$���8==�{����_�~��}��d�z/:""j�r����)C!��z����$I��?8�T2��hs����$�,#�ۋ��!�B��wa�
$�X\�q�,mK�e�8qb����v��}S/} ��}����C�;���6�}{�.�/~�%�KKKLЉ�,HUU,-."�Nc`xN��w��q��#X��13=���D�/�#y}>apx�%�صT�e,��"�N��R���M:t~��[�&��p���z	���;A������2:m�_�җ����u_l&�A�P����;DDd�b��'�'��GwO`��,���ߏ��~d3���"6��,w��ۍ��~����zK
���X�����	""j@�������iv���O�^l���@EDUUܺuK�3���x���	�Vщ�ȺTUEln3SS(��P�,^��ęϼ�W�xc��[���t��n�ٻ/�z���~�rɹR�`afs�Q&�DD԰OU%� 4u3�lP�Hx ^z�%ݏ62� nܸ��_]�3_���駟�sii	]�/��`��c�z#�B�X��������؁Ȧ�X�ǑX\Dj)�9�e��$	��n�"a��at�-��e%�B|~��;Q{;y��Ƌ�\�)�'�2~ }}}����m4A�~����y���W�Wun�f�ls'"j�� >����2���r7�w�,^�^�{��P�T�ZZBbq����l����AO8��p=����o1�R.��03�eDD�#����D"o�ͭ?v��簺� ^~�e���{[~�������~f߾}8}�4.]�Tw\Vщ��K!����It�� ��l����4�l6�"�������XN-#�Lbey��%�;�B+I�>��ݫC�zz�n�o}+����%,.���@DD;V��������$AO��4 �y�f�n���t:�w��ud2�|>�Ͻ���LЉ�:���H&H�� ����Un�۟V�C V��Ȭ� ���L:�L:�t:�b���+��p8��������ߏ�@dٺK��2��P��[})DD�!^=��旗 4�F���3�Cz���9��߹��;A/����O��}N�s����˿l��=��74������\*an:
�'�ށ�<��o�$I��<`(�JȬ��ϭ����r��r(��(
����r���xV��������C���
���u	%IN�>���j�ܴ�%�2>��� "���ۇG�m�Q����$�s��m���ٳ���*.\���`ii	���u����%��azb]� B}��;���q8�z �<sLUU�J%��E�J�՟���\���&��r	 �(*���m�����vH� Ilv;�N�����f7u�>�RA"G�{��:�P(��vo�\�bu�7�ZE�JзkW�U�:t`u�{#	z<g�ND��TU�r*���
��z��L2%I�����l���U]����mӈ�� gΜ��2��?��}M�z&}�3��z���y:�|]m}o��6���)�XYY���DDd]�� ����$bq�"@U��Lb��C��晜��jr�_��p�������ӧ5�U�$	^����x>��s###�Ul""�J��D,�I&��Zb>?3�R����!"��p8p�ԩ�7����"t����^/�=���F��ϝ;W���������d�Oԉ�:PeS��_���;��"�X���&�DDd�^x�����g�%"A�������*F�C��?����ZW���u�J��ŅL�?@|n�:w��Q)��_�����昘��j��\�iL	z��k/�֡����כ��A����^C���ND��EA2����G�}2�\6��K�*����c��C,.,�\.�����h��*N�x���؉y�����^Ьf;��&�޼y�L����ɟ�I�q��=�s�\C�!"����*2++�NLb����ˀ	��� ��l:���)L>x�d"�9DD�R�,����ja�X�w8x��5?�H�{�R��˗���o��oa�޽u�XE'"ڍ�榣xt�>b��(���֪ʥ�j�����z�l����DDDF�b@���{ ��^����T�F��/]�T��dY���7;�'�DD���(H-%����<z�Tb�,@U��R�NNab��j;ח�����?{w_Uu���ϐ9d"��1��@��*��*ʠ�� �u����,��j����:�j�S��U�jm{�U�e�@�<���#r!��9'����~�|��\�^�$�Yk��u�_��L���rҤI�f�5������c.\h����'""���PXP��)ؕKž2�]i�+{��ٶa�s���+n"""N8����pg�@w������3p��V����aF���t���s��'wx<��={,����4M*��(��eۆ����Eyi)����;P��u��uYi�>��7d������PwV�
t���7N:��'t�,]��u�VJJJ���W\�� ��Ք��Y���������2g'��K�ݺ(+-�`W.[��T���HD�8qb`��8X�f�^|�o�tb�:X��?��O��Μ9���dK�߽{���""ҳ��IeE�lߴ��6S��OE��·�4M���(ڽ��[��m�&��5��iW���D�O81��1�{\�Y��Ѽ�?f̘þon�=�����cccc-�����QSSc)FDDz���z��4�o۰�]۶S�{��4��{�}>U���#�m6��}%EE������t������?l�0����]��{�/���;vl��bbb,=��
:�u�]����vi]DD�0M���jJ���߹�m7�c���峯����jL�{����R^ZJa~>;�leۆ����Iq�^�*+��@DD�������z�>��U��� l�A�6�O?���AVt++� �bƌ����)**"++��o����e�uu���AiS�0�^/Q11DEGEtL������0M���������Z�jk���m?VDD���x�A������@�0��^�7�4���������m��ׯ���7�`�@7M��{����iy.����I]]uuu����=����m�������˅��]oBcc������������������P_��q���0N8!��s��	����.��l*����ða�شi�!�bbb�����#�m�ƞ={�ӧO��8��7n��{��۷o��f��H�`�&������S���2.��ǃ����vc�\�������0����Z��<p��3�&�飱��@A����_���H�1|�p��ӛ;�x��_���S�*�h�n��=66��:�_|���o)�n��9s�tx|}}=��Ť��Y�GDD$�|>��:t�����sZ\%~�-f��C��.����أ�ի־��ˉ\p�0�R����Z\%�?4վA�����G�Mjj�!C,=�N���zY�|�����j���,�%""""""�S�޽5jTsG@�L�)��m�M��M�2���і�B�ꫯ�����ȢE�,��k]DDDDDD��N���u�|��b�P軁/������� +�sMM��,'����-Ŕ��Q]]my.�~ZԴ���'T:���rܸq$&&2��6���~�V*7�tn��RL~~���DDDDDD��HLLd̘1��n���@�����x8��`�@�����~�mvv6ӧO�SRRBUUwވ�����H�7i�$�^o`��C5W(�m���Fk��Z�B�TRR�����V�t�M�c���l�%""""""�C�Z�i�uC"�:��K�'�x"QQQ�IJJ���u���J夓Nb	�b���g�`:�|111ב!���.�]�����1~��C�$''[z�[o�Eaa��t쬢���ښKDDDDDD"�	'�@lll`W��/`����6�^�zY:������^z�V2�f��?������rJJJl�'""""""��E�X��B]��Ɂ�קL�rH1n��m�/���iZN��rq��Z�������Y�����x�8qbs��|z���@�枔��1�sȐ޽{[z�x�]{��Ϙ1�q��Y����e��ݶ���s�q�ѫW��Wh��7Mz���SO9�����DGG[z��?l+�0X�r�市����l�)""""""��E��=�svE��<����N��:tZ���}���_m%t�Yg1e�K1>��]�vٚODDDDDD"����SNi�0������@���LMM���?dHZZ�aXz�C=d;�x��|%%%���ڞSDDDDDD������q��o�bޮ)��/�����8��Cx�^RRR,=��w��������N`޼y��rrrhll�5���������5�N������
t&����r
QQQ��۷������]w�e;�Gy����;���^w�������tSQQQ�m�[��5b6tU�~�6�^�z1aC����Z.�?��C>��[)��ۗ�n��r\aa!������5q�D�;\��Usw]�_�t�; ��vz��222,?��[o�u/:�M7��Ga9n�����."""""�ʹ�U7��Uswe�N�6��S�{Ȑ^�zg�_}���������x��'-���Ց��ckN	?���L�8����7]9��[bcc9餓Z���e�ѷ�~;>��S��>�l�̙c9������b[s������Hx�2e��ɮ�E�е:|��7Z;� ))���xK���oy�7l'��SO���n9.''���:�󊈈���HxhQ���ﮜ��t0�W�y�>@�~�,?��{率��VZ�{��G��������m�)""""""�!11���̍�λJ��4�"9�>@bb"�����a�^~�eۉ]v�e�v�i�����ٽ{��yEDDDDD�Y'�|r�u�&t��vp�@����8��s;��*�ʕ+mo97�_�����Z���ͥ���ּ""""""���W�֮���,s����۷�a���$''[z�;X�n��������O?m9�4M�m�f��:qFVV�{ls��KN��L�� � .��s�9���z��N�fϝ;��s�Z����f׮]����w޹��r(��p`{;8W���{�a�:066���<^x�N%���2h� �q����zMDDDDD$B��r��`��8U�����_8�Q�FvhVV�a��y�������^RR���/?E鰜�jkkm�-""""""]�c������jWs�@�w	�T�s�;����h���,=����g�y�vr S�N��o�����֭[1M�S󋈈���Hh��E� p(G�:��+��<�L���;833��*��?Lyy��iz���c��WUU���EDDDDD�Xtt4��zjs��o�^��,��ռu !!�ɓ'vhTT�{�����{����~~�����Mll���={�PZZک�EDDDDD$4N9��;\�moo��Y� ��7���M��V�	��ǩ������ȑ#y衇l�n߾����"""""":-j���s(��~���Nhs����Z^E/,,�瞳��~˗/g�����>������H��ӧcǎm�0X�\6M�/���@#�':@߾}-���]�����	B������/8p�����J���;5�������Ϲ�X[6 �8�z�q����<���ҧOK�����/�N�/55�7�x��k9�����������H�����v} �v(�¡@?h+��A�8��c����ak����^~ƍ��ի-Ǚ��Ν;;=�������t�����h�_8�M��(���|Z1s��6{<˫�۷o�>��\K?��9묳,Ǖ��QRR�DDDDDDĞ5g�C�$\
�:L~�o�zꩤ���ЧO˫�?��Om%ג��⥗^�_�~�cw����|�.99��S�6w���>.:��������;,�Ή�|��7o��b���t^y��n�����z'"""""��ӧ�o���c{;�S�[�?��f�j�8�~��i�A9,�o����s�=�����Cuuu��������gv���P:��~���̻λ    IDAT#��y��v�·�n�:�����׊;ѣG[�1M������ """"""�k�p����P�U������߳f�j7 ==��������{�;��ó�>��jK-i[+�ý�P*�
�������O\\��I^~�e{��I'�Ă,������8�.���p�����­@?�8����aq`}����c�޽��;�G}���4K1���59T8�~����RSS-��^WW�k��f;�֤���z�j�q�w禮�6������������7-��!�+��(�C�;�����r�,�m� K�,a���bL�d׮]A�EDDDDDD��7�����0;�/<t�=M/�p�������o��6m��X[\.�<���KKK)++j.""""""ҤEM���C��)\�:L��7&O�LVVV�			DGG[�$����;�8-Zd9n�Ν���|DDDDDDz���,&M���a�av8�_����Y��V�/���vCRSS-M���KMMM����.�}1.ׁҷ�_�7�[��L��7fΜIlll�V����w|��w��kCjj*+W������k�DDDDDD�$&&�i��3y��ש�M8���i������}��m���&>>���ZE���5j��������C�������HOs�y�ѫW��?q.���w���7.���]�fū��j+����n}�Q�q{��ѵk""""""A��U�/��;�J��{�F�*��!C8�������nh��������_�<�L�=�\K1�ij]DDDDD��ƏϰaÚ;j�p�:���+׼^/			�&��ok+��x�',�._\\LMMM�2��Z�Z�J��"�@?�ʵ)S��{�ZJJ��	^}�U|>����1l�0�-[f)�4M���B�������Hw����ĉ�;~J�	�a-
tp�<�3;r��m�yyy|��g�J�-��s�{��SRRBUUU�2�.������j	��EF���W�͘1��+�<����&�6���dV�Ze9N��""""""���ŵ�Z�5`�c	Y):�x��e�^�8����n�4�7�|���z{�u�UW]�СC-��۷����e$"""""��̜9��ۀZ2�EN��t�ځ}�s����vvprrr���v�ݻ�?��O�J�-^��+VX�۵kW��<s.���1�O�ұ,�
t0x��eVV��z�a����/��P݉�7w�\F�m)�������e$"""""�}�q���۷�#����U��;������y��m�o��VH�7s�\�{ｖ�rssC�������H�2������JŖH+�M�7�<�HƎ{��IIImn�o�������s�c�̙�7�RLee�V�EDDDDD�p�	'p�G6w<��%dC�� /�t�< �ο��].III���_��vba+W��WPP�lDDDDDD���a.���B$�Z~�o�)IV�����;���?��:�,�L�b)���L������������Ou�%dS$� ?*����W�^x<�?�����_~�S�uĚ5k,���W�������t��-<��������z	&?�79�/�a$''[z���sL3��*L�8�3�8�RLII	���!�HDDDDD$�deeq�i�5w�<�s,�N0B]��� L� ^����7<������`Æ���'�Xކnէ�~�ԩS-�dddп��$$A|>uuu466����t:""a�n7.����(K�
�H�������K��z�;LɶH.���+�����i�QVV������[�B��/�������_~���n��ѣG�rE��{LӤ�����2��˵�DDD�&**���z��Err�
v�����;��qqqM&/�b��Y��U�������8.�����ݻ��G���lٲ�~nt뭷Z���HQQQ��	?�����7߰u�V��ݫ�\DD�������b�o��7�|CNNuuw��H�4w����L\<�d>��:||�o̝;����V���Ю��F�z�N'؞��?��#GZ��aq�S�ٳ�������NGDDz ��Gaa!�}�yyy!?�HD�KHH`��ف]�|�P:A�:�������^��0��c���u��Q\\ܹ��a7�p�������n��ظq#;w����""��4��������-�05gΜ�h�s.�������o̟7?p��A�ns������Tr1w�\˹�ٳ'Dو8���������r�S�������?TVV:���������v} �ݡt��;�`���eRR�f�juX�^�������'�|2� ��Ʋh�"K1���ӧ�����ֲq�F��'""a����M�6QUU�t*"���ٳ�!mp�s�O�(��S�/�ƥ�/%::�Ձ}�����={�����w*��X�|9^��R�Vѥ;��|lٲEŹ������F6o�L}}�ө��x111̝37��O�g�Tݥ@�5�/���8���[���f�~�G����\~����b�̙�b����~�t999!��LDD�3���ٶm��i��x�f�"55��#��tݧ@������u� �0,����/t:��\w�u��766��;��PVV��ED$"����w�^��鱢���?o~`��'�d|ݩ@��_��Ӈ��;��a���\�~�?�p���>餓3f��ms�� 77��DDD:,//���t"=Ҍ3^p5X�X2!н
tx���q����x<�r�ݤ��[zpnnn���_{�������5�h���:tGDD"J}}�V�E��x�t���]�>r(���n�A�虙��s�9���Ȱ���j�*���׹��1g�222,�h]"�~��H��_"]o���dff6w�L�
��W����w�Ƣ��z(���|�xaa!<�@�;!::�����R̾}����	QF"���ب ""����u��H����+����iu��t������=�o߾�Wџ|�Iv��ѹ۱t��V��E��J$*//�4�Շ�""҃���;��H�q��|��^���9t��-�+�˯ &&�AvV�kjj����;�`[���ϬY�,��ݻW��Hĩ��t:��}L�k��Ʋp������Wϡ��f�i~�{�梋.ju`FF�aXz���������N%����566RRR�lDBC�f��H$��1��1gΜ����N7\=��[�| |�o,\�����CEEEY��4M/^LCCC��<��'r���[�),,Q6"����DDDB�����D�����������C�\w.���.��III̙3��a��������ox��g;�_;�-[fi|ee���������t
"""���B�Л?o>�z�j����]��g���������v|\�}�����v*��̙3���4K1:,N"���H��c"�����r��}��9�N����A�'$$$��������V�kKYY7�xc�S<���,X`)���X��"""""�\� �5es����Z�/���;��%�\r���A�~�,?���_�>�T�mY�x��C�tX������D�V��7uuW=�@��4����[���LBB���/Y��}��u*��>|8S�N����DDDDD$���*۷���n�g��&o�^x!���ou���-_��s�ΐnu_�d���UUU:,NDDDDD"R�~��1cFs��+�z��B=�@� ^���K��:,66���ˏ_�n��~�R<��3gZ�I��"""""��]~-QQQ�f=����_�)�a&/�g�y&#F�hu`ff&��і'X�x1����3<���(.���m�����DDDDD$Ҍ9�SO=�����f��b=�@����Aӡp����և�\0���sss�я~ԩgѢE�\�����(**
I.""""""�p��7�r\����̧����`���3f�&Mju`RR)))�'x饗x��W�gxC����O��m�""""")N>�d�9�����ݎ%䀞V�<��7~tݏp�ݭ0` ���K�.e۶m�<������PVV�<DDDDDD���v���e�]��S�㘞X�W^p?x�`�O���@��kk���}��?>��lŴi�,�վgϞ�� """""l\p����w =�j��X����߸z����ŵ:055���d�|���^��v���x<,^��RLYY���A�CDDDDD$X����ʫ����C�8�����o���2o޼�4h����k֬�O>����,^�8�ʁv���Ut	[,$55����ǀϱ��St�����7.�)iii��x<����|>.��R���m'�R߾}�5k����{�}�������Hg���3w����? 9���zr���Ut��U,Y|�C�RSSm��k�.�.]j;��,[���A|>{��j""""""�u�ҫ����7}��d>N��:����3f���#�<��A�Y�^���o�n�:{�bҤI�3�R̞={0M3h9������t�QG�y���a�+��
=�@w � .���o���C�n7����ay�뮻��7�N��k���������n���0n��-�\J�J\��dN�@:���c̘1�v�i����@߾}-ORYYɅ^HMM��,[�7o����b���."""""�;��=zts���4�}ޣ�@p� ��߼�����=����L,O���r�m��?����-��^[[KIIIP��#&&�eWT�ls(����Iu�a\:���6���l�n�剞z�)~����˲�e˖o)&???(s�������q��W�+��& 8[�#�
�f���, ++밃���8p��IL���+�d׮]������e�]f)���F��"""""�~��1����?o9�N�Q���z����/�fy��SSS{wz[����?>�����t�7��x,�����]t�r7\C��X��k0�O��������3�8����xo_�}�駬Y��z�-6�K.��RLMM�����[DDDDD��Ǝ�ԩS�;L��u*�p��%�E���7�x����].l��իW�駟�?�w�y������󃲂/"""""����M7��U���N��T�����ƑGɌ3����o�}��illd޼y�ݻ�z��:�(.��"K1tj^���袋6lXs��],�J�{������e$%%�зo_z��ey���\���N�~�w���ߚ={�PWWשyEDDDDDڒ��ʒ�K��~�P:aMz��1���HNN�G���ݠ��l�^����y��x�	�q�F���ٳ-��|>���:5������H[����/f����s��T�އ���ƴi�8����x<dgg�z��[n��>�����'::�RLQQUUU��WDDDDD�5cƌ���n�0y�ر�
��\�0�[o���+���Ȱ<UCCs���������,_���p���͵=������Hk�^/��v{�f.~�dN�Nz��1X�o2��s����EBB���v��������|�c���NRSS-Ŕ��QVVf{N��.��R����;� �mT���i�kc����n��ٖ�>���Y�zu�#%%����r�Ν;;}P������@ff&�/�<���s�1T����%� &&�o��ݠ��(lk�U�V��GيX�lC��SSSC~~��9EDDDDD�n��-�����>�AõKz������S�2y��v����IOO�<����K.aǎ�c��Á���r\AA555��8��S�4iRs��3��K(��@�(���o��-��ŵֿ��O�:����y��Q__o9`��ٌ;�R�i��?����o
�*��=N�iT�w�>n�7���˕W\�n���b�С��G��_��m��f9�ރ��G-�UTTPPP`kN�ٖ.YJ�>}�;n JK(¨@�����7o�<��nPtt�����q~���ي�<y2ӦM����Gee��9EDDDD�g>|8_|q`�G����T�[cb���x<�s�=�\��6&''ۺ�4M,X����-�<��Ӗ�|3M�m۶�ب3DDDDD�}n����+p�p-�:�S$R�n�FL�7F�ѡ�����g�~�
f͚ž}�,�4�{��r\mm��G����K9�裛;�68�P�R�n������ͥK�2`��v��`Ȑ!x�^�Snܸ�ٳg�Zվ���3f�帒���."""""m8p �-���5��T��S�����/&&����0��z�dggwhlK~�!+W����xx���mT���kk�^DDDDD�?����w�MTT���q�T�`ZK�}_a�1f�fΜ١���D233mM�f��~�m�q�<��r��9�m�Fuu��X�.��B�=����ǀ�;�P�3L�t:�H��7�P���J.�}{���P�M�(++�<iBB_~�%#G�������I����/-���z9ꨣ?����SSS�t"""��\����o߾����������a�@WB٤�Ω�``���s��wt88;;�V�k��8����/�Lbb��9���ٴi�cEDDDD����Ƿ�&�Qq�)*�;�cL��'N��3��P���aȐ!�����72�||>���aÆ���O[�����-[�X�SDDDDD��s�9�ɓ'7w�����&�+V�p:��g�)p)��1���{�v��(���(--�<�ƍ1M��O>�R�1�CNN��׿,�YWWGEE�����	TXX�]""�ð}��H$KNN汵������L@�.v�VЃc������xÍNKK#==���k֬��^���s�1i�$[sVTT�i�&��������@���RRR�;� �W�*Ѓ�-�㬳���N�p��HHH�<�i�\y啖Wã��x��Wm�[QQ��͛m��."""""���O�3�h�0�-��c	u3*Ѓ�i}��y�-����ڱP�`Ȑ!�������������~YYY��w�#::�� ���lܸQ[�EDDDDz�޽{sםwv��z���T�����������?�6y�^�j�и��fΜImm���	&�_��֜ UUUlذ���:[�"""""��.����;��V	�M*Ѓ�mL^�7&O�̴i�:ǀlM���s�5�X����y��l�	M��oذ�C�≈���H�9s&'Nl�0y	xӱ��)��
�I c����G***:GCCUUU�����IIIa	��&L�@MM��_-�	���HQQqqq����z��<:�]DD"�Nq��"++���������rqq>:�=贂�\	� ����s�=����=4��o棏>���p��ۚ���e�
m?CDDDDD����{�%..��ebpP�`Zݖ
������cǎe����̡q\|��lڴ�R�a���,X���~�i���Cnn��g�����Hx�;w.�w\s��3�K��S�J.nT��]{C��pxg�+))aڴi��Z����r�n�:.��2�s*((P�.""""�����z�Ձ][qq�S��*�C���@#4�=�r�J<O�����mM�a��Νk��r�>�|[�����өg�����H�s�ݬ\�2�Jf��ڦck�-:$.�vb���I ����7����_w���� >d.��͛������O��r��9s&�����/��<�_UU���$''c���H��C�DD$��8��]����:����!�9�QϠ�+�?`:�0��1|��W�޽�ÏHLL������%~���2�������ଳ΢������/�����"]ZR�.""�L�tW#G�dŽ+_�]��y�~p1mq������A�v�իVo�!���VӭZ�d���5k���c�u��.))a˖-��i�"""""Z���<p�����b0]��%T�w��1����ׯw�y���\.�f�v���fΜɮ]�,��p�����?  طo[�nU�.""""�n��6�l-�0    IDAT���;n�ϱ�z�]k-�q��s�9�Xz@TTC����]PP���ө���p����ӧO[� ����ܹ�v�����������9��3��<�P:=�
��ebp9P�����8p���$$$0`� [	|���\u�U�W�Ǐ���Ga+��;�l"""""�c���|�́]{�����]Hz�۳�H7���5����z-=$==���t[	�������0t�P��0z�h��(((�tH����������a��������L� `aQ��
tg�����#F�x�b�0` �����뮻��o~c+ ##�?����񶟱k�.���lǋ����H�-�f9�F�j�0yxϱ�z0�Nqq�/s���7��#�`Ȑ!DGG[����q�e���3�X��KKK�O�'N���;vPZZj;^DDDDD�?~<s����W���ҵT�;�]A4�о��$''[z���aذa��n�	�|>�/_�m��f9֯W�^��ly�D���ɶmۨ����������X�����+�;��`6�R�1*Н�on�7����=w�c��������m'��C�x�b���m����������ӧۊ��|lݺ���"""""b�a��w�{���G�KJT����1y�ߘ<y2��ͳ����$���g;�^x�3�8��;���Ѽ���zꩶ����زe>��V������t܂8餓����C��~*�Á�����/�f������Kjj��4>��&L����o+>::���z���~����ر�V������t̘1c�z�Ձ];0�ʩ|��
��P��E@4�W��Z~`РA����Nd��͌7�W_}�V|bb"��>#F��_\\LA�ns	���T֬^x�U=s��T����ap��ѧO����:��r1t�P������`Μ9,Y����:��iii|��<������:�]DDDD$�\.�V��O�>͝7�;��Dzxy��w? 7n�_~��x�^�����T2?��Ϙ4i[�l�ۯ_?���?�?�۶m��F�G�����ˢ�1a��7��JGZ�=�����8P/Y�����[~P\\Ç'**�S	}��W{챼��˖c�<�H>��[[��'���8��;v,W^ye`�f9���Nz�)�`PM�PV�ZMzz�����0|�p���;�Pyy9�]v��ͳ��|̘1���K������&''�r������4KKKc��5������|��iI+T���o�GOMM�5�Y~ **��Ç��^y�F����o)n֬Y�Z��֜EEE��~���n7>� iii͝ˁ�KJKz�z���ǌ��%Km=���2|�p[�·���˹���ٳ)..�pܝw��ܹsm͙�����EDDDDlX~�r�=����ߢ��Ö
�p�bp�R�2q�D{���{fffPR{�75j��N������s[w��}t�N���������{��Lzx��?z%4���w?��ٶ�������m��R~~>�>�/������111���[deeY�K����tܠA�Xq����+��w^�`Z���o=������Ѓu��4�:�N��`�&/���G���?lw|VVo�����늊�(,,�������H�����ck#!!���鶨;��t�
���kL��7���U�;�
ǈ#��^:��;8��3;�n�رcy��Gmͳs�N�'ɋ������ap���0hР�N�G�WKJ:Lz�pq3�9e�.���N=��v3t�P��������M=zt��/_��/����M�d۶mTUU�MQDDDD��Z�h1��rJ`ןpq�S��5*�#G���ѷ�;�.YʤI�:����̠ܗ����ә?~�W����:���}>[�l����3i�����t+�'O��+��ځ������"葥�Y@4wߚ�:uh�_||<G}4����~��o~�F�ɛo���?OJJ��^���@]][�n�4�Φ)r��N� ""b�˥�%|8�U+W�wY���q� �S%���%�F\\�<����~���&;;���l<O���{�n.��"�=�\�n�z�??��X�v��gWTT�s��Φ(R�.""�,X?/�tV\\�>�h�C���XRb�{ŊN� �}�I�����=��>�((���%--���Zjjj���M�6��/����0a�A��ƍ��������*YUUETTT�N��TVV�<�X���A�}(b�a�Y���;����1v.+�K+���M���7�qh\ ���СC����*guu5��s�G�>�Ä_|���:��ssrr���u��(66��DDDl��1	W]u��zj`�Ǹ�թ|�sT�G�������t�R�N��IRSS9rdЮcظq#g�qӦM;�E=))��������3MS��E���D�S�M���i��r
��Zؕ����P���=����|���1bDP'�<8����5�'�|������y��m}]__�C�"PLL111N�!""b���>�}_�.6|�pV�X�C���k&@tt4k]K�>}�>QZZ#G�$)))h�,++���g�ر|��L�0��^z�ֽ�l߾=h�I�HKKs:�RSSu��8�w��<�����-���8����T�^��~#==�����ʤ��eذa2$�'���_�⤓N��.cʔ)�y睶�S\\L^^^���KOO�i�""Q��b�HG��z5�d�ǒ��Q��]���W�ͣ�>��+V�Z��F�AJJJОi�&/��2#F�`РA�s�9������޽{�������u�����SRSS���8�0��^F���&.V:����Y�N�N�2L������C��MJJ
���TTT�����ܪ�*�y����())��ܲ�2]�A())��A癈�Hx�x<6L���ˮ^ƅ^����gR��nB�t/�� �d�E�q�Yg�tR�jz��%^�~���4M�o߮��a��;""����D:���Ooy�r���ʡ�$�z�-��_�x���:�,]·�~������ɡ��&�suTVV���N�!PTT���DD$l�g
q��ѣy�����`"��%!��������%QTTĂ�(((�Ħi�{�n����4h���N�"�ػw/;v�p:��dddп�Ӑ(33�_��W�����|�~�`Z"*л��Ow߸q#�/����K&���c�Ν���v�|�1���������I�^]]MQQQQQ:ݵJJJؾ}{�|�#""=�adeeѷo_�S�(11�_x��C�6w�<�XRR*л;/����\{ݵ���uY
���#''�K�lOjj*���@ӊmJJ�����)..��������C�	�)�=Muu5۷o��J�U���3���<x0			N�"=����'�bܸq͝&���减�H������#`�����c��t�{��G~~>�w���y'::�Q�Fx���r���Brr2���m�iR]]Myy9eee�����kr�\y���Ǉ�ҭ���޽{)((�xDD�{�x<dddЧO`*�0�իV�<��c��CQ7��gH�h���֭�ٟ>����Ԑ��Cyyy���ҨQ�ذa����JMtt4n��ۍ�磱����Zjkk;�!���娣�
<�Cl0M���R����+�DDD�� >>���4RSSU������:.�����?�ġ����@�9�c�p�t��y��_ݑd���ٵkW��qW������ccc9ꨣ�>H|>������P[[Kcc#���N�%""��!|TT111����~�M$�f͚���ؕ��	@�C)IR�޳�`�Jz4:��z�|�#�466���GaaaXl{��������t""""�&M���G�.�a0���iIR�����(���Z�^v5�|�c	UUU����e��;����� �0�NEDDDD�Ј#x��牍��w�cp.�iIӞ۞�c.Lhz�����1p�@����㨣�bРAx�^�����z�F.""""��߿?O<�D`qnb��=�
���V����<��Ӥ��:���ݛ�#G����-W����'99���|�����~�XR��=�*L^�7�����G�~j���M���9r$III��lN� """"a$..�'�x��ݬ&�8��8JzO�b)�{�?�k]W�EGG3l�0�8�bbb�N'(t�������y�^z�!F���.�u*'q�*������?��ƍc��UaSL��Ջ#F0`� <���tJbb��)����Hp�\ܷ�>N8���ap1�m�=XxTa�
����8�Ӹ��{��=p�0�ӧ?����ʊ�;J�n7qqqN�!""""3�;n��SN9%�{#�Z�é@���l�w�w�y�xÍ�e�
��Eff&�F��O�>�?@�z���ݻK?�HLL�<DDDD�9�.��3fv���t`�C)I�=�h&��;������W�y�d]]yyyӑ��].���dff�v����dǎTWW�4O����G�mޥ{���
�]�,���I��R�0�]Z��'@
�i�<����w�s6�6TWW���OYY������RRRHOO?�u�4��ϧ���CE�$===$���p�p�m�v����JI
ti�	�|��|>��.>��C��j_]]UUU466Ettt�N����e׮]���5�������SN��<���3��8���!�r8�a�;�Mwx�xӍ|����Z���PVV֩�\.HZZZ�2�H4n�8�x���E�zf�9���)�Җ������	VWWs��k��oN+����),,d߾}���u8��r���JFF��9��9�~��O.������%aL��g&�����,�f�ׯw2��0M���JKK���#..���D�n7555������@}}=�a��xp���|>������&111��k��5j������;n �p,)	{*Х#��d��QVVƲk�����ɜ�����-[�PY��Փ���$&&ү_��w�DDDDDq��G��3ϒ����ipp�cIIDP�.��>��7��˹z��ݢH���aÆ444�;6++����.�JDDDD"�G�s?}�����N����ٹ�$R�@�������%%%,Y���[�:�U�mڴ�CᲳ��+��؈i�RVV�ȑ#;t2����o��ë��=���$2�5L
��*Hm5E��J�ViU�:�^P�T�8{[Ǌ�h��j��^�b���8Q�9����CM��I����C��u�y�����^K�T��k׎	�'�Qp�m$���R:q���^�KS�GoԨw����;F��w�u�֝�ynn.�7&++��>���Z�hA2�dɒ%u+I���j۶-��_>���#��J�ƀ�}�`!w�7n����}�����mڴi���֭K�V�v96++��u���W_QXXX�I�$)�iӆ���MӦM�.�L!��K�����W!	�!dbi�q�ƌ�s�n�m����:t �H0x�`.��R>���[�la��� �Y���{�$IR������s,���_C�%�0��Gt}!	�&��B����xZ�le_�,�^�-Z���E2��[nᦛn�K.! V�ZU6v˖-Uޫ$I��%77wW�g��L Q[Jct}[E$�-0��P����͛G�־�W�^ٹ��_����{��˗�j�*ƍWv=5��͎�$I��J'�ʭ"�I�)�o����]l/����B�6m�8ab�̤AP�����Y�h�7o�V�Z4lؐy��m�6
ٺuk����]�$��jٲ%'L�M�6���	��s}t}W�<]Zhٲ%�O�u������5kFNN�7o.�'�Q�F$��{�]�v���srr��OI�$E�M�6L?�����%EԖ�	�AWE�$d:pbiaժU�}��iqNzQQ|�6l ���(**b�ʕ;�o^�N�v�Z�%I�T3�k׎qw��qC��p�`sDm�1��"�"ɽ%K{ X�z5�{~�a�}핢�">���5/�v�����Q�^�*�L�$IQk߾=��G�f�R˳Jn�t�\��V�$S8����W_qι���D��^[�v-_|�6l C�999dffҼys�?�$I�a���{�X5j�u1�!��9W2��2�"�D~[ZX�n#��;�e_�$C��$�jՊ�I�$E�S�N��s,6��� 	�b8W�&ZU�"�A���BNNw��N9�(��'A�%I�j�.]�0�q���D���\������`!w�������{��Q�%I�$}��={r���w<�'�N�$#kL՚]�)$�y��ZZhРc�ˑGe_�$I�n��Ջ;n�����]����#�Jc@WeI0��kJ���㖛o��?�q�}I�$I;�����NVV��Ő�&�E�U��$NU'ɕ\U�e2�u�_��?aS�$IR���.�ݥ$)���'���d@WU;��;(Y��!���L�:5�$I�T�2���5� JK!����5��f@W~E�=@Fi��{��αw��GI�$U� 8���:thj���a�=��ʀ���@��^iᩧ��k����(¶$I�TS$	.��2N<����� �FԖj0��t4!O egW����/�?��[�Fؖ$I������su����0x!��T����	yhVZx��Wu�(6n�a[�$I���ի�M7�D�>}R�+8x#��$�b�3!�mJ,`䨑�Y�&¶$I�T�4lؐ[o��C9$��o��"jK芏�%!�Siaɒ%���|���%I���e˖���?Ӯ]���p�YDmIe�<D����_��֭[3i�$�v�a[�$I��u��_��K�p�*�0�+&芓<SZhܸ1��O�~�"lK�$I��#�`�]�hܸqj�o�+#jKډ]q����2��P�^=n������?��/I�$�������~��dee}]��u�5&���+�~Gȍ���ӧs�-7��[I�$�I;sÇO-��\M��"jK�#���7%������~�k����۷Gؖ$I��*##�+.�����p.|�RS�����	��^y�.��%�_�>¶$I�7YYY�xÍ��8_O�/I��H�#����y
h^ZX�h�ׅ�X�"¶$I�͛7�[o㠃J-^r���%�57�S�x��#������<��;�c�$I�D�N��g�=���{��\i�t�������6mʄ���Ϗ�-I�$E���L�<������%��Q[�>s���Q�L$���B�L�:�;����$I5D�v�i�{ι$)s�!����Ț����U \B���������Uc�b˖-�u&I��J����忿��N�Ǩ�:J;t��_r/�UZx뭷u�(V�^a[�$I�,6���G=����f� ��-�;3��:�I�@��+9j$.���$I��n<�@n��VZ�h�Z�����FԖT!�$N���%;��^Z���e��	}���%I���ԧO&O�\>��/y/h8W�s]�I}B����$w���iӦ�y�$IR���fp�0�#jM�PtU7I�$������?�5�^æMn�)I��N�������Xݐ;H�_@2�ƤJ`@Wu�B����E�q�%�t��ے$I��jݺ5��8��S�[L��-��x�����������Ǵ��8�#"lK�$I{�O�>L�wj�p���b8W5����f�� ~XZH&���k,S�N��tI�������s	��ED�I�΀���6I�%�w�E�K�$I����,��Õ{�;^�@���H���]5ɩa2�A���|�E_�}�$IkӦ��8��R�[8�Q[R�2�������S�^�߄ax�����<;Ѱaò��֭c��G���/Gإ$IR�շo_���Z���S˟�s<�\5�]��g���%A\ ��k�����a��ܹs��0�:u*c�K2�I�$IUa���D�Ix��j���=b�    IDAT�3�<s`����H$8qЉ��;�_{�5~��Y�jUU�)I�Tc5jԈk��f�v��7?�IcR��V\�aÆ��B ���Gu�9�����ڊ+��Ѽ�曕٪$IR�u�a�q�u�Ӵi���F��FԖ9�����?��ƍgA��}y\�6m�ϳ����ܲZQQ�'Of��I.y�$I� Ap��'s��P�v��K�J��/��5)�Jf���o���u�rک�ѫW��/��"W^u%�֭��>%I�j���ۏ��\M߾}�_z���k#hK���7��/''��o�6o�̄��v�4�o�^V�ׯ�� �rH��)I�Tu�ڕiS���[��������aÆ W��oߞ�����=Q۷og�����{+�e$I�j���.�����>%�����J)�Jk%g������mР���o�޽��ٳgs���QXXX�/'I�T����p��/�c�)�	~|U�]I��w�����+��p�~�z�{'��NQQQY=??�x��;��_R�$��8�C�o�}���vB�p"�si��AW�:��ӛժU��~e�N^^��FÆ�j�d�iӦ1��q;ܳ.I�T�ժU�3N?�3�<�Db������QkRZp]i�v�ڧS��`ѢE\}��,X����D��C�2i�$Z���	|I�������3���>�|8���a8���]i+�S��
�s�L�o[�n-�|��<p���UՊ$IR�{�<p����3���d���/"jMJ+.qWZ:��3�A�8��nٲ%Ç�i���g��ƛnd�ƍQ�%I�T��ԩÈ�Fp��'�P_�~�����Gә���AWZ
�`��@�ʲe˸���x�v�0�iS�ѹs�:�$I�:]�v���)�ϛ7�+�p��Υ}f@W����C*϶mۘ��t��=�6��۵kǔ�S8��S��{%I�T-���3y�dڶm[V_�~=c�˔{�PXX�-���U;��o��� �׿���ŋ9��3��� 33�ο���G\5�*>��ӈ��$I�-[��+����م2y�d֬YQgR����U��(�z�j�t���t��d٦ݻw��`Ȑ!Ae��$I���������y2���'����n5�K�t��J?^m_�a�/���%K�]4�@@ݺu5rG|����V�\q��$I�&77�+.��#�<r��_|��)�Y�xq4�IՐ3�JW����p��m�$�& YZ�۷/3g̤�� ��$I��M~~>>���<C�̙õ�]k8�*�3�R��D�K�لL� dgg3�����՛o��e`�$)��������0`��իWs�_�a�u&Uo�������LȄ�b~~>3��~�����$Iڭ>}����v
篽�c�c8�*�3�R�ZG����r7�иqcn���<���v�mFۥ$I��rrr�����O�C}ݺuL�6���=�\�lΠKU�Q--A��~�3f͜�1�ak�$���ׯ���S8뭷�����Rq]�:_P �T2���I�&��M�͋/���7\ϗ_~m��$��hܸ1^p�N��7m�Ĭ�g1gΜ�:�j&gХ�7���ө���\��)I�TN8�f͜��{�����+�`8�"���%�@�l�X��~����c��������/���KI�T�lْ�.�l�s�7n��Ï<l0�"����t*��{�>}�5sC�%��SI���A@AA���S8�׸����RĜA���U�N�O2hP�n]F�7���ŵ�]˿���h��$Ii�C�\q�t��}���ի����Y�`AD�IJ�ԜOЕ�;�di��C��1�dffF؞$IJ7u��a������;��0�3gW���p.ň]��u$������K��k�f�С�xh}��=I��.����q�}�3|��~���_r˭�0�ilڴ)�%��w)�^"�0��!�BJ�_mݺ5w�~�?�<��z+W���MI�7͚5c��Q����PO&�<���<��l۶-��$�3�R|m$���K�пf͜Ő!C�DN�$�H$(((`��Y;��ŋsÍ7��#Υs]���N%�f�)@�5r�q�p�����oGۥ$I�L�Ν�����֭���7�ēO�����0#�N��2�K�!��In ` ���1e���׿r�-7�v��h;�$IU&;;��������wXU�!/��23gͤ��0�%���^V��� !w]�xIۀ�ݻ7w���}�YK.IR5�H$8p #�A�ƍw��l�2��>>�������mХ���� �!�Z�@ӦM�z�՜�˓�����I����]�rѨ�v:�|�֭<��s<��3l߾=��$}t)}mn'�aBn~^z�k׮L�4�g�}��︝U�VEץ$I�M�6e���4h�Mb,X�>��|)�Х����_ �J6���裏f��IL�>�][%IJC���2�3N?������X��3g0�����T�<�I�>#�sɹ��J������/���t�$I��޽{s�}�3�����ŋ�{՘��R5b@����e�]� $K/�mۖo�����Eǎ��P�$}��m�r�m�s�ػ�СC��I@�뮿�/�����T=-#�Y�^K�P���/������ړ$I���~�1j�(f<4��}����
G0�,��$U2�T������(-fdd��_���}��C����a��$)##�!C��أ�1d�j��a���	8��#�FԢ�*`@����J������^���a�y#x��G)((�iGXI�T��  ??�Y3g1j�(���S/o#�:Î��I��|7.�HpU��鏧^h޼9�/�_���vXD�I�T���ՋiS�q�7ҪU��!�	. e�WI՛]�y�'`P�2��R/t�ڕ	�'p�ػ8蠃"jO���}���xÍ��k�;w.��&����')Bt��z��~��0�B�FrW����M�FԞ$I�K�f�}���}�o�p0'��$ŀ]ғt#`$����H$0` �<�g����$I{)''�s�>�G~���jժ�zy%�L�x�I5�]�V�Vڗl$���BVVg�qO?�4#�A�����R��4R�^=��c�>�駟N�z�R/o-� � ��K���R�/�H.��	@Q酬�,���=�СC�S�N�mJ�_�أ�1����^��t.� nM4]J�#��]YB���<�z�aÆ;�V�VI�j���N:�$�x�	F_6�&M����0�$�%Ŝ]Ҟ�A����_H�������F��r��I�Tc$	���9c&���w4k֬���%;��0?�%�	����2��/�^hѢ�/������O"�?+���!�HпfΘɍ7�H�֭���p��.i/�6UҾx���|Bn+�СCn��F>��c�z/��_)**��3I�����sÇ�cǎ��� 3��5IiΩ.I��l�Wr����;vd�Ucvw��$Ii�v��8�l�|��=�ù�o��.��
)>C�0~|�z�U�V��l4�<��"###�&%I��233)((���a�Uch׮]�!p*S�=�\ҷb@��]�pPɮ�S/�jՊ�9�>�(C��x6IR�H=.m�e�iٲe�!p]���d�w)�:1�K�(I��u�V����ԋ��?�F���'�d�Сԭ[7�.%I����cȐ!eǥ����C	�& ۫�KIՑ��I�hI���?�H��@�ҋ�7f�y#��)��1k�,֮]Y��$�jذ!�O����iذᮆ���k��p��J`@�TY���<L����/�ظqc��ϳ9��3�={6�&O��O?��YIR�ղeKNr
���
�7	����\R%2�K�
�	�E�������0��?��s�2�)���[�u*I�1:u�įN��w��N�K�M��Uܚ�ʀ.�*�D���ф\ (>S�_�~��׏W_}�i�Mc޼y�����}���SO���Րx��?s��;I5�]R����"�y����Ջ^�z��2c��z�)�n�]�������A���z��]�_����Hp�N�'I�]R�> ��M$������J/x����l4g�q&3g���Ge͚5�u+IJ;�7fРA��h֬ٮ��!d<	� `YU�'I���`	~\�A�H�m����\�=�\��9�9s�p��{��$i�:u���~����S�ή�|Q�o#���J���8Y�N�]� B.�Wz133���|���y�����t�{�9�o��YIR�~&Gu'��dz�a�K��*lO���]Rmf0�O����@�t@�.]s��=�\��KRרQ#N<�D~��_�����!I�Y� ��G�I�)��8��x8�$�J6�kT:���Ts����������BB$�m�{Uܞ$�3��t�	.���̪w+�X~����=ʳ�>˦M�"kX�T�233��~@��{Z��!����_.)��%��B`�c	 �Jt�҅.]�p����s�1��Y,Z�(�~%I�C��0��~��!I��%�؟�e�Ґ]R�
���f7���ׯOAAΪKR�����e��Va{�T�蒪���倫̪�:�tV}�y#x��gy��G���#iV��gyyy�8�D~�РA��{��	��Va{�Ti蒪�B��7|�$�	������f���<����3{�l6l�YӒ$hР����� >���+�-� �^��IR�0�K��^#�k�(�7��:�{��t�ޝ�]�;�̙�3�>�ܹs)**��aI�i�ݻwg�O���z���n���j���tS�	��)��٥Rw����/y�x��'�XN�*I��������p�	�l�rwÜ-�T��%�$���,�"�g�O��:�Y�f�|�ɜ|�ɼ��[<���<���[�.��%�������㄁'Э[�=}��)ϖ����$)�j��Y�.$9��_�Sr�!r�!����̙3���y�y��}��H���t�����G���ׯ�����!�H0x�
[��X1�K���#�e��>$9��SH�X.u	��u�x饗���l�W��](��<��|�;�85j�����'	�<K����T��%�Xx�/�98J���0`� �ڵk�;w.O=����*aFԺ$E�K�.0���|�6m���_o���IR*�$�l0����%��S��~ea���?�o��=����LI5C�.]������ߟ�͛�i�G)K�?���$)��%i�>"�U���$�%���nѢ��v��v�~�)�=�/��>���(z��J���Ǳ�ˏ�cڶm���K	�A���+_�E�$�]��N�L��)>[�IN"����Fm۶eذa6�e˖1g�f�0��L&��]���D"A�N��wT?�;�8ڵk���	y�3�rI�gtI�w�����,Y�K`�ԁ-[�,;�m͚5���`���7o۶m��wI�F��{�4k�lO���DI(�+��&Iߒ]���"�� 9d�lذa�=륻��������c����.I_�[�.}���G��~��������y�d���l��6%�Z3�KR��<B�#@=�8��H�	@�ԁ���o޼�y��1�s�;w._~�e�K��rss�۷/}����#��N�:{���'I�(�76UQ��Tc�%�rl#�c@-����D@�:u`ݺu�я~ď~�# >��c^|�E���?�׿������)�b��Oޯ_?:w�L�q��/	����%�j�%��_߭$���ܱcG:v��СCY�n���
���
s��a�ʕUݻ�4��~�ѫW/z����GM�&M��!��̔��VA��$��wH�pp0�3BN z�ԁ999��瓟�ϥ�����~�����/���^�N��;w�O�>��(�v�J"���C�(>�)�1�]�D��h�%)Zoop�8�$���?u`��ݻw眳�a�ƍ��������+���{�Eѿ�hժ�����ݫ7�{�&''��x�������ޤ$��%)>V3K����$��l2w�8����E���o�V�\ɛo��+���K/�Ċ+��IU�Q�F~����՛#�8��-[����-Y�>�?�~rI��$�S�:	^�x)|+��p�	��t�QӦM˖Çaȇ~ȫ���?_�'o��7n��o@Rũ_�>�zh���M��R�����3�2��KR��%)=,&0��]�{������F
���:��:�SN9�d2��ŋy��7��`>���:_|�E���J�ƍ9����ѽ={��[�nԮ��o۶�	�]2K>�Z��J�*�]��O��:�N�M@Ч���|v�>�H��_PP �ҥK�?>o��7�|�O>��0t�f)
͚5�G���՛�={ҡC���!�8%�?�u�\�җ]���F({�М�7�;h���jՊV�Z1`�  ���K�x�ޜ�&o��6�-�v�ddd����!�B�=�ٳ'M�6�ۇ/.	�/ V�%��0�KR��x��|�8�$? �(�ӮԬY3���O���غu+.�w��w��w���>��o@�NڶmK�n��ֵݺu�S�Ndff����"	^^>1�KR�e@����c�cL-�:�>I���^�Ni!33��X�R6l��?,�����f���U�=Hi�A�x����у�=zr��ӨQ��}x�>!/�`.�?�grI�9�T� �$��%_gS|�Q� �����~����у=z�Ֆ,Y��������>`ѢE,_����)r͛7'//���<:u�D�֭��)6�2�d���z�$�\tIR!�	�+���8�$��8H����[��u��{�e������G��{���'������u�J+�ԪU�v��o�ء#]�t�[�n4n�x_��cB���:�*��@.I*e@�$�W����,>8�>!�z-w�4�i�}�֭|���,Z��O�G}��ŋ�����=^��H$����С;v�C����q������O�x��� ���qIҞ�%I{c����OJ�h�&���� Z��	233�ܹ3�;wޡ�y�f/^�'�|�'�?a���|��G,Y�����J�fT�ծ]�֭[ӱcGڷoO��С�۷�N�:��)�o2��QȗVhӒ���.I��� KH�HJ��A�P��(	���ϛ�u��2�o۶��>��O>���>��%K��t�R�,Y����I&���-��H$4o޼��֭ZӦMڷoO۶m�]�[��N��o�`>�f��J g�%Iߕ]�T��fS|.{����@ϒ�~0Ѝ�0�[���v�ӵm۶�l�2�,YR��tI��K�.�^�"33�� ^�K?oѢŷY��j�!o����qIR%2�K�*�f��}��6s��n$�J@7�+О�lHW*##�v��Ѯ]�]^_�n+W�d�ʕ,Y����U_�l�26o��ݿ3U�ڵkӨQ#�6mJ�V�h֬M��|޴)-Z� ���_����.!��]��_x�pV\�T�蒤����ݬw�X�/��F��t�8��n�+/''���:v�H�޽w��L&Y�z5˗/g���\����|�W_}�ʕ+Y�f_}��V�b������T�ФI5jD�F�hҤ	�5�aÆ4k֌��\�7oN�&M�
K�����y���)>�� .I��$)n
)>~��]̣��4�'9 �HP���d>U"��iӦ4mڔnݺ�q�֭[Y�f�V�b���|��W�Y������~�z֯_Oa��_�aÆ}���O������&;;���g�l5jDÆ�Cx�����YY-}Iq /≒?�?�(e�$Ř]��N>/�xi�=���hC�6@kZm)���s/33���\rss��q�d�,��[��m۶�y�f6o��֭[ٰaEEERTTĆ���lڴ�m۶�=W����ׯ�鈺 hР�Nc���w����Ƞ^�zԭ[����gէV�ZdggS�V-�ׯOffy� 3  	�IDAT&u�֥nݺdff��+`i���F����XJ�O�πO(�΄K�Ҟ]�T]��(���]�	`��zk�5I�-	hA�|3�iE4�H$ʖڷj����T��
`%!��u�^B�Qe�R<^�m�\�T��%I5EXV�Qlד���f�ܓ4��hB�&w���Y��N'�(�[��c5!_�I���e�+(�_�|l/{��[�T��%I�Q�r�ρe�=��CqPO��HҐ����! �����j��Z/�� v^�^��S����(��|;�Kŷ 	�X��:`;	֔�[S�cmɟ[vzC�$I{̀.I�w�X^򱳊�];Aq�/�!_����\�ZJ���õ$IUʀ.IRzHR<{]ޮj�$)U���$I�$i��$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IR�%I�$I��$I�$I1`@�$I�$)�$I�$ŀ]�$I��0�K�$I�tI�$I�b��.I�$IRЕ��Q7�+AĲ/I�T��a�-�v'�HĶ7)��JW�n`W� (��I�T3�a��C �d��Dҷ`@W�Zu��:�$IR͐L&�G���$�Q� �#��R�D��n,��I�T3�s�=_ k��cW���¨{�ґ]i)��Q���n@�$�(����]�jݺu�D݄���JKEEE�u��ߣ�A�$�(�{���͘1�(�>�td@WZ�2e�g1�E�h���.�$IU����Ѩ{(/���$���V�Ӣ�!U�S��A�$�,S�Lyx5�>R����|$�&�te@W�
�� .Gxl�pR�MH���'�[��!Ÿ�c����7)��J[�&MZ�9�>JL�<y򲨛�$I5O�V�f oG��'7G݄���Jk[�l�>����2�H\q�$�����+��9@q+�8qbl�f�ҁ]im�ԩ���R�?~eT�/I�4q���0�#��]�6.+��e@Wڛ4i��A����1a��$IR�Z�j]̍ॗm߾���&}wtU�Z��x�*_3�'��EU���$I�3~��m۷o?x�
_vM��/��5�j+èoU�*�Yg��QTT45��+���0|"++k�wܱ��_K�$i_�}�ٹ۷o�]�/�4�L�<y��J~��0��Z	� 8�3��`4��B$���u��]�2.I�Wg�uVV2�� ���^b0x�ĉK*���ɀ�jiذaǄa89����K� 6ag+�9%I�*Ͱa�~	�
����� \�v�ڛ���*�]��ȑ#�^ \4�O�&�[�n�zsɮ�$Ii��s�m�e˖�A��~˧�L�]����ƍ[Z��IJa@W�W�O� G���aE�KAL߼y�4��$IJw�~�M�6 �q@�7<d+0x,�'M����{�j:�j������D� ��m�3��0�,�%���CH�$UWcƌI�����H$�%��@�d2� VA�E2�\XXX�`ƌ[��U�I��_D�5Z0(    IEND�B`�PK
     ��Z�c^��  �  /   images/edd00682-873b-4230-8bb4-282089490c70.png�PNG

   IHDR   d   s   n1�w   	pHYs )� )�;d��   tEXtSoftware www.inkscape.org��<  JIDATx��]\�U�����@43\�����
�����̑[��Ie��ܳ4g����L-7KeȺ졌��x	p^.W���z��}��=���s��ʨ�QXX���/����'R��p:s�M�>��ܹS�Oip+�V�۷o7���w���S�R�fef�����?x�@���@\���z����}�:��z�rC�8SS�++�6ttr�Ӣ�֭��x�bj׮9::R�^�i߾}Dj�OM�F���),(���X���k�(.>N���ѡ�ݻw=gϚ�9s��|�]RR�~ZZegg@���ED�<C�;T�����JCC�D:::dhhHfffLF������ٝb2N�A��\�Іf��(6&��RS�b�J:D�biﾽ���+����hݺu�y��}�֭�111���T����|1r�pGW�7����ĒE��M��M����]�6�I	nӺ�a[[۽|��={��0�L[�)5J!���'�#�Q�t��	;g��~~~��z���q:�L1͓���RƒB)))����q��U�#G���ܹ�M�^mӦ�6s�;xv�\�n9�8Ӄ�D[�!5�J��z�n�N���x���G>�ƍ�/(8�099Y��Q�(��ZZZ������B��}���{�� �={��`������=y14$�\\](�A�hguSm= 2�̝C�ƍ��={�_��r����F�ٗ/\#++��I(ؓ�Djkk�����1P�h�O�>mx�ҥ�G��R������������߿D�U�hlBb��
\����ݤ��fy�=�z�uYNN��pt��!�?���I___87n�@IOOO�����`ǂ4BBB�:y���ɓ7XXZ,hаA�-�^�����Q(!������h�z3�f�'M�4�ܹs��5E�C�,(�	o
��i�_��xݤI�;w.-[����&�fY��Q|}�����;v
,�,�5�k�+�m
!�.#=C�������ŝ/��C�u���V"JC��z��	r�߿O���4t�P���o���Ӈ���͛7���	;v̔%ƿ[�n�Ə?v���Wq�i�id`h�o�	��
	!�D�.��0���Wl3ta�U����@�ڑ ���_d ����t�R�ѣ͞=[H>T.���>|�T��ﳳ�E(¶<!h��ի�7� mm�m[��X�`���b+/���$@�M�2EHΈ#J��ԩu��QH��_-���]~^��܎�݇]�4�ų�ReB${q,�\B�%K���o߾���*-OTp7�5��H�۷��/ )�+W���n��'�����ɳؕ*U�޾};q��a���;9���hS��h@20����hƌt��)��㏩E�%��@�AEϛ7O�cǎߜ�5s� ���|ҐU^CT��@"�U�VQ�={~:��O�<��$�6�g��1�@��������ԵkW��,--KΛ0a� �G����{���O��j�_>���J�T�IM�\����ӭ߼����|^U�� %,%��ޢa#J�W�^�ꫯҘ1c�&{k�fL�1p劕�||}*��*L�d��n�
��5����Ґ��$ =߼ys;vl�s�☏��޽�Ο?����E�gϚݟ���CW��W�|!��ѣG��G�ӦO��E'�4������Ed�8�<V�X!�d��'q ���_����w;z��K��V����/�~�:q0D��4n<mڴ�l�t^2 ɮ888ЦM����^�� i۶m��w�^:q��B��LLG&3}XR�J�mY}}㯾��'��,���B�(�������I���A�v�Z�������f�f;�|:�CFzF
��ix"!�`����M�����f҄��
)�G�#�^PmFFF4�|ڷ�������: }�4�뱄H����t�̙I�.�/%_f�S���R�q"X,�����B�8p�v���}�d�,-OT]��ݘ��~�:5ukڊ�⢨;Q�2ٍ'�ԩSG�Z|}}���@�*偈��?�����=���`[�����Qx$!R���H����.ԩ%�,$R0<~�xLj��K.��q������'z���O"�DU-^L��z�ÿ���jQ �ᨨ(Z�|���1x�`:{�,���O0�-_i9����I�G���A
6̮���#-P+�+��׬YC��Wy,Y�D,u
�={�����o~4pP��<��0=��3���2�/��0`�A����N �����`�֭�2��R#	ez������w�� ,D����RWv�����pvv����~������挋�K��J����p�גQ	�[[[���/ń����C����_����ܶ}یѣG�������B�a~����V]U�POH��d =u�T��������v��i,�� z��t�[�n�V-�����˗�����{�s�C^�ĉ�k��	#F�8]ZJ�z����~���?�[R���t����HB>����[$ 9z���Dߍ����`f�R�͇���j�JG�!M�^�x�`�7n��9�۷s+���Ρ_�t��,OOOqL&��o���6�IK*kQuHű��,�v{��O?�s�Ͻ7w�܅�V�=��y�gSϓ����[��#f���t���9�{����޸�����#�y0!,�-���w��v�yI��l�)�a3E�O5�
��\������9�����>}�t�_�rK�d0�[�lљ���.X����J"B�N�{�ZZE�jE���]��NɃ���u�x�&�A;1'�Pbǎ�����9xǮ]�օ��a.�e����]�[ᷜH�!M���446"==A���t>?����Ρ��4JKI�L�ZL��]�D�
���mۊ�F���NY�Y�"""��0)����:�����paz�d�zYO__�KOM���22ҹ��s4��utuɈ	321!K�dbnF)ؤ��$$F�҂6a���͛"�ׯ_���@Թsg�R��_g_���l��1����=����nyH��Eݺdja.^G߹Cw��!b%N��-6�}F[G�,�Z�m�damM�L����l�J�����4k�L,��y�f�1c�,���9�wÒHU�������̄UO*�
�d� �=I�ssr(2�6��Ē��� ��}C�a2�32�F�� � |i Ղ4UdT$�+�VW6�b�(��g�d�R������>w�z�*>�`�C�Rfz�4iL�Xg߽!S�F��BLR���1�����J���dmURW�l�M,,Ȅ�Ƥ��v���ԫ`�Ԋ�����[S��zt7"R��2 m�;y�$���P�F�J��M��>�@'(0��,**�	쇪,�sլ�ͭ,);+��X���>\���H���ۓ)�ĸ{JS]R�#�@@(A��������%��� �Sh`eef*���5޾Ff��
�(U�"T�2��;�����E�i���.Ā���.2�\n��
�����p@��!.&�48�q�|wYR\�6�Lҽ���j8v�!:���#ޓb(8U����E�JeV� ���o/�]T4R��z��NBCGd�9>),�~�&�w�ok�$BDa*� p!���2VV��
���z���DR���+���C*K�;H�(����]�z��=i�#�eee�rssuIE�ѫUG[tv�V�*�ŧ��r�X���e�7��B"�R����	\���i���H�$
33�KZ��
�	��5�2�J�#P�X̓u� D*���Z���0EP/v��aU���EG`*�
CE���!�^z��/u�MhWͻX$RQE)%��Ջ�)[;Hv�����ui�j{1�H�jhTAA���ji��R]�U�^k��K�e ���Xك�]�T�p!�����7j� L(���S����%tj���c0����Ҷ\�t�u��oCR ��t���rp��)8�55���XD��s�+=(����`.
˭�|�����%�zP�l/��efiAV�����>S�c	IM���lB��+$1"������(��pW�W�t2�D����RH	�u�O07
���	H;����M@
s-333���J�j�����ř�������kk���--)eg����f�i�f,��Bfmm7�F)oT��y�G�p,NH��kie%rN�7Þ9����А�7� �X������}��Dl�ƵAb�����K���qall�2�H[qGԤ
�o��Ƒ��69��_�NDdI��� i�֢�ȸ�EGS���� %O�����& �-�9���`Krk�tx@qw�R�vԨiSֳ�q�VI5�� �+��ͩq37���R)I�5N���0�H�S������A�96(�?Ɔ��mM���gR4K��m}�g213LX���EIjʔG �˖mQ}V 1!&��T�V�����ѲF~P�N�w.0�ŚS��I;"���;�#Ȝը1��+��<9Y�Ę�3RP���.F@�o�O��bˁ�a�D��.u�f�����m
2��^dgk�gÆ�a	��������`)dM���@̩�ݽ+�TH����PCP_пy�5�%B8��1D���F3q�j�?�M>n����*GY�W[����_�5J;��!�/Uٵk� �PE� +#C<�h�KI���\�9�81��_���Ey�B�T� ��@�q�xΦ�ɘ4��ҥK/���.\u:�l�"��H��)�ԩ�9�b�n�Z�6D,�-vً�qL]�� ����z��6{b�����>GG�ΨH����w�+�TU�PD��#^�)̣��2$uղe˽�7mo�~���z��AOO��7lؠ�ſ(����N���q�*��k,�^�p���k��	PE�8b_�zu�/����O���8?��#��P5Iy��עE� ���ev�BT�;F��m�{xx�D�ˇ~H{����%Dq�t mҩS���{p B *(�8Զm�&�bl(A9;,��-�P�^Q�K�9���9 �ݯ��J����!~��@A�VG�l�s�t�j����{��E��L$T݄��(��-��K<Liu�"!�Fa�X�a��� ���Q+���ǡ
����v�:y���Q�`ذa�.9(�����И��pq�U�(��T��@]�j��n�6b�-�C$�)ٷwE�D'���{ف��DG���H�F�mHLU�d<d �1�T����L���;�X����ԧ^��-�Yf�*l���+������>��3��o���Ġ����6��9s�C]�k�.��W�zC�y�2�@J�\��������]���?�]? ����w
��$�"�,����~}��߻wo���ʙ�9�M�Q��a@�Ã���@�-�CMA�e��EJ^V�����Ǚ����e�)��D�,�`����|���lе���ؒ#G���)�"�Z<��lӦ�����N�ܥ3��S��������1͞5�����°��y�Ӏr��ׯ�lP���jIy:�U�Ư��^g͚u�6�1]�HB�;��_0/w�w�^��Q[U@JӦMkIy�B��z�:�f�7�C,�x\���nL��b������q��Ӊ'�ɫ_�Ư�J���j-!�y׮]�YU�bg)OWG��Z�}��O��,/�N�N7|}}G�]�u��I�3g��}�� 60���C_�.��f�4n�����q3�&M�4���y"!"\\�������޳�)�Xǅ��K�.��*�n��`P�� �Q�yx�(q�RUUS�	:��=z�,V��q�i؍g�� +�׮[�N����?��aRǈbQ ) J���TLyR$}��Xn��j�HkT�� O#G�\��>�;M�����B�Md�2q{���ddf��+�/�i����X��Iy��HE�UR��� �>|o�~}}��3���Q�6T�ɋ����6l� f|�ƍ����	�`V�I��q�ʅ> H�6������|h�F�.�#�������~���;6n��s%PaR&�et���0��#F�x��"�Ҡa�J�_*U�It4�����.��/��6nO��e#���6c��^��H�x���D��+��t�,�y�"M�5��z9|�p��5k�����I��, �.���[�N�w>0`�pX��W�&�U�X��Q��`��ܺu�S>�b�ᙳg�ZUu���aR�վ}�_��}��Y#�$)�l��T9K\�r�Ad��077�w>4�������KG��֋Z�R���n�L�:uk�saaa���C�����\ӯX��GD��+f����?��		Q����fMY+P�:���<�s H:�:���*�(��>�~�j�ՙ�W�.������ǝ��pL�9YQX"�+��:t�@F�F��y�B1���7�/ER�VA233e�6o:8gΜV�yL����	�.]ҕ
5?/�HD }���!o޼yBxx�KPp��Np����+�z��)�\��G���bŊ�[6o��G�^AAA��U����ܛ��w��駡C�Ng����fWgm�j��F���ү)*2*���gz�͛7O:u�T?�/u`��V�U��}�1�Q�F�����������?����Y݃�Z����+R�HD���gҤI�����ݳ���_g�m0]���Х�ɑH�G�rIM�4�n۶�O}��Ycllܦu���G�����ɒ~1N�N��GEE�:}�%K��]�r�ۙ3g��]����۷���G��%�A�K1�X�����Oe��D�v�7w?4y��W_}U���)Vn*�STZ)k�R��l���ע��Rbbc�������۰��x��n�>��u�a|B��ւI�U�o�|T�_z.}o�b#,�v��mmm#����jѢš�-[�s��zHLQ��h�� M��eA��Kw F�[]��&O�G���n�~���p+����s�εd�i�4!>��<En�����Տ 	j���E#^]M]�I��[Y`���� ���D&!��u�@��c��!Ӹ�^S
�7�m���i�%A��SeP���K_4TZ��ݩ{���lv/�DGG_�����9�B���i��i�V���\.7���4B�BV+"%���������Ke���������D�Ç��{`! 11t�ʕ�;�T *S}���6�ɉ��O6l���$d��di�:�B��\����i,c��u�3�h��#ϣOU�2��GE:�qi~5��#�|T����y����&�ED-!*�ZBT���j	Q1��b�%D�PK������Q���~��"�|M�Dz�P��oL�C��[�"����~��8�"���ѝo�c#?�)��L�c)p�I    IEND�B`�PK
     ��Z?S�2� 2� /   images/da48ab5c-24bb-4ba8-ab59-39208c7b2ba2.png�PNG

   IHDR  �  %   ���   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���   �����
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �ك     ��FPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU&��M    IDATUUUUUUUUUUUUUUUUUUUUUUUUUUUa�ޟ<+;�?�9���/s��f a *�K e'�P��xvf m�T�w�����a��j�T*��$f�V�4j,%� 1\gg�/����y�/�*�9}y�~���~<���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ��Ū    �jkw�yIou������h�g�R��e�qQ��c��,�RY�Y�"�zL�ʲ�~�u+!OE�N)e�,���w˲lǔ�B)�!�����t�
)���\J)Ʋl��/e�8Ƙ~��S�Ն?��$�X�B��̲l�S�;�1�1�eE�qc��,�Gy��2���eEȲ�"����s���hƸ�5���x�ޙ�Y�����k��      �>�   ؒ����p�g4���c�UŮ,�]�t����L*˙�,gBJ�4�v��e��R���l��hƲ�������B�y>IY6y>�Y6.c�dY6�Z?fY?��/c�Y֋Y�k��)��q���Z�|Q��Z�����?      ��;    �IǏg?x�ˋ�bJ�EqIao(��yY·��+�r.�L*�nV�4���tڊ�m�h)�k�Q��)��1�7R���Zm=ĸZd�jȲ�!��!��b|)��ԥ�_�B<~���     ���!     LZ\����WN���8�.Eqi-ƽ�(�Ĳ�U��{�-�b&N&�4��չ�R)��T���<�Zm-���S���<?7M�l��?H�کZQ�`_��|\Z*��     �)   ��]wu_8�@=�ק�|}*�KCY�e9'�=i:����0ͅ���{���Qj4zY�����)�{)���Z�T-�_HY�Bʲ����T�
     ���   �`iq1a0�:��`*�+�x��T���$M&{�d2����X���[a��y>I��Z���b�~����,;���,;���g�����     ���   lc'?��+C���,���drE^��䒬(v��xw�L:n\��'�X�z���e������<?���z���d�ԁ�z��N     ���   la�...��7���XN&cQ싓ɞ4�K��X����W&�X�fs=��gC�~>���P�=_k4�N��w�e�w��Ҹ�N     �ׂ�;   �&�{�߿&���N��_��q2�4����pxI*�ZՍ�ŕb,c�������8����z��㓡^lay�LՍ      ���;   @�N�v۵�,�K��~z�F�ݡ(�U�[L�6L�湬�x)��_L����,{���z�ɪ�      ~w   �����Ņ�`������`6_�����p�'�e��>`g�1��\���h<j��k��ө����O|��U�     �   \ �>���j]��F��S��r<����p��M��������f�ƩT�?�'S������?ZZT�     ��    �Щc����五��x|m����eq8�R��^b,C�������:j�'k���Ӣ�ځ�z��<     `{q�
   ��X\�,�ظ)��[�h�r4�<�F��dҩ�`3��F/6��S��B�����E������SU�     [��;   �����b�����drS����+�h���]U�lIy>
����n?j�'S��x��|����sU�     ���;   �c��﮿x��i:�1N&����W����l2�K)yO�J!��l�f����h<���;e�����f���I�}     ����   ؖ֎�۟L�^����h��0\�KSQԪn�'b�E�j�d���E��O�f�Q��wW,-�Xu     p��   [ީc��R�F7���8]�����h4�Vv��)Ƙ�Fc5�tN����E���q���+�����     �זC^   `K9q�o���o����a8|S��x}�N;Uwp��(��gB��Lh6�����{�;�Ǐ�U�     ��;   �i�c�~��0����`�y��F�kqi��:     x��  �M��m�][�͵���p����EѬ��-(�GY��´�z��h<2��o/�'��     ^��;   pѭ�y�%�kk��drc>����!��Uw������9Z���������XZz��,     �g�   ��G����77��w���-�`pU�v���� �2)�����v�ټ�z��j�Þ+���x�=���     `'s�   \P+G�^3�ߓ&���~�-�׻*��W� /'�X�v�L�v���oO���^y��OT�     ;��;   ���ƙ���b8�9�F�Q�`���. �`�����>S�Z��z���w:shiiPu     lW�   ���s��~is8|�n��ᵡ߿,E��. �XR�Mb��b�t�(k������,,/���     �w   �Z9z���dr8��
צ~�> ~V����'B�����������U'    �V�@   ���w���b0�a0�!��o���ު� `˩�7b��L�j=Zk4������/��    ����   v�t����'O�'���-��W��Uu l;�Z?t��+��oN��W��~%.-Ug    �fd�   ;DZ\�ό��*�Û�`pS���h� _ʲq��(��G�F�s���/�    ���  �6e� [��;     ���;   l#��94>�7�^��Pͪ� �W�V�n����~���?w��?�p�I     p��  �v��[�.Cx_����ׯK��l�M �V��c��tj�nt:˗,/�S�I     �Z1p  �-d�ر������~��ac�m��_��	 ��Z����>;��;��KK��N    ���   6�G�^�l�R���-76ޖ�����< �bL��9��GC���݇--��    �Wˁ8   l2���E�wkn*�ׯ�EѨ�	 �b�OC��|��>�7�[x��/T�     ���;   T��ѣ�&Eqx��0���#��U7 �D����'b���h|bay�L�I     ���  �E��66�c�N�7��n������ ��-�Xf���C����l~f�����TT�     ?��   .��n����ht4���kko�I��& `���qf�43���K��    ��  �k��w�u����ol*{���-� �fc
���0;�������n�b<~��:    ����   .�s������}�~��qu��4�V� �4kav����|��h|lny�l�I     ��   �+8u��u���C���C�׻*��W� p!�,�����N���n�c�[^~��&     �/w   x�N9r���7���+�SJ���#��g���7R����o| ?^V�    ���    ^F���K++�L������x<Su ��P�������y��t���}��U'    ���  ��q�����C�׻9�zoHEQ��	 `3KY6N������~��v��KK/V�    ��c�   ���#G~=��76�^�`H)��	 `K�1�n��43��N����[U'    �5�  ���>r��t08{�76.O)yV ��R�}6��}5k6?���_��    ��ˡ=   ;JZ\�O7���
kk���U7 �(��J���Vj�>y���Ǐ�U'    �y�  ����Ɖ��;j���am��a2�V� @��X����v�ӗ^~����N�n    �Z�   lK���'_|�q8�=���3L&���  �%j�a��{<t:.\s�G�=���N    ��3p  `���Q����өQ; �Vd�    �c�  ��� ls��     ;��;   [N��?n�y�M�׏d��ׅ�hV� �EP����7c��Ʌv{9.-U'    pa�  �%����d���� !��h����7R���7��@<~���	    �_��;   ���#G�އ���o��x��  6��j���ه'�ֽW>��#U�     ���  ��>r�P���nX]}OwW� �֑��a~��N���g��    ��1p  `S8}�o���X���'{�� `��1ř������v�-,/��:	    ��g�  @e�]\\hnl�^\]�%�zW��<� p���47�T���|������ݷRu     ?��    գ�w��j
�ޱ����R^u  ;H�����c��yp������4�:	    ��0p  �5����-q8�=�?S�N[U7 @�Նa~�S���x�����$    ����  ����#G�^�����o��x��  ��Z��a~�˵n���oU�    �S�  pA=����\[�HX_�@�����  ^�N�T97�7i~�O�XZz��    ����  �_Y����K?���bu�����SJy�M  �+������	33���_ť�q�I     ۝�;   ���#G�އ��ʻ�dҩ�  ^+�����o���??���~��    ����  �W��m���)VV���uU�  �Ŗ�����gF��zpi�T�=     ۉ�;   /+-.�/�w���_���%��U�  U�1a~�;���_����?�/�n    ���  ��N�v۵i4�H<w��a<���  6��h�����ess�,,/?^u    �Ve�  ��x����z�����^�ꔒgG  �7J!�lv�{a׮�?�������A�M     [��   !�N9r���>Ο��0���� �-/�Ga׮G�����O}��U�     l�   ;�ڱc{{��nK����{  `ۚ�9����?p�%�=��_lT�    �Y�  �@'n����`�ùs7��hV�  ;ƿ�����������U�     l6�   ;ģ�w���VV~'��_Su  �x33'���]���?���3�:    `30p  ���=����������ɤ]u  ����7®]_����YX^~��    �*�  lCiq1i8�c��򑸶�����?  ��R)���^ص���]����{'U7    \l   ���ѣ�l���5;�����;���.�|�<�h�,ɒ��q��)KK
��=m;Rb�
n�a�f�iKSZ�����2���4t:�-�;�q�b'Mo�mg���8޴[�%Y:�<�7��[ ;����~�o��_��}~
��{  �g��j&Y�����ʛ7��{(v    �R1p  X�>�=���.LM]�����  �i�fIS�w�MM���K.�J�kW9v    �b2p  X���oo/��^�NL��ͱ{  �EVS3����bC��o�����9     ���  `��<;��tb��\���  ,�4����Uhh����u�_��    8��  V��mۚ�O��>LN^��<�!v  �<���cIs��,���{�l�    �3e�  ��Mn�v���쇒�ǯHJ���=  �2UQ1��_�?��՟ٴw��s     �-w  �eh����03�3LL�,	!�  X�4͒������}��{b�     �.w  �e"\}�ГO�+LL�5��97v  ��54Iׯ�rg]�Ӿ�B�    �Sa�  ������������B��.v  ����L���{MM7���7;    ��1p  ���UW]R9?}:>��e�{  ��-�r�t��of���=�����    ���  ,��ۛ��Sir�]���ܗ  K*$IH���[����.��+�]��M     O3�   XGz{[������oJO�l��  �$I����l�    IDAT���;�r�ʻ�    `�  ���tw?7�������+�R�&v  �3���K֯�����lڻ���9    ��e�  ����/33;���˒r�{   NE��Y����|C����{O�    `�1p  8K���H��ޖ��u��  8#��L��������t׮r�    `m0p  8C����n��ݙ��]��Ϸ��  8�Bm�h��z[W}��}}��=    ��f�  �,Mo��:=;�������Ph��  ��Қ������uMM�n�뛊�    �N�   �i`���$����ؕI�U��  XR��'���{��}j����    Vw  �S4��7]�MNސ?��P.W��  �)�狡���Om����    X�  ~�����'33�$!��  �g�4͒�뿕54|f�]w��    X�3   ~�cW]uu:=��dj�y�[   ���$!mj�n���s�����    X��  ���ۛ����剉����c�   �HG���?�|�+�K�kW9v    �r�  $Ir_oo���ٝ���u��|K�  �� ��	--�����Ҿ�B�    `�3p  ִ���[�gg?�ߞ
�{   V���f*kn�j]Sӧ[���b�     ˗�;  �&l������G���7�YV�  `M���K[Z�ַ�}����b�     ˏ�;  ���������b�b�  G��
ik���kl�x���#�{    ����  Xzz�K��>���_��"v   �4t_hi������b�     ��  ���֭�I>j�  �|�    O3p  V��ۏ�,�ˆ�   +��C�BSӮͷ�>�    Xz�  ��2��s~yn�F�v  ��+�狡��k��    ���  ��@O����ڰ  `u�ǡ�����n���?�    X|�  ��6�}���ӿ����&	!�  ����    �w  `E2l  X{���kj~�cϞ'c�     g��;  ����T��|${M0l  X�B.WL[[�   `2p  V�v   �����u��}���;���    �9w  `Y��y^:3�+���"	!�  ��'�r�|k��曚vm�����=    ��g�  ,KGz{�ɏ��Zz��e�\���  �����������5�v�X�    ���  �ʑ�ޖ��ԍ���5I�U��  `��8���7vtܔ~�K��s    �Sg�  ,����n����dl캤X���  �ʗVU����u56~:��+��    ~4w   ��ۛ���Q~Z(4��  `��=��������q�kW9v    ���  Q�]�rC�������������=   �~��~��������=v    ��� �%7���������\g�   ֠��#���Ϝ��G�    �_2p  ��`Oϖ0>���ĉ�c�   @�n����}��{����-    �?0p  ��5�\Z���1LN^�   ���$!���H��������=    ���  ���5׼�rz�?&��JBp�  ��Ҵ���<�����{�<�    �*  ���9/���X:6��!�|�   8U!�+���_�56~�s���=    ���  g��������'��㗅r�"v   <k�������H�����9    �V�  g,\}����b2:z]R*���  ��%TUͤ��_�jl����/��    ���;  pFFzz�\�Hz�d[�   X,��n0ݰ�w6����    V3w  �Y�<>��dffs�   X2MM�+Z[ol�㎇b�    �jd�  ���[�^�;yrW8~�U�{
   ֠��崥偤��ƍ���c�    �jb�  ���mۚO��ޔ��^���=   ]E�|hk��X����{�    ���;  �C��������'���N����=   ����L�6|���/��t׮r�    X�� �h�������/�����-   �܅��c��哛����    V*w  ��8����tr�tj��c�   �J��iH��Iׯ�X�w>�    Vw  ���tw?7?;{S2>��$�   �,��\)���uC{��o�m,v    �+  @2���trj�c���4˪b�   ��QQq�����s��>���b�    �rg�  kX��������;�B�1v   �Z���Ӷ�[������)    ��� �5�ӳ-��07��   ֊���{Ys��7�u���[    `92p �5�Hw�s+ff~;���$���    �Z�������56~�s���9    ���  ������w��ӑ����rU�   X�*+g���?�jl����/��    ˁ�;  �G�n}sz����'O��n   ��PW7�۰�7�����    �� �*6�m�K�������n   ~��$!���ºu7l��?�    b1p �U�-[�+�>���t'!�c�    �(�_(o����ټ�7�/|�;    ���;  �2�[��3�p��o��   <;i]�p�����ٳ竱[    `)� �*q�������O���ύ�   ��4MC���Hhj�������{    `)� �
7�m[���ٛґ��B>v   pv�\��nذw4M?��{�    ���  V��kWn��_�p2<���X���   ,��������{�~)v
    ,w  X�uw_V9>�+��97v   �Ě���ZZ~���;��    g��;  � O]{mW���o'cc�KBp=   kT�˕{WT|��w�=�    ��  X�C�4�5ɲ��=   ��������[�ٳ狱[    �l0p �e���W��jj����sb�    �TS��bK�Ϲ��Gc�    ��0p �ej���i~|�w����IB���   ��4�/���=]�{�G��}n!v    <�  ��l������I���   XYҺ��dÆ]]��w�n   ��e�  �ȑ���V���v���-   ���$����7tv~����b�    ��2p �e �����%���#Ͳ��=   �*QY9�tt|q�޽7�N   �Sa�  �vw��|��'��ٍ�[   ��)45}����Ϲ��Gc�    �c�  �Ll��|�ĉ�I��.OBpm   ,�4�/���=O57�xi_���=    �L�h   ���[ߙ���BXXh��   �-i]�H�aïw����    �5w  XBG����NMݜ��zQ�   `�
I����:;?�x�mc�{    �i�  �Booձ����##oI���=    I�$Ie�l���ō{��;    ���  ��-[ޘNN�f:;�1v   �3	MM�ͷ��b���ߎ�   ��f�  �dh�������&cc�KBp�   ,ki>_
mm{�jn��Ҿ���{    X��l  `l���td�áPh��   p:Һ��a��7����   ����  ΢�����cc7'Ǐ_�   �YK�r���w���}x�wL��   `�0p ��d�v���%�bm�   ��!TWO���qϞ�c�    �6� ���9?LO�&&^�   �lK�4����������7�   ����  ���UW���JJ%��   �Z����ut�fמ=}�[    X�� �Y�ܶ킓�㷄���n   X*O�����|}����c�    ��� �i��S�>)�jb�    DQU5]jo�����-v
    ���;  ��C�\���o	���.v   �r�67�[hk{���o��   ��`�  ?Bص+7x��7���w��rU�   �e��r6tv�|Ξ=_��   ��g�  ?��5׼(����p�ď�n   X����}���������   ��e�  ���S�ӑ�w�,���   �"TVΕ;:nٴw��c�    �2� ��2�m�K���φ��ͱ[    V���y_hj�����ñ[    XY� ���ުcSSϏ��\Ȳ��=    +ZE�\��y�ƽ{o��   ��a�  I�_sͥ���O���c�    �&����������?�   ���� �5-�ڕ���ӑ�w9�   `�TV�̵���y��;   ���� �5kl���FF�09q���-    kA�ܼo��c��}}C�[    X�� X���jg�p�eձ[    ֔��餽���{��E�    �w  ֔���ۓ��ϗ��_�   `�J�4�������Ë�w6v    ˇ�;  k��֭oMGF>
���-  ��U\pAe~Ӧ���p)��SS�$��Y ,C��v,��|d��w-v    ˃�;  ��[�4�W(ܒ���.��  Y��s*�~�g��ai(C���,����Yyx8ˎό�H�$	iZN�����?���/|��   ���{  X�F�n�2�d��o��  kE��'�@S����g�aa!�'&�?zώ-����K�	�2S_�����w��P�    �1p `U
��U�������\�8�  �\ݛ�ܐ��8������Ѭ4<��GF�lp�������|������ƿ��O�n    C  V���ݯʍ��~27��  ֪�W����Kj���'�lh(+f�GK���YRv�;�����x][���;�x"v
    K�� �U#�ڕ���ӑ�w�,;��" ������+j����l��P*���X�����,;v�����UT̅��Ϝ�g�c�    �t� Xƶo~ad��'Ώ�  $IRU��{���4]���!���d�<8X*d���,��w��Җ�o֯_���ݻ��n   `�� ��^u��00��$˪c�   �������Z[�K�{��\�<:��JٱcYyh�2�w��,���
�������-    ,.w  V����ۓ��ϗ��_�  ������ڪ�(����T
ah�T��ǎ��c��V��$!ݰ�o�ji�yi_���=    ,w  V���[ߚ,)�c�   Ϭ�yϫ����w�B(��e�#GJ��å��Q�w�$���6l����b�    p�� ����ު������W��g `YKr�~wc�)�Byp�Nx0xX�\����߶��{?�   ���  �ch����CC�Ofg7�n  NMû޵.]�.��t�R)���R��އ��$��Y <���o/tv�������)    ��  �[��?��$˪c�   ����+�*~�ǫbw��P,�0<l��L����iG��:ﺫ?v    g�� �e�-[�+nIFG_�  8}�/zQU��X��l
'O��c�J���*�*���r�&�5/M�I{{Ws�i__;   �g�� �e�Pw�eU##���[b�   �N��%W���5��XL�ĉ���S��'��ѣ���UD�n��l����uׁ�)    <;�  ,;a׮ܱ��)?<��B>v  p�4iر�1����NYYʃ���������W��NwXj��'�6|j�=����)    �>w  ����^�)7:zk25���-  ��Q{����_�#�p�D�9R*>\*<XJ
��	`-H�4����}��e�}}'c�    p�� X6��6�J
���-  ��Su�%�կ~um����P(�)e�����,v��WW7�l�������N   ��� ]������dd��$ר  ��Ttu�k���u�;������������ҡC��Tr�;�"�\!tv~~�=���   ��x ��ƶo~ax������b�   �$�Kv�lJ+*<��A�,�KŃK��/���r�$��&mnޗ����s���-    �`^&  �Ж-�-�R�eձ[  ��U��7��6m��ݱB���hV<x��<X̆���A �EZS3�tt����w�    ���;  K�-[�+nIFG_�  XU�zUM�+^Q�c%
'Ndŧ�*eO<Q,9RJ�w8!M�i{{Ws�i_���    �w  �����W�����'On��  ,���<��v۶��+��|�t�P�t�`�x�`))B�$��*]��\s�{;��y2v    ��� �%3x�CC�HB��n  �Xee����oLr9ϥϖr9�JŃK��/��G�����j&�踩kϞ��-    �/  Xtl��x�����Ǐ�d�   ������\{{E�U*�������W,8P���� �*MC���ծ��Ҿ�,v   �Zg� ��:���򊑑?LN���  ���u���z�K�cw�剉�x�@���c��䤱;�)�����߾���c�    �e�  ,��-[�[��$�X  ����+k�l��ݱ�������D��������c�    �U�  �u_~y��,�������n  ����&mx��Ϧ������G�)cw�g��i�ut|yӽ�~<v   �Z�%  g�@O��������sb�   �O��߾.�ܜ�݁�;���kiy��a�{�����   ��� p����-;v�cI�T�  X�j/�����ϯ����T-��/(�'���VS3:;�?�_���)    k��;  g,��Q9x�����թkL  ���|��j~���bw��lh(+}�������0?bĖ���RG��ν�[b�    ��G  ������҉�?���.v  ��嚚r��xGc�NA�|�X������ŤX4vֶ����jk{��}}'c�    �f�  <kǮ������'C���  X9��ƴ�>��SB��S������Ť\��G]�P��㽝w��H�   ���� ��v���ﾛ����3�(  8-u��u�.�����fg��'�,���B6<���Xr�Ig�omܻ�K�S    V#w  N����\��ѣ�975���-  ��T�җV׼����;8s剉������03�Xw`�H�4���{�.�����P��   ��� p���__�l����  X��6�����u�;8�B64��{�Pؿ��
!v��hhx*�~��:��y2v
   �ja� �)غ��tp�!�*b�   +\�&�{_SZ]��*J��=�d���c���å��`w`�����uv�j�]w��N   X�<  ��
o{[��c���]�  X=�o�ϟw^e�W��+��/y�P���tV�4-����l����]��   p� ������Eax��07��  X]�_��W��6vK�<:Z*~�ۅ£��R)��Xis�RG�;�����   �R� ��zz�%ǎ}2)��b�   �O~Ӧ��7��!vK/,,��'
�}�
��p��l����6���/�b_�   ���� �c��+>��ޓ����  �Ni>�4|�MI.�9�V��Ȋ��������S݁գ�b���y�y{��;   `���  ��{����7��99~��[  �կ�-oi�wvV��`(�Cv�`���#���å$غ�@�����wν�~$v
   �Jb� @�$Irt��Ӊ�?Kgg7�n  ֆ�׼���e/���������w�[,~�;�0=]��p����׶��������-    +��;  �PwwOyp�SI�X�  X;*~��*k{z܇��B�C�J�o�P:x���m݁�+��N���ݹ{��c�    ,w�  k��W|4zw!�  X[������oL<��Gss������C����TQq2�����={�b�    ,g^  �Q_~y}{�pkU�  `�����ZZ|p˩)�Cv�`���#���å$��E �'Mˡ��+��{�Gb�    ,W�  kБ������tv���-  ��V{�e�]T����<9�{�P|��BXX�tV�t���u�������-    ˍ�; �3��}Y������  ���ϯ�������\�Xف�·�Uț���    IDAT�Ʋ�= ���n����m�w?;   `91p XC�l�p:8��P.W�n  H�$I׭�5��]>��(���
?\(��_��;�TV�:;?�yϞ=�S    �w �5 ��V��.�"v  ��V��w5�֭���`�'O���=V(<�p!LO�c� �0i�fiWןt�sϧb�    ,�  ���k�ݔ�Rr����[   �I�-u^X��U(��>\*|�[�ÇKI�� ~�����jk{��}}'c�    �d� ��ݲ卹���&�Bc�  ���⋫�������n�����C�G-�,������ׯ{Ǟ=O�N   ��� `�:r���PȲ��-   ?L�ښo��u�;X��|��装�C��= �FU�L��M7��qǽ�S    b0p XeBoo~`|�������n  8%i�4��ј���b����ˡt�@���o.dcc�t��4�+�:;o9��{n��   ��� V��mۚ����<LN�0v  �騽�����ϯ���ڔ�
���B��'�I�s �$I�4MChk���5�ٙ���/N    k��; �*q�������/%ss��[   NW�O�Du�O�Tm�ֶ05���+��+$���;�,������_�ʻ�   �� V�����'CC��º�-   �F�ƍ���^�4,a~�\|��Bᡇ
��	�&х��c����:���n   Xl�  +�ѭ[ߟ���e�[   ��4�Ov�lJ�yϭY>��P:p�X��7���,v������\g����ob�    ,&/
  V���_��th��u  �
����6��9�ǻ,K�G��\(>�T)	!v�F��|1���[�{��Y�   ��b ����[�yt��&��/��  p�T_ziM��_^�~���xVx����c��r9v��iH:;���/���b�    ,w ��k���-����  �l�ؼ����kbw��(�8Q.>��Ba߾BR*9�Xz���u���#��+�N   8�� V�����%�÷&��-�[   κ��t�Ν�I�zv͊��˅}�
�\����J��n����ݻGb�    �-^  �#==o.=��$˪c�   ,�����!�aCE�8]�X�����}!�̔c� kHm�hn��wv�����)    g��; �
0t�7f��;�r�[   S��P[u��>�e�*�C�����̗''݁�QQq�t�9�z^��S    Δ�; �2v�|�?HFG���  �*/���f˖��p��q�>��o,��ǳ�9�ꗦi6n��ƻ��l�   �3a� �L��m��y25���-   K%��K������kV��:T*|���Cw`Q�iB[۽]�y��t�.E   X��   X��n�zan|��&ss��[   �Z�;ޱ.mj��-;v�T��7�K��b� �[�ܼ�P}�u������-    ��� `�ٺ�����g�b�>v  @5W\QW���U���R.-|��'�(�nV�P_,��v]g���-    ��� `9v��!7<��\���  K�EU�\vY]�Xl���bKkj�r]];;���-    ��� `�8z��H���K]�  k\��9W���7�R*-|�����\!ٸ���ٻ���-    �";  `��v�v��OFF�5n  H�0?�.��*��t�Ě�64�*/���r��0?���M�ꑆ�ϝ8�_�������{    ~/  "z�������NL�8v  �rR��]�������݁Ő�i��_��W��[    ~w �H��vV;���33ω�  ��T����5�}mm����X6�MWK˻Ӿ�,v
   �3��  X��tw?�jh�+���9�[   ��4��򢋪cw@LiCC����*7o���<1Q���ss�g�����[�����9    ��� �ر��������C��.v  ����%;v4��՞c�?ʆ�J'�gK}��rW�����ۏ�N   ��  XB�W]�~3�2�  �u�^[�?������d����ώ+�nV�P[{�z����v�~,v   ��� ���֭�O���$�|�  ����'���������U�����������p�X�*+g����o����N   H�$1� XG/������$��n  X)�\.�|��bw�r�66�+/���bÆ|62�����	X�������_|�ˎ���Gb�    8� `�;*��x��0:���-   +NEE�n���$��,~�r9���/���B��)��V�4M���s�S�޽��n   �6/  �×_^�6?��tr�ű[   V�����!��Y�V�P*��}��}!,,8�8-i�����Ս�W?�   X�� �S�^�U=<��ω�  ��U���5U/}iM�Xq�>�Px��BR*��%mm��ζ�w�}}Y�   `���  Xm��o�(70З��v�n  X�Ҋ�����bw��SQ�V�{ne�_X��J!͒`����'7�f�O���w����-��   �'� �E#۷��t���B�!v  �j��Ԥ�{_c�y6����dVx�����݁S�독���l�����[   ��� ��d����ţG3�2'  �E�o{ۺ\K��H
gAyd��p�}�C�J�[��!��=^��|�s����-   ��`� pl�zC8v�i��-   �M�e��V\tQu�XM�#G��w���X�X�Ҫ�������=�   X��x p�����ñc�K�ĸ  `�����.����I��)_y��U������P�
!v��eYU��ܖ.����|7v   ��� ��c�_�����u���  �h��|�z�K��g_�kk�W^|qUZS�f��YR.�n��*r��?�/{��g�;   X�� ���kWnG>k:2��  `�+B�EU�UU>.�E��ri�����/�JJ����d���e*�\z���>������'�;   X�� NSر�r�������&v  �ZQ�ٙϵ�z��(��J+�?����~�"LN���ӎs�I��w��u]灦��g�&� 1H��8�3�X�5q Ip��Dr�T�+�S݊ɝ�z�0�VwUuD٩NuW�R�Tű%C2)S�%��Xq�x��XII  A ĝ�9g��.ٚ8 �wx��Z������|�;2�����ͱS���6     ��n   n�O��-�d���L�    @%q���w_�tPI�˗�o}+LM1���-Z�R�_��o��      �w  �4��Uo���zf��-    Pi��+���T�� *Nh���|���.��im:@Z��[������I^�     ��w  �p���fgd�Y�J-1�    IJQ}�D�����"�rA�G?�~�Ü�}�5 �LP_�K-zDvw�M�     ��g�   (v���r�ge:�d�    *���j��:�l[�K�:Κ5��dt01��f ?'3����?��5k�����=     ����  �]�~������n��,2�    �Ώ�=�@����Vx��X�C��-� ?����/N��vu՛n     �M�   (V�zЉ��/�yQ�-     !��;��Ue���i�B�[���lV��Pt,Z[��vw�n     ���   o�Jg�Qgx��f�    �G0:�	�g�(�^�ƭ�g���ݺ5$�� !S�u����2�     J7�   �dh���p��2�    �o��t�7����B*t�=���W[--�� ��L�A%ώ=��t     (=�  ������+GF~_c   ��##�� o�jh��]]����Q�I�= ̒�|�78��cǎ�m�     ��t   @�ٷ�##�B�     -��p��5��I��`9�ׇD���Z�n`J���́'�o�?���g:     ��  ��{���"�xT
�v1    (bA:�C۷����߀"&m[��펳f�����`j*0��� �e2���[�^�Lo�k�s     @�c�  T4}�:aY*��:M�     n��{�JWE�|}(2VΝw�vs������X�T"�-53s�۶͜���G�9     ��1�  *���FΝ�y��L�     n�Z�Ȳm� n�����M�\aY2�f��@J�����֭����     ŋw  P�tW�5z������n�-    ���\W�+W��; �$���d���y�����`j*0�`�I�L����nu������     P�p  G�8�~A_���t    ���lV�[��Mw �52R��5��x�双�"�g�;PY�H&w<�ys����M�     ��À;  �(��	'q���brr��    �-*��n�#C!e:��SX�ƍ��R�##��̹D�Tj�[�ԝ��c�     �� @�Џ=y�/���ͦ[     ��jl�UCw�@��JI{�R�Y�����~�L2�T)��͟�뮆�����t     (\� ��𝮮��������`�    p�d$"�+� f��F��~�k��(oh��o:	���2���M�ZO]��u�1     �8��V  P�~�wolY"qZOM�7�    ���g������u�����jg�j^`*����޽�1�     ��  ��]��]�N?/���4�    �=��d����t��'�Q��E��ɚ�e�K$��|��5�     ��R  ��ɣG�r��i}��J�-    ��$lqʘ���T}����Ν!�x�T���}�     n @Y�<z�.36vF�̬0�    ���o���,ڽ;{�j���2�`���~���h:     �À;  (;�c��GG�"��e�[     sǏ���T�p�����"{�D��J�= ��3|����'O�<    �
�   (+�c�����J��n    �1�D��>V+��n���t:�}�;����M� �c~����Q���W[     � ��  ��@WW�?2�<��    P!�@�[܁
#�Q~�h��3*c1^p���į$��?���,�)     `�0�  �B���v�ʕ�2�n6�    �?^<�FW�BY+V��G�q7mrM� �;�ڵݣ��ݺ����     T� @�=xp���xNf2�L�     �W����`2����F��ɚ�{e*�vmk|l�!w     *}  ���;;���ǟ��L��    ����q_�6��,��͉���W��6�BJ�9 怜��+1:��~챐�     0�,�   ���#�D�"�]`�    `Hg�
GVU���pҲ��|�c���~<��l��_�r��6&�����]���o�     ��  �$�;�ڎ�?/��:�-     ��x�7� �xX��v�#�vw���(C�����v��    ��ŀ;  (9����^<���1�    ~<�W �Ȳdh��H���R��<ʌ��ڐx�guW�k�     �>.�  @I�8�=�3���[     ����t�⣚���#��t���PN������h�>q�1�     f7y  �d�;;���ĳ��v    ���lV���� E�M����� �GNM�5���y����m     ��  �$$�[,�ǿ(2�E�[     �'�L7 (n��Ѯz䑪�=����,,P6�]��z����I�}    P&8� ���8vl��H��t��    @q�}� J�R�ݺ5��_���rʄ��ؕx����!w     �w  ��]������J-1�    (^:���-!� J��F��a�+��Ȉ/�6��ve2�f��7>50��     p{x�  �ɣG�f._~��v    �{�ׯA2�� PB���ݻ#���*UW�33�ȫWH<��4�     n�u  �(]��͌����d��    @iFF<� J�jj���<R�n��np����=�={��t     �u� ���ݎ��\<~Z$��L�     J��3���HǑ���F��ɪ*���nt�H����2�     nt  ��|��+�4���33+L�     J�?4�n Pڬ�6'���T�+W:�[ ܦ���=�3     ��c�  ��tuE�%�����-    ���OL�"�Lw (m2V��c�C��2��{ �:kl�ktϞc�     �� @QЏ=Z>:������t    �Di-�D�-� f�u�n�#���.�M� �u��د����/Mw     �g�   �'N8�7��SSM�     J���Q�ҥ�� �A�B�Y�֑��
�\�֦� �<)S�͏o�R}���oL�     ��ƀ;  0J�8��/\xFNNn1� 7E)�l�RѨ
&'�9   �9�[皎 PV���h�+W:�訯S)�܁�#��̖Om�b=�����c     ��c�  ��������brr�� �Vc���9�օ�+`���4   � ����CBJi:@y���r֭s�eI?g�;Pb�R&�;?�m�~���{�{     �;c�  �O�T�s� �]�i� n��d���x "��,!���%�����(L'  @ka/[��je:@�R�K��βe�?8��\�)w��H=3���[��������     ��p  F��e���z�n� pC����n��ᘽd����@e($���;>�?   �Ԃ�ji�Mw (_��J9k׺:���W�= n����߶m�To�+�c     �[1�  �]|Ϟ?cc�Mw ��P��*z�@�ټ9,m[��?W]�dM����Y�  `��,a�Y�� PޤmK{�J�Z�@y�/{"`�(!J&��>�cǕS==�M�     �_Ā;  �W#����H$~�t �'ۖ�]����QY[{Cg'����\�'�\�  ���m���/� �\P��j���N���P*�V:�|��۷��ٞ��9     �a�  ̛xG�'t<�1) ���z�9|8�,_���P���f��LO��  ��ΪU��F�� �A���Y���'x�(Rk�J��~b۶|��g�t     �).� ��9p����2���ɪ*�쌆;:b�����KJ�ȁQUW�y  � /�L7 �0J��=�D�ǎ�d,�P*
���H���G��3�     ~��5  0�F����Bk��8I)܍]��#�qf�LM�駟N�\���  �Y��� P�t&d����w�/� �"�T��ǛΞ0�    @�c�  ̩xg�^=8��2\�- �v��+��C��h�����gΤD��  �� c1Y���y�� M�_}5����}�- n��FGessg���c�[     �d�t   (_��&��?�p;��d��ݽ;}�᪹nBk�R't�����  ��t*���� L��ƍ��?\���x&� �N7cc��G�+0     d�   �)��y�=:���P�2� ��^�Ԏ9s��R�闭��f[��A06�p  �<�/�UC�� ����r֯wu*���qΆ@���$���ܵ���x���     ��  0�❝mbt��:��1� o&�aٳ'9~<����m�)|�}����*  �y���� B�82�gO4�T8Μ�h`LO�M��}Awuq�    �� ��J;�X��~Id2�L� ��9�׻�Çc���B��0���^��)��D>����  P�<O�w�2� ?�,w�j��u:��(f�lKJ�ͧΘN    �Ұ�  ̚k]]�zl�[��M�[ �gdU��9?�PT����@2U�Çc¶��  0O���@g��� x3Y[kE~��ٸ�5������������     *� ��Џ=���=-ff�0� B!��Mn��3f-\XgU;v�    IDAT�*��Az{�[   *���b����  ��?}��Z�@y�.y"�]�h�Rw~z��EO���t
     ��K}  p�tW���x�Y1=��t !���U�C�bΦM!iYE�1]-X`	��?<�n  ���Z�mm�� x;���rV�r��!_d2�t�w�Jm���͡�����t
     ��w  p[�ɓj�ܹωk�v�n��mmwv�T]]ўw��VKOM��+�   �B8�ׇLw �;���r֮u��L\��9(NR�R�?�m[���0    @�+ځ  P~ǲ���z�~� ���T��ᘳqcH*UT[�߆��-s��O��l�  �CA:��m�J�7"�
&-K�+W�VM��/_���!)gfv?�m����s�c     (g�t   (]�={������ P��Ν�أ�V[�Ͷ�%m[���h�A+  ��B'�� ���u���j����P�����ȿ�z��C�S     (glp  �dh߾�Y�����������ъ=Z�^�
)K�G2�VK��?�g;  �ܑѨ���l�@	���r���׮���T`��/�Z[~*���۷�3==q�=     �#.� �Mڿ�7������$����}{(�kWX(U�����|楗Ҧ;   ʙ��QΝw:�u���e��R�󯾚Ͽ�rF��� �D�n�]����ӧ{L�     PnJ~  ̯xg�^=8��e8�[ T&�p�ݷ/�-�M�̦���M����Lw   T��ɲ׭s�U���6��揌x��~5��I��EFG"�VK���ӧ�L�     PNp  7l��������E�5��I)�-[B����,�����:{�l�00��N  �Ҳ��l��]�X˗;e�;@Y��l�}饴w�gF��TW\ji9�+���)     �.� �:~�����f�M� �<��V���Z��e���-r� ��3�`r��|   �L���^��u֭s���t ���:���fs?�ANhm������5�w߇�ɓ��     0��  ��ZWW����L�� FJ�n��;;c�����/�-��v�;� |�t  @e�<$~��W󅾾��<m-X��m�(@q�RZK�:Vc��_��qn���d�SW��qj`૦[     (\� �w�O�p��?���֙nPYdM����Q�������gΤD��/   ��e	{�J�ݰ�U����N@�����/���S�@�--���`�    �RW� �m�����,�]�n�@eq֬q���d}�m��U[k�PH��/{�[   *��"��
��
��t6��:K�B�0J���Y��&'���5ގ�E2���[��������     J��  ��<�п�cc�Mw �2���{�V{{�mm;ٿ��t���;   �&J	{�2�ݴɵ�����4����r��}/+�6�@!���%K>����|�t     ���w  �F::~O��� ��^�����Ѩ2�R4�@gΜIy��lr  (B��Z96��M�������B�k_K�\�)w��v�[��mg���t
     ��w  ������W���К�� �m�н��ݍ]�孲� ����`z�O�  )iY�^��q7lpUk+[������ٳi=1�n ���Tc㱦�gL�     Pj�d  ���#�\���;�[ �?���
�������bLL��g�I�B�M|   EN��+g�z�]���/��W�Pйo|#]��)�n ��FG��K.��f�    �R;  ���~p���ӢP��nP����Ю]a���]�Xȼ�BJhf�  J��Jg�z�ݴ�Uuu��	`>��������Yΐ�y����������Λn    �Tp�  �B?�*����|�� �M�֪ȑ#1g�ڐ�����,�����L�   ���	���+�`d�S��TuuJ�x�ܓ��%���ly��}�=@E���;N]����     J�  @|����mj�"�j5���9�׻���H��,rkt���҅����<  @	R(g˖��v��ob �A_��gΞM�W�2����x����O��     ��� �
�O�p쑑g���J�- ʗ�Fe�����ukX*� ϭ�ֲe�劧S)�3  Pbt6������+y��h�p�%]��� ����n�����`b"0�T2�N����͡�����t     Ŏw  *�����L_���t��e���ѣG��ŋm�-�@*%�+�BOOA���  �"��Ȉ��J.���UM����2��<I���j�#����g��`R�R۟ض�����4    @1c3  ,�g����#�; �)���kW8�cGHH��c����~�٤���<  @9��,�C;v���v[pw`������/f����4`��,O��>�|���L�     P��$ �B�vt<����֚� f���Q���������9�]��ϼ�b�t   f�Z�@9[�����]�gv �.����_�rJ_��n*��Tk�5=����S     (F\� P��<���>���L� (?���N��""R�[*A�o�6���s�;   0�d,&�M�B�]w�d(�]>�Y��� s�l�O$�,`��D&dKKG���c�[     (6\� PaG�l���(
��� eƶe��{��ƍ!�)FgΞM{/L�   `��t7lpݭ[C2�%R �'t��HΝ�<	"kj��������     �	[[ � �~�!;8����jM� (/VS�;~<f��9�[*��W�p��O���t   f��d�/��'9��j�B��� f��Ҿ�G!�x�3�T�\�>���S�.=g:    �b;  B?�Xh���3"�j5���H)ܭ[C����2a��!Ҳ��|�]8w� <f   ʒ��O$|�Wr��끪�W2�78��%��V�Z�Py��=@��d�>�eK���M�     P,p �B�N,�����f� ʇ�e��3�l�R�A�0
)���*\�P�E�   eKk����W^��㾪��T4ʠ;�ۢ��-����
�P0�T�dr��m�6�����h:    �b�
   �w��$��� P>��f+��S��������r��f�t   扔�^��	��R�ۦs �6�J�^H���o��4Z���|�o.>}�oM�     `�  ��������%���� n���ݲ%z���B)��R�r��V:����Mw   `I)��˝Ю]��-��t����^_�܁y&��i��x�����-     ��@
  el�ȑ_�\�s���� �O��2������-xA�3�?��\�L�   `����v����E�tp�t�������ﳦC�J�c�x������{�t     �0� @�=xpE0:����M� (}vs��舩�je�7(�R�<����)   0�no�ݻ�X�� �����g^z)#<O�n*���{���ʓ'��    T$.� (C��訩��|Nd��[ �8)��uk(�T����ۖv{�]8w� |�t   ����k���q�Z�В�(���U_o9mm�70P����rd���k��O]����     L`� �2�O�T���y��*�- J��e��3�l�R���$#e54X^OS   ,��
���ד���h��˫ n���RΪU�w����Y6��D��k߶M������     ��  ��a��^OL�c�@i�Z[����Uj�"�tn�Z����-�+W<�-   0+��򯼒��d�/����"+�"C!�^��$���C�����m������^�1     �'.� (#�>%��~�t���n��>���P��B��ٯ=]8w�M�   B!-K8�׻���a6��Q��t���^?�K`��v�Z��W�{��)     �V  (�VCC��Z� ��uet�ވu���́ Йg�Mz##��   Ǒ�-��}{X:� �7�u����~����R�Hd�ji�h:}z�t     ��j  �@�ȑ����3��[ �&U_�"��Ԃ�$S�t:��~:�gf�-   (.2����v7lp��<; �򯾚���_g�֦S���kjz[������     ��+  ���?ܐ��|�� ��Y�։>\�b1e�sK:��[[�¹s0�  �7)�?0�y����J��z%X��]X����h�*\��q�����H������M�     0�p ���.wrx��H���nP�������;*�bp�B�XLYuu���+�n  @�љ�.����AO��[���a�#�`�e/]j{���y�s��'���Ol�\s���e�-     �%� (a����_���f� J���V��Gc��U���?�p�%�@��o�   �)��х�_�W��vS�%C!��-U]��ի��eOg��tP�R��>�m��gz{_3�    �\aK#  %jd߾�GF~�t��c/]j�;:�2a@����/���~6�  �]I����nh���9G x{�l�~ᅴ?<�*w`�i����֏��=�]�-     �� (AC�����֚�� �qR�Ў!�}�)9@�BAg��Ť�*��  �d8,�;B���!�g
 o��:��250"�	����t����     f�  ���C�Vى�i��W�nPBGF��X+V��SP\��� ���3:��3�   �!j�~����wp� �VZ�췿�-���9�)@��uuo456v��n�     �
[_ (!��Gc���/�lv�� �C�թ�?Xe��8�[P|d($���;>/43�   xo:�Յ��B�Hx��Ŗ�D��& EDJi��;�u�?8���Z6�(i��.^|�t
     ��w  Jȉ�?'��ך� P:�����ѣ1Y]�o�#U]�dM���   ���tPx�ռ��	�K�6_��sVs�m��)���/TsG��k>�m[���0�    �la� ��ط�cc�; �)��sg(��CQa�lS�{�,��~"�'�  pS��q����y
Ik�bKHɠ; !�����-���A`:(WR$�;o׮>y� �     f��  ���>�����К!U ��qdt����b�k:%Fk�9s&�]��'�  pK��F+t�}���6��x�##^���S:�c�;0Gd8|M.Y�����1�-     �.� (r��Y�='
��� �O-X�"��T}=_k­����O'��)V�  ��H)�ի��#�����!��]��gΤ���M`�蚚ޖu��?����     nC/  ��vt��_������nP�����ȑ#U����:ۖ��e�w�|A���   ��`b"(��Z^h-��fKH�����HD9+W�ޥK��f�����-L�r+N|�t     ��w  ��>yRٽ�ψ����[ 9)������>����n����h�U�p�m_   �uA ��!���-�*YS�3	���PH9�W;�А�S)�܁9 3�U�ڼ�{����[     �U\& P�~�q�P\���� �MZ����u�+$�`��F��Y�q��g�   �Mg��p�|A��VK�ŋ�@e��#�;�t��q?��
L� eH�Lf�v���S.��    �V0� @>p�a�H<&V�.du��?����-(OVs��S� �M�   ����~����"�Vc�%�� *�TJ:�W;zj*&&rf�֖�f��]/<u��u�9     �,.� (2������2��x�--V�С��D���� Й�Kz�8C�   �5֒%v��"���E<@%�Z���L��W�S�r$kj��֭��'�-     �.� ("׏[荎>#���- ���v�9x0&]��v�=)��b�S��-�\N��  @y�33A���"��֒%�T��<@%�R�˗�B)�y�s�����'s�5�^0�    ��`� �"�O�TW_��L.7��HI)�ݻ��{�
�?0���Hk�R�p�\A|9   �DkᏌ��
V}�Ruu<� *���,�e8,�+Wrf��d�xb�V�T_��M�     p��, �H|̶�H^�v�� E�ue�����aC�t
*��F��Р
��|�   �+�Ӆ����u�Z�Ė���@���l��N����0��L�v~z��ן��0    ��`� �"0|���GF~K
�\ o���T���*���6݂ʦ,����f�   f]p�jPx����F�Z���P�TC�e56Z^o/C��l�Z�L��Ƿm�ʩ��i�9     ���  0l�С����_�g+3������ȁQ
)�-�?љ�|%�����   s�^��=�@TUWs*�?<쥟>%
�܁Y$��/6�����y�-     �6� `P�ر�2�xF
U�[ g�7�T8(&�^���<�N3h   �9LM�W_�K�VS�%�daPATM��[[�BooA����|��f�Z�����M�     �np �}�J�;��L��nPd������=�D�@1�JIk�rǻp!/
,r  �	�_��������b�H���
�����l�������ʆL�W<�m�>���=�-     �� 0���kq�ꃦ; iY"��u7n�nލ���d��?��E�   �;zf&�^{-/,KX��ls*��Ŕ�|����x��=2����;~�TOϐ�     ���  0���!�\�c�5/��9YU����Q�x�m��Q�����K/�Mw   �2X�Y�}��j�B�T�
LM��/})�gf�-@وD��mm�wwO�N    ��q �<�8�.FG�\�~�t��a54X��ǫT}=��QRTC���y$��   �?�Nk����¶����6w�B�pX�+W:�ŋ���1`6x^,�zד�.=c:    �_��  �HwuY���n�N7�nP<�e�����U*U�[�[a���zl���ؤ  �����\��A�Z�Ė�0g)��PH�+W:��K��2����4r���S���6�    ��1� �<:�����ڵ��� P<�M���}Qi�lD�R�˖�^?C   �7�̌�^{�m�@��+�ի��eO�Ӝ?�Y S�͟ޱ��'{zL�     �3\� 0OF;;�._�W���B�D��"�ƍ!�)�l	�����O'�\<   ���bG����Z� � �2�?��FF|�)@Yp�����K���M�      v  ̋�ǎ��_��%�y�- �������Q���1��6p��>s&%��t
   *�m�н��ݍ]�����\Ng����{�[��P[{���ȓ'��    �&  �~��tOϳ"�[h��y2��c�bVk+��(K��֒���/_f�    �+�?0������fK�a�(cҶ��f������4�����f�]kz���o�N    �w  ��oUU�����h��y��N�>��*��`�n���d�L&�GG�T<   �]05.\�[Z���� @�JIgժ��OM1��&�N�{|��˧zzΛn    T6.v �C#��}�t ��+r�x����78*���n##~p�:   ���(�?_��d`���R)���J)�^�A09��=R���~b۶�����    @��B �9r��s�58��2\�- �rV�v�{�F�e��Eg2A�駓�!w   �jkUd���jj�kZ@9���W�^�t
P�.5/Y�Wvw�M�     *�# ��G�����ݲP�6��,w��P��#�m��@�q���fΝ+��w   ��s9]8w./�vK�%��|�#)��r%�܁ِ��%-�S/~�t
    �21� ��DS�����J� �R��w�C��+���P�d4���-���z   0Gk�y��o����u9��蟆����LM1���N�||۶ԩ���n    T� �e#����;h��9ҲD��#�n�2��`�%��Аg�   �M_���C    IDATxo��WuuJ���(GRJ{�*6��O�Tjקw�z���L�     *��  ̢xg�^9<��!�� f�pXF������-@1��,���dLL0\    �|_x���Lv{�-�b�;Pn�i�;C��m�����]7~�O��r�s     ��w  f�@WW�58�_��GL� 0CVU����U��Ŷ��I{�
ǿr��ɤ6   ��~��߳[[m��� (7���P���6<50p�t
    �r0� �,�]]Vfd�9�N/1��U_���P����76�N����N��� �y��  `^&�o�Q����yY(7��B���oۦN�����    @e`#	  � 15�o���Mw 0�nn��]]U������{�Ѩ�<��   �Hx��}��׾���@�QJF��+V8�S�R&GF~g�Сݦ;     ���  n��ѣ{�ß�BH�- ���n��������UUJ��*���`�   ��`b"���
Vk���Q�x@9�R:�V9�ؘLM�"p+��D>߇7mz�O��r�s     �w  nC�ر�~<���"�[ �?g�:7�����.�MR��<폌��[   ���٬��x#/"i56ڦ{ �")��z�\�����@z^�:�����i�-    ��ƀ;  �ᓍ���d�� ��ݺ5�������v��mmv0>�`   �������L`���R)�}@���&w�܁[&���Ol��}�����[     �w  nQ|���U��0�`�I)B����}!C�����?0��tZ��   �,����Z�Ԗ��2�`��l�}l���rn��d���]����[  ��ٻ�8�����k�}�[7[2�dI�d0&��l|� _t�`
�&iZrNZ�6��4�$GI?INOj�i{.=9-m� �)���KJBp�M��E�-K��sifϞ�{�u^�$�o��ѳg����|~oF�k��� ���, ��c�w�7�?�8ϒ$��uW�|�u��)�/�R)���[��UF  �9��h:�яNw�|r>tp%I\۽�Qܴ�:�4��GG�����/�N  �?�� g(���c�>��ϯ��G�b\߳�Q|��ˡS��ĕJR���B���;Qn�;  =&ˢ�Ov���x��(I΄~�$q���K�i~�M�p���WMw:��w��C�S   �?���ϫW8?y�Bw �Q�7��6m��H�re!����ȑn�  x!��H�=�-\zi)�T�C?H��x�e���g�y���5��|f�?��7����'��  ��b� ��Ў?k6�v�����ո���7�����+\|q1j����LC�  �ɧ���c��.����\��X�K�yM�����hv֐;��8��ݾ��z�~���>�  ���� ��b���˳f�Cw �O�lYRX�\|q1t,����Vܸ��  =+o���'?93��#�(��B?�V�ƽ�6�/���P<?�,������~   8gl�Ӑ������B� �G�re�x�;ɪU~3���qi˖b�СN�n �7�y�=��FG��-��P�C'�L\*���.+u�Dss�G��sskf&'��w��WB�   �����pb|���N���8?�ի���e���!�j5���ۈ�eCB  ���C���>v*��LC� �\�lYҸ��F�l�o�p���~�����Bg   �����qbϞ�������QX�����hč���Pr������(6� @o��ǳ��~t�{�H't���+V�4�j�)��<�剉��V�n  `� ^����c��c��VC� ��qc�����R1�= ���B\,F�ѣ��-  ��4�>�D'ʲ��qc1�"����ŵZRܲ��}�N��H
�+�v��8~�}G����-   ,n��E�&�o}��|ffC�`�_��RmϞF\,B�RX���OMe��h�  ^Nz�x�OLd�-[Jq�x��E,�ד��s�WB����jm���^���SO}=t
   ��w x�/�Fccw�� ^鵯-նo�G���ŭ[Kٳ�v���<t  ��ll,K���l)ŕ��LXĒe˒Һu��Ot��#)���պ�g��������  �┄ �^t|��[������ ^�u�+U��p;��$���w7���=� �(���i�#9��8���2Ɇ�ھ}��`o��4�����>��*�S   X����0���th�cy��,t��ʯ}�z��(��C��K���aC���c�� `q�v�����+V$�5k|��E,Y��PX�&�<��M�p��Ng���٭<|���[   X|�P���������ׄ� V��kʕm�jQn�E"n4�ªUI���:�[  ��y�=t�u�yq�Ƣְx%\P(�Xwv3���������~��'�2t
   ��w ��;v�è�|g�`a�o��R��zd��d��B�eyz�D�  NW:8�f�fZܲ���Ea�J.���JQz��!w8q�I�}�?�����c���  ��a� ��Ğ=WD'N�z����-��)�xc�r�-����+n�X�FG�lb"�  �+���:G�tK�7�J%	���ºuŨ����A��t�i9Nӛ�;z��C�   �xp�(�������Q�}Q�`�Tn��Zyӛ����l)�G�t�V+  �mv6�|�;�����d�rC�H7m*�33y6<l�N���E?s�u���z�C�   �8xy
 Q�����ԩ��;��Q�o��o��:87�R)���ۈ��8t  �����g?���Ȯn�Z\���Zi����i������ׄ�   `q0���wlϞ�
##�
�,�8�jo{[�|�5��)���,_��v�l��� ���i�>�Pk���Q���$���v5
�\b�NC�e��������R�   z�)  ��|`�<=4��h~~e�`�qT��Z��C�JV�H�+��C��-  p��cǺ��t^ܼ�űۉ`�I��x�e���g�y��
�������ݵ<t��S   �m6���NL|(��Y�X ��a�(]qE�|�5��  p6:���O|b&j���-���+���o_#^��wW8I�y��۷��   ��y������]�����;�`����[�R+n��Zx  ��������O�SSi���ōFҸ��F�h��^F�����}�����  @�*� �&��_�7��%�vk�[�s�p;,Mq��n-v�z���ۮ� `��������ƍŸѰ���RI�6;�?މ22�K����t���#G�  @o��%ivj�����Bw ��vX�*���o_#�Tl� `Q�[�|�f�g��n�\�W���5�c�r��ѻN��yo�   z�w ��;w�'�9tp�n�(JV�*�v�G��]  �n7o����t����)��+\rI��}{=�����GQ�����w�{M�   z�� ,)��������o����-�9d���ʕ��T�ңG��[  ��y�=|��y^ܸ�:83Ʌ
�F�=r�s)��n��Ͳ7�맟�x�   z�w �����ߊZ���;�s(�����f��>�u���L���[  �l�Ǐ���LVܲ���A�b���U�(����qC�����?}�����|�OC�   �;����q|ǎ��''_�8��8��}w�x商ہ��~{��~���  ,j�o}k~���mEi��n�L妛����v�(�����ܵkk�   z�w ���.����~����v���W�H��$���w7���=� ��u�z�3��OLG�v�83�m�j�͛��;��u������3t   ��G~ �^>0P���(Mmx�>R��Z��]/)�Ւ�޽��X�C�  �+�=q"����g��iC$I\ݹ�Q��"7��K��z����,t   ���; }����/G�Nm	��;��n�����p;pZ
k��;vԢ،;  �[>6��x`:��LC� �/.������x�
�f�%d��ox��kBw   ��( ��c�w��� Νʛ�\-_w]5t���n-�o�ѿ  ,z�ɓY����QC��zR߷�W*N_Ë���������_
�  @X���o��@e���>w:+B� �F�曫�n0�
����|r2��Ʋ�-  ��t:Q�;��֭+�+V���D\�%��������<t������:��?x��B�   �� ���o��ĭֺ���Q���J��e���+w�Y/�Yc  �ů��[���L���N���֯/V﹧��ËI���qd��m�;   �G} �����{�E�����]W��v[-t���I�l)u|>� `�����S��ʕI� ',��Յ(���رn��QI)Mo�;?�C��  `	����gw��h����ө�n^���W��۶�"V�s$�T��%�����+� X��<�>܉k��p����9��)n�Pȧ��ld$�=��i4��-�>���)   �I�  8�.N�峳�Cw �\����;�0��s��k����  �<������o|�:8mq��;j�K/u0^�����}���  ��g�; }ex���i����aXX�J�_^��uW=�c���H.�������Аmy  ����n��yq��R��4�q\��Rz�H7o�\1�g��7�{�Ϳ����n�   �� �?���Fub�7�N��xe��7k;w6�$1�,��M�|x8�&'��-  p.�Ǐ���\Vܼ�Y=/.��e��:O>ى�����t��ō�>�P�   Ο$t  �+k������5�;�W��iS��g��v����z�=��< �7�����/}i6�"ò�čFR߿�W*އ��slǎ;Bg   p���@_ܽ{[wdd{���)�[W���m�8�*���w�A  ������|�󟟍�ܐ;,Ʌj�vգ��[x�<O
�����)   ��� �J��顡ߎ:��[��WX��P��q��+p���jR���B���;��  �D62��'Ofŭ[KQ;�	=.Y��PX�,�>��=��Y65;����|�   ��! ����_�[���;����Z��hD��ߧ@0��K�7���  Υ�c�uf?�V�eNr�"P���J��km��Py{s߾[Bw   ����ݻ�-������ً�/Ojo���^���|���__�  �R��!CTo��Zܼ��zM�������)t   �:  �V>0P����Y�8;q���wY�r�ߥ@�(^zi1L��'��-  p�dY6<��.���q�x	q/���9��[-S�{ĝΊ����>���-   ,[2X��&'%n�օ� �N\�ĵ�%\`��-IWw��+Vxf ��t�~�;���36�C�K���wo=�VH�P}����ׄ�   `��X������7���Bw g�X����7
k�nzR\�%�={Q�d�  ��b��x��Bm��F\�
�W���tx�C����   ���! ,:��@afx�������-������wo�p�%��- /%�ד��Յ�OvB�  ���MNf��pZ���R�uBK�/O�+��C�M�{�ϯ���\~ߡC_	�  ���D3 �Ή��_���7�� �BG�;�6m2�,
ŭ[K�n���  �s�������?m�;,�+�(�����zM�l��yｯ�  ��g��E�]��OFF��8;��n�������LTn��R��
s  �;�#G��"Q��jq�VϦ�=�,+eCC�4�   �g
� �t��ّ���ss�n�\��+�n�X���-����n>=m� ���MNf��HZ|�kJQǡ{��qq��Rz�H7o�<��_���`����}O=���S   8w�d`�<y��O��4tp�JW^Y��|��v`�*�ڞ=�x�2��  ��Α#����^+�sC����R)���S��U�Q�{�CCw����Cw   p��0��0t��U���Cw g�x�e����V��ȇ7`Q�����kW=.� ���y�N����C��W�(���mx6�����:  �sǛ z^~�`2��o�v�n_�83�����{Q�n�B�lY��\�t�z��  εll,˧���֭��Au�Y���I�bE�=tȳ)|W<7�槯�.�逸�8t   ��w zޏW��"�3tpf
k��4�RɭA@_I֬)D�n���[  �\�FF�|~>*^zi)t��
k��Nǳ)|���k~��o�̿~���)   �2�� �i���_5�����d�ʤv�@#�T���R��[��͛��;  `!t}tn�k_����ʛ����W�[�O��P�   ^9G �����FiZ	����Z�k��7�z�oM��q\ݹ�QX���h  ��������7ڡ;���qm��z�j��p�]����w����   �2^v гN����xr��;�3P,Ƶ}�ɪU>���Jqm��z\�ơ[  `!�}����G5���RIj{�6�rٳ)|Wwx��&��_�  ��g���4>0��{��oD�n5tp��8���U/l�X
�p�ĕJR\���y��N��s  ��K���/���.*�n^X\�%�/L:O>�	�=!M+����9���)   ���I����{�nۮ�He۶Za��r���-ٰ�Tٶ��  D�G�_��l����C� /�p�e���X	��"������Bw   pv��s�xs::zW����o��R~��}@����WW�ox�C>  ��<��=�J�}�vh�a�[n���lq�DQ�yR����|`���   ���9 zJ>0P898�[�����H����T���ZEq�����6���4;y2�  �\�G�'��7m*&˖Y��).n�\�>�T'o���1Z�鬘.�k�:�?B�   pf�����<�s�������)l�P��uW=2�EI�v�'�Vy� �?u���>5�ML��S�Q�$�={Q��}DQ��w�&t   g�Gw zFs׮��������x��B}��z�$>���j5���ۈ�e�6 З�v;o����d�N��zTrᅅ�]w�Bw@OH�Jiz�_��   ��p�gd�ӿ�i%t���e˒��}��R�{�$\P�m�^�b3�  ���ԩl����gg�C�*��5����{�Qe���5��y_�   N��$ z�;ߓOL�!tp�帾#Y��oI�Qܲ�T���j�  X(��d6�;�3����[�V���jq��b��ݡ����;V��   ��J �?ޱcE4:�OCw �!I�ڎ�d��B��^W���J�u�+��  ��������~v&�2C�Ћ�8��sO=^��7a��xnnե���  ���e �m������^�xy�m�j�͛k���z���u з�G�v۟�|+�"C�Ѓ�j5���ۈ��8t7:�����7��   ��p ��{�ޚ����xy�믯�����`QI���{w#^���7  }���t���ڡ;���^]��uW-t���y�01��zO  ��l� �|`�0�l�V<?o{;���֭��w֢8��	�ťR\ܰ��y�N�e�s  `A�'N�q�.���x�d��B>?�gCCi�j~~��ɓ���z�C�   ��L ����MOo������;v����䢋��� ������������������%�8��7�?zb��KCw   ����О=[������ ^Z�lYR۳����^��嗗�7�P	�  &ϣ��~��uC� / I�ڮ]���𮏥�ۭf��}�3   xq�"=y�CQ���^V.����q��7#�9R��j��J�;  `��i�~�3��x�x��VKj;v4��+?��d|���v�|g�   ^�7 �w'v�|O<1���KH���cG=Y��:����{�֬��+  }+���[���L>3��n��p�%��7VCw@h���?����F�   ��u :h>    IDATΫ?ޱcŊ���/NS/ϡ�Un��Vz�kˡ; �Q\(ą-[J����:��9  �0������n�+�q�ġs��Wܰ����Ԕ�(,]�nm:�6�w��C�S   �~6�p^m�t~5��[�xq�k���������%˗'�ݻq��s  �W�l�s���L��y��y�����x�rߋY�����G��!t   �� Λ�����GF��� ^\q��b���ܰ p֭+V�m���  ���9r�;����<_\�&�]��_���y^(ML�j�   ��w Λ��ؿ��ܛr�QɅ&����Q�6�<)^uU�|�5��  ����5�x��⋋�[o���%-?y���w����   �� ��w�|w<5������ո�wo#�T�>8�*��V+n�T�  i�K_�M�y��x���VJ�_^
�!%���h|``e�   �c�	��G�dt�gCw /"I�ڎ�x�J7, ��$qm��z�j�gt  �W�E��~������S��+w�QOV��\ʒ��ͭ�NM�  �s�� `�m����y�}a���U�m�6m��	 �J%���׈+�8t
  ,������O�䳳Y���ŕJ\۳���KY����=C\�   � ,��.�FG��� ^X骫�嫯���  ��U�
�]��Q�Q ����<������Di��n�_�zu��ַVCw@(y������   � ,����_���fh�A����o��� �o6n,Un��0  }-J�_�B+�"C��c�W]U)��u��d%SSW�ع�=�;   �:� ,��{��O��^�x�d���[�]9�c��]W-]uU9t  ,��w�ә��7�Bw �W��z�zu!t����t����    /& X��@yvp��y��,t�����w,K�/�[�G7o.fǎu�S�l� �o��>�-�Y�$^���8I����c�u�,��_�[?�n_��Ç�:  `����q|j���V�U�;��Q}��zr�>��$���w7���=� п�<j}�s���x:��|n.O����s�/|��~�V�e]�d�##���_�  `��C �N��yi48��(M]�=���7W��__���IGG����OGݮ�  �V�bE�x����ժ�p>��e��D����Y��f�f����Q��������җ�:  `)2��97t���gcco
�|��_]���U��XT�Ç�[��tˠ  ���aC�~�@#J�-��[�,I��f��i�����Y�.X�8ΣM�~b݃���-   K��� �S����9w��o��=%��¤�����T�	���k�s?<�  R��k+շ����<ϳ��,N���4{n���vZ^�z}h�ƍ��<��N  XJ�� ���@�ıc�d�zK\���}������7W��������-  �P:�>:W\�:)^ye%t��������4���neφ��yj�ιVk��'�YE�:  `)1��9s�{~.|��{�qT߿�Qش�:�W&�v����NGGM,  з�B!����
k�Z�Q峳Y6:��V����٧��(��Λb��^v��6>����)   K�w Ή#k+�)�t\!=�r�m��u�UCw pnd�Ne��}�T�j�d  �oōF�x���ǍF�Χ��ʲ����l���p���>7�_t�W�����p�  ��; �������󑑷�� �F���K�;��| }%��~��Ӯ� ��֯/�ｷ%����<ϳ��,N���4���ǻy��03��8��֭��-=���)   K��� �b�}�nI�~���<�Q	zDa͚B�]�Z�~����w�3?�{��
�  �t��[���H�����4����4m6Ӵ�L�n�0;,6˖]w����ݬ   ���� X�ґ�_1��#�V��޽u�� ��x����p�y�ѹ�-  �P:�>:Wxի
�+�(�n�ӑ�����D����Y��f�f����Qn���������'�(�w�S   ���' ^���;2;v�Bw ��Q}��FaӦR� X�����9��  %.���޵,��"K��)y��e##i��L���4M��)[��ߕ���-o����S   ��w �������#G�0��_�xN�[��n��� �<���f�:��0D @ߊW�H����ˢj�-��y�g��Y>>�v�Ʋlx8M�y�e-;,U�z�g��?:  ��p��}��w���� �Sܼ�Xۻ�ű�x KH69��>���|n�p  }�x��ھ}�{���,Ϧ��bN�f3M��4�v=o#�����{.�ԧ�:  �_y	�Y9�s������4-�nl2X��g��>�ə(�� ��U~ӛ���nrs�F���##i::�f##i�l���d�
8�<r�W����   �ʀ; gep۶����7�� �(.���޵,��b� �ѹ�?����  �`�8�8�(l�X
��ⒷZY62�v��4O���,K��bv���q��6����\�  �~d��3vl�g���(�m��P���Z�u����  �������_̇�  ��W�q�=�Y�,_��$ϗ�y69����iwl,ˆ��tp���Z&فs��8��{�<��  �s̖O �X<9�K�ۡ7����l���Rݶ��MLd�c��-  ��v;�{衙ڽ�.���"��,��lj�!���4m6Ӵ�L�n�0;p~��lh~��?E�o�N  �7^�pFN�������_�DQᢋ
�w�kYT(�M�_�gg���}l:?y��0  �V��*�[n���������lb"MGFҬ�L���4I�4�,u���ȪU���s��	�  �Olp����ğ��?6I���j\۳�n���jI}������OG��ͅ  ���?�ӹ�ڵ��֭��-�[y��e##i:6�f��Y�l���X�o��n�ZE�KE?:  ���ഝ�瞟�����8����5
�^�. /*=|x���O��  Я�J%n��������[8y����Y6>�u��4N���n�jy��Ba.}�������C�   �� ��g.,>�?�N����ʍ7V�7��
n ^�������v�  X(�u�
�w�cY�$�y��,˳��,N���4m6�tx8u��/�.��K~��,t  @�(� `qH&&���v��aC�|�M�� ,�o��i�;��n ���L�_�j����X�+��tt4KGF�ld�����i�e�� L2:��Ğ=׭��GB�   �� ��c;w^��c����qm��z�6�p���wֳ���th(  ���sō��-[J�[��������;1�e�f�5�i:6�F����Ғ�y!����(���n  ��� xY�۶}<c�X��8�8�(l��C- g,o����~t:���2 ��W�q�=�Y�,_��n�Wy��e##i��|n+��P7��1��=���|�wCw   ,v�xI��woˎ�p�T�����7�����+�>���<�� ��Tذ�X��n�{��,Ϧ��lx8M��Ӵ�L���4�t�����8���{�<h�   �+P @o�'&~�p;�Uܸ�X���J� �d��b����=�
�  !=v�;��:W��KNS�����X������h���e��P��X���̬���"���  `13���:�k׏��>��;`)�������.��u�kpN�}�������\�  Xq��wY�K,y�y�����iwb"˚�4k6�tl,�r��Υ�Z�Z������o΄n  X������G��ή�KVG���K�S �+�����wB�  �B��/O���=ˢju�.�[�,I��f����P7��1�p��_|�%���?�  �Xp���_����KY�[���`!�N>�_��t::��n ��P���RuǎF��ey65�e��i:<�fcci�l�y�m� �<I�7޳����n  X�\���8��g����⥗�7�P	�@�K���{w}�#�����  �w:O<�)n�4W��ʾy��w:y66����i:6���f�u�ԹU�^gY9o�FQd�  �Y0���'O�r���Bw�R7q��{��v X@�ʕ���Pi��ߜ�  a��_n7֯/&\P�r��V+�FG�td$����SSY�;�
�X䣣�5����O}�B�   ,6��>C��]�?��>�@ q��jI� �_��+� �[�n����k����eQ���"���ʲ����l>7��l���t��W(ϓt|��(�:  `�1�������<��F#��7��R���R� ������k��P�  B�l��_�z�|���o���<����z#���s���}# �jj�;w޻����o�S   ���V��7|���;��f�Da��B}`��7���������??�  LG�w�cYa����)�t�|r2��ǳ��[ٳ��n�:[
���Ɖ�������A�s   �&��k���_0���Jqm����v η�嗗��|����	 @����ϵ��}��T:��^��tb"KGFҬ�L�f3M���(��(�gf�=��GQ���-   ��* �(���v퍟}�߄��cG�x���� ,M�/~�������  �t���w�_��G�je��H�m6�lx8�FG�lj�F^ ^Z�6�nӦ��p�  �i���(��(������T����l����W^Y6� @����_Η�l).������y�MNf��p������X�?���mk�8s��NO ���N  X�5��y_��3�Cw�R�\pARٶ����+;u*��ַ� �$�~���u�q������w�y>1�f��Y:<���f�6�i��f�����~���-<0�  ��pX�������;`)����}{=.��- ,=y���?��\�ߘ�S�c �4��v����Z�M����H�6�i69�E�Yv V�n��r���DQ�/C�   �:�T Kܳ۷�d�ĉ�
�KQ�o�������%����}tn��G�m�   8�J���֭�\��S�S   z�� KX>0P|�	�KQi˖b��kʡ; XB���G��{�����1�   p�u:�٩�E�?�  �˒� �3x��?���Cw�R��q宻��t 8�n7���7���𩹇�3�   N<2��鷿}]�  �^f�;����}��=��L���W��z\�9h������c��}m.���B�    EQ�V�'O�|E?:  �WpX����~>��_�����P.n�\
�@K�y����Wf��	��    =&���k�֋?�á[   z�w�%h���W��<�?t,5ɪUI��[k�; �_��P��կ���ǻ�[    xaq���V��(���-   �(	 ����<�Q�[�KI\(D�;�q��n��d����>5=s��ӆ�   ���ۚ�����   ��w�%�Ğ=��g��ۄ-�_�o�&�z��^ �[�v6�'27��o�EY�   �Ӕ�y!��(�B�   ����V��,+�΀���~}�|�u�� ��4��y�}��>5��#��   ���76��%t  @��E`	yf߾��~��<t,%�R\���Z�.N �\��C�:�����IS�    �Y������EQ�;t
  @/��`	)MM�b�������\���W,�x`���O��   �|r��={v��   �%6�,G��!:z������.��T��r� �lz:���?nw��/�C�    � ��&���:  �W���D�����(����I�lYR���Z� �4��~���O���v   ����:uٱ�;��  �WtXF��3���2t,%�;�Eժ�Z ����g:��応�����y���   `���8?x�w  �(��� Xx�����y�����W��^Z
��Ⓧ���/y6=v��   ��'��Y����,����  �ӿ }nh��=��S��"^�"��v[-t �L���}�˭��|��v   ��)��|`��   4��\61�S�`Ɉ�v睵�Trc �+�>�x��0��Zy�    gg�4���nd�;  �����ǎ�ڵ7:ujK�X*J�\S)l�X
��␍�����}衖�v    �(�򉉿�<h�  X�lp�c���O����#Y�*��rK5t �/����~�=��o�EY:   ���Z���?��(��C�  �P���S�v�|g>=�9t,	qU﹧�q� zZ�}������͓�<b�   �����}[� ���w�>ON����T�o��RX���* ^T61�������رn�    z[�j�z�����á[   Bp��ݹ�������;`)�W�.T���j� zT���<�n��o�2�   �i�q[� ��ʦQ�>T�������ąBT۾�%I��ޓ?�m��ﷲ��,t    �K�j�y��E�
�  p�9��gN������)���<(�pC��fM!t���޽��Y�w޿�u�! PP!�B�A@��TZ�l�(ۖ��ֻ7me�N{ߏ:?�o�{,�� �L*��h4*2:�z9ه�ֵֵN�����-�������_��e�\;�}} #��-�_�z���-�v    N�`~�/]q  ��� &;�i��a��S��tS=v �e����:O?�	�/�   �Դ�����$I���N  XM� �ȶm$�]�&^���v��k�R��$ $I�$E�Yt�~�=��/�[    ��7�����  �2��
`�,.>;�A������  I�$a��������q;    �-Ͳ�ٱ�Obw   �&�,�	�����������n]�~��3�; �/4�����38xа   ���t�$���  �Z\p��c��� /M���|䴤TJc� Q�������M�v    VZ�e޶���   ��w�	ph��������IW���z��<?L�b~~����=:��   ��HJ����   ��w�	P^\���0�Jg�Y��r�L� "�������}Ӹ   �U�e�{�w  `J�@
0�^���'8�!vL�4Mf����RIc� ��\m   `T\q  ��� c.,,�M��t�-[����׋� ���v    FI���жm��  ��� �ء{��pz���!vL��]�*�o�u&v ��X\v��m�1l   `d�?�$�bw   �$��X9���B�&�̇>�&�V��L�0x��n���2n   `�Z�_ݱ��   +�w�1��Ν��WZ��ʩn�T�\rI5v ��h�����������-    �V���_'I�H�  ���;��*?�&�};���^O���kbw �:�?�Y����5��   y���#۷4v  �J1pC�}�c������0�f�c&=�4�J .t�!߻��~�v���    �G�����   +�h`��?���z;������ʕW�bw ���C����>���r/v    ���h\��Ν��  `%Tb pb����N8x�f�Eae��rR�Ї�$I�%�IU������}��OU    ��|~���$���   ��w�13h�?��J�Bj��:S:��r� VF1??l?�p��o�q;    c-]Z��Ў���   Xn� c�q�����?�&U��s˵�[�; X�����=�pk����-    p��$I+Y�cw   ,7w�1�<v�����VB�&3wݵ&)���) ,�����_�:_�j;�m   `b��o:�s�U�;   �S%v  �煻�^[���f�+��eK�t��� &��ȑA�_m�f���    �-�Tm��.I�O�n  X..���w��_�^���0��3�(�o�u&v �(���z    IDAT��w�������   �d����Gfg/��  �\��@x��j��0�&՚;�I��4v ˣh���#�d��~7O
�v    &[+i��w�;   ���;�8z��'y~v��D�K.��7l��� `y�?����ȑA�    X-a~�#Gw�>/v  �r0pűc�.vL��\N�wܱ&v � ��ݷ/o?�x�<��   �U5և���;  `9����gg?�������v��3���*�� �Ԅ,+ڏ>���>O�m;    �)���<�6v  ��2pq������ ��t�Y��7�cw pj�C����7��b�    @T��iG^���   ���`���cǝI�ui��D3��TJcw p�B�o�������,s�    �$I�(����Z  `����F�oC��̪�6U���Wcw prB��/})�}�{�$ض   ����uG�����   8� #굏}lsXZ�6vL�Z-��~��� ���ѣ��s�k^ye�    F���'c'   �
w�5���O������>��]�`^~��y�Vh���-    0�B�y�/�o��  �dw�����������&M���˵k���� �Ą� �O=�u����0v    ��Z��W�   N��;�*�����P��%M��}hM���`������o��~�    ai��C�����   8� #�q���&��w��IS���Z���+�; 8~�����=�p+;�l;    ��4I�R����   '��`�,���g���&J���o�u&v �-�~�����Y���1    0����[^۾���   '��`�|{nnMyaa[��4��n�IO;�s�8(������>�l��v    8Y!�r���  �Dz����CI��6vL���sʵk���� ���,+�_�b���˽�-    0	���]߹�w��   8� #�XX��� �f�w�$�R���7<zt�=�psx��0v    L��`�%!|:v  ��0p���~<�����IR��jy��j� ���嗻�Gi�,�[    `��{�؇   c�/0 #�����`�T*i����� �m���?�����	C��   `%��ιo��_�  ��e�0^���)i4.����~�-��gx�U�n�y��o_7v
    L����b7   /�/�Pi��&M�4vL�ҙg�j[��cw ������_h�n   �i�6W�2;{S�  ��a��/?����������~�k�R�K# #h��+���?�*���-    0-Bi��z(v  ��0p���l~6���0)*�\R�\rI5v �?����җ����1    0m����~�я�'v  �;1p�腻�^���$vL�R)���kbg ��Ð����'��    bH��:�j}&v  �;1p���4}(�����IQ��z��˱; �5y^�{,������)    0���an��  ���DTZZ�/vL�tf&�y���; ��B�1̾������A�     I�^�]���S�3   ގ�;@$���q_h�ϋ������$33�m FD��k����V��P�n    �������   ގ@,��'c'��(�[W�]}��������=�H���    ��B�y��ٻcw   �w���yUXZ�:vL��;�X��Ji� ������Od�``�    #*m6��   �V�"�6��1	��A��+�.���  	���t�~���v    e������m��  �1pXe�ssg&�����TJ����� S�(B��S�޾}��)    �;KC(�{��  �1pXey���d0�����z�u�Һu�� S��-ڏ=���~�    �������X�  �7���tq���0	ҙ�t����� �f��f_�Bkx�� v    p���5G^���   ���`ڶ���>/vL���7�$33�e ")^{m�}��b~���    ��tqq.����-  �H�K
�**�Z��� ��t晥��͵� �j��_��G�B�b�     ���y���}�c�3   ~��;�*9�s�Uai���0	��>��Ji��i�{��n�'�d00n   �	�O�n   �u� ���j�M�A.���{�S�\vY5v�4���y��;IQ�N    �IXZ����][bw   �w�U���w�Mo����v�mk�$���
���t�}6�    ,�4IҢ�|(v  ��0pX�T�"�����qW��j��+�; �J!��N�����N    VF�������   Hw�ձ����	0�J������� �*E�j�_|�;    XA����7����   Ib���^���&Y���0�j�^[+�}v9v��C��_��?�i?v
    ��J����   Ib���*ͦKp��մv�ͮ������c�e�_�r�    X%���C�����   � +���ܺ��xS�w��n��k�xnX!ϋΣ�����   ��I��S�   � VP��x(k�;`����^�n�Z��0�V�h���oc�     ����xs���ύ�  L7w�����=v���[o���J�`�������*��-    @a8���2v  0��V��;fC�}A�g���.U��ҷ  ��b~~�~��,4��    0����{c7   ���`��f�`���v�L����������/~�Z-�v     	��y�����  �^� +���܅aqqK�g�.(�7l��� �d�Ç�#�d!�C�    `t�f�S�  ��e��j���IB(��qV��f�$q�`��w{������    ���..n=87wa�  `:�,��gO�XZ�;v�����W)�_�z;�
<��<�x���)    �
EQ�6���  L'w�evd߾?y�.v����n��� 0���   ��1�����+  V�_D �Y�����0�*�]V-]pA%v�$2n    �W��ux߾�bw   ���`-�ڵ�XZ�*v��4M���z;�
0n    NT�����  ��1pXF�,�i>[�$U���V:�r��Ic�    ����t��;.��  L#L�e��j���]�;`\��rR���z��Ic�    ��J�<���  �t1pX&��Z�Hz��cw���l�\O�8��v�ed�    ��tq�#����;  ��a��LB����`lU*i���\oXF��    �r��G���  ��0pX��ڵ�h46��qU۲���Y�`��    ˩h4��   LC2�e�o6J�$��c�ZMk7��z;�2<�o��?���   �e�h\~t��kcg   ����}{nnM��p{�W��[k�̌g�e�/��d0�[    �ɑ&I�f�_��   ��1�)��v���`�&v��Z-�o��z;�20n    V�pa�07W��  L>w�ST,-}4v���֭���v�SV=:h����    ����׾�e;  �|e ���ݻ7���e�;`��zZߺՕ�ST;6l?�x�����    ���Zs�  ��g�p
���CIi�G�믯'��g�SP��ۏ<�
yn�    ����t��]bw   �ͨ�$�={J����;`��zZ��:��NAh4���ˌ�   �UB��e�g�  `��������a��g��qT��&��NA�j٣�f��*b�     ӥXZ�;����<  ����I�f��n�q��̤�͛�; �U����c��h�    �.���׾���;  ��e�p��]�,.^��Q���i���� K�n�y�Ѭ��7n    �ɲ?��   L.w���.-�e��ƍ�� �`8�/�=|��a�    `��o����;  ��d�pʍ�ݱ`ծ���v��Q!��lx�� v
    @Z�����   &��;�	:2;{wh�Ϗ�c�VKk�7�bg ���?�t���_�    #c��4�  �L� '�Ȳb7�8�m�ZO�u� '���o�����    �ץYv���[bw   ����|{nnMiq���0v�մ�e��� '���ۿ��    �j�?;  �<� '��,�D2���㦶eK-����p/���>�\�    ୔��n>X��  LC3��l �&-��ږ-�� �dx�@��u�b�     ��^��#��;  �,� ��ȶm�Fcc�7�뮫�����8��>h?�d;)��)     ��n��n   &���q*��!�܄���I���]o8N���<K�}��   ��P,,\wt���bw   ��P�8���ߋ� �z�t�Z� �!�y��җ��n�    �#�r��|*v  09� �á{��ph�Ϗ��$-�������� �aȿ��XX(b�     ������  �� ǡ��>��M��+k�3���NB��Of�#G��S     NJ�u�+��7��   &���;ss���ts�+i��n��;`�O?������     ���n"v  0����v����?-v����WKg�U��0�z�����^���     8U����ܜ�  �����FcW�7��w����^�����     ˢ�{��Ngw�  `��������[n6����r�ŕ���Wbw ���7�|���;    `�d�}�  ��g��6���?Ea�'�v�������,ڏ?�%��u;    0Q����s�=��  �7w���j�~�'�w��\^��K! o!��!���B��    'k����   ƛ�;�[8�m�šټ4v����7ד$Icw ����?�c6|��a�    ����Z��  ��f�����ϓ|N�q*�uV�|��� �*��7:�_�r�    `E--m:87wa�  `|n���ټ+v���M7Փ4u�����G���/�bw     ��B����g�;  ��e��[��kזR����0.ҵk��W�bw ��������vbw     ��V���	  ��2p�-Y���K�p�j�__O�e?3 ��XXv�|��E�    �U�f���;w^�  O� �Eh4~7v��Z-�^}u=v���v�Η���n7�N    XM!��Ȳ?��  �'w��ptǎ��N��0.j�^[K�u��~]�󕯴����   ���l�;  O� �a���Q��RR��Z��Q���7;��;     ��t�9�c�]�3  ��c��k��\9YZ�5v����W�3�(�� %��^��~��^�    ��  N��;��9���N{��cw���m�Z�� 0J��G�7�щ�    0
�KK���9ǒ  �b���Z���N�qQ~��*��ϯ�� ��.�O>��a�    ����z�����  �x1p��o�ͭ	����0.j�_�z;��(��?�DZ�"v
    �()e�#c  �	1p��K��O��`&v����g�*��;���J��ot���t;    �o(--���j�;  ��a��+����xp������4v�(��b��⋽�     #��_s�w  ��$I�ؽ��R�yu���LZ޴ɕ�$I��G�g����     e�NgW�  `|�$I��v?��J��뮫��������v�~�,��S     F�pqqkx����;  ��`��$Ih4�� � -����ͮ�E���?�C���)     �.kG���(v  0܁�wdv�������AeӦZz�i����}�|x�� v    ��(�Z;b7   ��@�z!���$��p\oH��/~�������     �$4���[�  }���K��ñ`����J��*�; b
KK��W��NB��    0V�pXI�?��  �>w`�ڶmch����Am��ہ���y�v��Y�    ��J��~�  `���m0x M�4v�����K���; b�~���ocw     ��F�ʅ]�Ί�  �6w`��Z�;c7�8�m�\KJ%/� S������܋�    0��pX����cw   ����Z��vm���bw��K��z�5�� �����3�tbw     L�f��	  �h3p�V���D�$.R�;�l�TK׬�� L�0�ΓOfa8��    0�ͫv�:+v  0��Հ��l�;�Am�f�ہ��}��v1?_��     �a8�tz�?��  �.w`*��}����Z�F]��ﭔ�;�� ��K/u����cw     L�4���   �.w`*z�O�I���QW۲��v`*����3��;     &R�q�®]g��   F��;0�J����`ԥ��^�l�P����B�:O<�%�A��    0��pX�v�s�;  ��d�L�׶o�4�Z��QW��ZR*��`�t��N��P��     �h����	  �h2p�N1>��`�o�TJ�W]U����?�I���˽�     �n��t�w��]�;  ��c�L�f��	0�*�^Z-�q��`��Fc����;�;     �AZ����\�  `��S���܅�պ$v����ͮ��%��?�T;��B�    �i�f��n   F��;0Uj���I>��m��:�T^���`5u�>92��    0U�k�ܜ�K  ��a�	L�a�uW�u�͛�I���; V��ȑAo��n�    ��3�β]�3  ��b�L����3�V���0��r9�^ye5v����󕯴���]    0������  �h1p�F�e����FYeӦZ:3�� ���uB�e�    IXZ�!����S  ���05J��ݱ`�ծ���`�^z�7�����     �j���o���o�  ��2p�B��g����ձ;`���=�\���r L��h;��f�    �$t��c7   ����
���gK��z�e�-[\o�C!�v���)     $I�l�?v  0:܁���l�� #�VK�7�S����wG�cw     �+y~�k;w~ v  0܁����I��%v��ڦMմZMcw ���o{��n�    �k�e��n   F��;0������kcw�(�^}�����+��}�v:�    0rZ-� �$I܁)P��{c7�(+�{n�t�y�� +-�ַ��oZ�    ��v��;w^;  ����xi�uc�e�͛]o&^q�P���ucw     ��jy~_�   >w`���kז���FUZ.'����; VR��C{��NB�     �F�e��  ����hE����0�*W\QK�u��D�>�l'4E�     �^�ټ��{�f  0�ڀ�Z��n�QV���Z���T:���R/v     �,�Pnt�s�;  ��܁��ˏ~�=!�.����t晥�{�[���RB��{�v�b�     p�J��]�  ��܁�Ui��OB�9o��ys-I�4v�J�~�[��h�;     8�Ƶanη �3�&V�ݾ3v��R)�n��?��5<x����{�;     8A����<�;  ����Hߞ�[S4��bw���\zi5=�4��D
�n����IB��    �I�d��;  L�J� ��pI��N�Cש�-Ԯ���0���=�	�f�    ���e7�N   �q��Hi����`T�kצ�.�0��G��/�ԋ�    �)�t�9�}��;  L)w`"�����`TU�����i�`��!߻����    �ST��?�  ����8������{W�U�M�j� VB�;�ɋ��"v     �.d�-�  �8܁����;FU��ʥu�ʱ; �[q�ذ��vcw     �<�V뒣�w��  X}���)e��Dŉ    IDAT�`TU����v`��{�a8�]    �2IC(%y�3v  ��܁�Ҹ��s�,�(v���\Nj�_^����z?�Aw��k��     &��]�  ��g�L��јKC���EeÆj23���(aii�{��<v     �/4׆={�}  ��_�����n�QU���Z�����0t�    `"��k��w��   V��;01��\9i4����(=�r�E�� �i�ӟ�bw     �rJ����  ��2p&ƫy~W�﯍���z啵�TJcw ,�n�ȿ��N�     VX�}S�  `u��#Ϸ�N�QU���Z����[yh�C�     VX�����܅�3  ��c�L��jys~���K�S���\���:���ǽ�     ���j�},v  �z܁�pdv��$���FQ媫\o&GQ��׾�I���     �"d��  ��c�L��߿/M�4v��4M�7Vcg ,�����p��0v     �'4�W��9�X  S���i�s{�E���+�ڵ��&Bh6��}���;     Xe���W����  ��0x�^س��6��bw�(�n��z;01�g�ɓ� ��      �N�b'   ���{�|��J��bw��I��|饵� �ax�`��cw     G����  X��ثv���n�QTٰ����i��SV!���;�3     �'�Z���}^�  `��c/Ͳc7�(�^qE5v�r����-��     DB��v  �<w`�5v�>'ɲ��;`��ji��܁�W�ZE�{����      �R�sg�  `��c-�v�!�cw���n�XM��4v���>�L'��C�     �Yvm�  `��cm���� ��v���co��+��?�s?v     �!���Gfg���  �,w`��ͦ7��7���^*]xa%v�))��?�L'v     �%��gc7   +��[Gw�6�vϊ���z��$M�� �����b~���    �h	Yvk�  `e�c+����0��7Vc7 ����E���cw     0zB��ᅻ�^�  X9����tn�� ��t晥�y�cw ��������;     =iQT�]��A�  `��c)<�`54����QS��j�$i���U;6��R/v     �+�v?�  X9��Xz�С����FM���k� NE��g;IQ��     `�����  ��1p�Ұ����0jJg�Y*�{n9v���������     ����~��ݻϋ�  �w`<����N�QS��j���V!��7��     ��J���;  X���	<�6�Z��QSݸ���d�^x�[,-�;     �۽#v  �2܁�s�ر{�ʱ;`���>�T:�?�x�v�޾}��     ���j]�  X��ةt�w�n�QSq�c�}��!�C�     �G��{h۶��;  ��g����e�c7���n�X�� p2B�9�����     ��R�b7   ���+Gw�>/�t.�����n]��n]9v���>�\���     ��<�@�  `���%�w&!��3`�T6n��n 8�k�����cw     0��ͫb'   ���+�n���`�T/����d��>�'!��     `\�z�ؾ���  ��2p�J9˼���t�٥Һu�� 'j�����bw     0�j����  ��2p�Ƒm�.N�|]�%�ہqBȿ��<v      �o��   ,/w`l�!̆��0J��^j����O~�ǎcw     0�B�yyس��  &�|`l�y~K�%�g�J�_��pB�"���N7v     b08����  ,w`lYvU�%��.�&I�[���{�^h4��     L�r����  ��1p���]�<_�FI��K+� ND�vCo߾<v     &�o��   ,w`,4�|{�%��LZ��Bw`��~��n���    �����Þ=60  0!<�c�����FIeÆj��i����������     L�������?v  �<܁�eW�N�QRٰ���Dt���&����     ��r����  ��0pF��]�<_�FF��V.��;�x�V1����v     VN��;  X���k����0J��^ZI��4v�����ycg   ���ޝ5�u�w^�n���Z�,K�d y����WQU��>� �9�;�ӥ����Y6�<)��{�5=�I������꽮���~Z�� Xb�ѣϥ�7�`  `	���r>�Vt���gW� �V��qW��Ut     K�i�����  읁;0|�۟�N��(�l��3����U�����     ,D1����  `�܁A{��߿��f'�;`(&�/O��U�7p t�u��/��    �B����  ����6�N��Rʣ;`(���W� �V����    ��<y�\t  �w����U�������'� O#}�a[ߺ�z;     �W��{7n|1�  �w`؞<�RtEq�D�?^Fw <��/̳���     `d�����  `o܁�z��m�����ɳϮD7 <���a[����     ,\1��et  �7��`�m�|���S��&ׯ����?v�    �����  ��1��N�.��"?|8//\(�; >M��q�ܺ�z;     !���ԝ��K�  ������ӯF7�PL�_�dy�Gw |��'?�����     `�RJ��ɓ�;  ��3p)�������������+� �&mow�/~�z;     ����o�  ��3p��W_��Զ�����&W��� ^��s��    �����  `�܁A����`(&�.M��Uo60hi:�^r�    �x��>��:�  쎱0H�|����������OS����iRt     �)�����;  ��1p)=yr-��br��$��OI�y�]o    `@�l���  ����������Y]�Ew��Eq�D��Կ��<�箷    0i>�rt  �;���4��?D7�P�\��z;0l]������v     %��t�]  @~���Ͽ� CQ>��Jt���ܺU�Ǐ��     ���9�����  `�܁�)��?� �PYy���p���/�8��     ��s���1�  �9w`P|�{�i:=�CP^�8�WW���OҾ�Z�=x�z;     ���f߈n   v���Y]�s���M�e���5�ہA���'��    0Xɷ� ��dD
J���&���|晕��Oҽ�V�޻�Fw     �'�NO߻q�7� �c�J�Ͽ� C��������i`��/��z;     ��gY^����  ��0���"��jt��ڵ�,������}�A�ܾ�Dw     �����_G7   ;c�Ɲ_�f�4G�;`&�<3�n �$�O:�R��     �O��S�"  ��;0������<��+W܁AJ�Y�ܺUEw     ��ȟ<��n޴� ��/��`t��ף`&�ϗ����h`���^�R�Fg     ��i��;/����  �����oo6����v`��.�/�4��     ��(�ڷ� �b��ϟ~��N�Fw��W��D7 |��W���I��     ��(��?�n   ���;0&��O)��-/ˬ<ޟ`���?����     ���f��  ��g�B]�� CP^�<��2�� �C�;Mz��6�     v���>���_��   ���;0E]9����zu� �q��t�      ��R*/=��;  ��c�B���Lt���w`p�Çm��Mt     �V5��Vq  8 ܁p�n�8�f��-?|8/N�.�; �P��KU�Rt     �Z;�}5�  x:�@�j>��<����6�zu��?���m���*:     ���N�G7   O��7����n�!�\�:�n �C�+�Ti6s�    �-��N޻q�lt  ��܁pyU}!����r����g?s�    �/��M��  ��3p�mo_�N�h��cE~�X�𿵿�mӾ�^�     �����*�  �t�@�����gRU�Gw@��ի���S�����     �7U���  ������ot���w`P��v׼�j�     �f:���  p �����ztAq�;0(��[Uj��     �7i6;����9�  ��܁X����c��͢X_�&C���^��#     `�u���G7   �1k:��3z��ˮ��Ҿ�f�>�;     `��M�[� `�܁0�����YU�Gw@���;00��    ��|�8  ��;&ϲ��n�!(.^4p#=y�5��^Gw     @/��g�  �?�����߈n�h��cE���=���/���3     �EU}k�|t  ���0��~�lr����p���_����     ������өo �3p�t��W� Zy���;0���Mz���v     �Z7��Et  ��܁o}����Z��h�K������z;     cPV�o �3pB����n�h��F�ol���f��}��:�     ��M��D7   ����V�ף ��ʕIt���oݪS�Fg     @��lv������  ���!��~.��M.]r���嗫�     X�<��v{�o�;  ��g���g�����x�w`��������o    `4յo ��2p�߿��c�l�����������Pߺ�z;     �R���  ��gX,��VW����Gw@��ҥI�e� ��6կ�RGg     �"u�ٵ�  ���7�N�"���/�� Y�eͫ��i>O�     �Hi:=���|f  d�,\�4��n�h�ŋ���,˲�嗫�     X���V��f_��   ���;�pi:�� ����3g\� ¥��s���     �y��ut  ��܁�J7oi:=���s�&YY�� ��~Ue]�     !���+�  �3p���ϯ�m{(�"�/��B���ut     D���g�  �?f�,T���o�^y��$��{���}�6�     ����rt  ��܁���W�1z�.���[���     ��W�����K�  �G��5���7F���,�#G��@�T���ut     D�L��   |���P�|~1�"��.M� �;w���Q�     ����	  �G����_��|~"�"M.\(� �W^q�     �,����E7   e�,̛|+K)��H���.���.տ���;     dY���W�  ��2pf��� �&��8y���j�x�Ϊ*Ew     � L���͛>� ��:�8��� Ry�|��o1 Bտ����     �?�v�������  ����SUע Ry�|� �[��T��Z�     CR��_F7   �g�,L>�]�n�Hw X���u�4)�     �$��_�n   ~��X�{7n���z=�"�g�N��q���:�     �&o��D7   �g�,F]�uJ)�΀(�ѣy�������]{���;     ��4�^�n   ~��X��i�� ����]oB5��V����     ��)��3ik���   ~��X�|>�ltD*Ν�b@��׿v�     >Fj�ɻu���  �w܁Ũ���	irႁ;&�穽s���     �������  ����f�s�&ϳ��w L���uj��     �n>�Bt  �;�@��ݸq6����R?^d�{s�0�o~SG7     ���Ms-�  �c;�w�i|��V^��z;&5Mjn�n�;     `��|~)�  �w�u����T�=;�n ƫ}�:k��     �6��N7o��  � ���]^ן�n�H�ٳ.�a�����n     �������/��m   w�w]U=� a�<+O���1�.կ��Dg     �Ap�,�<�  0p �f� Jq�X���zo����MVU)�     �����   �=����#yU��(���et0^ͫ���     pP�U���  ����3��7����a��3g܁(�y�w     xJ�|~9�  0pzV��E7@���Yw D{�^��<I�     p`�fg�   w�g��>� ��ӧ܁�믻�     ;Q�k�om���  ��3pzU������ol��#�Z D��Mt     4���7�  `��^u�����R�=�z;"=|ئ��o�;     �Y�/F7  ������OD'@���R�����     �u}=:  �������|�3YۮFw@܁(�k���     p U���  ;w�7�����T�>m�,�|�5o��;     �BQU�  `�܁ެ4�� J~�p^��{g��k��i����     ����N��7}�  ��B�&U�g� Jy���@��7\o    �]ʻn�ß��zt  ���;П��� Q�ӧ܁��}��     �`����   cf�����E'@�����X`�w�m���]t     dE�>�   cf|�"mm��|~"���N��,\�曮�    �^����  3w��7�s��&�"ϳ��Iw`��^3p    �=Ju})�  ����E�4_�n�(���E���Gw #3�w�{�     �G�|~>�  ����E[U_�n�(��Ӯ��ܹ�d]�     ^1��H[[>� � �@/��y&���N��.`�7�p�     �AJ�|��>�  ce����k_��hMΜ�׼���;     쓕��bt  ��Џ�:� Qr܁�<hӣG]t     ,�<��F7  �X���f������eV?�}�y�-��    `uu}5�  �� �w�����y������e��yt0.����     ��ʺ��   ce��Y�})���O���Ȥ�Z�    `_�Uu6�  ����w�R�ltD)N���ݿߦ�<Ew     �2ɫ�dt  ����&Ms-��'O��,Ts���     ��������tt  ���;�ﺺ�� Q\p�y�Mw     ���G���   cd��4���n�yYf����V`aRӤ��]w     �A޶��n  �12��]WU���q��,�<ϣ3�����mR�Fg     �Rj����  #w`_����ײ�Z���S����B5o�m�     =Im{)�  ���W'VW��g�֌R~�D� �K��[Mt     ,����G7  ���jҶ��n�(���"�m���3p    ���Uu*�  ���_m{-:���,Rw�n��6:     �V^U��͛�5  �`~	�W�^�N�y����U`a�߶n    �����}�+�  06�x��Ju}>�"�E>����x�o��D7     ��+��G'  ����*����ar�7X��K�ݻ�     г�m?�   cc�쫼�ND7@����2���޽6�mt     ,�I�^�n  ��1p�M��:��z-�"����T`aZ��    `!����   cc���M�\���+�Ra�,P����     � y]��n  ��1��MWU�E7@�����`4Rs�n     �PU��  `l܁��ҵ����eV�����8tti6K�     0i>ߌn  ��1p�ͤi�D7@���2�sw`!�{���     ��]}�����  �11p�M[�� B���=���o��     ����s�  0&y���k��:�T�����.�    �"uݳ�	  0&y�����DtDp�p��    IDAT�X�٬�<�3     `Lڪ��   cb�쟪ڈN�����S`!����,��     ��m�G7  ��������=����2�����6�     Ʀk�s�  0&��������n�yYf��z��Cw�~�      cS����  w`_�������Yfyn�,Bj��s�     ����  0&������jtD(77���B���4���     ���֣  `L��}�������;�-����v     �ж�o�8�  ca��Զg� Ba�,H{;     �����n  ��0��E�4�ouF�8~�[
,��;     �Y��k�  0Fy�����	�w`!�.��c�     AR�\�n  ��0��G]�N������]��A�5M��     ��j��bt  ��Q�g�?\Mu}$�-_]����<�X~�;�4�     0fE۞�n  ��0p���o\ϳ�ȗ�)67���B4��E7     ����=�   ca���jY^�n�����Q`!�����     ���7�  `,�=���RtD�76���"���w�     P�4��  0�y����3pg�r܁H~�eu��;     `Ԫj-ݼ��A  X �x{׶g� B�;� ��    @��Ry����Ew  ��{V4ͩ��P;�zg�     �0��k�  0�y����=� r܁��y��     ���D'  ��{���ft,Z~�p�������s�     ��Ȳ�  0����u�� �V��{C�ޥ�KO���      ˊ�9�   c`��I�y���z-����p��]z�}��    ` ڶ=�   c`����^:��TFw����P�w�t�     ��Ms2�  ��8ؓIU]�n�kk�P�w�{��     C�4��	  0�y���Yv)�"�yt������    �@��9�   c`��IS�� B���������#     ��V�k�	  0�y��L��TtD��ּ�@��G�RVU)�     �om{$mm��  ���iwF���[���mt     𿤔��e��  zf��I׶'�`�����<:Xn�     0@���  Xv�����9� �V�����<�     ��Jy~1�  ���;�'e�nD7��ǎy?�ޥ>p�     �PӜ�n  �eg��Ig������O�w���     ӥt.�  ����'y]�n�E+�ͣ�喦�.��)�     �Ms2:  ���;�k�_�u%k����p.�=�<p�     �(%w  虁�kw�޽���5�S�����Uz�n      �X�4ǣ  `���֥t)�B=��zպ�     ����Xt  ,;=`׊�.D7@���܁^�>p�     ��mף  `���Vtݩ��;г��\p    �JM��   ��@ص���D7��M&y���;П�KݣG�     0Du}$:  ���;�kyJ���h�ښq;Ы���.���    `�R*����>�  ���ص�m�G7���kk�N�W��C�v     ��y~>�  ����{)mD'����.��j?���     ,�L�D7  �23pv-o[wF'?z���U���2p    ��S2p ����4k�	�pG�x;�^u�     0lm{::  ����{mk���kk.��j?���     ,����  Xf�����X8܁~�d�     ��u�  �##=`������ɏu��Mz�$eM��;     �O��t,�  ���;�+���u$��Jt,Z��j���{���v     ��m� �G���<��}!�"G���I~h�     ׶�Ft  ,3w`W�8� ��Y�;У��#w     ��mף  `����tݩ�X�|u5�����Mz���     ��#�  ��܁]9����X����v�W�Ç�     0pE��n  �ef��Jj���h��;г�ѣ�      �i�mW�  `���R��Ft,����M�W�w     ���  ze��N��N�E�]p�4�uY]��     ��n�o[[G�;  `Y����n=�-?|���M���q;     W��Tt  ,+w`W:wF�w�O�ѣ.�     x:+y~2�  ���;�+eJk��h��@��<1p    ����>�   ���ؕ�uG�`�\p��>~��     ��S����  XV���4��;㳺��z�\p    �#ϲc�  ����]��Ht,���@o����     p@�]�;  ���ؕ��V�`ъU���I���     ��Y��   ���ؕ�m-}�|e�w�7����     pP���;  ���ؕ�iE7��:d����R�N]p    ��H�ht  ,+w`��͛E��Jt,�d�gEa�����NY�o    ���5p ���;���h=K�ЗQ���<П'O��     �饮;�   ���ر���ft,Z~�Pt�ĺ�m��    � )��pt  ,+w`Ǌ��Xt,Z�;Ч��w     8@R׭F7  ��2pv�m����p����S�    � i[� �'����4�Ft,Z��j��&mo�    ��R:�   ���ر*ˎE7�¹��(�f�     p�t�jt  ,+w`��,[�n�Es��S���     ��Wt�Jt  ,+w`ǚ�ۈn�E�]pz��S�    � Im{(�  ���;�cyJ���p.�=��    �`i[� �'���)�n�E+&��`���mw     8HR*�֖+�  �w`�����L\pz��&eMc�     ���ٌn  �ed��X�����1pz�f3�v     8��f-:  ���;�c]��F7���++�	�����    � �ő�  XF���Y�;㳲�;Ћd�     R�u.� @܁�k[w�g21pza�     S[��  �w`�R2pgt����`Y�    ���V��  `�;�v��;��;Гn63p    ���2� ����Y�5��O&�	��JUe�     ��  �w`��3pg|VV\p�1��    �A�uG�  `�;�R2pg\�"ˊ���E2p    �)O�w  聁;�c�w�f21nzc�     S�e�  �w`��&��H��C�@���     ��m� ���������e� ,��6p    ��K�Ht  ,#w`Ǌ��}w�G���     �]H)�n  �ed��X2pgd�ȣ���U��     p ��$�  ���;�s)����L���#w     8��]�n  �ed�
�X�:?;��t��O]�    �4�s�� @���X�g#��et��RJ�m�+     �]hRr�  z`�
�XJ��ƥ�<Џ�4�	     �.)M�  `Y�;�n�,2wƦ,��`I�u�N      v��2w  聑*�3��+���,��e�4�     p@Y�D  聁;�#��;� 7����"5Mt     �[)��  =0pv�j���X��s	�#u]t     �K��� �{��4y~(�-/}� Џ�iRt     �K)�   z`���z׹����e� ,'�    ��*���  z`���R�zҶ.�    ��R�D7  �2��v��:Ag|܁����N      v)��;  ��bؑ"����ɣ�����        a��HӶ~n0:)�m܁^��     W�V  ��Pؑ�����oz��.:     ح�|�  =0pv���2����I޶)�     �5$ @܁����F'7p����    �J�  �CU`g|�cTx.�~t�     p`�>? �^X�;���       ૠ ����������3>�]
��     p`%� ����<�N'��p�@_�.�      �=$ @܁9<�og�����    ��r�  za��H�eet,��@_��;     Tɡ,  腁;�#����\=�o    ����  z`��Ȥ,�       R��9  ���          �A0p          `�          w           ��          �A0p          `�          w           ��    �����-�m�gF��!�iYm����+JUbo�8%R%��  [�rve�>(vs�y��=�J��     � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           ���=       �r�<��45�w�i�z\�0��   �M�      ; �0��n�ǻ����5�����Ƚ   ([�{       p=~l�7�u�ɽ    >��      vDa>N�aȽ    >��      vHa:I�4V՘{    |*�;      옶��')����so   �O!p     �tc�,�W�w    ���     ��z�Փ�y�{    |,�;      찣�y�0�U�    �1�      �㞵��a]or�    �E�      ;.�0�t�B�so   �?#p     �=C���˳XUc�-    �G�      �'��')����so   ��     �9���ҫ�;    �C�      �g�x��i�s�    �$p     �=��i.�Y,V�w    ��	�     `O=k�7w�z�{    ���      ���^���;    ���      ��b��ry�j̽    �      ��Ɠ�NCU͹�    ���      @uc�SJg�w    ���      @UUUu?��QӜ��   ���      ��I�\|�X�r�    `?	�     ���Y۾�[���;    �?w      ��<O�lY�}�    ��;      �O���=�U5��   ���      ����"��uUM��    ��      �Z�8��ҫ�;    �w      �Oݏq�]Ӽɽ   ��'p      ���M�z�X\��   �n�      凶=��U�    �.�;      �Ѧ�(�    IDAT���e]�    �&�;      ��B��ry���1�    v��      �$M�IJ/몚ro   `��     �O��q�1�W�w    �[�      �g�����y�{    �C�      |�GM���bq�{    �A�      |����^�W�w    p�	�     �/��m_-�˽   ��M�      |���"��&�m�-    �^��  �?7�s8�n��so  `���&�1�n��tܶ���u�M�m   ��  P��86�5�7����  �~9j�sq;�c��<���v�ӹ�B�=    �.�&  @�Ά���w���v   nړ�y��i.r��������y�{    ���  P�a��}��j����   ���qu�4�r���{�4�y^��n��   ��!p �����ߺ���kK   d� ���Rru�k�}۾�����8�ɽ   ��A�  ������  �\��x�SJ�s�`�<k��]�-6Ӕro   �|�B @f��q�o���v   r9����}�{��a~��i{    �� @&�<������t��XU1�   ��2��$��:�9�vWa:n۳����[    (��  2�NS��������[   �_mË�R�΍H1�S:U��    H�  7�rқ���0ϋ�[   �_M�������ܘ�1n�o�7�w    P.A  ܐi���fs�O��p   ��U5�H�e{��QӼ��y�e;    >DX  7`��6��?��9��  �~��j:I鴭�m�-�����v����N�-    �E�  _�TUa��t����   ��擔Nb�so�gm�z�x5M��[    (G�{   �~�����  (A������c�ro����:��8��6�!�    �!p �k6WU��������<�!�   ���z�ҫ�1�s�ߋ!L')��U5��   @�  p���T���w�Ðro  ����i^?��*�������)����    `�	� ��\Cz�^��NS̽   ��iӜ?j���w���c�,�W�w    ���  ��4��|��s����[   ��/�6�E��1�x�x�x�{    y-r  ��l��6��?��9��   ���b���m����⻶};�s|7�wso    �;  |����j�9�Ʊɽ   �у/����;�s�ضo��[\M���    �P�{   �6�8.^_]��  P�;u���m_���+�0�tֆ0��   ��� �G���Z����fsg��{   ��e]w�)����[�K����NcU���    p��  ���T���w�Ðro  �I!�/R:���숶���)����    `O� �_���f������{   |H��b�<�!L���u:��{�ҫ�;    �9w  ��<�����e�/so  �?�j<I�t{|c�z�4os�    �f,r  �m��f���<��[   ���U5�%��m]oso���i��ߎ��[    ���  �;SU��fsЍc�{   ��PUӋ�^���[�&<k��뚫i��   ��s  �Rt�x}uuO�  @�BU��)�����7%�0�tֆ��:    v�� ��7WU�������<�!�   �3���R:��&��i1��d�<�U5��   ��!p `�m��>_�ﮇ!��   ㇦y}?�u��K��$���    ��;  {�rқ���v�b�-   �1�������̽r;���1�W�w    p��  �i���z}��   ��z�4o�4�E�P�1^=i���w    p��  ��vۼ^��ӴȽ   >�7���i����9j�w�u�ɽ   ��#� `/LUV��A7�M�-   �)���Y۾ɽJt>w���+}    ;D� ����qq�u��<��[   �S܋�꧔^��%�ǃ��ǹw    p��  쬹���}�\Cʽ   >�a]o����;�D��q�k�=ɽ   ��'p `'m������4��[   �S-�;I�4�0�������]�d�*��   � �;  ;�r�e�/s�   �ϑB�_�tZ���lƱ���NUU��   ��!p `g��T��&߹   �JMۓ��4�0����i�s���   v�� ����n�U����ij   n�XU㋔^6!���@i�i�?w��XU1�    �.�;  ��TUa��t����   �����EJ/ۺ�������뎆y��&   ��@  �Z�8..����v   n�PU�qJ����[�4�<�?o6G�<;n    �'�  �:sUU��~���{   |�PU�O)�݉�˽J3�s���l�ͽ   ��#p �V�NS}�u��i���   ���1�W�c\����{ܾ��e�-    �,�;  ���0�˾��&   ;ᇦy� ƫ�;�D������t�{    7O� @��i�W]w�O��W   v�QӜ?j���w@����]���;    �C  @�6�m����y�C�-   p/�4�E�P�����o��^�    �#p �HSU��fsЍc�{   \�ob\}׶os�������w    ��� ��t㸸�CW�  �%b�|�қ�;�Do����0<̽   ���  c���}�/�Ðro  ��t���?��*�(��q<�m�ͽ   �2� (�0�q���i���   �u:�����r���q��]�8�    �!p  ��aH�}�̽   �۲�������[�4������Uro   �w  ���^u�A?M�K  �9m�IJg1�)�(�zۿ��   � !  Yl��f���<�  ���j|���Ec�-P�~��t�ө���[    (�� �5UUXm6�86��   ��PW����^6u-n�0LS���滱�b�-    �I� ����qq�u���  ��ꪚ^��2�8�����s��뎶�v    ��� ��n���}�/�Ðro  ��%T�|���A�}�-P�q��_��i?�^�   �O	� ���q���?�N��\   �PU�O)�݉�˽J3�s���n��ͽ   ��	� �j.�!]��2�   �ڞ���~���;�4�<��vݓ�4y�   ��"p �ڍ�T_t��0M�7  �y�5͛�1^��%���_N�A�    ��#  ��f�mV}0�sȽ   ���Ms��iV�w@�~�oW�x�{    ��� �k1UUXm6�86��   �M�v�x��i.r����߼ǻ�w    p�� �b�8�/{�����m�$�����HJ��������'�h�$�*��?�d�I�;�$�I�s�!�-pq:�^m  স�-��Kw@��{��l��    �j2p �O�M�|���4��-   ��	���ߔ��Lӝ7�ͽ�    \]�  �)SJ�|�6�J�   �ײ�u��˓�P�w�t�izX�   ���� �?�b���8�Jw   �״��y�Gm���-P�Ӕ���ǥ;    ��� �di���aؚ��w$   7Jl�q?ƣθ~�CJ����   ���0	 �O��l��q��9��[   �kZ��Z���K�@m>�_�nngF    |�  ���iڳ�zkL�/�   _[h��|�:Z�m*���Li�¸   ���� �kLiq:�^m  �&�fޏ�pٶ��-P�q�/�awn��t    ׋�;  �����0���i��[   ����q�*��t�f�9�^j�P�   ���� �_�R
�㸵�g�   �Hm��g1o�0�n�ڤ����zo��=#    _��'  ���4ŋq\��   ����xr;�u���/��1�t    ח�;  M���l��y�}  ���m߿����P�9��`v�9/K�    p�0 �p�ͦ?ǭ�s[�   J���w��C��͜s�rv��K�    p�� �PsӴg��֘�_J  p�������?+�5z5��/�y�t    7��; �4��8�m��  @�<X,�����t���0<:Oi�t    7��; �s>���i�;i   h��^O�˷�;�F����iJ�Kw    p�� �SJ�|�6�J�   @nw���OJw@�~��o7���;    �y� n��i��*�   ����w1���Lӝ���^�    n&w �k,�ܝ��[�<��  ����vx�q׶�t���fs�izX�   ����	 ��Zo6��8n���-   P�e�N���Qh۹t��4����q�    n6w �kfn��l��S�K�   @MM��W�C�v���V?�q;    �� \#CJ��a��j;   �Zh���a߶�t��"���0��q�   @q�  ���8n��iY�   j�5��<ƣ�T�js���q;    1p �⦔��0l����-   P��i���BK�@m�y^��ݹi�+   Pw �+�b���8�Jw   @�ڦ�Oc<��P�j3�s8���4�t    �_�  WPʹ;[���y�=   �Ɠ�?��e��Mʹ;��)ggK    Tǡ ���l��q��9��[   �V��7���c���/��1�t    �+�  W��4��z�5���   ~�^߿{��Jw@m��ð���e�    �w� ��!���0l{�   ~����t���Jw@mr���aع��X�    ~��; @���qk=M^�  ���~��,��Kw@�����U�    �w �JM)��a�N9w�[   �v�B��{�oKw@�^���Kw    ��0p ���4ŋq\��   ��`���O��7�;�F�����fs�t    |*w �������z{��P�   ��U��c<��6�n��Nӽ�����    �G� Tb����㸕snK�   �U��q߸���i�s<M�Kw    �e� P��4��z�5�ԗn  ��bٶ���B�Υ[�6�6�[?M���    �g� 4��8�m��  ��M���VG��M�[�6�)m�8��Kw    ��e� P��8n��iY�   ���i���m�)��9Oi��0�   p�� |eSJ�l�S�]�   �Jڟ����-P��)��a77�?   p�� |E�/�qU�   ���i���BK�@m.SZ�0n   ��0p �
R���z�=�s(�   WM�4�i�ǷCX�n�ڌ�x1�s��[     ׂ�; ���l��a�.�   W������.Kw@m����0쥦�    ׆�; �27M{�^o�)��[   ����w��C��Mʹ;X������   p�8� ���gð�snK�   �U����w���t�&���ޘ��    �v� >��q�ZOӲt   \eB8�����P��s�rv����	   �k�� �3�R
gð�r�J�   �Uv/�Ob|[�j�sn_���y^�n   �/�� �3���x1�.  �/��ǧ1�)�5z5��.�y�t    |I�  Aʹ;[���y�[   ����w��I������,�[�;    �K3p ��֛M6ۥ;   �:Xu��<ƣ�ms����q|�>�;�;    �k0p ���i���1��t   \˶��c<���7������n�    �Z� ��!���0l���-   p�m��_�C�Υ[�6'�t�x���    ���� �����z���;   �M��c<��6�n�ڼ��[?M���    �� �SJ�l�S�]�   �.�����x��M���YJ[?N���    P��; �︘�x1���   p��M���x��X�j�!�իa�)�    �� �i���a���s(�   �I�4�i���!�[�6S���Nn��t    �b� �O֛M6ۥ;   �:z���.Kw@m�)�/�awn��t    �d� �iڳ�zkL�/�   �ѷ}��~Kw@m�y^Þq;    � 4M�4CJ��a��9��3   |�}��a�(����9�^j�P�    j`� �x�ͦ?���   p]=^,Nw���t�&���ޔ�;;    ��� 7^��7   |!��o����;�6?��wǜ��-    Pc.     ����œ��m��Mι}1;�y��[    �6�     �gw��.��\�)���e�~9ϫ�-    P#w     �Zu��,��ms��ͫq|t1�[�;    �V�     �g�v܏�3n��x=��R�U�    jf�     |˶��W��жs�����������    P;w     �/M���x�h�T�js<Mw�l6�Jw    �U`�     �%]�����p�u��-P���t�p���    ����     ��ڦ��c<�!L�[�6�)m���G�;    �*1p     ���i���BK�@m�SZ�0�Kw    �Uc�     �am��1�a]�js�R�~vsӴ�[    �1p     ��o����.Kw@m.SZ�4n   �?��     �C�������t�f��ŋa؝��   ���p     �d;}��qߟ���L9��Z��IMJ�    �Uf�     |�����^ߟ���lr���Ƹ    �2w     �?�o��w�;�6)���0�9��[    �:0p     ~ם>>��M��͜s{0��y^�n   ����     ����n��ryR�j3�ܾ���<��-    p��     �Ҫ��1�m�K�@m^���y�*�    ׍�;     ��m���:�v��W���<���    p�     �ҷ���ju�v.��y=�NS�]�    �+w     ���I�1�m�J�@m~��o7���;    �:3p     ��i��i���]�)��9��;'�ͽ�    p��     M�4�Y�G���-P�w�t�izX�    nw     ��ڦ���xt+��t��t����ǥ;    �0p    ���1��	a]�j�!����    �U�    ��m߿����P��)ŗð���-�    7��;     �P{}��a�(���Li�¸    �0p    �h������Y���8ϋð;�G   �"�    �� ��?-���rð��&�n   ����     n�{!\<��m��Mʹ;X�����[    �&3p    ��v�]>��t��q��s_�    n:w     ���n�]�ǥ;�6s���0�s^�n    �    ��[u��,��ms��ɜs�rv��K�     ���     ��e�N�c<m;�n�ڼ���U�    ���    ��
M��c<\�m*��y5��S�.�    ���;     \C�i�?b<�θ���q|p����    �o�    �5�5��<ƣ�T�j��8����-�    �k�     p��M���x��X�js2MwN6�{�;    ���     ���i���o�0�n�ڼ�ln�4MKw     ���     ��'1���t��4����q�    �?3p    �k���{?���;�6�)�~�v    �"�    �����w����t��"���0��iK�     ���     ��ǋ��nߟ���\��|i�    W��;     \Q�B���r��t�f��ŋa؝݅   ���P     ��;!||��P�i���0쥦	�[    �?��     ���[�\���ڤ���a؛r^�n    �w     �BV]7<��m�\�j�˸}̹/�    �y�     pE��n܏�3n�_�9�/�ag=���-    �_c�     W��m��1���K�@M~�_��t    ���    @�BӤ��ѢmS�������b��Jw  �/K    IDAT   ���;     T�k�y?��e�nJ�@m^���Kw     ���;     T��yܾ
a*��y=�N7�ۥ;    ����     *�6M~��Vc����4�{���-�    |~�     P���xr;�u����4�9����;    �/��     *�m߿����P�w�ͭ���a�    ��1p    �������}��t��,����q�    ��2p    �J������?+��9Oi�jvJw     _��;     T��bq�����;�6S���nn��t    ���    @a�B�x�\�-���Li�¸    nw     (�v��xR�j3����0���    �Fq      �lw����Ҹ�ɔs8���4�t    �u�    @����xܵm.�5I9w��ޔ�t    ���    �W�l�i�:
m;�n���2ns�K�     e�    �WԷ�f?�C�v���s�rv�9/K�     ��    �W�&��x�w]*�5�9�/�a��<�J�     e�    �W�5��<ƣe�mJ�@m^�㣋y�*�    �g�     _X�4�Y�G[!��[�6?�ó�n��     �`�     _P�4�i�ǷBJ�@m^���)�)�    ���     ��'1���t��p���l��     �b�     _ȷ}��~Kw@mN����4�/�    ���     �������?��ڼ��[?M���    @��    �3{�X����Y���YJ[���Q�    �^�     ����o����P�)�^�Nn��t    P/w     �L�p��ߖ��|L)~o�    |w     ���n�d�|S�j�N�1��{)    �8H    ��h�u�����ͥ[�&c΋�a�3n    >բt      \e������7�yð��&�n    ��e     ���l��y�G�m��-P��sw0{S�[    �w     �BӤ�1-�6�n���<n�s�K�     W��;     �A]���1.�nS�j2�ܾ���<��-    ��d�     @��}�T�j�j��U�    ��2p    �O�6M~��Vc��ͫaxt��v�    �j3p    �O�6M~���֥[�6����iJ�Kw     W��;     |�o��7wC�,����q��v��[�    ��    �?���w���P��i��f��W�    �>�    �w������?+��y;M���A�    �z1p    ���bq�����;�6�)m���G�;    ����     ��{!|x�\�-��9Oi��0<.�    \O�     �O���i�oJw@m.R���nn��t    p=�    ����u��˓�P�˔�/��   �/��     ~���y�Gm���-P�q�/�awv�    |a!    �i�e�N�1u���+S����oRӄ�-    ��g�    ��׷�f�:m;�n��lr���Ƹ    �J�    ��BӤ���M�[�&)���0�9��[    ����    ��k��y�Gˮ۔n���9�ð���e�    �f1p    �Fj�&?��h+��t�dι}9;�y��[    ����    ��m��4�����-P�W���b��Jw     7��;     7ΓO�pY�j�j���]�    ���    �Q���7�C�X�j�z��t�t    p��    pc�����}��t��������n�     w     n�ǋ��Nߟ��ڜLӝ7�ͽ�     Mc�    ��`�8�f�|_�j�n�n�4MKw     ���    �k�^O�˷�;�6�Ӵ��4=.�    ��    pm��˧1���ڜ�����    ���;     ��V׭��x\�j�1���0��iK�     �3w     ��ض�����ͥ[�&�)-_�    3p    �ZY��Z���K�@M�y^�����    P1�     \�i���m�J�@M�yð��&�n    �=�     \]�����p�u��-P��sw0{S΋�-     ���;     W^�4�~��1��t��q��s_�    �S�    p��M���x��X�j2�ܾ���</K�     |*w     ���i���o�0�n���9�/�a�r�c�    �?��    �+�۾s7���P�W���b��Jw     �Q�     \I����}Q�j�j���]�    ��0p    ����������t���8>8M�v�    �?��    �+��bq�����;�6?��������     ��;     Wƽ>|�\�+��9��;'�ͽ�     ��;     W>>��M��ͻi���4=,�    �9�    P��[�\���ڜ����4=.�    ��    P�U��c<j�6�n��|Hi��0�    ׊�;     Պm;��x��ï\�_�nn��t    ��d�    @�����VG�m��-P�˔���    �ue�    @uBӤ�m�J�@M�y^����    pM9�    �*]���1.�nS�j2�s8���4�t    ��b�    @5~��B�J�@MR���0�M9/J�     |I�     T�m��4����-P�_��c�}�    �/��    �*<���N��P��s�bv��,�    �5�    Pܷ}��~Kw@M~�_��t    ��b�    @Q{}��a�(���~_��V�    ����    �bv���Nߟ��ڼ�G�)m��     ���    (�A�{}Z�j�z�n6�Kw     �`�    �Ww/��'1�-��9��{o7���;     J1p    ૺ�u�Oc<)��9��;��t�t    @I�     |5�]��.���P�w�ͭ���a�    ���    �*V]7<��k�\�jr��֏���t    @�    ��m;=��8��\�jr����0��     ���;     _Th����mS���ǔ��ð���-�    Pw     ���4�1�]g���:���q;    �o�    �EtM3?��(�0�n����8���=    �o88    �k�&?��h+��t�d�9�^j�P�    �F�     |Vm��1�
a(�5I9w��ޔ�t    @��    ����xr7���P�_��c�}�    ���    ��������c��Iι}9;뜗�[     jg�    �g��������P��s�bv>��t    �U`�    �_�h�8�����P�W���b��Jw     \�     �%�C8��r��t��axx�ҭ�     W��;     ڝ>�=Ʒ�;�6��������     �j�    �S��n��ryR�js8M��n6wKw     \E�     �a����xԶm.�59��;��t�t    �Ue�    ���q?ƣθ~��4��i���     ���    �d˶���x�v.�59Ki��4=*�    p��    �IBӤ��ѢmS��ɇ�V��a'7M[�    �3p    �?�fޏ�pٶ��-P�˔���    |6�     ����q�*��t�d�R0{��    ��Ɓ+     �V�4�Y��[!��[�&c��v    ��oQ:     �z�=Ɠ�!�Kw@M�yð��&�n    �n�*    ���m߿����P��s�rw��="    ��    �{}��a�(�5�sn�aw=���-     ו�;     �����w���t�dι}�?��X�    �:3p    �=�|��OKw@m^����*�    p��    �4M����I�oKw@m^ã�Kw     ��     4�C��4Ɠ�P�����4�ۥ;     n
w    �n����-����O~��o7���;     nw    �lն�����ͥ[�&��t�d��W�    �1p    ���m;�V���O�N���izP�    �&2p    �������x�v.�59Mi��4=*�    pS�    �0�i�~��}ץ�-P�)�~�ǥ;     n2w    ��k��y�Gˮ۔n��\�_�nn��t    �Mf�    pC�M���x��X�jr��Ҹ    ��     7@�4�i�ǷBJ�@M�y^���ٝ	    @�    � Ob<��e��ɔs8���4�t     ���    ��������c���&�p�^�M9/J�     ���    \c�}��a�(�5I9w/���1�t     �f�    pM=^,Nw���t�dι=��u���-     ���;    �5t?��o����;�&s���a�Y�s,�    ��f� �?v�"���[U3Y�$��h� ���3m@ԍ��Ƭ֡��g�VT�f�繱�4�?�Û�?_   .�k��\,�=z���������F�     ��    \ �9�����y�����էG�^�    ��'p    � �伺�X��Rꣷ��|�Z}�փ�;     �cw    �`����b�c���w���ߵ~4z     oG�    p���{�ʏ%�6z�����������     �=�;    �9V"����)�:z�ɓ�f��fs}�     ��;    �9�#ڿ�vsގ�s�t����f���     �yw    �s(E�����R6�����z�[q;    ��%p    8gRD��X��W�z����Z߬V7zD�    ��F�    p���~k��頔��[`NNkݽ/n    8��     ��W;;?T���0'�֦��Ս�    ���    ���bg��';;ǣw��lZ+�V�/jD�    ��O�    p|�������2z�I�=�[����>��    ��!p    ��O��苝���w�����׽��    ��#p    ��k�,������;`NZ���ju㬵��[     x��     3uX�ɭ����;`NZ���j��ik��[     x��     3t5糯ww��s�p��층��;     x?�     3s%�՝��ǔR����j��Q�WG�     ���    ��"������,n�7|�^�փ�;     x��     3����Ε+?����-0'������~4z     ��    `JD��X���R����fs�x��6z     ��    `���.?������f��h��>z     ��    `��o/?^)e3z���Z�~��|6z     ��    `��o-?헲��dY�oW+q;    �%$p    ��b���RNG�99�u�`���#��-     |xw    ������Z)'�w���ֺ{_�    p�	�    >�/vv�\��Y��s�nm��Z�h�]     \j�    >�Ϧ���;;���s�i��[���e�     ��    | �L�ї���7z�I�=�[����>��    �xw    ��Z)�������0'/��u�;��     0w    ��l?��[����;`Nz���j��Yk���     0w    ��h/�ۋ�O�w�����O[�2z     �"p    xO�伾�X��Sꣷ��|�^v����     ̏�    �=�Misg�����Fo�9y�^zT���;     �'�;    �;V"����)�:z�����'O�ۃ�;     �/�;    �;�#ڿ�vsގ�s��fs����G�w     0ow    �w$G�����R6����<�l�l>�    ���    �)��^,~�+e=z�ɓ�v��fs}�     ·i�     ���띝��)պ��zO�ED��"Z��Go��Z��[�?�    ��C�    �7�,eyѣ��_W���_�
�s��SD��z�����ܞ�}Q<��Q�W�V���    ��"p    ��Q���9o������Dk�A������׃�H�G�=��zD{�c]Ϝ�Ժx�Z}����     ��'p    ��n�|�iΫ���WyĿ�����u��{�=�_��g!���]:�u��ju�E��[     8�     ��9��(�l�׼q��s�u>���������󿾈�?�l.�ukӽ��q;     ��    �O�$�՗�����W��
�{yv��e����^xv������z��^�/����˽��QFo    ���    �	��������?zޥ�H�ڛ��_�/B��_^}���Z�D�B�=�;;�bӻ�     �-�    ��~J�[�t|	����"�Dk�zŞ�G������%�)��,~o��grμ��׽��    ��'p    x{)mo�����=�����o�^�g���>�������Ӄ����wGo    �b�    ��ED�3M�<z���?��Z����<x=�O9���Y ߃az���j��IkWFo    ���    ��݈vwg�<����RD����<~�GN���zzv齥�[�xq��?����z��qk{�w     p��    ��)��)�h��NJ)zDN�G�^"����Տ��R�)���[DK)�Q�/�oW��Ժ?z     ��    �7��~���ݜ��-�%)�^����)�E�-E��{����w��������_���w     p1	�    ~%G�;�-�����9Z�/����s��{J-Rj=�ų�����a����v{m�     ..�;    ��|]�r/�:z\����_��=��������%�o6�?m6��    ��&p    xͭR�9oG�`^RD�֦�5���%|���?�l���    ��'p    x�R�������2��Ժ��f���     \w    �������9�G��b����)�9�x��H����f�/k��p���G��[     ��    ���yΧ�����-������ߏ�.��T{J/���;_8�u�q;     ��    �Ԯ������;��^�����}�)����{��"|���׭M�W�-"��O    ��#p    .�k)��*�d��/R���KDD�="RD��[���뻌�7���9;��F�w�g    ���    ��aJ���t<z���_J��2z���=�\SD���\SJ������˽�ꋭ�    �A�    �������iZ��C�I)Z�^�qO���)��R��kv���?����V7ֽ�|��     ��    ������뜏��\)z/�����{D��R�)��/���ӽ���Yk�#    ��    �4v#��iZ����?RJ/��xv�G�oj=�    0w    �R�"ڝR���^��p�=X�.n    `��     �[��wK9�͹��s�#����/�v     fD�    \h9��)�h!n�7��v���/F�     ��	�   �+G�ۥ,�r�����<�u�߽_�     ~M�    \X�JY�����qk�ǭ��    �%�;    p!�*ey(n�7����G�^�     ��;    p�����k9oF�9y�������     �G�    \(7r>�4���0'�֦����     D�    \��|v����;`NNZ+߈�    8'�    ���IJ�/K9��䴵r����Fo    ��!p    ν�RZ5M'�w���Z��k=�    p��   �sm?�ͭi:V��+���Z��      �3�   �sk/���R��vxe��o�[�  �[�    IDAT    8���     ��ED�3MK/�R#ҽ��pQFo    ��·    ��ٍhwwv�JD��Gă��`%n    �s�    8W��v���I�/���A�'�{�    �\s�    87JD�[��n�m���k�_��3z     �]w    �\��N)Gq;��#�����/���     ��    ��ѿ.e��s����v������     ��   �ٻY��A���;`N~���Ͻ_�     �%�;    0k_�r�QΛ�;`N�������;     �]�    ��e)'�s^��s��G�^�     ��;    0K7r>�,���0'O[������;     �}�    �s=�ՍR�F�9Y�6=��`�     x��    ��\Ki��i:��䤵�    �K@�    ��AJ���t�F�9m�ܯ��E�W    �O�    ��~J��ӴT��+����Z��     \w    `�����vxӦ�t����-    �Kģ8    0�nD����c%��}�o��    p�x    ��"ڿJ9�r�\Ԉt���uD�     >4�;    0D��w�����ۃ��    �Kj=     �|JD�S��"�6z�E�=�zpһ�{     .-�   �*G��KY��\Go������e�;��     �Hw    ������~���;`.zD|��^�����[     `4�;    ���*ey n�7<�u�I��;     `�    ��RN�����Z���ڕ�;     `.�    �{w#��Os^��s��O���     s"p    ޫ�s>�Q���0'OZ�}T���;     `n�    �{s=���vx�/��|W���     0Gw    ླྀ����RNF�9Y�6}+n    ��J�    �s)mnN���0''��oj=hi�     �+�;    �N������^9m�<��P�     �O�    �3��z;�eN^xa�Z�_�A�    ��    ��nD�[�єs��b���zX��    �[�    �mSD�#n�7l#ҽ��p�-     ޚGu    �o)�n)G�9��[`.jD����#��-     p��   ��,G�;�-���R�������     �4�;    ��~���^�u���q�I���-     p	�   ���f)��9oG�9�v��_��3z     �W.�     ��R����G����է���     ��    ���e)'����j�{��b�     8��    �[����g9�F�9���+?�ve�     ��    �[���ٍR�F�9y������F�     ��B�    ���SZ�����;`N�����֫�w     �E"p    ~�G)��9M'i������|W���     p��   ��j?�ͭi:��+��&q;     �w    �7��=MKq;�r�Z��փ�_     x�    �XD��9/= �+g������    ���}
    x���r4��Go��X����zP��     �^	�   �����/q;�a������M     �;��    @DD��~���ݜ��-0ۈto�9�zO    �<    9��.�h!n��jD����#��-     pY�   ��U��j�u����l��g�v     ���    p��*ey��v����ۃ��wFo    ��F�    ��W�_�y3z�ɷ���R�     CL�     c|�����ףw�\���֫O{��     .+�;    \B��|�y)g�w��<�n�����     .�<z     �a]Oi�����c�W~����     p�	�   ������i:�����?��7z      p   �K�0���i:���Ik��[���;     �g�    p	짴�z��i���ek�w���     �"p   ��JD�:�cq;�r�Z��փ�;     �7	�   �ۍhwJ9*9��[`.N[+j=l��     ��;    \P��}��K����Z��     fI�    P��wK9�͹��s�n-��    ��	�   ����N)Gq;���H�k=�z    �Y�F     ޝ�o���˹��s�m-ݫ�pQFo     ~�K5    p��*e���v���Z;X��    �\p�    .�[�,���R�=�zpڻ�p     8'\p   ����\�y3z�E�����/{��     x{w    8�n�|�iΫ�;`.zD|_��_z��     �s�    p�}��ٍR�F�9yT�ޓ��w      ��    ΩOr^}Y���0'�j����+�w      ��    Ρ�RZU�I=f�qk���v     8��    p�짴�5M��vx�Ik��j�:z     ���   ��Ki{����^y���w���     �}��    ��YD�;Ӵt�^Y�6=��`�     ���-    ΁݈vwg�D��[`.NZ+߈�    �B�   ��M�N)G��^:m�ܯ��E��[     �wG�    3V"��R�vsn���\�Z��k=�    ��#p   ����N)Gq;���=߫��z�    ��     ���o���˹��s��H��ۃ��m     ��|    ��g)��9oG���fs��(��      ��    f查_�y3z�E�����J�     �4z     �ʗ��|��z����{<���w��     p	��    3�yΧ����G��Z�����     |w    ���9��(�l����o�W�}w�     ���   �`�RZU���0'��۽'�/F�      >,�;    t����4��s�C�W~����     ��'p   �A�S�|=M�4z����?��7z     0��    �Ki�u���vx�Ik��j�:z     0�4z     \6���4-KD���ik;�պ?z     0��    �M��4-'q;��lmzX���     �xw    �@JD�[��nJm������7�v     �9�;    | 9��)�h����;m�ܯ��E��[     �y�   �{�#��R�{9��[`.V������    ��	�   �=�U�r?���0��ҽZ�7j     �W|<    ���V)�Cq;��}�o�O     ��    xO�Q�ɵ�7�w�\Ԉt���uD�     �'�;    �7r>�4���0="l�+q;     �;��    ��,�����s�{�����M     �].�   �;�IJ�/K9��G��Z�����     ̟�    ޑk)��9M'�w�\��~���Kﻣ�      ��    ށ��67��x���G��=�}1z     p~�   �o�Ki{��e=f�Z���ڕ�;     ��e=     γED�3MK�$��ǭ-~jmo�     ����    ��݈v����Go��x���Z���     �Ow    ���v���)gq;<�Kk;�պ?z     p~	�   �O*�n)G�9��[`.��Mߊ�    ��I�    B��wJ9Z��ᥓ��7���4z     p�	�   �-��u)˽���-0������    �wA�    o�f)�9oGX����zP��     �;"p   ���U)����b���zX�3     �    ��,��z���;`.���fs���     �c>>    �︑��g9�F���fs��(��      ��    ���)�n�r6z�E�������     xO�    ������4���s�"n?�}�     ���    �+���9M�i���o���e�;�w      �K;    ���6����R���۫O{��     ��\p   ���R�ޞ���^yT�ޓ��w      ���    "b7���y��^���+?�ve�     ���   �Ko�h�*�hʹ��s�ŏ���     \.w    .5q;��'��>����     ��#p   ��*�v)�ݜ��-0O[������;     ��I�   ���#�ץ,�r����\,[���     �Hw    .�[�,�sގ�sq�Z��փ�Fo     ./�;    �έR���vx鬵r��Cq;     0��   �K�R�����b�Z�_�A�     3 p   �Ҹ�����ףw�\lZK�S���[1     0>Z    p)|���R�F�F�{�v     `f|�    �»���q;�T#����pQFo     x��   ��Z��J9��G�7�����     �!�;    �AJ�����s�#��v{p����-      �E�   �������4-��!0#�n��Kq;     0c��    �-"�����\���۫O{��     ����   �����r4��Go��x���=�}1z     ��   paL편��c�W~����      oC�   ��P"��R�vsn���\<im����F�      x[w    ν��r���KO[������;      ��;    �Z��KY��\Go��X�6=��`�     �?K�   ��v�������w�\��V��     ��   �s�f)ˏrތ�sq�ZyP�a�H��      �w    Υ�r�^Z����zP��     �9&p   �ܹ���9�FX����zX��     眏    �+��|v����;`.��~�[�     �0�     o��V_�r:z�Ŷ�t���uD�     �]p�   �sᣔ�����4z�D������     ��;    ������4����{<���wo�     ���;    ������4-���L�����/{��     �]�   0[��z;�G,x�G���^�����[      ��   ��)��-�hʹ��s�ֽ'�-F�      x_�    ����%n�7<�u��֮��     �>	�   ����r��s���qk���v     ��   09��.�h!n�������֫�w      |w ����	  <�u)˫9��;`.����]���w  ��wߧ  �?� �ܶ۝Tk= ��[�,rގ�s�lmzX���  �L�;Q�UGG   ��#p .��s�lv��  �Y����k9oF8i�|#n .�֦�nR�;��    �4�  �Z��Z飇  _�rr=���0�������M��*��v/r�"�H�s-   �� �4z�9m�S�  ���9�~��j���Uk�~��v �Rhm��6�i:�����    �G  �R�S�lvB$ 0�SZ}Q���0���Z�w[ �I�o6WS�W�w�   �� ���b���)�o#  sq-��W�t2z�Ŷ�t�փ�� ��RJ�[ۍ֦>Mg�5w   ��|, .�����n�� 0+�)mnN���05"ݫ�pQFo ,�k�   p�� \D)m����������]{��9sΥ)�,K�H%.
�E���rR�q#�%Ҭ�ʲ7P��j�p�-��iP�j��m�4Ha�H� TFI�D��%)R"E�佤$�"M���g��sESI�眵g�������9��g�γh͏�  &f?��;f�3�*p�Eĩ�O\4n ����}���B�Tz7   ��� �,��i��7�v ��ٍ(�����p���r>q�5�  �������   ��� `S���6��%  ��ED�y>q<���^��'J�?�ڼw �T���RQ����H��n   ���M����� 0i��z�8�83n��8�����^hmѻ `M���~���;   8znp �Y��gɭ�  �5F�w�㋋ap�"\�T)��Z3� �:)j�i��b6;���   �-� �zjmH��<�� 0YCD�y_�1n��<]����  XW)bL9���[   ���w `�Rf��ѭ�  �5D�����rJ���gj��n���   ���1������   �A��u�b�����; ��v�8���ܻ��ZO��׻ `��:�Zǘ��GJ~\   b�  pEJc�Z�q; ���8�gn0n��<_��[����  �PC�y?պ�;   8� �����r�G��< �~bϽ~V�;`*��:{���;  6Y��V�N�V�њ3p   Xs�� ���0�V��@ `-�y���a�ػ��\��i�v ��4F����y�   �ڹ	 ��Tʬ�:��!  \�7Å7���0�k/�zp�(  �'���1������   �f���I�Z͛ ��x�0\��q<߻��b��㥜0n ��y�:�lv>R*�s   �+7�  xI)cZ��a �6^�ҥ���9���U��Rn(�� L��r�O���   �����RD������]�  �c?�Ս��Y�v8�/�۳q; �d��h����6�#%��  `��  }�6�j����] �F�)���q;(�Rn�1�n ���Zg���ڼw   ���� t�J��ZG��  ����r�lv�/�@��S9��h� 0u�弌a��0\p�;   L��; �C��j�� �YD�w��/��^�z���kͳV �uQ�<j�lv!�Tz�    ��E[ ��j��i���q; �ڙEԛ��řq;D��?�'r�?�ڼw  WmL9�Z�C   ���V! �ؤRfQ�h �~ƈ��q|q1�wLA��o���BkQ  �+�Rv��1��B���5   L����R��V��; ��7D������vx�S�,��u�w  ���y�y���6   L��; p�Z�j5o��� `�q<��һ���Rv��u�w  �'E)��ڼw   l;C3 �ȤRf��E��-  \������aȽ;`*��u绵.{w  p$R�y�,[k�k  @'� �QH)�y���\ �������aջ��ZO��׻ �#V�<��Z�   :0p WkCZ��5g  �����7å�0/�:�V)��;  86c�y/�6�   �f�;  ���Y�ul�C  �.o��o���;`*��:{Ҹ `���2�a�p!R��   ���; pR�y��v ����a���q�л��\���RNԈԻ �Nj�GkC���H���  �Mg� \�ֆ�Z͍� ���S���q<׻��|��Rn0n  Z#���ڼw
   l:C4 ���Rf��{  ��)��>����Sq����RN�w  �S��L�����   G�� �)�<o���C  �~�)�n���Xg��UDz����  ��V�"��ͦ   p4|� �NkCZ��� l�eJ��pָ���juC�� ��6���[k��!   �i�  W��1r���' ���(7�fg�ah�[`
JDz|���R��U p%R�V{Q�n�   �$~M \�����v ��1����g���N�|�q;  W!�Q�"Zb�GJ�c  �u2R ~���¸ `s��������:n?ךA  �6��"��֚L  �u2T ^]kCZ���z�  p8��v�8��3�wLœ9�im޻ ��7�����-  �� ���1V�y3n �CD�i�,���n�)h���omѻ ����j��Zw{�   ����] ���<�ֆH��  ���xfr����JY>��N�  6KJ)��E�6�0���Z�&   X'np ^.�ju�� ��r�8�9a�/��Rv�u�&  G��Y��Z{�   �:1^ �6��j�m �0?1��^?��0�Ժ�G�.{w  ����^Ժ�   Jm��    IDAT��� �vp�̼� l�7��?;{w�T<W��R�zw  �UR���J�!   ��� @g9�Sk~� ���4�<�zw�T<_��[����  `;�Z���x.Rj�{   `��� `{�X�a� ��ސ�ŷ����0gj�� �]kc����S   `�� `�:��j�w
  ���)]z�lv�wL��Z�ӥ��� 0C��.z�   ����I�̢�Y3�  �H'RZ�}���P��x)7� 01)J�M���  ����  �O�y�Z�7 ��L)�cϤd��j/�D1n `���-�C��H���  �)0p��b�Z� l���r�lvf0n���X՚-��(  SW����  @D8����ڐV�y�� `c-"�;���1�m9"=f� �IC��Z�v   �� �`��1r�7�v ��5��7�㋳a0n��(���W�.E��[  �*��y/j]�  ���`C�Rf�V7�  l�1��s_\C��S�"�t���� XS)"���T�n�   ��� 6P�y�Z�C6 �6D������v���q���O�mm޻  �W;��}�a8)yc   [�� 6K��ja� �ن�v�8�YC��S�"�ۥ�1n `��:k9�g�   l_�`S�6��j��`
 ��z�8���ܻ��;9/��u�w  �1D���5og  `k��h����� l�����êwL�wJY�qk��;  ���y/j]�  ��`� k.�2K��� `�e���vx�3��<[�q;  /ED���J��/   � �X�y�Z�5 �-��a8��a�ػ��ZO��׻  �S;��}�a8)��=   p� `=�X���  ���p���x�wL��οU�~�  ��Y�y?�   ��|��5�Z�j5��o$ `��>�K?1��{w�T��u�D)'zw  @O)b����ػ   ��; ��ֆ!�Y3n �
�K���g������jO� ����y/�6�   ��� �E)c�<7n ��)�n4n����u<U��w"  x�TW�e�u�w   w X��Y�:�� ��X��o���X�����r�� �I)E+e'JY�n  ��`( S���Gi  [bQn�3� ��Z+��  xm��#"�a8�Rj�s   �Z9�	K9�ø `k�"��g�`� �#��9�Ȟc ���u�rދּ��AZ�^���>���  �i�4�X�nn �����r����Kc�  X3c��8���ع�~���  �i|���Ii��G��U  ���n�3�a��[`
ZD����E�v  �V�呻����O������7zw  �&1p�)imH�ռ� l�!��c�,���n�)h�ũ�O�omֻ  �\���Rk��!��Ƈ��'~�>׻  6��; LE)c�l� �en�3�Ð{w���x���38  pXR]���֝�!����]�����w  lw ��T�,ju;! ���q��`�q0n�v){/����  �$����T�n��dCk���Ώ�����w  �;w �-�y�u� ��z�8�}�0�zw�T<U��9�J ��i�.���֚7��I���_�˿��G>r[�  Xg� �Q�y��< �2?>��8�zw�T<U���Z�&	  G��Y�y/���ȤK�R|����'>�3�[  `]�@)V�E3n �:?6�l/�x�֝g�� �8���x�褳g���������-  ��|a���j5���  l�7��7n��<W��R�zw  ����}��j��?޹��nw�1��  ��� �SkCZ��͸ `�~.�u��x����J���  �*E��y������o��������  �uc� ǥ�!�<3n �>'RZ�}��8S��RN��   ^��a����#7����+�;  `���1h������ ��~J��f�3���jO� �����^Ժ��jv����c���N�  X~� G��1�2�d��b�R;���"��q(�- �i�R�q6;�/A8�kMO׺\D��- ���)��&)ED�y7�c�q�ػ6���o{��[������w  L��; �V�,�:���Rjo�����|�z�|�� �f���9gzw  }|��ݧk]�� ^YJ)�֝H)�0\���&��/|�~����s�����w  L� ���Rf���w     �+e�J���(]���w������'�|�  �2w 8��Y�ո     X;��E+e/Z�Z8d�����]w�l���N�  �*w 8l9ύ�    �u�j��Z�F�p���|�ĩ/}��;  `������њ�W     `�Zg������y����~�{w  ���!h)V�E3n     6��r�OF�p�ҽ��������  Sc� �/��j�     'E-�}o���5��;�����G�Z�  �_>���     �`�����;6J�i������O|�gz�  �T���jmH�ռ�     �!E�{F�p�ҹs������O}�M�[  `
���ֆ��̸     �2)r�k��z��&���w�_��ý;  `
��j�6��     ��J)�e�á�x����]��  ����j��      ��&w#w8d���'�����  =���jm�����      �Z�{��y��)"��_�����ڻ  z1p�+qy��;     `JRDԜ�Qʢwl�TJ��{�W��{�  @� �#�Zg��      �,ED�u7j5r��r�ܘ����祐|�w
  7w x��E[�<�     x)"Z�F�p��yf�z衇zg  �q3p�W�j�i����      X)���{);�[`S�<���/�w  'w x%��4_     �JJ)�֝��p��:�����  p\���Zw�V]     �Q;8o�\8����7���n ��`� /�J�us;     �!(ea��#]���w����v�[z�  �Q3p��R)���E�     ��Q�"�b��`x��=���  p�� ��     �J������江��{{w  �Q2p�R���      G�����������  G�����JٍZ�;      6]�uF�p�Z��K_��S�����S  �(���J�us;     �12r�Ñs����㛷�~c�  8l� l�Zwø     ��պHF�p��/�<p�  8l� l�Rv��v     �NZ��T�N�Xw�O��������  p���.���     `Z);�#w�N�}�������w  w �F�uǸ     `:Z�F�p�j������?�я���)  p����4G     &�պ�q��\�8��������^�;  ���; ������CQ     ��j�9���ax�ٝ�����;  �z���R��v     �iK)E�y������#o����  ��a���uQs��     ����Ƚ#w��{�y�o��?��  �����T뢕��R�]     �J)E�u7�6���*���_��O}���Z�  �� l�R��;      �j)"j�K#w�v�ܹq8y�K�;f�[  �j��QRk�V�q;     �3r��7<����?��{zw  ��2p`c���5�q;     �����=Zs5\����������w  \w 6Bkm�rvs;     �I9/��;\���X|���ѩ�n{W�  �R� ���Ɣ�2.?�     `��tp���;��ŋ�p������E  X� ����9�q;     �&K��^�f� �`x��S���}�;  �J����J�%7�     l�9�5#w�&����������  ?�/} ���R�y?|�     l���M�.@���Z̿�����m���w
  ��@ �Ok)J��c      ['EQ��;\�t��0�<���g>�ӻ  ^�a  륵�X��S      褵�������3����so�  x5� ��Z�ɸ     `륈1j]��u4���������Ի  ^��; 룔e�:�     �D�:�R���j��w��}���w
  � w �B*e7j���      `bj�G)��3`�\���w���O}����S  �����Rv[���      LT��T�N�X7��gw.=��=�;  �����T�"��     �Z�;�V#w�J���+�}��w  |��; �Uʢ��u�      \���˓�*������O}�?�;  "����f��ݔR�      �DJ)Z)��ڬw����ᮻ�y�  �0p`�Z#�i;      W+ED伌���-�N��|�������  � LKkC���=     �5H��^�fW!�<���n��ӽ;  �n��0��f�     �������\�Tk�����ԧ�Ի ��e��4��"��	     ��3D�{��������ɓ'{w  �����Z�1��      `���,
�B�#����_����w  �����JٍZg�3      �P�΢����V�������ʿ�; ��c�@_��D���      l�ZQ�N�Xi�J����Q���� p���&�6o�z�     ��h����;`]������?���{w  �]�袵6k9��!      l�-��hm���b�����?���;  �� ��ژr^��3D      8N)rދ�l&�J��]w����o��w
  ���5 �Wkɸ     �ξ7rwfW �=;�|�w��  `;�p|ZKQ�^��     ��������?~�~����  `�p|j]Fkc�      �l�Z��#`]���߸����� �f3p�x���Zg�3      ���:�R���J\���<���3  �l� �T�N�:��      ���y���;���䓯��#w  ���; G*�6��z     ���Zw�5o$�+�8y����Gn�� �f2p��6��wS�      �RDD����ػ&��Ծ���ÏB  8t� ��R伌��     `���2Zs�?���3�O�����  lw ���}/|�      �~�Vʞ�;�h�����c�Ч{w  �Y8|��F�W7     ��Rk��3/����'�O>��7�N `s�p�R);Q�w      \�Z�֝�0u������{;  �� ��f�C>      6D-e'Z��K=���>���ݻ ��`���hm����w      ���6�n�Ik-Ɠ'��o��-�S  X� \��R伌���      `����2Zs�!�93{���ٻ ��g���9���      6��J�kF��o~������V�  ֛1" ק�݈�JF      6ZjmLgc��i-fw�����_k�  ֗�; ׮���u�;      �E��(e�wLY:{v<���_�� ��2p�ڴ6k�zx     �Vi��Dk��0e�o|�������� �z2pવ���y�z�      �1K9/[kc����b��W��ß�ԛz�  �~��:����2.?�     �-tpf֚33x��g˯~���  �w �N����      ��3�U�=���>��;zw  �^�r��F���      0	��R);�3`�Z��=����O��w
  ����+�ڬպ�      SRk݉�\�"���셓'��� ��0p�Gkm����w      LL���y��`��~�'������ �z��
���Z���q��      �CR��l�9S�W�Z������O>��7�n `��xm��F��;      &��1���`x�ً_��zw  0}� ��T�N�:��      k��y�u�;�j���~��[n�d�  ����W���J��      �B-e7Z�dx%�F����; �i3p����R�ˈH�S      `���h9�Ek����g�Y���_�l�  �����J�k>#      �����J���S5�{�O�~����  `���>���䕉      p]Rkc*e�wLQZ�Rz��ܻ �i2p�%��y�uѻ      6A�u�Z���)�x�������w  �c�@DD��Ɩ�$      ���w�7(�+N���o�~���;  �w "ZK)�eD��)      �aR伌֜��H�΍�G�|�  �����Z��3      �D�R�ަ�`��#�8���f�  �Ø`˥Zw��Y�      �d��y�uѻ&��H'O�WO}����S  �w�m���J�      �A+e'Z{w���'�N}�w  �`���ZK��2"R�      ��弌֜��|��8}���� @� ۪���9       �*E��ꀗI������w  �6l�T�"j���      ��T�<j]�΀���N��=��w  }�l����J���      [���h�n~�x�}���'?���  ���6i-E�ˈH�S      `��ݵ��^�������w  ��l�Zw���     �T��Vo_�0{��<u뭿ڻ �>��Djm��{w       �պH�9ǃ��5����  �a��ZZλ�3      ��rލ�l8�e��O�?����N�  ��/G ����,#"�N      ^Q����5gz�r��{��گ��w  ���`åZw���w      �ơ֝�0%�a��#��w  ���`�����E�      �G��,��Y������y�[���  w�M���r��      \��RD��֚=|O�1�����; ������y�w      pUR*e�;&�g�����; ��a���R�;1��       �Akc���;�d<y���?�?߻ ��g��iZ��]      ��j]Dk.���xqH=����  ���l��Z����w      p�R��9����#����������  �h�l��֝��v      �c:8""����{w  p�� 6DkmVKY��       O�u�Z����{�����  w�M�Z���)y;!      l�Cλњ�@�l�կ�������w  G��`Ժ��m      �EQ�n����f�����;  8� ��E�:�      �Z�5�p���?��G>�ӽ;  8|� k��6D);�;      ���r�m��z@D��*�G���;  8|�� �����zg       �"�Zw{G�T�������O��  �p���RvR��;      8F�μ���b���C�  ��;�j��Q�w      �A��֚˰ "��O�?������  w�u�ZJ��FD�      t�R)��5g���������zw  p8��M�;�6      �n���֝�0�����O~�w  ���`��6k�.zg       ��Z.ǂ�׾�3O~�#?ݻ ��g��&Zk)r���A       ""ED伌�#���j�꣏���  \?w�51�^���     ������0���O�~����  ��J����Z�w      0=��E�6���R�Q|��� ��1p���R�띂      �+I���+���'�xã��ٻ �kg�0u��D��      �W��8x+4D���׿�7zw  p������y      \�V뢵��,�����.O��}�g�  ���;�����      �J)���0�W���������  ���LT*e'"ܮ       \�1�a��^������w  �2�    IDATW��`�ZZ���      ��u�ل������蓟|K�  ��/3 �JYFD��      ��g���҅��G�l�  ���;�Ԕ��Z{g       k��1�5����W���ZU�w��v��l�I"d 	A�@0�0c�顙�p��bP��%DG	QB"R��"AJ�H�3�� "!{<���az�O�ϻ�֛��V��O{�z���<R��.vZ����]e��+�s�_���  <9w�U1�	      ���l_��aئ�:~��?Ύ ����Bjk�K)5;      Ѕzg	�6~����x�9  x2
� ����hm�      �G�6q�4��Z��_���  <w��2����      th6�W"�$͠��{ߑ~%;  �����\�      ��ܞI M^y巳3  �x
� �"&��Iv      �c�m�sI�����9p�+�1  x4w�DQ�tjS      �x����fi��R�/���9  x4w�D5b_�,      �cT#6�C@�����<������  <�R%@���l��      �41�m�}m���_��  ��ya�2��w�      �d���?;�z��w{���ώ ��)�dhm��2Ύ      Pk���2կ���3  �`
� �Q�l�/;      0\m:�_"\:�`�.\�<��O�Qv  �2w�%���+��P      ����;�K��׿�\:4�� �_���L���fv      ���f�g�,�K�6N|���� ��H�`�f��V�      ���R�t�?;d����OǗ��6 ����,��>�      �3.��[��z����7��s  ��)�,CD-��(      ������Q3X�W^��-�  �C�`Z�_���      �bꝙ&R�rer��W�gv  nSpX��Iim#;      ���l����e���?��?  ��)��tj�      ��j��N���s@������W��߳s  ���X�mV�Z      `=�kkJ������8tȌ  ���D���fv      �'��f���9 ��ҥ���'�5; ��)�,Jk�K)>�       ���ΐM��͟��  0t
� �1��6�c       �Tkm3"��9 ���ō7>��?�� 0d
� ��~��     �uTK)#[����/��� `���Fl�Rl3       �V�6)���a|�������9  �J�`�"��tj�      �����%���R}��/eg  *w�9��m�V      ����2�s��~����� 0DJ� �Q��;      @b6۴ŝ��x���� `��極��v      ����ھ����=�����of�  w�y�Gk�1       歵����a����� `h��a6�ou;      УZJ���@MN�|����� `H���Fl�
      ��Ek�1��KQFG����  C���5�S�
      ��M��K�˭�ё#:���?�� `(�����Y<K     �aՈ���t��v��e�  
�L�݊�q��      01�m�����^�맟���s  ��;�.����R|�      ��ޙ� �[��ӧ�Wv �!Pp؍�Q���      `٢����9apꫯ~��/|�d�  蝗�ݰ�      .[����룭7����  �Spء���      ٝ-����l����q��$; @��v�����v      `�j)e��fvX���59����Av ��)��Dĸ���      ��Ek�wh��+�eg  虂;�N�f��#       �3T��;����>��9  z���"&�       �#bn�fp�����  �RpxR���       ���ff���������3?�� �G
� O���R���       ��׈���T���g��^v �)�<FD�2�mf�       XU͍�����?����� �w�Ǩ���{^      <D-edqCS����o}�d�  ��&��DԸ]p      �jk�Q�s�2�_{��eg  荂;�#Ԉ�Z�0       ����b��ҥ�ѧ����  =Qpx����      xr�m[�����Rv ��(�<Lk����       ;Q��Za0Fgμ�������9  z��� ����      `�a�;�Q�����1  z��� ��v      �ݲŝ�>����/���  =Pp�_D��      v�w�f:�����  =Pp�_���       {Sk�fvX��k��@:4�� ����Q�lf{;      ��l�i�;CR�^����sv �u��p��lo      ��Z[�ŝA�8|�`v �u��pWD-���      0'њ-�J=s���z���d�  Xg
� wԈ�b{;      �<�b�;R#���''; �:Sp(������*       �f�;3:|��g���wf�  XW
� ��v      ��ŝa�yst��7�Kv �u��`{;      �BEk�a�;2>z���3  �+w`���M>�       ,H-�V[����Oy�/d�  XG
���E��      `ᢵ�b�;QK)�';; �:Rp���v      ����������>��=���s  �w`�"���      �g6�ŝ���n��+�� `�(��5���      `�F�wd��?; ��Qp+f3M       �,f37m3�s���x晗�s  �w`�n0�      X>[��v��gg  X'ʝ�0�X      �&�S[���c������ �.܁���I�g�       ���-�1��w^����1  օ�;08�5�        ���/;,������  �.܁A��q�f��       C�٤D�0o���Ƀ?� `xI ���Yk͎      0x�V7p35�LO��w�9  ց�;0��f{;      ����6J�-e����OġCz  ���GľR�#       ���[��k�����O'; ��Sp�!���l#;       Q�f���3�ȑ�3  �:w`Z�,��      ��Z#,,cF'O���/}�oe�  Xe
��0��c      ����l3;,Cm�\;r��s  �2w�{w~��y      ��F%b��at��eg  Xe
�@�b:�K      ��پ������~���s  �*w�kq����       <Z���]ar��W�3  �*w�k�5��      ք/C1:z����K��� ��܁~E�b6�d�       �ɴ�6"B���ݼ9:���!; �*�B t���Yk͎      ����a�;�0:~�@v �U��t)"j����      ���6J�mft��:���{��G�s  �w�K�v��      ��Sk)���hu:�������  �F����       k+����������  �j܁�D�K)��       ������6:{�]'�{���s  �w�?��%?      ��3�eZ+��g�Sv �U���%���&�1       أ�&%�fǀE;�w�3  �w�/���      �����3�ܹ�Ǟ���9  V��;З�6�#       0'f�@-����;; ��Pp�1)�k       =ݙC�FǏ���  �B臫�       �f�@���8y����s  �w��hͯ�      z��$"t\�^;q��  ����Bmm�f�       `�j�=���V��Xv �U������md�       `AZ�(��ѵz�����>���9  �)��/b����>       }���IvX�ӧ��  ��;��f3��      :��fvX���?�  ��;��"b\Jg�       `���q��u�k�ڵ��<���9  29�kmԚ��       Pk-�5[����ԩ_��  �I�XkM�      `8Z�dG�E�8��  �܁�1����       ,ͨD(�ӵz�����_�� �E�X_��      7}3 qꔂ; 0X
��z����qv       ���I�p�7]�'O~Wv �,
��Z���,       ����N�F�/O?���9  2(�k)Z�dg        ��;0:}���  ܁��1��      @�q��{�k��'?��  ��>�v�_�      ��it������� `�܁��Us       �lfvL��o���  ˦���Q)�RJ��      @�ZJ-���H�ӧ�;; ��)�k%lo      ��j�L���N<��g�  X&w`}D�hͯ�      (���MJ�[��WDi�����  ˤ����6}�       ��F��N�N����  ˤ���p�       ����,���Μy������k�9  �E�X��      �_6��qvX�:��o�����9  �EYX��      ���IvX�z����  �E�X��      ��lfi]�:���  ˢ����W�y^      �0�;�e�R�qct�g~�W�s  ,��(��jk~i      ��E�-ӷs�~%; �2(����Iv       V�lf�L�N��Dv �ePpV[�$<�       x�Q�g��E_��y���$; ��)�+���      ���mdg�E��=���3  ,��;����       �PX�F�Μ���  ������I)�f�       `m�J�8;,����wŋ/>�� `�܁�e{;       ;e�LϦ�z�ԩ�ʎ �H
���ru       ;
�t��;w ; �")��)bRJ��1       X/��zg�]�9��  I�XM~Q      �.U7�ӱz�������  ������Z|l       `��R5zQ��ʎ �(
��*�Rjv       �V�����ٳ?� `Q܁���       �Q5{�c��7ߟ� `Q܁�Ӛ_�      �7f�t�^�>:���(; �"(�+��q5;       k���qvX���ۿ�� `܁�R��      �y��Ȏ �2z�����  �
��jQp      `^f33h���[O����d�  �7w`uܾ�s	      �y�sh�Tg�z�ԩ�� `����Qmo      `�Z�Ȏ s��g�#  ̛�;�2B�      �93��g�����  ��������c       Нq���!`!.^�<��ߝ `�܁�P#6|M       `�����ӥQn�?���  ������1      ����̤�V�;���  �I��QKk��       t��I�p�8]�g�~8; �<)��`\n�
       �P��l�3�ti����Wv �yQp򵶑      ����&�`jke���d�  �w ]��       ���Mӳ���Tv �yQprE�k)5;       ���qvX���o8; ��(��Z�Ȏ       �0�[���ŋ�^��_�Xv �yPpr�u<       K���;]����s��yv �yPp�D�hM�      ���R�%�f�E������  �����Lj��       �娷���N�Ξ�Hv �yPp�Dk>       �Tf��jt�¾#/����  {���im�      �a�f����R.^�Jv ��RprD��g       K��"Bɝ.���"; �^)�)j�+�       HQ[3��K���#; �^)�)B�      �<6�ӧ��ʎ  �W
�@��|,        Gk�Q�c�����z����g�  �w`�"ƥ
       �R�w:Uϟ���  {��,]��dg       `�jkf�t�^��3  셂;�t�G       ��f�;]��ν/; �^(��QK��       ��R�%�f�y�[[�>����� �[
����}        ۝ٵmt�F���˿�� `�܁���M�3       @)�3l:.�Dv ��Rp�*Z��w       VC�6]���ǲ3  얂;�<5|       `EDk�Q�s�ܝ?���  ���,M-eR��       ��Zk��L�s�����z��g.; �n(�K��(       �ji�M�t���K�8; �n(���        +&̲���Ofg  �w`9"jDx�       �R��q���9`�.^|v ��P6���2���        VK-wJ�Йz��f<��� `�܁�p�       +jd�M��tZ��f��� �S
��RD��       �$��U�|��3  씂;�xU�      ��e�;�]����  ;��,øf'       �����6zt�·eG  �)w`�Z�dG       �GRp�C�K��eg  �)w`��Un       �:w:Toݪ�<�Lv ��Pp�z�       ��,o�S�[[/dg  �	�S`�n�½f�       ����m��.^���  ;��,Tu�       �c� �mt���3  섂;�P��      ����̸�N�x��  vB�X(/�       �3n:4�y���쳟�� �܁ŉ�%�s      ����KD���y��/dg  xR���"�k��      �z��N�:S��~ ; ��Rp�Fx�      `���̺�N\����  ���;�0��      ��ѧ�?[[�ʎ  �ȁ�	�j      `ݘuӡ��˓8xp3; ��Pp#��Rjv       ؉(eT"̻�J�V����9  ���;�(~�      �ڹ�lש�;uk��  ���8��M�#       ���yӣ˗�Nv �'��,��       ��̛�ԭ�eg  x��b�6Ύ        �ҚNݩ[[���  �$Ɓ���Q)�f�       �݈R�%�ܛ��+W&��K��� �8
���U�       �؝f��7]���7����  �� �]�gg       ��0��G׮�tv ��Qp�/³      ��f�M�.]���  �� �]��W�       �5�o�t���#  <��;0_5��      ��7����nm=�� �q�P�y���      ��W�n�]�:�C��] +�a���6       �`Nof�z����d�  xw`���=       ��Э�;׷�?�� �Q�j�s      �.T�:4�r��3  <�C80o�+       t���s�3�z���  E��QK)5;       �C-��۳p�Ǖ+�͎  �(
��ܴR�r      ���Y8��r��  E����j6       :S#�k�����q:�� XY*�<y�       �w�3����g?� �a���i�3      ��D����Nm���  F�'�       �b�;�]���  �����B_�s       ���aNW�W�~4; ��(���y      @����˕+�͎  �0��\TW�      Ы�qv��+Wޑ �aR��Pp      �cf�t�^��G ��r��"<O       蕥ot�N���s�}ov �q��5�       �f�th����3  <��7�w�w       zUK��`ަW��Pv �QH�,Jy�      �c�D��Еɭ[��  � �����:       �gCW���fg  xo`�ZgG       �����δk�ޓ� �A��=��      ��Uw:3�v
���    IDATmv �q��,<K       ��8ݹvm#; ��8x{ךg	       }�p�9}�ys/��Tv ��)���%      ��E��ЕQN]���  �s��$n��+�      лj�;��u�Əeg  ���;�'�s      ��0#�+q��'�3  �ϡ�W�      0��ћɍ��  p?�n`OB�      ��h͌����Wߟ� �~����Rjv       X3r�2�~���  �Sp�$�:      ��]zs��fv ��9t{b�;       �њ9]ݸ1��  p?w`���      0�6�e{��4 �rP�݋�E�      ��wf�Ї٬����3; ��܁��      `P¬��lߺ���  ����Z�      ``�����͛ߟ �^ʩ��Ek�!       �Y9��y��  ����^�~�      ��T�r:3�~�#�  ���^��v       �Ŭ��ܺ���  �Rp��K;       ��6��ƍwgG  ��7�{�)�      0,f�t�޸�Tv �{)�{�      ��(�ӗ76�#  �K9ؕ���      �A	}:3�qc�� �^��n�Z��      �ZJ)�ё�uK� X)'��TW�      0P��ӓ:�ַ���wg�  ��a�-w       ��̜�ܼz���  �Rpv�Fx~       0H#w:Ӷ��'; �]
���D��u       )Zӹ�+��>�� �.�m`W�_�      0\f�te|��G�3  ܥ��JxY      `���M�y��  �Rpv��:       CefN_f��eG  �K�؝ּ�      0H�sCW���{�3  ��얂;       �f�tet��;�3  ܥ�얗u       ���ә���?; �]
����5:       C
�t&n�ڗ� �.w`�"j���      �Z������Fv ��܁��      ��)�ӓz��8; �]
��nxI      `����h{[� X&���:       CW���HL�zd ��p0vl�%       �u6� V��;�s^j       4��ӕ�J:4Ɏ P��;���       f�t�o}�C�  JQpv���       �2)��  JQpvA�      ���֌��ʾ��gg  (E��/�       ����y�և�3  ��        ;V��p������  �(���-      �A��s���  �(���       �/���fg  (E�؅hM�       �#m6{Ov �R�       `7,��+u6{Wv �R܁����ػ��F�,=��8�KDV��=�G��XcdR���"�� ��� +KU]y	�q?��Y������       Б� !p.�w       6����Lӗ�  "��xI      `�2���.�; �w        �T)��ѕ�ֻ�  "���#�       l����V- �J���Ru;       @gjݵ�  !p.4Ex�       菖 X%�E��}�	        \Y֪% �C	p��xt�       �3%���  !p.Tw;'�       "J�ӏ�; �J����s       ��l= �h�	 A�        �q��]�  w�B;�       �S25! �"�        6�F��E�).�       tgp� X�;p�����       @ojՄ  �����n�z       ,Cq𚎸� ,�����e       �?� `!�� ���bl=���a���Vc(%[o    X���r����-�)|� �&p B�\����<��C��+    0�/�0}��Z� �k�10})~��e���׺       �n ��܁��K�{       ""2[/  ��U��LӮ�          �$p.R]p      ����z  �H�
\�n�;       ���  �K�\�m��       �z   tH�\��7        ��  0�*p���          ����Ȱ���       �w�R�< �A�
\�8���7       @k�� `w�"%��       hM�  ���2Zo       ��2[/  �.	܁K�{E      `��wzS�H � p.�9x�      `��  0�;p1/�       l]I�N_�D K!p.Vjm=       �� �,���Jq�       �#�� ,���\��      �M��� ��        p�R��  f p.�;       [Wk�  �%�;�w       ��g����� �A�\,��      �u.�ӛR�� ��;��
�      �:���?� �R܁�e�w       6���Ng��A �e���      �q�g�  0�;�^�      �4��� �B܁�yI      `�|v  ���Z��       `�j2��
  �H�X��wR      �Y%��;  �B�\N�      ��e� o �y܁�MS�       �L�:�����u ,�����       lX�,w  ����XN��      ���L�� �L���J��'       @Kw�R�H �!p>$k�f      �6��  ��2�kt       6�Q8  �������      ��*w  ��@�_�      �F	��N�# ,�����u�z       ��w  ����/�       lTN����� ��܁��      �QC��'  @�����      ؠR�w:��  ��;�!9M��       ��2b()�3ŝC `9���LS�       p{�C
� `6w�C�8��]       6'kB�  ��3���:       [���m�Kq� X�����      �M)�>+ �	܁+~�       �1w��; �0�T��2�      `Sr}V  3��|X�u�z       ��49w  3�Vj��      ����M�# ,�����&�C       ،���4��W�w `aĩ���q�;      ��"���z\�� X�}�����w       6�ֺ�;�q� Xח���y��      �fdwz�' X�;�a�V_S      �v��cr  ������u�z       �B���З�o6 ����|��w       6"��g�  03������       �0��]������Ӵk�       nB�  ���R���;       �+�1M�g�U�� �	܁�9��      �{�+��g�U���%�������      ��M�.���w `�����q��      @�2u6t'U �y�>�K<       ����q  ����e���       `Neu6  p��ϛ&�;       ]K�;�)�� �_���<_�      @�ql=�K� ,�(��<�]p      �[��]��z  l�������       �Uk݇��Τ� �B�R�O+�s��l�       �Pj����; �P���ˌ�2      @�j���  `+��U�L/�       t�����; �P����iڷ�        �G�  ܈�o�*r]p      �?��8�[���r� X0�;p�t��      ������ ��	R����y��#       �ڦi�q  ��;pe�z       zSkݵ� ז.� &p��dz�      �+e�5t���� \M��u       :�糾��� ,�p�jr��7       �5��Y	  7$p���N.�      ЏZ�1M�W�u�� ,�����q��l=       �!�i�cp  �%�;p=�X"�      ЇZ}�9�q� X8�;p]^�      ������?w `�<�W�Ӵo�       �B�N�� ��y�k]p      `�JD����;)p N�\��(p      `��4��4��  �#p�*ܳ�       ��R�o���v `��U�Z#�n      `�r���G� ����iڷ�        �r:	� ��;p}��      �U��IWCwr�c ,�'��N'�;       �U�~��+  `�����CDd�       �9M�L{ӡRZ/  �Cw��Ʊd�7"       V)kݵ� W'n VB�̣�}�	       ��t� @#w`�(p      `�N'���� �J܁Y��$p      `}jݕ�Y	Lwr�� ���Ey�ED��       �u���n��6 ����8�Kz7      `e�8��r��E� ����M�&/�       ����k=�N� ����M��w�7       �%�񨧡?w `E<�����_�      ���c[�  �M��y{�gD��       FN�>���th�� ����M�5J��      `��7�ӥ,� `=���r�Zo       �?�x� @cw`Vy:	�      X����񨥡?�� +�����>[o       �?P2�1M�g�ե� X�;0�r<%B�      ���4��r�T� ��܁�e��'        �v:�ZO�Y�����;���'       ��:u4t)� ��x0f����      ���Z�y:��鏸 X!�;0��a���3       �WM�^L�� �
	܁ٕZ#3w�w       ��G�iӥ� +$pnc�ZO       �_���o=f!p VH��D�w       ��:��QL�� �
	܁�8���g       �߫�t���l:$n VJ��D�ޜ       X�qܵ� �� +%pn&���       �{y<�[o�Y����7���]�       �7��xT�'�; �Rw�v�}Fd�       ��E��W�,R� �����2�^�       X��}�0� �bw�r��[o       ���x��'�; �bw�����      ��j��]L�r�� ��I���p�GDm�      �m�i����3`.� +&pnkK��      @c9���  �&2no�[O       `�������� 	 ���ps��v�K�       h%k���XZ�9d� ������ᮔ2��      �6�i��t��N	����7Wj��ܷ�      �F��>��_w `��@y:=��       �F���ZO�Y���܁6����}o       ��4��tR�'�; ��;�Dy�EDm�      �m��t�z�%9 �~�h�62#�O       n����`6.� ������       6����^�>���Nx`�9�JDm=      ����>����� ��h��ϥ�=      ����y�z�F� tBX
4���C�       lCy{�ӭ�` @<� m���ED��      @�j�����5}r� ��h�翎��g       з:���7�l� @G�@S%3�V�      �Y�����`6w �#w�����![�       �g����d�V
���xp���R��z       }���>km=�#p :"p��R3��g       Ч<��Zo��0 �/�n�exh=      �N��:�F�\o :#p��p���      �u�zWƱ�
�M
���܁E(�㐭G       Н<��Zo�Y	���܁�Ǉ�       �Kw�5ȿ ��x�#���p�      ��uW�G���� @���b��a���;       �C��}�0+��y��#3rZ�       ���]�	0�R"[o  ���X�<�|      �Y��!�޴1����  f�!X��׻���g       �n�o�w�� 蓧`QJf�i�q       |Jy��3]K��N	܁�����l=      ���u��AC��� @�<���//�����       �)��>�i5:&p :&p��1M�*      �ɷ7�9ӵd_ @�<� �T��#�      p�����a�z��w �cw`�����0L�g       �2���s� 蜧`�J�Q���;       X�����`V�� ��������      �?���î��S�� t���X��r���;       X����Hw���� �܁�*�����z       �oo��7��� �܁E���1"�y=       ��֡Z�6� ��X����O�;        ��>����-]p 6@�,[f�8>��      ����'��\o 6�S�x�����      �J�C:��z; ���+oo;u;       ������ޥ� �Fx�V!O���       X�|}�o�f�z; �!w`���}D8�      �?�Z���]�K�\o �ē���N�      �?9�\o�.� "p��x|l=      ��y}�k=fU�� ��;�//Q��z       ː������o�v `c��z�NCd��      @DD�����`v�T �O?��Loo_��       ��Z����o��.� #pVex~��al�      �Ʀ�>jm���z; �A���u��R�g_1      �u��ώ�� � O@����뗌��;       h��]������  ps��)���"p      ج<�\o��v `���*�����       yy�k=f7H� �m�����c�2��      �m�4����5�K�; �Q���u:�KNӾ�       n�pxh=fW� �]w`��/��g       p#����k=f�z; �a����ʗ��(���      �m�8>D������$�VɌ8�[�       �6�����])�� �4�;�j���K�p�      �w�tW���z�-]o 6���j�x��2      �������	�; �q���իoo_|5      @�j-���o=fW|I ��X���t_�al�      �y�4=�Z[π٥��  w���<�}      @�^_�[O��� ܁>��˗��Z�       ��j��ۛƅ���z �"x��P�}��      Н|l�n��v ���=9�FD��      �Ք|z�k=nB� w�#����0��      �u��鱤;gl@).� ����F�5�x��z       ��Q���[p� �o<]�?�f)��      ��4���TZπ[H�; ��x2�R��R���       >'__[o��(�� ��	܁�L//_��o�      `�jݕ�W]���]�	  ��E �����o�      ���ǣ��l��  �@������       +Tk)��w�g�M�- ���Х|zz(�L�w       p�Ǉ�|��F� ��'$�K�����W�      ����}�	p+YJ�	  �#p���Ǘ���g       �'M�]���Y��� ~��$�_����Z�       �Oz{{h=n%�  ��Sе|}���z       ��!_^��g�M���?  ����Zyy�+���;       �}y:=F�_�F�� ~���^=~
W�      �������ݮ� ����+OO1c�       ��<�b�Zπ�?{��    IDAT(ŕ> ��!p�Wk���C      ��Ɉ�����;�V��v ��%p������w      �����!N��z�L�� �{��6�c�����       �Qy}�Y.�1ȵ  ��'&`3�?e)S�       �U�w���_a3R� ��<1�Q��!���       ~V_^��� 7S���  �]w`S���OQ[�       غZ뾼�jW��� �OM�������>      ����[O��Zx���d�  "O`�������R      �H�u���}�p3�,?T��z @��ؠ��r�z      �����K���p=�]��� �R܁mz}���       Z(���0��������Rt �"܁M����      �\�_���3�v��$Z�� X��<=\WɌx{s�      ��2#���[π���Z/�S�pe ��;�Y������      �v���2��W�픲��{EC ,��جRk���e-/�       kW��Zo�[ʕ\o��Մ� @����}��e�s�       ��q�/�si�n���G>�A� ,��ش2���N���       �OO��w�M�K�� �"��)
�������a[�       ��4���Sa[����z @�� ��\�tz�g�       ח?~��ζ�YJ�q X
�;@DTW�      f����z;��۵^p��; �^ ��+�y:=��      p=�������]o��(�ݩ� ��;���o?��      p=y>����+��/��z @���o�8��      pE����v6'w��>f�w� X�;���o�~\q      ��:����=k��e� �"���
`eK=��d��      �����v�gŁ{�c�  w��߾}-��+�       �z;�TJd)�W|X� �E�(�X�w      ��p���Z�����2o�7  D�~ݷo_�0L�g       ����lT�<p�axo=  B���~����;      �e������������� ��;�o����0c�       k���P���z��꯷GD���o�  w��6�����      �Y?~������������ ��;�������;      ����!N�*_��n�z�u���  !p�}�X�x��      ����xzr���)%��������O�  w�?����p�      ෝN����E9��_������ ��;������_�w      �_���C�	�DG��������  "� J~��%K��w       ,M���ir����(n/�]��w�n ,B?OY 3*��//��;      �_e�%�p��M�ݮ������o� C��'���os       �_�_Ku'���z{DD��I" ����I`^���/�;      @D�P~��k=��-p�� �bt��0���r�~w      D}}���3TJd)�W\����z �/D� ����_"bj=      ��Z���y�z4�۵^puywwn� �w�K����4��=      `����k��D���#"��N�'  �B�������a��\      ���4���9a��N����ZO  �E�O\ 3;��<�3��      ��zzzl=Z�N���� �����o?���w      `3�|~��w�	��i��wwϭ7  ��ߧ.���c���O�;      �?~���f�n�z�|���'  �B��?~|�a�Z�       �[=���\Z������/_��� �_���0�Rk���_"���      0���ZO�VJ���#b*�?Zo  ���ೞ��0�     �n����R},�FCd�3����n� �w��ʌ�Ǐ���L��       \]�C|�~�z��C��������  ����� n�����4�3{��m      `K2"���O�w@3����s���� �_����?���ײ������־���3���!Eʒ)Q�2,+p�H2$Y���YQ-ܦA�(X�@�]((�-(3R,�I��i#������k(��N|��h�\���s����#�C�C���ۗ��'5|�2:k��ٿ�����z\�      ��L&�tpP�΀b����n��G�x�F� �0p8)��U>:�ǭC       f���R�(&��pz{�zM� ��������U5)�      𠚣�~/���`No��ȝ��� S�����������      ̬�4)����;��E9�="R�7*�  p;w��6ts�b|�      ����Rj���[���#"��;,�  p;w�Ӱ���S���       �gMS�`�.��,���M��_� �v� �a8��x��9�.      �k9"�`�\���lR��n�N  �݂]���fss%���t      �]��qxhO��J)�ܛ^o�t ���j���85+q�      ���#R���l�Qw:�)�  p�Ż"8Ci{��      �,�y4J�3��E;�="�i����  �[�+2���s4����Ҥt
      �5M�۝�PT]�.(����t ���NY��k�ɤ����     ��#���[�4Yp�xz{���^��Kg  �n�� �^��\Ku=*�      �C�������j������G�ۤ�^;.� p;w�3�F���Kq��      ���#"���Kw@q�xz{D4KK��  o��Wf %ln.GUMJg       �i8���q*�%-���KKG�  ���������E��;      P^�T���-��-�����=(�  �v�{uP@��m7�I;�      ]΃�rdO/Yp�|z{DD��S: ����X��\����       W3���p������������W: ���
���8����єN      O�H���/���E?�="�����	  og�P@���5�t      ������dR��J)b�Oo������  ��U@!ys�\��q�      `�4M+�v�(θ=""�n��n  x;Wj �����9:�GD.�      ,�fkk�t�Rd�Hu�������  x;Wj %mn.GJM�      `���q*���.�0���I� �wb�PR�D3�E��;      pz���[[��P\J�~��tT: �������y2i�K�       s(GD3��g�����4����  މ�;�4��\����/      ��F�txh#No�����	  �ć�i0�|p�M�      `~䈔����;`8���r����  ���`J���^��      ���9G��_J/�����~�_�N  x'� �ds�\��Q�      `��J�A�tL���������  ���`����j2.�\�      �q��˥`*T����&G�vοY� ���L����H�)�      ̮��p9F#�^��5p����#o�q�t �;q�0eR����SU�J�       3�i괽�.�S��";������N  �w�i4����R�z+      �]��lm���i��t�tZY�+�  p'� S*ol,GJM�      `v����t|�j���L��$���,�  p'�� �T�9������ƥ[      �闛����ۥ;`Z8����KK��t ���L�ttT����$      pGyss�tL��wW/-�^� �;1p�ryss9�d�      �Q><\J�Q*�S�2�z7���_J7  ܉+9�)�r���q>�j\�      �BMӊ��N����*�0���|��ם� L-w�����8:�G���     ���[[˥`j�t�w�WVF�  ލ�;��h66�#%w      �M��p)���y��t��kVVK7  �w��r�fs�|�4)�      L��i��v�tL��";��=嵵��  ���`����GG��p�;      ,��#om-�΀i���~W���*�  �n�fL��\����      @9�p��ǎ������ߕzy�wK7  �w��r�fc�TU��-      @MS���N��*No�k�^�WK7  �w��������rD8�      L��\)� �$�u��3"w����_�f� �wc�0����R���}L     �E�#���_��(�n��R�@ݵs熥  ދ�;�Y�s����Tף�)      ��L�i0h�΀i�[��	3%��J7  �w�Yv|\5{{k1)�      ������r��*)���]�kk�)�  �^�f\����ɤ��H      ̟�wvVRӔ��t��I���,�  �^�����ZT�S�     `���~:8���U����ø��ǥ  ދ�;�<�LR��}>�d�      �i����΀����{��*z���t �{1p�i���݈ȥ[      ��#"oo/G�n��ڃ�����FO��/��  x/� s$ol�4�#      �����ȶn�RD��}9~�t ��p�0GR��"�I�      ���ɤ���ۥ;`��.�0��s�]� �n�̙t|\僃���      3*���R��:)����YY���	  w��`mo��i��m�     `��ȃ�J��V��6No0���_/�  p7�����ZU���      ����ǽ�߷ⅷ�*��?�V+_{���t ��0p�W�q��윋�I�      �.�\��f�tL#��?�|��qz�5�� 3��`����v�;q�M�      ����lo�����]n�J'̼|��v� ��e�0�66V�)�      0�rΑ��ph�o�ҭ_<�ɹsV� �n�`0�&���QU^5      Өi�i{�S:�Q���	s�^]�?J7  �-w�����fww5Rr�;      L�Ԭ�/���i�����'d�����  w��`A���;�:�K�       ����ժiJw�trz����~�~�wKw  �-w��66VsJ�     �h��ph��ĸ����K7  �� Hj�����"b\�      Y�L�i{�S��RJ�+����z軥  �+A�Es|\�����$w      (#�����0����OTu���]� �^�,����q'"r�      X4ykk55Σ�wTU)���+yu�WJ7  �w����W��     �l��å�5��������n秮^���  ��&��r���8U5.�      a2i��v�tL+����<��0���]  0S���q���E��     �iʹj�חKg�Ԫ���JW̝|����  ���`�������ND��-      0�����8w
����"�?�/J7  �+w "���dw      8��p)�6p'u��)�Ν��  �O D�9bc�|Tոt      ̓<��c{�S��VJ�+�S�j�'�}�(� p�\p��q����&�'���׿     ��)��/��i�=�>5���k���  �W� �)�4u��/�z��T�t      ̪yss55M��^U�R銹�.\�^� ��a��[�kk���W��ou�_o��     �Y�#"����ё]�IJNo?e����t ���A
����r���^���~��[�W��      �{���{1xc2����W]��F� ��a����G���Ո�$彽^�����g:����	      w�i괱�+�S��"��Ч)w:����z� ��a���:/�q�.�hT�ᰓ������N�h      L��4�Y__)�S���y����  ������H++��Ї����ѨU_��z��L�7�     ����;;�i2�P�M]G.ݰ.^�v� ��e�@DDt�_����ٶ����z�����?�:�2      �n9"���r�0�ݤ����L���n� ����H�v�?��;��yw������J����{W      �&���N�tL��r��Y�;�ߗn  �_� D�������U��Ij��zQU���O���V      ""��N����0�r]G.�(VW'�~�+��t ��2pXt)E祗�����f8�D����S��F�      ,��4)ol�D6ۅw�R��L�4/n�n  x�\�����Cw7V?<lE�T��s��S?�7       X`y0X����P�^�t�B�/�a� �a���:��rO}�9"�W���O~�}JY      0�rΑ���������|�,MΟ���  �-�V?�xԗ/�󝄼��M)5�_l�_|�um      0��hԋ��A�{I)�7���v;���~�t ��p	��:?�c��/�LR��׋���'?�j]��}r      ,�����f�t̂\{�|�&/��^;.� � �Tu�\��{���Ѩ��a'�:�?�v}钟)      ̵����J�\:�^��t�/�A]��g�  �1"����rDz��	���<שӉ���v��w'      �K9"bkk5�c��ཤQ�%��/^���  ʕ$�J�n�?������n7"�Z^����I�����      0Er��_�����B���	�)��}����  xP>x,���/Ft:'v�D3�"�\_�T�>�َo�     0/rΑ�å4�J��,�u}�w�\s���ʗ��G�;  �"�����\�~��gӤf0�GJM��պ�?�w      �C�tbk�[:fBJ�@��.]�Q: �$��X0�| ����]~2Iyo�)5��~��~�E'X      0ۚ��7o.�΀Y��t�Bky�wJ7  �w��y����G�*���R���'[�k�ܽ      `&刔76VRΥS`6����)�:�˥  N��;���~:�G=�;
���<������ϴ�K���     `�ln��xl�w#�ȕG�%�s�FW^��Kw  �W� �{����&��ur�)u:���N����      3!GDV��Ȧ�V��ޥ�G�Y� ��0� ���~�3��5�A/GDZ^N�/|��:�3�{     �};<\��}k]�[u99󬸋���	  '��`At^~9"���*��#���""ח.U����N�}      �X������&�[)E�̏��������  '�&�HKK��Ї��o<�����M)5���u�ӟ�o�     0��ɤ�76��;`��V�t�WW�׾��,� pR�@����V�̲|4����nJ�i?�\����h�      �;ɹ����s����=5�#�l�n  8I� �Պ��/�m�����󱏵:ׯ�?      S!G�fcc55M��U�2;��.�~� ���J`�u^x!��r���o��ߎ��RD�}���?���      �#"��W�hT�y̐����rx���(�  p���YJѾ~�tś����#"R��_�K�֕+~     PJ����qxh�����ӤY[?���s� ��dX0�Z�<�ŋSs�D��<�rJ9WU��s���%?�      8S9��GGKi0h�n��RU���<�&"���t �I3*�c�W^)��Ú&���U�D�����ک���     ��������0SR�\{����\��OK7  �4w�9U?�h�W�L�p|2I��n?Rj��r��j'z��l     `�L&����/��Ƹ}
������t �I3p�S���t»J�q����H��.\��^}��Z��Y      ̳����7WJg���u��Y6m�GϾ��?/� p���PZ]��>P:�W��Rj���z?�S���h     �4M���WRΥK`����N���cV� �4���C��_�������pX���vD��3���O}���      �����%s�    IDAT�jL&D�=���=������  ���`Τn7:�H�{����y<�SDn}���'>�.�     �|�[[�q|l��ȸ}z���;��Q� �4�̙��?����͹��N�4U�ȝ��[��^r�     �����#�^UUx���j.]:��o�(� p|��'U���KWܷ<tsD�������:/�P�n     `6�����i�3'�W)E��љf�c�}�t �i1p�#�矏t���~�>ED��Ӌ��SJ����v����5     ����p)�v��E���or���X� ��̑��/�Nx`)�Ȼ��F�U����t�}���W      ܵ<u��V�t̤��H3{��B��~s�k_��;  N�� ����z*�'�����Ij��z)�&�u�}�s��O��     �{ʓI;����;`&���hv�5O<�^� �4�"��pz���x���=Z�����;���ǀ     ���4u�ys�t̪�j�N�n<���V: �4�́���h����3N�hT5��ݔR�~���zm��     ��4U����r.]3ɸ}F����Y� ��d�0:����|��ú;)�&���ޗ�ԩ�����+      �%G�fcc5M&�S`6UUĜ>r�7���_�f� ��d�0�R��^(�q�[��q;"ru�\�{��N�tJW     0rD�ki<�΅��R�.]�]ʏ?��J7  �6w�����"����Y��ߎ񸎈\?�H������.]     @A9�ț����x����ii�Jp�G�j� ��f�0�Z�h�c�+�L����dR��\?�x����;�I      )GD��YMGG�p�r��tw-w:�����7�;  N�y 3���FZYY��(��n7rN)"�W�Խ�~��g      �&����C�!������P��gߓOn��^;.� p�,fX����	E4;;����{�ڵ���O��x     X)"7��+�����WJ��-{�L{�J7  �w�պv-�G]�Uw����)"�����_��F�      s.G���`%��-0�R�q�,��Xz����t �Y0p�Q��_.�PT�[#��u3��`���B�l      �%�1.��τ�4�V8<l�4�>�����[�*� p�fPu�R��{_��RΑ�7G�_lu?�q�u      ̣��~lmuJg�L�*���<��7K7  �w��y啈[���4)�������~�ݹ~��     `�4�ǽ����R�.]�}j~���n  8+� 3&-/G��,�1]&����{��D�����      ́<u��F�t̼�s�fU>~t�_���  g��`�t�_��k����d���^/���R�'��~�y#w     ��'�vll�Kw��k�n��Lj�|�OJ7  �%w����h�c�3��x�&{{�H��U����t���sF�      ��iZq��rd�\x U99Cm�=���.�  p��fH�������.�h���^���{��5#w     ����nn�X1n��R����Y���|�G~�*� p��fEJ�y���a4���A7Rjr]���~�ݾz��<     �Y�4U�ys5�Ãk�J���˗o��^;.� p��� fD�����CNo�[GGu>8���{��\���S~�     L��4us��Zj��)0�Z��5�ٗ�|��n  8k�~ 3���+�f��Q�|�$�h�R�_贞|��>     �)����7o��Ã�u99?m�۹�r寖�  8kF~ 3�~��/_v��~|�$��G��c���     0Mr����q;���"*�D�A��[O���m��  8k�ff@��/�0۾?rO)5�餥/~�S?����      ����ɤt	̾�"�Z�+8!����*�  P�q���Ν���ϗΘ}GGusxxk���W_��/:     �����͛�1{n(ED�u�NJUE��c�Q� ���\祗"RrC�$�>r��S�K_�֗.�Y     PB�Tycc5&���4�Vd���F�����Ϳ�ǥ;  J0��b�ۍ�G>R:c��6rO�~����t��     ����Nn��QU��s%?��7J7  �b�0��/���q��i�~���     �B�Ta�''��u]���S�������  ��L������+���G�_�R��     ��}���l�'&�Z�8i�>����)� P��;��j������;M�a�;F�      g���v'���1n�O����� �B3p�R��^*���pؚ�Nr     8])on��I�����I)ң����  %�L��駣z�qw"�H:<��p�$w     �ӑ�����<��RU�+��y�}t����v� ��\�L���/�NX8��e�     p�rӤ��͵d�''��u]��S2~��+�  P��;���~8�g�-���~0r#w     ������Z�=o���R�V�t�$��K��j� ����L����n��[����I�?�3���y�}      ܋���͛��p�>ߚ��{�+_��Jw  �f�0E��R��GKg0��������Rj]��.     ��j�*ol��q;���jE$��ڕ+�S: `�L���>�j�#1�����N     ��i�f}}͸NXU�ϻ���C���  ���`Z�Z���GKWp��������     ܅������4��.���R��K��]���Ͼ��?/� 0��D�G4���O�Ѩ2r     xw�iZ͍��x�'*�ȭV�
�@~�Z� `Z�L�����K�+�#w     �;�LZq��Jʹt	�'�/�T�9]����;  ���;�h=�LT/:�}��F�dw�o�     ���d��7o��q;��V+"y��&�/o_����t ��0p���_.��]H�qjvw��-     ��ɤ7n,��)�������|��n  �&� �U�<��O���n��)�����     ,��n�X*��(WU�ʤgQ�N'��z��/� 0M\����#"|�~�L&���     ,�<u�͛��pR����������}��~�t �41p((��F�G~�t�c2Iyw��k7    �E�s�||܋��~��K)En�JWp�&�/�R� �ic�PP祗"����j2Iy0�EJ�     �\������-0����N^Y�\�����  �������F��Kg����="�[�v     �M���R��4n���jE$g�-����uz�q� �ic�PH��"�]w(�AӤfg��sNF�     ������J�����Uב��ӓO�ץ  ���;@	U��^*]�	J9G���妩��    �y�#���[M;;��-0��*re��������W�t �4r�P@���"�?�+�s(�f<���     �a9"���j��m�n���R�.]A!��O�t ��2p(���+�8M{{�||�N)5�S      �U�H����-oᴤ���#��b���?[: `Z�R8c���Q=������A+���;�9�B     0�&��͵4y��ȸ}�5O<1x�+_�g�;  ����sz��ȇ��|x�u�;     0�������pʌ�IW����  ����U��G���/����a=����     �,7M+߼���q;���jE$�Y�t���O�{�;  ���;���rDr�bѤѨ����#"�n     x�<���ƍ�h���)׵q;�\��g���o��  �f� g$�z����KgPH�S��u�;     0U�hԍ7�#;�NS����L��橧���  �Ε3�i����/��$5����    ��rΑ��{���/�s/���.]�h.\8~�׾�s�;  ���;�Y�JG"n��wv�NA     
�y8\���^��{)En�JW0-����/�  0����7�ǿ�;V�D�9���^n����     �����W��v�t,�v�TU1y����t �,0p8CG����7�a�L��������
#w     ����`-�v�X���._�����~�wKw  �w�3v�[����}�f"""�<�RJM�     `~5���\����t,�V+"��L��k�\� `V����c����?�#wn��o��F�     �)�)����ё� ���jE6n�v++����ϖ�  �>���s��?�����;�[y�g�     �������w.�Fֶp�������3�����kǥ;  f��;@)M���1�ַ�ܹ���ʻ��d�     <��s�ɤ�o�XM�Gp&�*re��ۤ͓O���  ��U5@I�I�������ȝ[������	     �䈈Ѩ7n,G���DUE���L���'׾��,� 0K܁{Rյ�N�F����.r�d����~���     �9"��`)66z�[`a�d��姟���  f��;pO�Ng^�v��h���F��3)��;;�f<���     �Ky0X���N�X)En�JW0�r�ߴy��-� 0k�T�{��:��O^>:���=��~ט�?����GG픒�'      w�#R��\K�����3d�λi�y��{�~�t ���P�K�눔Jg̝|t���F���a�9<��     �$�\�͛kqtd gȸ�w�#b����t �,���o��2r?F�n��zF�     �[4M��qc-�c��,y^�{y≽g����W: `����t��F�����ǭ/�     .�F����D�|8K�Պ�99�a�쳿Z� `V��k�NǛ#��o���s�qʃA/r�d�     �*7�a?����C`�ԵC�xOyee��/�;�;  f��;p"��OG>:����w��y��I��N�i���     NnV��V�t,���\���ޚg��fz���  ��U7p2R�0r?Nr睤�������:�佣     � rD�����.����۹;U��'���  �̕7pb�����á�;�(��u��î�;     ̷�i���~.��-�p�*r�w�y���+���{�;  f��;p�rJ>؟�<����J47n��V�a������    `NM&�t��Z�R�X8��ܫk׾\: `��'.W���)��Nr7r��F����ӭ7�     �/7�ǽ|��J4ι�3��q;���p���/��^� `���"WUD��bNC>8���}-��~׈���LR���o��2r    �ٖ#���_I��-��R��j��`�4�<�ۥ  ��)pjr]���<�:��;�1b�-RD�`�ͣQ+��(     �Qykk-�����۹�N>�x��*� 0,O�Se�~z��Q|��1������!y���F�     0cr���7ϥ��C6(!��v����g���_��o��  �>�.���� ��|t�_�zL��O���!y8�'{{}#w     ��I��qc-���A!��
_�g)Eu��X: `^�g"�ZF�$���ZL����gᇤ�(5�A?�)܋    �)����^�qc%5έ�R��۹O�˗w�������  ����1r?=y4��_���[����$坝^n���  ��g�^c-��3�?��־�SW0U`(�
0�.P��f���T<�(��vҶb;،4���H��hZ�h$^��h�%;�Q:qbn����)�!]��6q����c���U眪s�9g��Z�߼8U6v����ߗ�G*��T��bW�����g   ��%y������ ���}6�O���/��   0N(�(�Q��}�����3����˕��̌�        ���`���I�˥�Y�I�=6·o�����C�:v  �qB���q8�~�B�GU���Qr�k�2o�*��       ��=�ɓ������ȳL��5�Cx׻�c�   �e �<Mc�_�K��?O�oȻݴXY�Qr       `�\���䳳���j��g�y�J�+�]���9   �w q�����#���u���J�xC����j�d���       ��so��|nnZ��<��X�k^����h.v  �qC�@<���W������_�+��xc!������g��       ��|ii�����9�I�i�r;�_��/���  `Qp%����_���O=E�o��,�v�"J�        ���0?�Y�V;
0��TJ������/_�rf�b�   G��@|f%�u�{�u�qI���:��WVj,�       �v\��y9��m�<g.�-I�۱F®]�6v  �qſ����zG����%w��<��^��L|N        8_�������9v�Ky�K�F.��y��~�   ㊂;���frJ����o��I!p��7d���rŻ�k�        ��,,.n�z�; Qnǚ+�����   �w Å%�u����W��_����;�\���F�J�       ��B���M��p��Xc�ys������9   �� ��Sr_w�K/����R�G�o��O��rM���g       �����W|vv���b� ��X�u����qG;  �8��`(������*^yE��w:����B�^�Qr       �My��A'N�b� p
�v��j5�W_���1   �w ��L��a]ǎ�}���f��2ޔI���w�%3��        0L\2_Xؤ��R�, N�܎u���������/��  0�(�j�$���Y17��̌|a��;�Z���F�J�       �UB���M�v�{��v��2�/��3�s   L�=J��/��j:�0;K�o��O��rM�L��       �T�^U��T;�S(�c�k�y�ꙙ�b�   ���� b�y������x�UJ�xkEa^�WC����       &QXY٨�'��s x��D�s翌  `RPp0:Xr_w�����ʿ�=J�x{�F9�ZQr       L��p��fk4��Q ��v�3����+���s   L

� F�Sr_y������쳔�����ԗ�k��$>3       �q�!��>7���}���Pn�:sIv�5w��  0I(�9�� u�|R�������W��z��<5��       c�h46������`�Pn� �;�.��;  �$��`$Qr wu�~Z�#G\,s�x�Q�v��;       `l���'6'++Y�( ~�v�_{��  `�Pp0�(�F��Qu{L
��;�^�����$7�       ]�y^ss��߷�a �������<���  0i(�i������j��R�SX��+
�z-�y*J�       ������2�:��1@a��/��   0�(�y��#�%���Z���m�$5e�t�fb�       ���'~��f[Y�bG�(�c��t�x��ߍ�  `Qp0(�Fq�Z33�J�83�N��k��Xs       /�</���&�z;�7@�f�w%v  �IE��ؠ�>aqQ�C�����3S��Z��T��       C(4�4??%�J��1`�ys��n�\�   ���;��B�}0��T���U����8#&I�F�;���B�<        �b:yr�-/�b�&(�#�p�uawܑ��  0�(�;�$�,�c�y���W�����M�g��I}e�&ɍ5w       @$.����������܎|�Ƣt�%���  `��`<�Qr��y�Iu�z��2�\�[��k^�(�       "�fsZ��S�SC�r;"�ݻ��_�b+v  �IF���2�(�D�g����]!p
�3b�|e��NYf!v       ��!�'6��r)v o�Ӕr;�����֭��  `�Qp0��T��b� ��|G�/Y��(���u:�//�\���       X?z����nR���0�<M��:"ٽ�?^<3ӌ �n��    IDAT `��D `칙K�����Z< o�(*����^��n�d��       �AX^�h'OVc� ��(�#���m�   �L
39%��(�SkfF��IJ�8;�v�*%w       �ZpI^���m�f��"`�QnGd�u���Ew޹;   (��$��&,.�53��G?�䎳��'E�>�L�w        ��VkJssT;����r���k��^{�?��   �x: 0Y(��w:j=���瞣���b����w:e��       8K!�D'On���r�, ޞg�vDW���̎�~!v   ��	��1�(�FQ�����9�b�g��I}y�&ɍ�       ���z����w���,[��"�Z-,����  �L$7�J%K�w��:�KyNIg�(���Z��3c�       �&\RX^ި�'kr�#��@�C�����ff�b�   ��Pp0�\,R���z�y�ũ2�^�Y
�F��;       ��\���i~~�5����e��d@d>5��k?;   ~w ��������̌�ɓ��q�����ק�i��       0��;��fg7(Ϲ�F��*��=���_�   ?��; �C�A
��j�̨x�
�8k�._^�x�Sf�       &����f[\����q/�a�7�m�Xo  B��S�;�zH���Srǹ�tҰ�R3ɍ5w       �$�</���7���f��b�={��;�\��   �� �:�eR�_���j?��zO?��s����Z��3��      `2���>??e��02(�c��M���Xo  R�8�x�Rrwu�~Z�G��h��f�T���Ě;       �+�</���-�lf�� 8�����	��=fw�ы�   o�' �O�բ;"���Ժ�^��2�d�c�       ƕ�Vk���-p����R�ys����+v   �9
� �f�D��>0�ܜ��ޫp�%w���f������      `t�$/������R)v g)I(�cx�����   Í�; ���e���P��!��?O1��O�z}��<e�       F�{�5����s��YJޖ��.��w�7|.v   �5
� �v�$J�j?���O=�b�����F9�ZJ�       0\����'���R9v g�Ӕr;�Zػ�O�;��9   ��(��p3���]�g�Q��a)�)���u�iXZ�)_�       �a��n����&��YmFQ�J	5/���?����  ��Ǔ �)J�����W��L1�.��劷�e��      `���$��<����J�< ΍g��r;�\�{����   g�� 8fR���3���S��{������ay����>O       �{�W�c�6����UY��)��_q���?��;   �� p�\���7j����~�R2�OQ�/-U��)�5w       �&�����f[X�����y�ɹ7Ős3����wc�   ���� 爒�`y������{䈟~_)p�:��Ys      ��󼬹�M�v��F���~��?�u��}�s   ��q`  ���LJ��t�zG����/K�.�d���k��n�5w       XA2��7i~~�زF�v��4�p�U�;   ��L 8O����,��P����9���k���k�ƚ;       �������7��Nc�pN�ہ���\93�W�s   �����5�i*���RX\TkfF���O!�5w       X!�$,.nf�IB���\�ގ�<v   �=
� �F����^O�GQ���\,oc��5w��g
       ΙK�ݪ��m�N�{i`�%���0B��{�^=3�\�   8{$ �Z:�J>��c�����3j�+R�K!�(L���t�ƚ;       �w��-,l����XmF��)�v���d��_�   熂; �53��.�%5�W��INʱ6:�4,-�Ě;       �)W�[���7���.�eR�g�������/��  �s�S �3�TZ�N�TkfF��/SF���|y���vY��      �rI
!	'On��b%v k$˸��H
\н|��O��  �sG� ։�Ԣ�>坎Z_��zO?�buk��M}i��y�Ew       x=W�]���M��q)�3y�ɹ�Ĉ*n����;��c�   ���� ���E��O?���K�.%w��L�F94�U3�(       L6��p���묶��v��bǎ��=��c�   ���q	 �iJ�=���ռ���y��X;�^��)��T��      �LZ����h�>-X`\$��r{��9r3�����9   p�h[��x�Ji;��	j��(���v��F���$g�      ��p/������R)v k(IV�3��W_���C�   珂; �'��+�0P��}��:O<�
�"2�N���z����Xs      0Ƃ�bee���6(�Ym�I�Rn��+��ع�7c�   �ڠ� �frJ�Q��}V��7��ܱfL���R��Rk�       Ə{��5;�%i4�� ƌg��H0��޽��<t��9   �6xJ�̤Ri�gT��j�}���^���5eyn^�׼�-�5w       #���y��I��S8��N�q_���6�۷�j�   X;� ��"�F��++j:��3�Prǚ�v;󥥚B0��      `�����t��f��i�< �ة7N;������33s�c   `�Pp��<�$^�7x!���S�|��<�莵���r%4�U3���       v��H�ĉ-��X�s�	��S�vF�0.¶m��<��9   ��hT��4�������wԼ�n�'8������bqq����5w       ��%�Fc���m�~��+0��d���3ٍ7�^�   X{�`Xp�M8qB�����.%w�9���f)���N��9      04L
��%���b++��y ��$apc'\}�Ov�w���  ��G� ���Wb��U��G�y�	W�����|i��NY��      ��WX���E���8��o��8*��ع�7b�   ���� ��L*�V����}V�{���ܱ>:�ԗ�j��Qt      �K�N��c�6[�˝10�<��	�1~�{����=;   �O1 0�\��M���(�W󮻔���ܱ>B05��hT%����      ���^���o��b5v ��L�c*lܘo޽�Wb�   ���� C̳LbQ!
�v�~�u�q�@���O�^�y���5w       ��%�������`yN�gf����1�n����_�B=v   �Z� 0�<M�4�c2��w��Z< o4(�c�x�Y����%��      �!3��?���,v �,IVG��1.�l���l�   X_�`x���BQ����w�x�e��X?Ea��T�N�,�`�      �WI8qb���O�s��;O���,`\%��ݻ'v   �?
� 0"�ԫū��VK�/Y���k�c��N'��T��Lf!v       ��%�fs���nR�ǝ00<ˤ�?�o���/�:t��9   ��x��Qb���N�=����7պ�~y�A���ܥF����5���B       �^�^E��[ly�;�`$�k���^����  ���� #��Cl�+��y�*~�J�X_Ea��T�f�̂��        o�B�'On��'k
lf �r;&H���;��~;   �v$ �(OS)McǘX�j�����{�+J�X_�^R,.N�^�$� �#      @�ճB����ݨ^��_`R$�j�� �}{��Ç#v    0�<I$��qW��Q�ff��:�c�+��V+�����̘`      &[�^���j++��a P���a��L�={~/v   w qΫ�+�S󮻔���ܱ���|y��ͪ̂I|�      ���BN��j5㍏�dɲ�,`B�~���z��?��   ��S ���%w���nW�GU���]y�m�_�����T�vKb�      {~�GXY٨�ٍ��|L3�T�3z�IR���kׯƎ  ���b  �OS�$�����{N��j��']�	#�_��y��jj�o�R.w��      ���:�)��Uہ	tz�
�0�o��λ�~!v   ( 3������m�"��La~^����=�-#S�Q�F���9      q&/����jq�*����I��H��[;������  �8(���׭8L}��*�rK�D��{=�\�Ç]�.7�~?�z���nIf�(�      ��]����Yss-�yc(0�<�Vǭ�I�$�o���1   w Wf�RIJUn��j���T��j��_xA�;�T��S4��ۙ/-�B��2��       8s.yh��u��fu:4[�	�Y&�m�d*������{O�   ���; ��4�̔��cS����͛c'�8aiI���W���\!Pt�`�`j4ʾ�\Sf�     ��f<�K>;�Ֆ�ʱ� ��L*�(�cb�ƍE����`�   ���; L 7�̔l�nS����+��i��3Ϩu�}��EJ���0_^��F�*�O�       0$L
^Y��ߪ��ilU +I�Y�A>&��tӟn��?<;   �� �ͤ$�U�V��'T��ؑ&R񓟨y��ʟ��IV��x�^�N�,�`�     ���%+7knn����5�,M�i;�_q���_���;   �� �%y�HfV��V�}�#�R)v���ݮڏ=���în��1��IC�>��LfLA      v�P�C��Aǎm�N�F+0�<�V���	�Y��={~+v   �,v  ��y��ܕ��mS^��GQ��cǚ8�^Pq옪����]�2�ܥf��Nf��=�i!wN�     ����L�z�j��	0����@����ˮ{����9   0(2��r3�L���6���*۹3v����Ժ�~��~���f`���|y�VVjr���      ���E����V-.Rn %	�v��p��������9   0<(��s��5�j�j��_�|�-�1$>p!����j=��|i�[����R5�Z3�ӷ$      8O�!XXXآ���s�ȳL���c ��La����_�b+v   
�  y�HfV��V�}�#�r9v��T��wީ���R.F�nZ,.N�n��$��      �;���Fc�fg7[�˽, �lu���)৊����>���s   `�p� ��Ӓ��뮳��nSrᅱ#M$�v�y�	���U�N�r1�$��μ^�y��2�u�      �qw�Y�v{ʏ�j++�ؙ 	���?�7�={~9v   
� ��r3�LɅ��m�)��ؑ&V����'���i#�������$If!r"      `���*~����+G 8��t�����o������   Ç�; ����{�l��\�[oeI"o6�~�au���s�8��|i��F�$��       ��/�,��o�����" �N�I	���v��z��;   �OQ �7�I"�Y��[�����*�ؑ&V�����җT����O���z���vY�      Ir!�'�hnn��9k1 ~�L^*��A��+�=\}�Gc�   ��� xSn&7S��w���+��ؑ&V��պ�~u�z��b���^�׼�)�,Ew      L�{⋋�4;�Q�w� ~^�ȳ,v
`h�n���w:�L�   ^�  ޚ�<Id�7�ԧ?���M��{��ffN��T��:�4,.N�n�D�      �%yh46����餱Bi*O��x3~�%�]�=���9   0�(� Έ'���V9x�j���\�ibǎ�u�����ߺ(#"��v;󥥚���%I;      ��N�zh6��ر���R��	�p�,[�S�Ʋ����>;   �OV �3�I"�)۳Ǧn�M�EŎ4���W�?���O��H�q�`�l���Ҕ�<�Y��     �hswɬ�N��Ǐo��e�_ �13�TZ�������ϗ�}���9   0�(� Ί�II���m��[�ݻcG�hŏ��w��(k(�������nfbG      ΉY��(�����b�t �f�du�=v`�����+���[c�   �h�� 8k�SkU?������J��5���9rD��//s~����|y�R����]�     02�
��,��]���i��3�7�e�4��z��n���;��cg  �h�� 8g�$����{m�ӟV�eK�H-�e5��%��}��;���ii�Z��VK�|6     0�B!�'�j~~��9�v o�L*�V�|�m�����W�{�}�s   `tPp �7�̔l�nӷ߮��kcG�h����j?����
eb�n7���)�t��     0d��`����fg7�����[�4�g��
^ؽ�}�{�   -�  Λ������V���T=xP�u�Q���j�韲����a��^�Y0��      ��]RXY٨����t8����LJ�Y g,I�8��wtbG  �h�� �f<I$3+8`S���lÆؑ&�O�ܿ��F�"1��IR����ũ��Rt     ���.�oбc[��(�`�I��ꛍ��|߾�/��;   Fw ��r3�L�6}���v�i��/���w*���(ch�$��?-�[��     ��V���v g'I�Y�6p�|˖��{9v   �&
� �5�f�$�MMY��P��[W�-��Zj?��?쾲�,���{��8]Pt     ��sI�++��1�2y�Ǝ��$�����c��P�   �)�  0�<Id�V����\��}M�lƎ5��_T�WT����?�:��0�բ{��Y��[��3w�Sx      �,���i[^.�`ĘIu
�\���=�}��A�   ],� ֕�IfJ��¦o�]�Ν�#M<�v�y�	���e��e��1TN�C�>���Ew      �%���ִ;��r;���$���s #ʷn�m޻��c�   �h�� Xwn���>=m�O|BՃ%^�]�����/����1���K�f��;      ΐ�Y���;�5YZ*�9Np��L�p�D����_�B=v   �6
� ���$�̬t��M��J�l�i�y��Α#j:$_X��'S�Y
KK�     �F\?+�_`�z�b;��f&�J�o&p��n������c�   ��� (7�̔\r�M�~�J�];$����]w���3.��C�(~Vt���Ҕ�;     �ds��ݮ�S�v�h�9�4�g��y�/얯��c�   �x�� 87��D*���яZ��]V.ǎ5��W���Ժ�>�'8��p*
S�Q���EB�     `�����Ǐ_h�z�b;�s�e�wV ΋���o��|��؊�   �'5 @.ɓD2S�w�M�v��m�bǂ���Լ�n��1܊�|e������g�$�     ƛ�,�v�N�B�L F���TZep�����ͮ����9   0>(� �r3y�(��B���6��8L�/��}�)5�K�'?�4��U�f����B���,Pt     +�R�N�������Qlp>�T�e�S c#l�־�[���9   0^(� ��'���V9x�j���V�	��ܜ�33�<�ף4��u���KK5�     Ƃ��C�5���/��b�x�$��a&ϲ�;) k�Tr�|��;��Q   0^�Z2 `hx�H����.���bo?���W_���?���^R�C��]�bb�+S�Y*Z�RR���Z�)��%>�   ���� �ug���i[Y)��^_kg� �9Iy��N���K����w�}8v   �
� ��b&7�m�dS��[����Q��ߔ�"v��獆�_���k���>$��    IDAT۸�R����[�Rh�JV��V��l�2��-   p���~��)v ��J����%%��N����a�KF����,[����
;v,]��c�;   ��� %O)I�|�-6��O)ٲ%v$���������=��"	C�$������T�tJ2�s     0<�D.)YXP��?T��(9�7 ր��T����j5���;;   �w ��r3y�(y�;m�s�S��bG�)��s�Z��/_X�	C�$���|qq�;�2Ew     ���T��z�_�Zl�я�.-�N`����r;�u���=�\}�=;   �Ot ��$R�bՏ~T�UWy��'��~�T�T��wީ�����[n����N'�NgJ�ja�Z�$�;_�     �䢋T=p@�m�d�E��ѣ�cf�4e�XG��k_������9   0�(�  ��K�$��)ۻצ>�%۶Ŏ���\����Լ�.���"6FG�����Th�*2���     �u�^v��~�״�WU�-[d�����<��G>"+�cG0�du��r;�n¦My{׮���  ��ǂ; `t��͔l�fӟ�����-u��-)�Ia~^���Si����*������M�۝�J��Z�'3��      ��L�Ν��ۧҦM�<���휥ݻ�n߮�#�(�8!(�QG��$Q~�Ϳw���;
   �w ���$��Y���W�s�w\aq1v,H����=����Ty���t��$q��ѰZt�y��MM��,�=�4v,     ���$*]{��{�(�VeE!��[��/��g>��7������3�2j� ����]�g�.v   L�) #���I���Km�s�Si��ؑ�:��s�Z�)��{�<�ٰ<7-/W����,I
��     �+�T޿_�~�7��T*�V��g��+�>�QU�Rv �5OSy�qx@ؾ��������  ���W� #͓DV�X���3e;wz�'��v�X8�x�U5�[�o��> �J��ct���J�Ӵ�j5O*��BH��      ���T޷O�k�Q�.�K!����T>p@���j>,o6�6,��g&O���v �Tr8�)��^�(   �� #��d��k����.��7�����b��iE��ѣ�_zIՃ=��jN�1Z���l��V�d�jn�jO�&��     `���ͪ�ۧ�ΝJ���K�o ݱCӟ��ڇ�x�5��qI�Zn00����.���ñs   `�������{?`/����9p�*7�,���_�4���J%+�ޭd���"���o����Q���^avV٥�ʪ���\b��$�y�N�$)�R)73�y݋��$���v7�   �z2K�4�Ď �/پ]���G��y��6(Y�b��Y��Ҿ}RQ�������w0��L�$�S %\s��ˏ�9v   L� c�%)Id�Vڿ_��y�1Ǐǎ���_|Q��P������{��$�Ga�t:�w:S�\vMMn&�?˅Y��)w XgY]���G   �|�)ݹS��S��dy.�����&�*�ުd�6u�xB����	`���D�6���{oѷ�;
   &w ���Sk�Ʌ��m�y�o�F�o~�5�!����O?����W�C����(�c$Y�g��2e��Ԕ�e����&���� Xw�=O(�   ��J%���Q���Vz��#����{�ҋ.R�G�����Y&W��%���ϫ���WbG  �d��] �����k*��ʷ�bӟ���.�����S��!uܽ���y�sey�tyY�Ғ<��5!.]     ���iU��^m��'�a�efg�����\t��o�Mٵ�F�` ���@$�7��>���s   `rQp �57�'��w�Ӧo�]�86��?������=��+��YVJWV���R�O�     �����T��Vm�����UW)�s)�ر~�*�>�1U�x30��lu�@�⋛W��}�M�   �l< &�'��T�����v�������ш�㽞�O?��w��������I+�+%ͦ�j�+�jU2��e0     �O�)ݱC�={T޾]I�+�z�S�+8�d�vo>,o6c���(��y��a����w䱳   `��� �����]�l��ە]sM�Hx��I�|P�v_^f���]��(�ו4�r�~�     `X���޽���k�>��-������aӟ���K/���JS��@d.�x�{�rf�bg   xo����������c�����|�T.���zf�R�J�]g�ƍ*^}U*�ة����w�,Sz�%��c�4+
%ݮ,�W/kJ%%ժ��Q��%�� �^����?� �|�%E�Vb�  ��d�VU��M����nۦ4IF��sV�Xi�>��Qq�X�8 ����v�A������+�񍃱c    ��W� ��df*�p�eW]�'�T�⋱c�x���_��z����z�k%w�<�sY�!%�ljJS����R��U��x�6     Xf�.�L�}�T޾]I�#���S��$�ʯ���K/��O�{�؉ �OS����\�ݸ�=�T�(   �$��%�G�o�N����m�;ޡ�?��<v,�o���y�ɓJ/�TV����s�幒Ng�M;v�|��J7nTh4�V� 06Xp�5; �$�TTڷO���jW_�R�����1�\t�eW]��G?��۱� x3��åT������w�ɟ|;v   �4
� �
��C����$%�x����UX\TXX��
o �8����J!(��R)I�lc,XQ(�veE���U��z���B�s���{� 0�(���� #%ٲE��n��>��E)u����b����}

'OƎ�%�j��8������^��C�&v ���ޝ�u�w��=�9�^l$H Aw$�k��HN�I'�d��I�;q��+3U�L��j��K=USSS���Ju�����m'q�Φ$vK��ˤ�E�)S�
�$ @,�lϼ8HٔD�8w�~�P�i��S�s�{��� �V� ������!c�Нm�/M��;���wde;;����a�T&��}�2��7��m�l(�z��$ �K� P&� P����۫�GU������"�$2�v��`�6ن�gϲ< �lm*R�u���o�Ѽ�    ~���   Tg��s�n5�==n�;�Q|�d�c�6҉	�<���c�\�SO������Ԕ4=-[,���
{�*�я���Ѽ'     �44(Tq�V���L�$MO�=V�L��lG���˿���k�<v��&mk���{��Ky�   ��EX6�W6����Ww횢Ç��������QSL����H�k֨04���_����Ii�� P�� e�w �8^g�x@M�>��U��T&�[�[�+L08����&'��/lm*W��������W~��(   ���X��C�~�ɂ��v�ءtlL�իyO�O���(:rD���Y#��{��$���Lʶ��߰A��A�bQ�Ą\�=" T,w (w ���`�5>����Thh��"n��D�X4�ΝR�(�{�>X��휪*Rr��;��3�{�s    ������W�{�6��ǊO�R|ℼ+d������c����,v�}y��*��%��K
C�׮�=" Tw (w ȕmmUq�>5=��֮���1�0^[��ӧ%6�����@�K7m����߽/�9   �O��=   ��Y+���[MsO����w�<��X��+���?��i�kx�)�+�Q{�����7;+��
�����*�vM���
�C��ټ�     ��Z���*��)��C�̌T*�=UU�M���n���\��h�� ��Z9�{@%K��±���W�   �T��� lp�>lp/#cd��)L�m�ܫ@z���Ç�(���-y�j�IS�0�-�d�[��А�erׯ�MO�=" �� P&lp�%c[ZTػW�O>��u��#E�sy�VLS�)l߮���W��=P���T� p�����_3�Q   ��B�`Aܫ��"0F2FުU&رC��A*Y�*Vt��L�(o�j��	�,ǲ��2��[�Z��;��J�)��4�`��@����V���P�C���*/�dX��8|���2����9n ��<��k' *�;p�O���O����    ��;�!p�>m�U&�����'䵶ʶ�q\��ݺ��,[&Ӧ�[ݧ������@�������*�ܩ�'�T�ƍ
<O6e�I})����}}�O���(�y����v��$������=��   ��"p� �Շ�}���6�kה^���T�nfF���J���uv�47s|��9'E�Vwke׬QahHA�$��@] p�2!p��V~O�yD���j��8f[{Nlk�	�|����d�� �����lm��[�z�߳g��;t�;�   P5�,�{�!p_"s�ܷn5~W����0�{*|�t|\���r���֮��8A0I�mtCٖ�7��c[��<w (w �gs�ڛ>�95l٢ ���	߮���&عSJ%��y�T&c䂀��"�Xt�#��b�W�z"�Y   �� p� �Շ�}	#c��ʕ��k��J.^�{*|�tdD���R��[�V���5�ܲ�]��c�;�G� eB� w�Z�׫������*��ɋ"�(���{:�����M���7 ��KyPU�Q��ÿ����?�=
   �P�� �Շ�=�����ׯ7��@�X[�"W�$Qr��wߕmi���$��ǲ��Y�l�������r�Ӽ~�	� P&� � v�
��S��>��u��ރMW<��a���=+73��8@����v��U'޵������?�{   �n�X��C��c$cd�-3�ݻe�@���ld�p�TR��{JN��mo�]��cuä�Lfڭ�����l-P���L��3� Pa�5<���x@Ak��7��V��l
;v(�rE�իy������{
 w!��������o��=�
  ��D�`Aܫ�{β���==&ؼY���r��yO���&'=�txX���2��C�+&IdK%�0�ii��a���v�kk�C����2� P&� ����5<���T��U`��ګ��`pP��A�ٳ,0A�`k;Pݖ-KJ��߿��~�Rޣ    w�����W�
0�ͽ���vɶ�d�ܹ�U���qEG��MN����XB�qN&����i*��C�ࠊ[��46*���ü���D� eB� c��TT�O�q�.�����	�k�񺻍�۫��))��X<�da;[ہ�e<υ�>�;��g�   �� �����Wcd$�uu�`hH����+W�
��9��.):|X�T���-y��IS�0�-��bQ^o�
�v��꒒D�k\�P���L�@2F~O��=���W��%?�eJ%�4�{:,"��j��A%~�S:Q���Ԅ����j�3���y�   �+w B�^}�+�12��
&ض��]]�ϟ�؀\��D�𰢣Ge
y]]��L?�Э[ݓDv�J�[���}�lS��Ԕ��L�S���@���cv�
��Q�SO��u���ٙ�l[;�)M04$��(�x1�q��`k;P3�m�����?��   @9�y  @�qR��y7���^7����a�qpSS���w<���;�f"w�-EY�n��bQ�]�TسG�Ȉ�'�<)7;���     �S,*ذA�֭�;;eK%�RI*��y���g�]�f��m9nr@5�<9�v�&���3M7������(   @Y������������#���߸������m�|\�̌��P�ȶ�ɶ�r����8ζ�G�̲e�ׯWq�.�k�HI���5n��6�@���@=0F~O���߯�'�P��W�1ٶ�8�{:T��i�-[��;'7=��8��X�mm�!�@Mp��i���?��k_� �Y   �r!p� �Շ��
���n�/7�]�d�Ur�!h�pׯ+:vL����V��ij�xC]3i*�مIf�J�7��}�lK���},9w (w 5�koWÞ=j|�)�mS��,of&����t�����oWz�ҫW��l�H���v��8k�>����7���,   @9�X��C�^E����x}}&ظQ�Ȉ��d�S��W�*z�m��Qy]]2w�{&IdK%�RI�}y��*l߮������J''��0�1�w (w 5��*l٢�GU�}�)X�Bލ��&��G�!�7��lC��3gX\����v�&%���0��/�   (7w B�^}ܫ�12�ȴ��`�.y+V(��(��p���Q��K33�e|��pN&�egg��w�����T��ٙ���	)Ms@�"p�2!pP<O��jx�!5>��
k��7&{Y�=��񺻍�v��S�8���bL����9�M�?����    ���   ��4���l��J/����!��T�8V��(:rD�޽���CR�H�(��n����)� ��鑿n�\)>}Z�ɓ�Ν#v    ���ѡ`�V�6��~v��ky�����/|����_(�p!�q 6�5̵�ϚةW_�{   `Q������������#���_��7*�tI�����J%�Ê��$yk�H�r<7�4��,*0F��C��-*n�.��*�JJy�Plp�2a�;�*c[ZTرC�O=��ݻUhm�W*ɖJ2�X�Eb�E��9nȅ���@sMM�;p�s}��?���,   �b!p� �Շ��##��l�]�d��?	�VՈc%g�(:vL�P��z�d�� ���q��L�[�F��A6l�mhP:5%W*�=&�*E� eB��
�BA�T<p@�(������q��x��`�x+W*9s�s�X:�da��yO`�X����u�׿���G   �;�!p�>�5�c���m��!��i�##yO��C�￯��	��f��vI��na����,<�"��fy��*)��	�Q� p�2!pP����ե�}���T���y���2Q$9����S�����6)9wNnz:�qP�<O����Ը���fݟ���   Xl� �����ט��M�`�͛��۫��%.�T73���	%�/��*�r%�(p&Me�0���T��U����CC�;:$InbB�� >�; �	�;�
㵵��g��zJ��
ZZ���dO�"*�ij2��ە^����ռ�A-�6��N�Լx۶3�{����    ��;�!p�>�5�F�n[[Ma�n��F%��<�ʸ������s�dW��mm�X>�I�R)��%��v�6�04$��MJS���l�p[� P&� *�ilTqpP�?��}��X!/eJ%΍�R��	e<O���@y#����yO`)tuM�{���w�Ey�   ,?�  ��s�J֚`�~�7���S��y��JΝ��7�!���{L^_�;�I�ˢ�R)�NU,�nܨ`˖��g�(:uJѹslv   �a�E�7mR�f�l����Jy�,�)<����k��_����T��Y+���˖%�}����Hg   ���X6�W6��	cdL08h��.%.ȕJyO�r��S:<,��]���c�4���q������vu)ؼY�;�\)9�tb��h@�c�; �	�,%�S00��}����T��U�����L�=p�lk�	�|����d���#[ہz.}���i�����=
   ���,�{�!p�#�H�Ȯ\i
{��X�����*���+:|8�;:݁;`���"��ٟ�ݷn�]�L
C�lG��; �	�;��f���x@MO<��u*44܌�9υa�E��)%�����A50F��%����%�<���?���#�Q   ���;` B�^}��1�����3�m۔^��t|<�p��qEG��]�"��!��ı܁���Q$S,���Va�66o�mn�+��y�+P/��L�,k�]����j���R�ƍ
�J2QDԎ�e����b��ӧ�4�{"T*k���pz�7�=��}���   ��;�!p�>�u�cdM�c��+�m�Q�Gu}    IDAT�d��訢Ç��Ʋ���2iz3v�c��F��^UܲE��I.�݁G� eB��\�6��ۧ�'�PÖ-
���vC�:b;;��a���g�fg���)��{ 9H׭����7�=   �?�  ��p�\�n�;Բe��xC��_��8��Pi��w?�`h�~X����X �2ׯ�Jr����f��Sq�^�k��:���)%##l   �23A ��O��
��e$�RI���]��4��o��g�U|�d�� o�H�'��v�~uv�Lm՛o�=	   �6�X6�W6�CR�{����La�6��)���yO����˗��6݁{`�D�T���ɶ�76���Qa�6�l��|��J���@�� ʄ� �44��~������'T\�^Ac����0dS;p+�7��lC��3g���N9ϓ</���%�Ԕ�~������(�Y   �<�� �:��B��6����+8s��~��J?�(��p7�$����*ر�zHf�
�z w���LJ�6���I�]�TعSnbBѩS�N�R|�2�   �3�e��[�`�y]]�I"S*�LN�=PL��l{���������{,k��@}�}>���n��?x%�Q   ���.��������?�F�n[[Ma�n��F%.H	KM���F��ޒg�;p�L�Ȇ�����kת�m�����+VHi���ubw���� ʄ� >��ޮ�m*>��zHAw�|ߗ75��T�y'`A�&ضM�����y���d���K��=	������o���?�Wy�   Tw B�^}�񉌑�5ޚ5&سG�c%�.lV+甎�d���lG�LS�>pL�Ȅ���l�y�(o�6oVî]�W���V��$7	�� ʄ��c�ut��}��xB��)��/�NO�����&��Pɇ�=��<��s� �^�g�[�>�sy�   T
?�  @���2������)r��=�dx8�p��St™�H��m���ò�Vq��G&�d�H��|_�X��n������JΟWt���3g�J���   ��3�/��G��u�֭�mhȶ��J2ccy��$7;�О������,n����?���ߟ�   @%!p  r�H��vu��_�u�8����+���{4ܭ4U����q�+8 �z5�;P&�e�Xvjj>v76�߰A�q���eE�N)���SSy�    w���{z�(X�^&nF�33y��,75���@ѡCr7n�G0&������k�i���z㍼G   *
�;  �猑1��[��߸х�����Kq��h�[�)>yR���+غ5������L�bwMMI���X���-o�Z5<򈒑�g�(:{V��h��   �g�--
֭��n���ket�V��2ׯ�=P����+����c���^c����	���q�o�ý_��d޳    ���  |��$ke��P�}�+����'���9E?���'���=$������DvzZ���6�
�:;�uu���r׮)V|���s�4�{b    �$ymm�����[�F&M�M퓓2D���scc������|A�q�'Y�� *�+����_�ڱ�g   *�;  �-g�d�L[�i����=�f���~�Qޣ�^�mt?yR^O�+>����	݁2���>=-Y+W((miQa��o��P��ΞUt����L�#   �#���uu)��a�lK�ǲa(s��-�Dґ������9�j�����=�Je��c��?������(   @�"p  �j.t���M�o���R饗�J��G�=J��5��3���D��[����ʛ�����Ţ����[��GUr��|잎��=1   �d������'S(d7熡�ؘ�\�#u#�|م�����8�j�1��v�iV �,����Y��o��y�   T2w  pG��2�	��?8�^Rx���j�|�z�
?��-[$Bw`q8'���0���/W,��v�|Pɕ+�ΞU|��˗y�   p׼�v���׭��ٙ�dʖJ2SS�ԡ��9����3g��F����w]����y�   T:w  pǜ�=Z����g���^Rt�Dޣ��˗5��.�ޮ�:�v�pEXL&�e�X����<�BA��M���퓛�Q<<���YE������=2   �
f|_�ڵ����['�l��$ٖ��	�$�{D�.%|�J���dx8�Q���e���3���?�{��y�   Tw  pW�������Wp��+=���˗�e���j��ge_~Y�p�Ν�����$��̌43#Y+W((-�oެ`�&5�����,v?{Vɕ+<�   �lk���>����֮����f�RIfl��@~\|���_Wr�R޳`1X��� pҮ��e=�Eo���(   @U p  w�#c�����/���	�^xA�ky��2H��5�����+*��+��-
���RHS��Yy���#��@i�(o�yk֨����NM):wN�ٳ�/\�ü�   �<O��5�Q�mk����"��Y� �J=���7����=����ۇ �)��M���@ߗ�<��,   @� p  ��I�1�1�ߺU�ƍ.<xP�k�ɕJy��2pׯ����
_yE�޽���Ls3�;�T��	Cy7"��rA �Ԥ`�v�8V|��s��?���՜�   PN��Y~���>y��2�Bvcl�LL��q�#(�\���
�������b0&��F,@CCj���k��=
   PM� @�8k�B�|P���.|�e�o�%�iޣ�\������*����ˬ\��`��8�╙�l�{� �{{����8���uE��+>^��07   ��Z��W���S00 �jU��q,�2SS�cw0P	���.��>���Z�y��o X ��.~���m�׾��y�   Tw  Pv�Z���?�9{����8��X(�8V���
��q�+>��lw7�;��dJ%�Н��
2��*�mwO%�����_������   �@��IAO���~�}}2R��D���$[ځ
���\x��Ç%���E��.9c�y�+����/�Y   �jD�  �1r�ȶ����^��3����JFF����'�<)���|P�ƍ�D��d~����������԰w�ҙ�,t�pA�ٳJyl:   �����]+��W^gg��q,�2ccli*Pz�r����qn �e�fq{�s �Z���?���3_�{   �Z� �E匑���n�i���r�*����k��e�k��g�^�:�V�Bw O���2�7oV�i���J�\Qt����\�(��9   `�x�V����>��%ߗ�4���T2�|��Jo���ܹ�g�b2F��$Nm����G�}�g�   �f�  `I�ݍ�u���]x���^��^�6$�/k�/�R��U��>��%�>W��
0��}f�c��MG����*��+E��K�+V2:��H   ����==
z{���ɴ��9'ǲ����$�s��9?��o(�ɔ���@��6\x��y�   T;w  ����R�`
>�`�n���·��q�5&��sϩ���*�����{�mn�{, sn��nuc���������+���Y�.d���<}   �,�'��k�����萬�I�lK��[ځj�.:rD�����u�� �(]�v��i�F��zޣ    U����D��ż� P��2������)عӕ��=ŧN�=���̨��+�}�u�mS���� *��vw)��{#x7
6mR�q�L�*��V|�b��=�tj*��  ��#��]~OO���-��Y��2SS2Q��� ~�E�+<xPnv6�q�Ȝ�I��=��V�*ŏ<���?�GN�   e��� ����Ԙ������yς;��_�ZZx�GesN�9%�î��JΟ�{"���ہd����U��>y9O��X+�2FrNJS���Y��ᇊ/^�ü�nˏ�)����{e���� �f[[��7�v�ؘ�ۈ��#��T���E�������I�5�([��</�Q Ԑt��8<pࡍ���   �� ��/}�m�/�5.4�=>�;�������)9s��>��ґ���B���<��vv��w��;$�U�Z�BAiHA��\�Ji�dtT���ٖ���	�Q1��L�Q�Lc����,h��]~�0�c�(��P� �F.y�}�*>s&�Y���<O܂���ң���o~��=
   PKܕ�_��F�w���r���,�t�F&�]|�J������G�=�]�>�,[����
v�ihXҹ �;���v�BA��7�i*%����l����/_��$�qQ���L�Q'L�(͚lK�ڵ2��12I"�ٖ�8�{L w+�\t������=�a;��.|��������=
   Pkܵ����;�y�\��s+�;���6���Q�^zInj*�p�>-p�c�ECC
��]�bI�P~�{�Y+㜌srQ�mw���,x��X2� P&�Q�PȂ��nyk��ko�<OJ�,f���nnr҅�):|Xnv6�q����;83	 w�Z��?��������{   ��n�=9��/������ffl޳���Q��7G�R��kr�R�ca��$p�g��͛Uؿ_^O�b�`�Y{3x����ǃ��_����e9�`b��@���F� ���%��[~O�����A{���~�Z�^���7�Tt�O��d�	�,c�<�ȟ�����ӼG   j��ܳS��_�υ�~��
C^S*�;j�IS��Y���%BȪ�������
��Q�}�e����}_.�G�;���;�dt�f�><�M(w (wT)������Y#��G~w�����q,{cK;A;PS\r��C���>�w�0&;�`��`q�������o?��   @-#xP����}�������C��Zc������p�W_Ut�hvA�n�9��Y�={��#��\�� ������c��sri��76��/�y�5w (wT	S(d�׬���-��s>h7q,C�Ԯ0t�ѣ
�zK�իyO�%�</;�  �,:����y�   �:�G es������;.UwԪ��=u��/+z�=.LW�{�����m�Tؿ_v��r�� *�1�9ke�w�^������-���d��J�@���B��F�]]Y̾f���v��d�D�ڣ��@sW���;���ꍵY� K ٴ�b�����{   �<(�S���/�x�a.UwԼ�c��n����=��D������߯`p��L@�2&��^(d?z^�&6M����%##�/]�6����T��; �	�;*�mn����uu�vv��}�x#f'h�KΜQt�����������K������/t����   ��ݙ�������[�w�#e��Sr�+����˗��X��}�mmU�w��]�d���"��s�,xwq�mw�t)��/_���w (w�Ķ����΂��n���匑!h�+�;�·�Rz�j��`�Y+y�x���Ҟ��e�?޿��_�{   �^<(;��oyg�����ו�, pG�1Y�����Uz�%�ccy�-n�>�
�oWa�^َ�E�����/���7=�4�sN�ؘ����tb"祝w (w,ϓ�ёmh�꒷f�LS��s2Ir3h��'��ҫW����cǤR������I��9����:��/�=   PO,��_�Rc���S������^�$�B�W^!t��R���߯`�6�G��ڛ�}?� ���Pra�����\��dtT�ŋr�R�Sc��@��c�bQ^G�|��wwK��}��f�(�I��G�甜=���a�?����r���놵r�.��E Ȥmma�Ou���|2�Y   �zÙ  ������
����ϟo�{�zF��z6�ŗ�=K��1--
v�Pa�>�e�r� @�n��r��}}HS�-���J>�h>xOFG���� P&�(�|�͘}���6c�$ɂ�8�	C��+����
T::���O�u�9�#l����y�����   �G� ����җ�6~��?�/6�=K�"p2sݣ�GUz���ɼG�+y��<O��-
�퓷vm�� � �� P�vPc~r����JFF�/_f�{�#p�2!p��og_�Z^W���.������e�(���GP!�+W����c�>�}�{�#lP\KKb}������C޳    ��3 ���ۛ��?bGG�y�R�܁�3i*�)���=p���z��={��
y��X�mw����Ƕ�KR:=�my�e�;�{� p�2!pǧ�Vފ����uv�����̶��i��=��(�ޛ��4U|���=��Op p�Q�� *ECC�<��������{   ��q� ��8��/�[������?i.Z��_~Y����Ǫi���1Ţ�m�Tؿ_��=�q Tc���F����nywN���|𞌌(��#)I��A� eB��[��fy7��5k淳�$�B��� n�]���w���҉�;��D�^S�TW(���'���_��W�   �w�) �d���o?f���	/�Y�	�;��L�Jq�ÇUz�5����G�I���3F��
vaC%O
 O�����cѻ�TF�K%W�(���}l�3�b��@���-YȾz��իe��d[Z��4I��}.fg;;�O��ӧ����>����A���8�w�O��?���;�Y    �Xb����_�������{�zA����R���B�EPс�-LK��;TػWf9���`m��=�<O��7��e_W$�8V26�tl�M�9"p�2!p���[�b~3��萷z���e���b�8�{ w���*>qB���JGG����{U3F�<��8[�nX���G�<��3�Kޣ    �p� ��;�����,���Wl��k� pf.tR���r��y�T�%p�g���>��g�;�q�'ݲ�}>zOS���]�*�v-��~#zOFG��8��k�; �	�{�]���)���V�$��c)��� (�tI��Ê�}W.���{�W)6��T�*=p�����~3�Q    �� �8�������_E�C���X���н|�.p��mkS�{���!��Ƽ�Pm�.��|���bw�>���݌�GG�\�R� ���@��W7k�\)��#���mo�bv�nne'fp�\����q�o��td����ܫ
�T2c�>��_���_}>�Q    |g ���?�g�6x��/�8�h�wo>tC�����^�+���*Us�>��l٢`�y==yO�����A�m{�q��'�wI����+W�\����%��J���
�@��Wk�Z�mf_�*����!���vǒ�p�ґ�s����{� lP���������y�   �'qF@�N��~����4i��(5���ws����u�o(z�-B�����v�*CC
v�b�;���������y�٭�/�0Tr�j����U�7>wlZ�D� P&��
���d�ڲ;;�����4���� �Ǌ�_���JΞ]�f�+���ۚ:��{�����/�9    �g ������7���$r_�@���F��_����{��Pk���mS�k���k�@�m�nL�ܺ�=M����o{�����!p�2!pϝij�6�wtd��;:dZ[etㆸ���Ɔv X,ɥK��Q|���/� p�PllPE������~[�s    �d�a PN��/����˿B�^~���0i*E���Q����_�{��V����lG���;���Vw ���,x�%zw�f��-ѻ$���ن��իJ����I$� P&�K�Zy+W�����.��]��%���F�n�$�ړ$��7;���w9�td$�9D�^Q�T�e˅ޗ_��{    ��3 *��_���^{�g������X\&M�$qѱc
_}U��D�#U�z��y��ѧ�    IDAT�M���!�z�ڼ'P����~��ݘ�M�\�~k�>=�dl,��>�_�"E���; �	���0Ţ��+�uvʶ�eQ{{�LHi*3��}n;;�� ,���%E�g������&p��d7]��Y? 5 ٴ�R���L�y�iw   T8�8 �(�闾Sx�v\�+w`i�4����Ǐ���J�^�{��RW��-��V��;eZZ�@r����s��o����ѻsN��D���g��ؘ��q������@������+W�[�Jv�*y���V�ʞ 5��}.f�� r⦧��#G�^���8C��3�v U*Y�������^��Ӝ#   � g T�3��/xo���!r/w`i݈]|�J/��tt4�*B��󬕿a���;�o��Vw ��5|w�/��	7�7iz��JJ''��}l�f�>>.W*��'Xw (�;�y�V��]�B^[���6�U�d�/�1&���2Irs+; T��9����'OJI��D�E���v Ṷ_�Qq;   PU8�"����38xp?�\�w�@>�B����Uz�%/�=R��>p��iiQ04�`�Nٕ+� n��nD�s�R�.I��������U�׮)W:5�ǟ��@���\Ⱦre��\y3d���F�$��(��s] *���Tt�X���ڵ���L�K�Z9k9��j��֍������   Յ3 *�������������+9sƕ^zIɅy����0F^__�o�"A���ͅ�l|w�fh?!|wQ�d||>xO�ǳ���5�(Z�?�; �I����緱��즭�fȞ�R���q��=I���JǊ�_ѱc�O����-�%bmvt�s �=�׭�'n   ����v������V^���;P�C��a��F���:B���L�(�&;v������`�͍�7>dm�1����w��TR:1�m}�>��Pr���$�2*�; �I��X�6�߈��U��˖�8���5��=Id☍� �N::��w=*7=��8w��}����������{��O��=   ����  >��#��8��q�ȑ�y� ���m���5�==J.\p��+~�}�ȕJ���wޑ]�\�ࠂݻeW��{4 �di��~Q��w����s[���wcd�56�����?��T���|�����1�8^�? ��Y+��2��ݶ�ʶ��[�J&n~}�5d�{j �'nvV�
�zK��H��R��!Ioﵦ��u��   @�b5$���~ڞ���O�ǎ��{�j�w�B9'�ґ�����ǫ�Q����`����CC
6o�|�MP����wy�܍�H�_��/����J&&�^��}���׮}f��w (�j��n�����Z[����5��W��iiɾ椩Lߌؓ��ߓ�CI���=��ԩ�z�c�{�i�= Ԋ���Z���}_��d޳    �{tF ���ַ�s��?��~�Þ�g�6�@���?��f�$yOUv�����V��!y��y� �b.x��)�����������I��o����SS�Ð� ʡ�wϻ�/_.�bE�/_.��"cL�ߺ�=�k*���I/_Vt옢wߕ���{�EA�^&7n8�Z�������t�+�y�   ���������}�}��w򞥚��ä��Ԕ��~[���r����L����
��l�.�Ғ�8 �4�6
�m~�6�2hm0ވ�o��=Me�_51��MN�t||��tz�0 ���X�]�,�[[���F�n��onb����f� u�MO+z�]Eǎ)�{�EG�~�ɢv�v 5���   @m�3PU��O۳/�x��uy�R-܁�2h(]t��Jo�!7Y��b	���������!�&�B!�  �܌߭�X?���:Z���<H�tb¥���]�����.��pnb¹��]29�j��* pW��߿�/[���˗���\���i��=I�� I���;��ԩ�|"�'!p�s�8C�F���ז=�غ�_��x޳    (�b �:���_<��w�z݈8\|��Jo��������/.S(�߼Y�������� �ʶ�;�y�</5֦�6u����l뻑s���<�qΥ��J''oF�nn���t��q������ڏ�7"���3MMٓ7n����g�����{�~眪��n����bSX$!��l�2f��xñ�`g�Or'y�ܞ之����:�Ƀs�b�%��g�	BHn!��[��$��ݵ��?NUwkC-����ޯ穧���:���|�Saxҧr  �p�>7mRa�&��^��8A��,lP�3�������   @ma5@U��}������;n߮�ڵ*����p9��Y��/V��K�M��z H4k���Yy���[šw+ϳ��"�y�'ɖ�:�:Jڨ���c���{O��Ax{�X���ciP�N�#��QިQ2�G�/7��-�hy� ������l`H�Ç�P�[o)z�}��8G�}</��+V� Ըpڴ�ŋ�/~��g   PY�j �Z����`�ƹ�gI2�@m0R0$����kUش�j!���&OV��K���b��f�� @u�<k=O��#���&�G������||9_�����zz�y� I�l֘�&y��F�G3z�W=��=Z��I^c��Jo���� p�lO���7���[
�y��8�B��Cx����� �vڴc�/�G�   �M� T5���u���֠����ipjO��]���m��7TذA�Pp=և"���)�=[���*X�@&�v= �c$߷2���x^Tn�����d�5F���O�g4ah��^EǎY��_���V��}���5�Q ���Lc�1٬1������Ƿ�@���T�(d�Y��&��Fy���d��d2�$OQdly
��vz&��7� *�PPa�67mRq׮�MC8	�3�� �b��noٲ��~���Q    rF ��mm�:V�����\ϒD܁��t�鱅u�_�V����X�D�=9L:�`�_���%: ����M��<�ʘr||����0��5���nz{m��km_��zz��k{{m��'���}}����ԊL��MM2٬Q6kLs��� {c�Q6k�lV^S�1�t 4Ɩ��xc��3�E�`�߀ERq� #%��ޭ�[o��u�l.�z��#�^b������DӦk������N׳    >�x �	����x�ŭ�ƍ4����;P��$E�T(�ʿ���#G\�u��d�Y�)�h��3�W�$�}k�Q��_��x^d���Zc�a��DQ���k���R.�����0|o�J���#�g����fM)�.����dLc��Y���7�������S
�{6�ʷ���0�h $ڿ_���Ra�&��n��T���lP��iӺ�/�������   ��b�@Ͱ��^��/o6l��}�@}1�Jah�[�*�f���d�pO>o��8�~���Lq= �L�A�R����qصt�1&ɫ?/�C�CY*���S��g��7×�﹜�������`|.gm>?�t �L:-�Ԧn�Y�55ɜ�uCCjoh�1F��z|_�Z���ˡuE�ܼ^�-�!�� P%�>Pq�f�zK�{��j�m���d=�U6 u+�1�H�d���?|��,    �+  j�mm�:^ziK��6��,IA��?F�;���ʯ]�b{{���	��ś8Q��/V�h��q�\� ���	>�z�5�P|����x^dJ���i�/3�Z��)*ߕ�٨tm���`|>](���|�@{<�����a�8���e��kl�J_��ֽ�k��e��NjXhZ76���q�QƟ�`�hZ��b��UؼY�͛������ZQww�� ����pp���?�p��Y    �VB ����u�^�!x��K\ϒ܁:g��������u*l� [(�����Z���q���E2�ͮ� ��8��R;����Ǥ�`�)�1�A�r0^�qX�,֡LY���!�BA6����@0>�����@`��,�WU���ˤR�!u�� ��`���3�54H٬J�������z�>�%��a]��d��� ��ӣ��o����
��!�^a�p��/y��1 ��h޼�3?��٦����   �'W Ԭ�[o]�����~�;�2ER.gmmʿ���#GF�gp��'�,�-R�p�LC��  	U�[cd��K!���r@�?_˗�O)oN�-�EX�P�[�K���
kˡ��>k��ds����^��+���
ih0~:-e2�d2R:m���L�(���� e2*�M�uj7��Zc��_�Zc����
��7�GQ�� �ӳ}}*nݪ���*vt�7�����YI IRq��wf�|s�im��   �:�����~��/�^}�[�'�	��H�	�(�ŭ[��u�����%�^c|_AK���.R�`aw ���/��cl�A>��wJ�gM�Քt����Sf���4(4�}���vx��'�rqS|.g߶�\��*o�m��m��xCCܞR&#�J�L9�2AS�RF��g2��:�6^&clx&�*�Y�;��)]�����4� ����Tܾ]ŷ�Vq�N)]�Tj2�N� N.Z�>���溞   ��� �y�w������zmr'��TJ��ZE��6�v�
�6[����
�̉����v $Z9��,_���j�� ��/=^~��Ue)D�r��V�ད���e��d�y�P�|^��s����V�|�-r9�(R����!�H���s���j�]����<OJ�=E���ϓR)c�LƗ$�N�A ���1ƤR�L��$y���1��{^X����oL:-�N�!v�7����5�
�[k��  $^���Ν*lڤp�N񦶑WSwϋ�� ��/�t[���/t=    w8o�.����N���g��ca	�8#ke�����_�6n)�� �^� �/\7�g2�'    ��E��ݻUظQ�m���p7�>�n����o> �$��7g��^�z    n�3P7v�u�㩕+�h�,�N��P)npC[ܼY�5k<X��M��v    T�bQ��v�oWq�Vٞ���j���m��i�W^���_�b��9    ��

������af�ʯ�b�n���c�d��ە��o�칟7$�^�L*%�\�-�?w�L:�z$     NV(��s��[���cM�	Uuwϋ�Y��3F�%������(    ��� ug��?��V����$�N��y�V�Z�Çm~�:6l�-���p
e�f�y�\x�Lc��     ��PP��Cŷ�Vq�6B�U�j�7� >�1*.[���g����Q    $9# uiח�Ԛz��?V>_��A� *�D����B[�򯽦�ȑ!�^�8%ϓ?}���.Rj�"��&�    ���S�ޮ���*n�*�ϻ	g!�wc�P;+a 04�����O�<���]�    YX]P�v~��z��?55r'��Ҍ�R��-ʯ[�pϞ3��8#c�_pAv_�Pf�(�    j����[���k�T,�	�(�w�� p֌����������{]�    yXeP�v~�k�������^��,Å�;��`$�Z�ZE��o���_���;Ζ7i�R*��by�ǻ    P�lo��;vġ��;�0t=* Qwϓ|?!� @�}^w�_�^��ף    H&rF ���{��{���u���z��@��H0Q$��i����):p��	��|�S�(��"ț8��8    ����TܶM�m���+E��Pa���H�'��lo �T����{s������(    ��� H��կ~�a���׳Tw #ɔZ�ý{ma�Z�m��;*�;V���
�ϗ?kVܔ    �k���*����۷+ܿ?��9�,g�r��U. 8w���������z    ��
 �l��ז4�Y��:�v=K%p���2��vw��ƍʯ[g�#��B�1٬�y���ܹ2�څ    N'���NjߺUkueD��ġv�` 篡!ҍ7�?������(    ���# �����e^|q���g�� \2R�Q�Qd�[�����
;:hRCřTJ~KKx_�@����H    �J*T��C�۶��r�'�##p7F�}Y���"lssX���{�>���g   PX���|��)��/o�w��z�J � )�����R��M�7��d4���ɟ>]���
.�P���'    ��ӣ�Ν*n٢�]R��z$$���=O����[@��Ə�篹����U�g   P=<�)�l����l�>��,狀;��8nCE�����7+�n��\��:�M��`�ȟ2%na    $Rt�۶��u���N>'�x���v 6��ɽ�%W�y䑷]�   ���R ����{S��n����,׳�� ���R�{�٩�ڵ*l�,��H��:b��̛�`�<�--2��    �����={Tܾ]�;���뉐p�{����Fx &ьG�/�h�~��z    Շ �����x����U���;��8�(�d�Ua��7l�=zt$�B=�3f(hiQp��Əw=    ��۫��#�o�&�˹	U���� �&\���Y7�<Ǵ��]�   �:x�!���Ϭ�x�S��K�@RyCd�E
;:�_�^�m�huǈ�ƎU0�����Ϛ%q�    *&:x0�o߮p߾��?p�)�N[; ��pѢ��/�4��    ��8 0Dw��f��&�\�rV�H���Y+Y+{�
mm*l��ǔcĘlV�����w���z$    �.���}�Tܾ]�-[��6T̐��ġv�� #���ju˿����G   P�<�Y���/������X���'w Iq^�A�UܲE�P��h���}�3g*�;W�ܹ�&Nt=    $R��7��ܩ���R��z$Ԡ3�ik���y��-�٬���Nף    ��� �Y���/�Q���D}}U�%� )*�!*��������ʯ[����J|g`ȼѣ�ϛ�`��--2��    ��(R�w��;v��c���]O�:pʀ;m� ���}����9wŊ{]�   �vx�s�q�=_�_|�ou���z�3!� )*�!*����N֯W�hu���<�ӧ+�?_~K��)Sh�   P��c*��7���%�˹	u渀;m� �V:m�o�O�~��?v=
   ���j ��-_��'�������)׳|� �bX7DQD�;�45)�3�?�n\�    �PP�o����
��vv�����l 8c���~s�O~�g   P{<�y���o_شr�:��w]�r:�$ňl�NluߴI6�������Ϙ�`�\s�ț4�F9    U!z�=w�R�k��{�HŢ둀8���R�� ��=�^�������,    j�
 8O;x`J�z�f��}��YN��;����-�,k�V�͛UX���98g�Ϛ���E��y2�F�	    $I6�W�{��۷+ܹSё#�G$I֘8�~��	��C���9-_~ìGy��,    j�G ��m�ߟImذ5ؼy��YND�@R8�juϿ���۷��8�7v���--��̑�d\�   �^X�p�~���*��+ܳG
C�S1c�v�;ݯ � ���ӻ{/^���G���   @m#� b[[��k֬�׭��䬯p�I��ׯW��g]��,̜�x�&O>��    �K��5h����u=p��P��_'g �H��rh�u�-��C]�g   P�� @�0����+�o�����WoHR� P�����E2Q$��H�bQ�]�TܵK9I��Q��Y
ZZ̝+3z��	   T�۫��#���+�"����ġ�ӷ�  ����>��E����z    ��J@ �w��xjժ߲Ţ��,� �"	�|[���{n�k��@�yc�����--2�G   �4���}���������d��P��}z��`����W����u=
   ��B�; �����R�W���q�    IDAT�!x����^�g  ���[�}�?�(JD,��R�~�
��K�'�d�3fė9sd2�#   iQ������q�}�^�H�*�˖�a�a� ���}^w�c-+V|��,    ��G 0�v�k_0+W>f��]�@�;��H���)���t�jP���g̐��   Ԣ��k оk�l.�z$��#[nk�l `�54D����9?���\�   �>%!g 5m�7�qU�WV�\�|� �"	�!��huG2���3����Y�&O>׏|   �Xt���={vt���!{�둀��8�><�G	��0�c��믿�Gy��,    ��~ 0����_���������ߵk��y  g�����}Y��6�Wq�w�PN��f�Ϛ%��8�>i�w    ��Ç�ޭp�nw���v=0d�M����M�ړ��߸f�#�lt=   ��F� F��?���k�wʄ�淃��9,�@v�"�(�ށ����*n٢�-q�=��7m����--�L!|    8uu)ܻ7��ڥ�\��c�� ��f��}o����=�P��Y    � ����o>x��G*9����f�� �K(�֦�瞫�7��5�����M���   ����ܩ���#g��r�4 @���^�u���_�z    (�� FX�3�|l�]w�Mvժ��X$	 �lp���q�{��
8+6�S�ޮ��]�d�iyӧx   * �ꊏ���U�{7�vT7ϋ���0 ���h���f?��-�G   �����z��;���M�^�/���[�#[
��Z)%kivGձ����L&�_p���3�O�*�Rn�   �(�����{�ā�={d�s=p^�1��� @mI�l���|��O~��(    p"� ������;�ws�������b{ ��)(mڣH6�d,����ds9w�Pqǎ�ϓ?yrz�1C���2٬�!   
����a�}��@{_�멀�F� j�ml�����'����Y    �T(� Ƕ�We֬Yi��o��?����f�� �K(�֦��s7@�Aw��1�ر��3�M��z$   ��lO��wމ�{�*�씊E�ca��߰���G
V �<D���|�ͳyd��Y    �th ����_����`��j����-S\� F����V�"�(r=PQW���.6n�$��f�Ӧɿ��--�L��   @���
��U��]�}��˨-���� �Bt�GK�^6��w��    >w H�y����������7�7�\l8Q ��Ԉf}��;j���Vq�6�m�$�tZ���-�\ ��:�   $�><�ξ{��#G\OT���@;�v �;т�f�|�<�ښw=    �	+W �0�>���W�����F���>����= 環!ʷ����\�qz��Q/��7aB��~��O�7a�
   ��ݭ�w�ۧ�wuv�
������P;1 p6�Qx�����/��    ��w H�9+V|q�����������<��  F��f�(���|�j���Tt�
6H�L&#oҤ���3d
  ���
�{O�޽�:;�߯��\O;k��y����� ��o�u�=9{Ŋ/�    �w H���?�����7�W��G����y  ��լ�v����FͲ��½{���a���ZާM��   C����w�UTnh?p@
C�c#�j�7Н«( �SQ����C�O~�]�    g�5- H�m��?/�r���}���=F�w������sI�������s��8?4����tZ����N�7uj|=q��   ����8���3~��=�ǎ�Q�
��8E ��	�pɒ[[{�W�g   �sA�; $؂�Ƕ����֦��mN¡  ������	��N�|���wI��Y��i�O�?}���Se2�S  `؄�����n�%:x0~#0Pg�0� �h���{/���>���,    p��J@�h�����^��lO��� )��!���S!��;V���-��ԩR���  �J):|Xag�����z�~�B��d�3����� �^z����?��9    �|q� �D�3�|���~����^���瓐 $�1���gwKawYށ:uu)��6n����'ާL�7q���n  @�ZE����}w ̞ϻ�pϘ8��� ��	k�����+V|��(    P	������'�g�׿��{��a�� �d�Nz[�݁X���w����>}_���q؝�w  �e������W�w�lo�뱀� � 8��94�]��f>��_��    *�` �B����"o��׼}����kG�w������sI�������s��p��;pfA �$yӦɟ2E�ԩ4�  ����Kс��w�%���5F���3aa J�ĉ}vٲO�z䑕�g   �J�� �P�~��>���=��ϛͦM3� $\���J�݁�)����w�hz/�ާN��ާL�?q��J��   y�PѡC
P�|��)�˹�H.cd	� �Q4o��Q�\�h�Cu��    *�L$ T��;����f�gL��q�$E6Du��~:�{I�&��	H<ϓ7z��I����ԩ�M�i:��   ���+:|X���q+{g����e�3�f����^�[@}3F��/ok��/�    �� P�f?���{����}���7�gE  gǘ�R:�n�h����E���.E]]*n���ih�7q���S���ԩ�&L��c   U���):x0�wv*ܿ_���|p� *&������<��}�G   ��D� j��'����޻*��+�ÇӮ� T��	w+ŭ�4�Cf���ݫp����L&3��>i��ɓ�M�(��  $L������+z�=����vw���J�� �fG�
��˿5��'~�z    n��F�{�៿���?���ڼ]�ƕ��"�D ��t"ޖ��Q�x(���\�л$����}�DyS���V��t  0�lwwd?xPQg���:$[(��j�� ��N�z,�U��{�6׳    �H � 5ƶ�z������ˍ��F�V��;�M��6�SI�������s�Ǩ~�JQD��4ߗ7~��	��{c�H&	[Q  Pml_����8�������q=P3l9��1�H�� ��͛�?{��N���9�z    )��@��y�]��W����E� P��\r	�} �$aD�}v��ih�7y��I�����	�&M��f]�  ��XTt����ST���'{�Pi֘8�N��%� ��x�UϷ<��'\�    #��7 �a�����^~�Auw���^�X7�,���I��pf�������k���f�M�4��^�75�  ��+:|XѡCq+��C�����cq â?����GA�E 5Ϧ�6���?k����}׳    �I� �ў{�Yf׮���ٙ��`�Le�C�f� QI��paQ4xw=PGL&#oܸ��}�e�& ���OQWWb?x0�]
��7�#[�=��(8B 5-?>�/_��^��#ϸ�    \��6 ԁ=��{�pÆ�A[�I�F�V��;�M��~ ��I����C�vwC�$���d���'L�o�'o�8)\� @]�G�(,��jf�==�Gꎕ�14���YQK���E�/|��}�g    �X��:�����"X��N�FA��M7)��R� FD66���8�N�Hϓ7fLx|�0A����t  T�B!�wu��Rt��l.�z:��3��N���pP{<O�UW����7�    ���: �3{����]�W�7s��/I�ŋ�p�M��38 �W62����nm|@��L&ny/7��[�Ǐ�R)�� �a8`���r�pb?z��t J�$c�l��Պ ���!�>��<��?�cף    @R$!g a;�����WW���,I��j�������a���*E� �44�;Vf�Xyc�����'�ɸ �aa��<��˗R#;�P$WK;��ZA�@͈&N싮��������Y     I��3 8����3�-[��ׯ�X��5J�;�7u*� �"	�U�vw�j�����}�Ō�\� �酡�#Guuɖ��V��.�Xt=!��0f ��W�"	 Ԅh޼����fѸ��r=    $�z P�������Uw�X4
e?�I�]��@�%a�B���E�@û�Y �3�������c�ķǌ�7j�� �ag{z� ���n��=J;P�hi�+�T5��6�t�?�����p=    $� ��}�+�Ȭ^��IJ/^���n�5���$lP��ke�H6��@����Q�d��e����)��i� �Q*:zt��}p����es9��c�vZ��w U�67�����|��?w=    $+~  IҾXX\��5ϞQ��Ϙ��;��W ��$lL��(k�(��V�vw���tz��}̘��}��ѣ�-���zD �H(}���#Gd��.5�����@�)�ii�wl�T�pڴnٲf����]�    IG� �o���gR�6�:hk[ k���wʛ:����	�:A�;P��@^��}p�;V^s��ƌ�R)6 �p���?�n����_�v�^�ҎSc' ��XI�e�m�u����֢�y    �� 8I��?�Cժ�+�7
eo�I����� p^��!�^���ox��@ݲ��de�LS��r���Q����Ms�dHO��)=*{�hܼ^jb�Ʈ"���Yc�vZ�qz�T�.[����~��g   �j�	[ �)����^��С�$�.�D�O}J���w 8'I�xpG�ݽ?��.�܇�44�����r�{�_�7N�d��k�D�}}ǵ���nE�ݲǎŁ��m�� ��v�=v$ ��3�PX��w�>���g   �j�J! ��~������f���$�de�Cf�X� �Z6�qke���]gp
��Ȍ-oԨ��}�(��F���MM2�FIA��]  ��\�FG�*:z���n٣Ge��[׻��F�����
 ���v�'^�H�h���ë��j�_�U��Y    �q� pF���R��v��Ec�i5|��
.d�$a�A��v7��5g8�Ce2��f����B�^S�LSS�XS�Lccv� �I�`�ѣ�zzd{z��z�v���>v,�
�$K�2�s`���v�Ҏ��E;��2F��/ok��/�    ��� �!���/�^zժ��=�KRz�b5�t�����I�Ƃ�;Ί�2Q$E����ܹ����!�l6�g�q��1����J_+�f��d����m)�����+���w CV
�[��>�P�l&��\��[�z��p=    T;V C����V��::�H�?u�����̘1�O �Q6�q^��?���TE��l�L6�ˁ�lv _�44�ߖ�'aw`�r9k{zd{{Oy�ʏ�������:w �c��vv�s=j_m��	vʔ^��+���G�z    ���  ����u������7�*�d�Yeo�U��9�S |�$l$��b��/�л�y |�����Nx?U�44H��J���y���닃�\����B�'�����=�~.�̖�쥶v`���=�d	-jO]tѥ�~���,    P+Xq �����I�Y�]����e�.U�dٷ 8�$l�c��[γIC��<�L&����4(���d��3�����$ ��C�6���x����@}�� {9��ñ=�D���-�ۖ��o��    j+� �s��w��pժ�:;��̜��g?+56�p�$l�cĔ�D���w�JAw�T�?�TJ&���oh�L�T������A�����8�0�*�6�|^*e��8x^(ķ�y�tm��8�^(�
���\|�P��pꇕd��oi����I±= ���ɽ����͹?�ѿ��    j� ��b|�iϳ���{�9�V��Q��n�?{6� �I�F��;�!�8E��6�L�л	�8���}��僠��^��!zϓ|?�?&<�y�mI&��`*%y��(��%Ɇ����?Tn4���E���_z\�|��
������ ��h������;P۬4���y��>�� ����K.ٞ���ߘ���=��   �Z�� @Et|����7��y�<e�/W��d�e_@R2<	�#��[��#��;*jP ��_
���Sih8�q���'�JCh"��\�k�W
�����F����
RynT'�@m����j�>�p¦�6��GZV��׳    @��| �b�}�_y埼����̛�쭷J�� �8�$���*5�Zg�aA� *��;P�hhG�����&N�+.]z����_]�    ��L @�\�����t�����[�1*�ءc�<���w9�  ���<��eS)� ����M    Α5F�������JI�O� ��-X�oԧ>5�p;    � �a����^}����j��F�����Pǒ���U�ځK%�T��2hp�ɘ�Ͳ��Q�8�02�i.Y��짟���(    PoX� �9O>���-�|�N�֣bQ}��o�{��|��  ��r8���T*ny�}Y�#b   Գ�k�}�v  �_4qb߱��v��    �i ����{���6n|�߰�Y+o�heo�M���L��4��fE���w ǡ� *�w��rC;ov8�0����Z���q=��z    �W�� FĎ����ի�7��y�<e�/W��ke�u#	Ov�Q$Y;z�w ���Ȳ�@��'����H�m�dɣ��   �{|N% `D�{��o�o���Ѵi=�"�V�RϓOJ==��  ��<O�}� �M��kϋ2    �*�[��?�WH�O� ������wn   �d`U 0�:��ݦ�u��6n�P��d���r���s�'5.	Or܁�r���R%��	'��2hp*Ș�����Pql�����7͟�x����Q׳     b�� �h�����Y���x2F�+�T�G?*�y움��'7w�CD������{��@�p�� ����0���L��� *�f26\�쑖+~��,    �㱊
 pf������ֽ���5N��)S���v�q��?5(	Ol��Y(���ZKv Ս�; Tw`h�4d���8o�ԩ=�W�y������,    ����
 pʶ�zo��o��_����1��27ܠԕW��jL��܁sc�8�^nw/��w ���i7�������3�y
/��m���/1��y��     N��V @"���W�I�Y����$�.Tç?-��쫀��'3w��hyG� � �A�(P�[�	��pl���ѣ���W�Q˓O>�z    ��c� ���{����-��6͖$o�eo�M���쯀��'2w`D�����ޑ ��2��Ycd��� �8�p֢��Å+��r���v=    ��X� $N�]w�(X��m.���Y�\�뮓���PŒ�&�8`��M��A]"� �A���;av �8�0t�-.Y�Ӗ���mף     ��s=   '���S_�喛�i�zEʭZ��'��zz8q @�1F�<)�TJ6��Yϓ5�T   �0&>&����4���Y}?>~%� @ճS���?���n   ���
-  ���&�}�jݺ+E2����r��9s�U(	O\܁��n����hp�ʠ���J��ׁZ��=�e�Qt�%[g�x�妵5�z    ��c �x����?�^y�߫�ۗ1J/Y���|D��؏U$	OX�@��?�n	��<p�� ��ja	���c{ ��U�.��9?���\�    8w�� �B�}�͵6���m�l$y'*{��&Of_T�$<Y	���JqȽv/�I/�    IDAT�]��@� *��;ɘ8�N��'�8����px�UW����jw=    ���� �*����W_���r��@�k�U�kd�e�$\��܁D�;���; Tw�d���� ��c{ �K�l�������3��    P��  8-+V�v�'>�);}�1�ʽ�����ǲ|�I  �Q�������T|	Yϓ5��  @�1&>����.��R))$ߧ�  �L�-�t�g	�   @ma P�lk���������
C�LF��~T��/g�$T��4�u�Z)�Z�]σC�; T���Fvk�i ΄c{ �1
/�dkj��+�?�p��q     ��:1 �����W��z�տ0��%)�p�n�Yjh`$L�����v��2�ۨ9��2��|Xi �N;��ñ=P�lccT���<����z    ��` P��~����7o�%ke�����g�ϙ�~H�$<!	��rȝ���A� *��;��0;�aƱ=P�¹s�3K�^;�����z    ��aU P3���ς5k��zz|��嗫����}�w@$�H��y��N�p�� �������r���% ���@���ղeO�\�⋮g    ?V� 5�o~�Q�����Ν�%ɛ0A��n�7y2�<��$<		��$+ɜ*�n�Z$w ��u��;� �ñ=Pg3?�-�̜'�X�z    ��` P�v�q��S���i
F������\{�,�>��$<��1��[ߝ!� �A��>�b�_@�plԋt�������gw�    0�<�  0���?����O�f�M;�(Rn�*{�	ٮ.N~  ��g��y��KA R*%��/�y�1   ���I</>F	�TJ
����8V  �ةS����o'�    ���i @M���ޞ7�x�[��*�I����ǔ��r���K�w �uB�h{�(��2hp�>V�1��Vv �n�5���-\~����^�ܴ�]�    p��l @]�}�=w��_�[��$s�*���H������'w UǖrQ����d9�w ���v�;�b j��@��&䢥K�9��Gw=    �-V� uc���gR;v��[�Ta(�Ԥ�?-�\���H���;��Rnz�V����"� �A�=��wh4��o�5�z���.k�}��KLkk��<     �X� ԝ�_��7��^��С�$�.T��7K��a��'w u�|����c��2��+�s�Fv �ı=PS���������?t=     9X ԥ��~����mU�~�劢�����ϟϾ&IxrpP��4�N� *��{��C���`�8�j�1
/��}��W^9�\�    HV� um�o�ֿ֮���H���)	O*� p����{�	�@ep?��`8plT9;zt!\��OZ~���z    @2�� �{��{�������Z�܁a��'w 8����VvP�ݖ� w ��`L��91��� '��*e%���?o�U�{��y     ��*;  %�_����~�tw�m�@�%�D� �����������; TF��K!vSnc/�-Xc�: ���@���aqɒ�w������    �|�� 0��o}kfj����ޚC�;PYIxp�v�����p�ʨـ�i�5���Z��=Pe�y��kɒ�g}��;\�    ��� p
;���S���s�(m�@�$��C� fp�|����1"� �P��rӺ\/]J� @u�����1�K��p�SO��z ��ٹ����N����$ے�y�dɒeK�m�1	�vf�vnJ�,P�܄I�i�;y��z�f�ܧ�3�tڛ���%�@I�L�i�df�4��$���"/1�"�����1a���H�����2����~�}? ������O�������{�[پ���������;�(���{��K���0�7ph���2\�v����a�ww?Ѽlٻg�y羬�   0��~ x?��_�<�ȯ�N��Dx�;�]y��1p�^��|����12���)��ꧯ_�{ �n9������Z���=�+Yg  `�r  o�?������kOs��/?,� ��i��+~�Mi��=�?q=�x��J��<J���;<n`��_���Y�  `tsJ  o��~������AOs��.?$� ����ݓ4}ipi�����'��$"R�u .r&�4�B�z��n��W�U�Y   �& �[t賟�\ڹ���lY����oR~@�
�!�$"ҋF��@������Ș�9�&I����V�Z=�_x&�<   �N �m:�я~2ٸ���O�""����|����?E~0�
��`.z*�K���t/4���5�i�D�Ҙ��_/�7._8 xM�4�@:mڹt͚ϵ�{�d�  ���a ��>��ɱm��Զo�K��H�����k��t�{,�J~(�
+���G�?���F����q�S�_c����!������Pl�1d()���˖m�\��dp�|�y   �F @�v��ˏ<�;������h���H&Nt������;@a���EO�y��^�c`��iOW�����Ju��  ����O�~vd��Oο�Yg  `ls �>�`����YiӦ�$�V��n]4�]�{.������
?���>�>)��^�����;�zOT�������5*B0�)�p�U�i}���1��+oH���  ���0 ���>vSy˖�G�L��(Ϛ��{_�f�rߥ���`�PX0�P鏟��'ƿ�(�H����c�W���όa��&�5%.����3��ܰ�Yg  �8F �%r����J7�?Ξ-E��+���T�)�<\�� �e �?ʿ�q�ϱ�+��{��{œ�)����������d������Ϲ�ޒ<T{ �ͭ.��VK�W��o�񍛲�  @�8� �K��g?�(y�o���Q�2%�o�1���N.zw��2�)�$""M_~��?^�����E��z�O�/����I�����Ͻ�яG��[���O�o%#�J�= Ŧ�%62oީ��E?3�����u   ��a \?�����q�'�ӧˑ$Q]�8���>��ٽ�����n�PX0�ڛ�I�O�'�O�o����P�(6.�tܸz�f͗ۿ��۲�  @�9� ����g>3��m�_U�o�4�dh��ڨ���Sy���
� �q�P�(6�-I��`���%K��y����   # �2��G>�l��[���n���twG�7F���̘������` '��b��)S��W��7<�/��   ?�0 2��������[��##IR�FmݺhZ�6R�gƨ<\�� �e �8y�� �~�P���K�~�㪫�K�g   .�0 2t�����eˆ�ѣ#"�s�ĸ�n�d�t�hƜ<\�� �e �8y�� �~��H[ۙtŊun��ͬ�   �kq 9p�������ͿgΔ�\���k�iݺHK%�jƌ<\�� �e �8y�� �~oWK���ʕ��������   ��q 9��m��L9t�[�]�:"M�4eJ4�pC���w�fL�Ål�PX0 ���j@�����I��G�.}��?���Y�  �7�0 rf�-��Jm���,=�TSDDe��h~�{#imu�fT��l�PX0 ���j@�����ӧ���bův���e�   �,� �CG?��q���v����%.$I��+���u�"M�oF�<\�� �e �8y�� �~oF��l����������   �[�0 r���>vMeǎ�KNK"�<cF4�xc���qg���Ek�PX0 ���j@����ꝝϜ_���l���Yg  ���a ����*o�|{r�t9�$��G�{�1n�{9�F.Vw��2�h�<T{ �M���"mmIW������d�Y   ��p ����}n����Uݽ{~Z�G��M��Gm��H���p���@���Pl�=�Z������ҥ���/<�u   x�F �(s��[?\ݶ��Kǎ�FD���"�o�1JW\�N���5p(,���C����{�H}֬�+V�J��~)�,   �(# `JKG}��ң�����K�$Q[�4���j���\�Åi�PX0 ���j@���iss�������o�ݬ�   @�9� �Q���n�r�з*�wwD�Ʉ	�|�Q�4M��ɕ<\�� �e �8y�� �~O�%I�,8~���g�{����   ���0 ƀC��zGi���.?�ĸ��ʼy�|㍑L��^On��b4p(,���C����{
�>k֋���i��N�Y   �Rr cD:8X:��W6o���ٳ�(���|y4�����{>���Eh�PX0 ���j@���Oss�����}�7�qS�Q   �rp c��;���{��ʻvu$i�ɓ�������O��p��@���Pl�=�Q*E���x�Zu]����   ���0 ƨ#��'���m�'�EDT::���"�6���L���3p(,���C����{
a���L}��;���_�:   \n# `KK�}�����;Ξ-E���ˣ�]V� .�<\p� �e �8y�� �~Ϙ�����,[���?��[��   Yq p���]�l��g�{ۣ^���%�֯�ڲe���>�e������` '��b����r9�00���d�{�}��d�   ��0 
��m��by��?(=:1"�|��|�Q�=['����Ef�PX0 ���j@����9#mmg��+om��?�:   �� (�#7���ɦM�&�OW"I��xq4_w]����L..w��2�h�<T{ �M�g̨���XqO�׾����   @�8� ��J��&m��畭[����V�ښ5�t�U��J:�������` '��b�����tx``�s��q�ݧ��   y�0 
���_[ڽ�����3#"JS�D���G��KO���pA��@���Pl�=�Z������{����ݬ�   @^9�  ""���>��J�>��KO?�Q���n�d�4}���Åd�PX0 ���j@����J�)燗/���>�O��   y�0 xپO��|��7�{��ܹR��Q[�<�����jUo���d�PX0 ���j@����*iSS:�t�_v\y��$����   ��� �q�������,����z$--Ѵ~}Ԗ-�4M�ޖ<\8� �e �8y�� �~��P*E�������Yp�۳�   ��� �:t��6o����Q��h��(͞�C���1p(,���C����{r������ޏw��׳�   ��� ��Ї�]�i�/'�>[�$���@4�������iy�X�
� �q�P�(6��ܪO�z��t����?�լ�   �h�0 xS�~�s�����S�Ǯ��gKI��+��n]D��S���p���@���Pl�=���W^��w�Z�����p�y   `�s �%;︣g��}ZٹsA��$��֨]}uԖ.�T��u���0p(,���C����{r#)���E���[�躙_���Y�  ���a ��~��Iv츻t���Ҵi����Dy�|��ה�����` '��b���\ig�3I�/̻瞿�:   �5# �w��/���Uٲ�ג��j���ttD�{�Ɍz�������` '��b���T}֬G�.�����Yg  ���a �������m��-o����̙r�JQ[�$���&b�x}���G�4p(,���C����{2QomNW�x��k_�%�,   0�9�  ��g>3��gϟ��n].$I��5k�i��H�e����p��@���Pl�=�W����o�0w��3��t�q   �F  w��x�ȶm_)803�4J��Q���-[i����7����` '��b��,�R)��wu���{�ٝu   (� �%3�K�tk�c�JCCS""�W\��]�y�t��Ûn�PX0 ���j@���\r#mmg�K��1��_�J�Y   ��F  ���|��)o����SO5EDT::����#�>])�<��� �e �8y�� �~�%S�:�|,[�{�>����   @�9�  .����G����[6Μ)G����hz׻"ƍ�I
 o��;@a� 4N�= Ŧ��pik�H:0��y+W�B288�u   (:� �e��y��\ڲ���ܹ$ij��ڵѴfM���n2����5p(,���C����{&��ґE���jk�qٽ�>�u   �%# �L�����Ν���s�IJ�'G���Q��4Mu�1(o��;@a� 4N�= Ŧ��%�r:��;4nѢ�ͼ��}Y�   ^�a ���;�!�o�P޷ov�i��M���룲p��2���5p(,���C����{޾R)���?���}h�=��e�q   ���0 ȅc���;~�t�XkDDyΜh~׻�4o��2F��4p(,���C����{޲4"��杪/^���_��W��   �>� @����/��l�X��gk���h��(͜���ryx�
� �q�P�(6���d�����E������u   ��q �N:8Xڶ���-7'�NU"I���M�^ɤI��(��7����` '��b��yS�S���/Y�;z�W��   �5# ��z�S�j9{��ד�[�O^x��r���k"Ə�cF�<�a� �e �8y�� �~�몷�ח,�fǊ7'���Y�   �:� @���gf�����Ҷm+��瓤V�ڊQ�ꪈZM�%��F��@���Pl�=�)7�����+��;3��t�y   ���a 0j}�]�}Wv����$7.jk�DӚ5��JzM���2p(,���C����{^�VK�-�~n��]�Gt<�8   �;�0 uv�r�ږ�������z=J'Fmݺ�-]�~�[yxc�
� �q�P�(6����H��t��wh�����g[�y   ��q �Z�n�������~i��+"M�4mZ4�_��u��Ûb�PX0 ���j@����FD��������ڰ�[Y�   �a 0�������s�o��o��(Ϟ��~w����ur$o��;@a� 4N�= Ŧ�TiGǳ�E�~���{��u   ��q ��?��]ڹ��QY� �֯��̙:O��M0p(,���C������7��H_߯w���e�   ��F  c��?�';w~��{GG4]w��{������@���Pl�}��g�z��dɿ���W~#�,   ���0 ��>���l�zG驧�"I������Ën�PX0 ���j@���P�5�Ŵ��7;x�_f�   ��F  c��|�?T�n�x<�tS$IT{{��k"�:U����b��@���Pl��V�6�\�lٝ<�٬�    �q B:8Xھ�K[�|�t�d�����ɔ):�e������` '��b��Ǡ��i�b`�K�=��Yg   ��0 (����C<�G�-[nNN��D�վ�h���H&O֍.�<��� �e �8y�� �~?��Ӧ��E����÷d�   �� @!=���O8�gσ�;nJN�.�<t_�>�I�t�K /��;@a� 4N�= Ŧߏ��S�%��   ��a Ph����#�<���ץ/�P�r9j�t�5���J������` '��b��G�tʔ��%K���k_3l   ~*�  ��ݴ���[ߓ��B9*�����7P^Dw��2�h�<T{ �M��҉/����+nN���   �� �����-G6mz��c�M����V��%�t�U���P^<w���І!    IDAT2�h�<T{ �M�E҉��/�˦����}�]/d�   F  ��tpp��ƍ���c�5ə3�V�ڊQ[�6��I�z����@���Pl��h��:R�����U�~><�u   `tq �:��ԧZ^<z�Ҏ7&�OW�����Z�U�"��u�� /��;@a� 4N�= Ŧ��X:q��ŋ��2c��g�}���    ��� �7��O}������l��3�s�U�Z-�K�D�UWE��S�	yx��
� �q�P�(6�>��I�./Z�������}�]/d�   �F  �/�w����ԩJT*Q����hiѭ^G^w��2�h�<T{ �M�ϑ�������+nN���   �#  ކ��;�G����+m���ɩS�(����M��E2e�������@���Pl�}ԧM;�,Z�м��%�,   ���0 ���'>1���?���yS�ԩ��C����d�T]�"yx1�
� �q�P�(6�>C������~���f�   �F  4@�����_��+[�ޚ<�TS$IT���i��(͜�sE>���;@a� 4N�= Ŧ�g`���L�x�o��W�Ϭ�    c�� �;|�Ϳ������㏏y�n]������+߼�;@a� 4N�= Ŧ�_&iD���Τ��������F�y   ��p p���Ї�E�޽�)921"���M�\�ٳ����M��@���Pl��%�FD}޼SI�?i���?�:   P<#  .�C������������H�(ϝMk�F���P],߬�;@a� 4N�= Ŧ�_*�R��۟���G��oC�q   ��r p���%{������3�^y�^��4M�|/��7h�PX0 ���j@����V*E}��'�}}��s�=��:   �� ����m�������Wݿn:2���ڢiݺ�,X0���y���
� �q�P�(6��Q������ឞ�ߵa÷��   �#  2r�c���o�]������pR�2%j+WFm��HK�1������@���Pl��;U��#������[��瑬�    ��� �����{�CC��w�Z��=[J&L����Q[�:�V3}-߈�;@a� 4N�= Ŧ߿M���##>6������:�u   ���a @Nl��'�O;q���Ν�%�=WIj��.YMW^��2�{[�w��2�h�<T{ �M���ɓ/��}�eƌ�ϸ���Y�   x##  r&�۲�K�k����Oע\�j__4]uU$S�������� �e �8y�� �~�&էM;�,Z�м��%�,    o�� �;|�Ϳ�����'N�D�D��;���*Jmm����!��;@a� 4N�= Ŧ߿�4"�mmgbѢ����2�<    o�� �Q��G>�b���MM�4�s�F�ڵQ��4MGE��CHw��2�h�<T{ �M�I���tu�0z{?�~�=�u   �w�a �(r�[n�8�ۥ�g��HR�1#jk�D��?Ҝw�<�3p(,���C��������ZZ���w���#6lؔu   �Fp 0
��k����Ҿ}]q�|R�4)j�WGu�҈J%�/��
� �q�P�(6�>"��u����7͝����/>�u   �Fr 0��ԧ�mHvﾦ��s�dܸ�-]�ի#Ə�U��Cw��2�h�<T{ ����>�2���������녬�    \
#  ƀ��;�C�������,?�ĸ�Z��%Q[�:�I�r�������
=�h�<T{ �����>k֋IO���=��-Yg   ��F  �1>��\=t��(M�4�Jww�V��rGG��/�����
9��D�P�(����R)������v���e   �rq 0F���_�<�ۥ���pR�5+j�VEu��H����<Ow��*� ���C����~����ឞC���Oum���    \n#  Ƹ�xo����]�V�/�PNZZ��lY�V��hj�l}0������� ���C����n�om^�౑���w�uב��    d�a @A���-G�l���k��M�~�)�բ�hQ�V��dڴK��P<�
k�` .�<T{ �mL��4"�Y�^Lzz�>wٲۓ���3   d�a @��~��w�m���[#I����ի���i�^�����i�PXcj ��<T{ �mL���\NG��N�̟����w߆��    �� �;|�-�[����,���.$�3��bE���#-���P<�
kL` r"��b�����>�`����Y�aæ��    ��  �_����۷�Sڽ����*Ʉ	Q������7�3�x���� �K�= �6*�}:e�����eƌ�ϸ���Y�   �3�  �,}����C}��o�/��k�J%�FӕWF2}�;�y(�� �5*0 9��j@���~_*�Ȝ9�����k���_�:   �h�0 ��t�[n>t�_T��##Iy��hZ�6*�ݑ��[�y(�� �5z0 ���j@��ߧ�ZZ��J���t���:   �h�0 ��u�;��RyϞ�ə3�ҴiQ[�:j�����o�O�x�V�0 �H�= Ŗ�~�N�|!���ދӧx�����    �V#  xS�v[sr��K{�|����㓦����EmժH�M{�^���i�PX�� �By�� [��}�Y/&==_��l�����p֙    F;�  �e��z�৓��鑦Qio��eQ]�0ҟ�1�P<�
+W�Q.��b�G��V�zW����_���/%�8    c��  ޶wܱ���З�{��NΜ)��L��%Q[�,���]3������1��P�(�L�}:q��Hw��������{ �,    c��  ޱ��;�G����|�t�xk��Q]�0j�WGi��$"������'��b����T��9sN%]]_m�O^��   P0#  h����*ǎ�F�o_Wr�|R�⊨.[���$)�3�f�PX� ��������--#���;����Ԃ���}]   ��s �%��ۮhy��/%{��Pz��Z2aBR�ڊQjm�$��;@a�4��S k��ߧ�Κ�b���[�Y�>2���^��_   ����  .�����|f�޽�zT����re�;:.k!5p(,w���w� d����VK���C����;���/��    �ͩd  ����������L{��X��1��b���4uj�V���%�T�Y�   �`�����,����'߾��{��:    �  \FOO�~�5��[+��y7��_�E���w��h�KOu�>=�    �e�JZ��xr����u}���6v��:    1p �K������:;����X�eK�n��n�JGGT�-�ʂ��JYG   `�H[[�G��vU���������}/�H    �w  2u��5N\sMT��:V8s7m���ϑ�Ձ��-]�ɓ��	   �hT*�Ȝ9�������t288�u$    ^��;  �0\*�zz�==�y�d�o��l��?�AT��_z�{O���   ���q��iO����ٿ�y��=6o�x衬c   �&� �;�'O���}oT��>V��s6n��o|�S�   ��$�3g�X���քi�n�q�ݧ��   �[g� @n](��{}}}}��쳱xӦh}�1Ou   �jm���Y�;�3����}{։    x� O�����h��ڸr׮���Q�Tw   �b*�����t̟����?f�   �1p `T9W��w�.�X�4�O���-[�e˖8���G��+��lYT/����   �5�I##��;Ks�������H<�H֑    h0�  F�#�'Ǒk���kb�ѣ1o��h�����w�����re��O�:&    �@�Z�����oժ���v��?����:    ���;  �^Z.Ǧ�����3Ϝ�e۶Ŕ-[�-�x�;    ������Ԋ��%K�j5�8    \&�  �)O��ķ׭�dݺX|�xt?�h����5�}��Q�:5�x    ���V�{zb��W�ޙ3��   @� �҈�1gN�3'&�tS�ؾ=�o�嬃   �
i�����qb������K��#   �!w  Ƽ��Z��ʕ+WƢ�0<�h�߻7��糎   PX�	���%�uŊ8>qb�q    �	w  
e��ٱk�������]�⊭[�z�xD�f   `�+��lgg]�<6wuE�i�    ���;  ��b��dIĒ%�v�Ll�S�n��ɓYG   sF�O�g��%K��㳎   @�� Px'ZZ�ĺu��Ţ'�{˖��{w$��e   `Ԫ�g-�+V�дiY�   `�0p ���jk�]mm����Ɗ���m�֨ER�g    ���8��GW��M���R։    e� �5��T�{}}}}�v�Ll�S�n��ɓYG   ȕ4Ibx��xf��xdɒ8S�f	   �Q��  �����8�n]�UWŒ�0�o���������   dfx��850ۖ.��[[��   �a�  oV�Ķ9sbۜ9�4<���۷G���##Y�   ���Z-^��CK�ƶ����    0� ��p�R���F����s�bٮ]1}�֨>�xD�f   �q��87wn<�til���R։    �� �:���Y�<b��s�T,޹3�l���'��   �L��ģ�̄	Y�   � � ���O��׭����?~<��m��{�Dr�\��    �P}8�xq�^�<M��u    
��  .�$�s�Ǝ�s������#Gb�c�E��g�   �eiSS���c˗Ǧ���R)�H    ��;  \b#�Rl��M��1���X�sgL߶-�'ND�i��   �"���Ů�8��[�Ϗ�r9�D    �  pY����;˗G,_3^|1�n��w��O�   �V���΍�/�����j։    �a�  �Ѹq��֬�X�&�:}�wǔ;��e   +�$.̜�,]���㹦��   ��2p �8>iR_�6b����я�w��hݹ3J�=�u4   `�I�$�gΌ��Ŷ��xr�#   ��f�  9s`ƌ8p��^���}۶hٹ3��?�u4    �F&O�3}}�cٲ82yr�q    �m1p �;0cF���H��.����;c=��=�u4    �'�龾ؽdI�:5�8    ��� �(��J���=���G��c���1k��h>t(���   \F#&��}}�wɒ�?kV�q    ��� `��P.��zz"zz�yx8�8m;wF��;   �Y�q��Ş�840��̉(���    ���;  �bg+���F�^���Ŝmۢ��Acw   �����������������r֑    ��3p �1�|���ccww4ǲ��m�Ncw   E�&����ű}��H=�   ��1p �1�\�?����5v  ��������1�xql�;7¨   �3p �1��   ���/tu�4joo�:    䆁;  ��c����Xz��Kc�C�"9w.�x   0��L��{{c���qh����    @.� @A��T�====Q��c�cѱsg�߷/J/��u<   F&O�3}}�{ɒ84uj�q     �� �)�b[{{lko��o���y���޵+&��ɩSY�  �Q#M��O�g,��K��Д)YG   �Q��  x�4"�Μ{gΌ�����я�gϞhٻ7*O=��YG  �\I�$�gΌ��Ŏŋ���֬#   ��e�  ��3fā3"��&�?�l�������SOEb�  @Q��q~��xf�����OM��u"    � �7�Д)qh������̙X�kWLٳ'�'ND��Y�  �K�����Ϗ'.���Ϗk��#   ��c�  �-'ZZ�Ě5k�����c���1s��w�`$��e   ���/tuŉ���2o^��YG   �1��  xǞ���{}}}}Q��c�cѾ{w�߿?ʧOg   ޴4I�>mZ�Y� ���ǁ�ӳ�    �b�  4�H����c[{{�M7E��~�{�F�}Q}�Ɉ4�:"   �R���΍������7~�Ғu"    (,w  ��:0cF�1#b������ѷo_Lݽ;����:   �67�َ��Qoo<��/T�YG    ��  ����0!�X�<b��x�\�������HΝ�:   c��ԩq��;/\���"J��#    �b�  d⹦�����#��#��'��ν{�e��(?�tD�f  ��.I��̙q��'�-Z��N�:    �� �̥�r�jk{��y�^s�{.��������##YG  `��77����xj��ؾ`A�ln�:    ��  �s|��8�zu���1~d$=W��������Y�   G�$���i�|GG���s�FZ*e    x�� �\{�\�M����7��'OFϞ=1y߾��8I��uD   .���)�͝���b{oo���%�H    @��  �ʑɓ��ڵk�Ƥs�b`߾��o_49�ٳY�  �RH��1#NwwǑ���5k���   �e�  �Z����""���'���}����!Ow  �<�    ���  ҈�;sf�93b��h�p!����{�D���Q~���#  �z�$F�M��;:�hool�;�S�   ��� �1�L���#��#"�����>x0&��MG�D��d�  ���9�͙�������8�ܜu$     c�  @!�<9��\�re4_�K�YĸC����sY�  (�$�3gƙ��8�`A�5+�S�   ���  �s�Z�Gzz"zz""���g�{���|�PԎ���  �#�&�َ�x��+vvvƩ���#    9f�  ޑ)S�Ț5k�D�^��'��yF�CQ}�񈑑�#  ����8?gN��ꊽ��q|Ҥ�#    ���;  �EFJ�������"֯�q.����c���1ah(�O?��Y�  ȏJ%.̚��Ϗ�]]�k֬�R)�T    �(e�  �:^�VcSggDggDD�x�������{��<�<���I�~'E��-[��6�3�2���v���ޯ�(�A�fQ��b�U̬: �`Ќ���lY2%^D�&�<�v<U�q"�<�>�,��C�whs����Ǚ�w/����  x�*���߸��w�ɏ�]K�応    �ç�   _���t�?y��$���qn}�q�?�8�$�ޘ  �x���\no���o��[�r211�I    �kJ�  ��������N��=潝�l}�I�|�i����p8�   _[}�J.��s��[�護�7;;�I    �B�  ��������v�q{;I21���lݻ��O>I{wW�  �n�2X_��[o���o����I�1�Y    �H�  ��6��pk+nm%��nf��|��O�v�^�ܿ����I]�{&  �&�t������yx�F~���A�9�U     w  ���i�����w�$3�~~kg'�w�d��O�8<L%x  ��v;õ����V]���lm�/h    
$p  ���v�������$���e���'Y�w/��y|�w  ��2��L��՜lo糛7���j�Fcܳ     �Mw  �BON���^��{I��^/�>���;��쳴R�Fc^	  �h49���zί_σ��Ώ��A;    �
�  ��y��+�~����ڧ��ʃi��&��X7  �1��J��՜]����ۂv    �!p  xE<k�����a������?���x�(��ƺ  �f�,h?y��ܿ~=wWW�=	    �!p  xE����xs3?��L�y�~{w7[��e���L��
� �U���bk+G7n��͛y877�I     /��  �5�o6�9    IDAT��V>��J���4G��up��O?���N:;;i���{&  ���������<��Ν��<���*    ���  ����F�����g�O�歇�r�~�>�,�Ǐ��p�+ ��3��Jm-�ׯ���빳���fsܳ     � p  x����������$�T��wvw���Qf<��g���vǼ  ^#U���|�[[9�����f�{    @��   o��N'?��N������$���qn޿����3�����IR�c^
  ��Q����Z�]�������ƍ�LL�{    �+C�  �s�/,���B��o'I������N�<��Çi��Ƽ  �0�����fζ���ڵ|������,    �W��  ����t�o�Nn�N�4G��<<�֣G�{�0S;;i�r�;  ��Q��zi)[[y����ܸ�'���    �Z�  ���]]����/oy��vs�ϲ������t��Ru�c^
  ����`a!����nme����Y[K���2    �ך�  �����D�ϭ[ɭ[_��?}�[��g���L����q2�q%  �r������r���������v�''�=    ��#p  ��73����O�?I25��ݬ��d���t���89IU�c^
 ��f45���z�mn����ܽvM�    P�;   /�E��mm%[[_����y�ѣ�=z��G�D�  �p�v;å�t76rz�jv67swuuܳ     �%�   ���v;?��N���<��vsco��y|<ƕ  �*F�Fꥥ\lm}�������4     ~Ew   �r:1�����yn>|��3��a�i\\�q%  �6j4R/.~~3��V>�z5�VV2h6�=    �߀�  ���OOg��w�w���l��2��������$��1. ��0j�3\ZJe%竫����G���l��=    �L�  �+�xr2�?w��\��{{�w �W�hj*å�tWVrz�jv67���r�Fc��     x	�   �6N'&򣟋�;�Q�f�ѣ�=|���ݴ?N��1.  �<fﯭ�rs3��������̌{     c$p  ��k4rwu5wWW�o;I����A�ww3������4?N��y- �k���`i)ݵ��oldc#wWWs��{     ��  ���7����F~�������e���g�ѣ�<z���a�GGn{ �::�������ի9X]������q/    � p  �/ON�x{;����3���A6��2���ɽ��Ӹ��R ��Z.,�������<Y]���F�Ύ{     �0�;   �+z�F>Z_�G��ϝ������n���r�� �Ǐ�<>N�1- �fԍF���|�������Z��ϧv+;     /��   ~���ٿu+�u����Os���,��e�� �Ǐ�><� 嫪�ff�_ZJwe%O��r���{kk�h6ǽ    �7��   ^�������$7o>w���in<|����L�sx���Q2�g( �FMMe�E�~����++�����Ng��     x�	�  �%؛��������_����\?>���^�2qp���'i��
��bt�J�KK�\[���J���`m-O��qO    ��$p  �1�7��xy9//?w��r��$�g�� �����I��ǩ��1� ��lf8?���B���9_Y���J>[^���ĸ�    ��"p  ���|���O�w�}��le�� 3����}x���IR�cZ �u����b�++�\\����쭮���r��Ƹ�    �!p  �W���d�77�����Χ��l=~�����f��0����NO�^oLk���n�2ZXHq1���./y��v{��     �'p  ���E��;�빳�������ţ��e�� ���T''i��cX ���2\ZJa!���9^]���Z�ͥv;     o0�;   ��~v�{~���$�8;���a��r��0GGi�yz��cX ����hz:ù��#����./���J�--����<     |��  �lwv6����͛ϝW�Q���e��(sO�d�ɓt���>9I��4U�7�� P�Q��zn.���tr������.-���\���'    �+G�   �������|v��!~O����le��(3GG�<:J��8���4�����k��t2��K~>�/"�ӥ�,,���\�h�{"     �V�   ��v<9����ds��k��zv�����no���yv����b �j�v;��l��9Y\����<Z\LO�     /��   x��f�/,����W��>�����i��2{z����tNO�<9I��,��HU�/8 ��zb"���ggӟ�Own.�ss9Y\�Å�<���D     �_�   /�E���++���W>��tq����,e��(�GGi�q~��ӧ�`�WP�f3�+W2�r%Ù��o`_Z���L�fg����Ӊ�q�     ��;   P�~��������$����|5e�ٳ���d��4ӧ��8=M��,���4�>M��Y��h�xQ�J��2���pv6ݹ�\���bq1�ssٟ�u�:     ���   �+�n4� ����/����YV��r�ѣ�5wxخ/.Vsy��Juy�γgM<�xԍF29��+MO�77���\����da!O��?3�~�9�     �K&p   ^?�Fffr03�76��������U/������F���Z��oח��rqq����˳g���e'Ϟ��n�!<�����pj*��t����Φ�J.��sq�J���r4=��+W�Fc�k    �	�  �7�;�����������~o�3�����w�����ŵ��r�������T..ڍ��f���%�x��F#��ff����gfҟ����l�gfr6;�'����     �!�;   �����ov���/����ѻ秧�9�ᷚ�ލ���J�����fsq1��ˉ��]]^6�^O�W�]grrTw:�zj�Wu:�É��LN6&'wF�Tw:��������������h��q�     ^ow   �d�/��$�*�}��x�wq��u�;������u���������J��N�׬��f��U�x��j4�NgTON뉉A&'/���g�N�i��ebb/���a�y����h�����_��ٸg     �<�;   �\����%�_<~%����ð�����6������F5,�۝K�;S�z�U����e��v������7|#�$U�Sgb���G癘8����t:������֏������_�     x�	�   ^�?������|��?��[9;����Ż�7��j0X�z���g�����:��lW�~3�^3�~U.��_GU%�v]w:���ú�֝N/�v/��E����9�[��F��_��{�Vk���|2L~��~�q�     �q�   �ƶ����&���|m�����|�;����ht���_�zk�3�T��T���כ�`Щ��v=6���f��F5$áP�WG�Y��L:�Q�l��f�N�3���~��\֝�eZ���9����<�;�Gu����nҘ�����      �5�   �J������_[���������7�޵�h���`u��5G���p8Q��s�h��`0Q�z4j�כ�꺑~��~�Q�uU���U��*�A��~1o�WKU%�V]�Zu>�n�h�F���j��u�5H�u�V�n6{�v�4������6:��a�qTU�Q�n�j�u���������q�5     �7��   �oT���$������x~py�T��z+Y�3�p8���ѨQ�kIR�U]���p�'�Ѩ��`:I2LV�Q����[��J��������_��U���r�hTU�����W�Q�W�����R�Z_��uU��tFIR�Z�TU]WU�v{�$i��uUՍFcX�Z�$���n�j������$I�u�h4��d�v�4I��:�Z��Q�O�����v�~�l�.������{��g���_      c!p   ���/��b���o����_�����_��u����쏭f�I?��ػ��~�ʕ;��[	�     (��    �Ak��Ivǽ      ^�q           �D�          @!�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @� �3�v,    0��z;�#         ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��         Y�A    IDAT ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��        v��I������tϮ�n7&��s�s1��v�c0���)�`�6�4���(>@���>gFZfd�Ekbq����	�cW� �1UƱ6S������'?s�v.��=����޿��|�  @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�      @'���    L��;      �	9��    �,w      �677�   ���;      �	�^���    &��      �G    0Y�      @'�R�    �d�      ��s6p   �r�      @'�R�    �d�      ]���     &��      ��    `��     ��xȱc��   ���      �q��w?6�   ��1p      :���?%�   ��1p      :c4=-�   ��1p      :#����    &��      蒧�Rrt    �a�      t�����    L��;      �)�~���    L��;      �)�w   �)e�      t��;   ��2p      :%������GFw    0~�      @�����Lt    �g�      tN)���    ���;      �E?SU��N   �)�      �E9p��3�#    /w      ��z��/E7    0^�      @W�rt     �e�      t�E+++O��    `|�     ����z/�n    `|�     �.{YUU�=   ��=      @�=z0<':   ��0p      ��e�    ���;      �u���:   ���      ]������    v��      輜�n    `��     �i���p���    v��      ��    ���      S!�|�k����    v��      ����_��    `��     ������������    쌁;      05J)�y�/��    `g�     ���s>�    ���      ��Y���?   ���      Sg4]�    ���      ���~Nt    �c�      L�+�    �w      `Z�|]�?   ���      S+����    ���      �Z��_\YY�$�   ��1p      �Y��z�>:   ��1p      ��/��gFG    pn�      ���9��    ���      ���/��    ��      3!缼���/�   �{g�      ̊=}�����    ���      3c4������;    ���     ���s~���ܑ�    ~0w      `�\���tat    ���      �5�����EG    ���     ���s��+++?�   �w3p    ��666F� 0f����������    ���    �s����� 0O>y��GG    ��     �S�y#� &���UkkkEw    �m�     ��h4r���TJ9�����   ���    pN�^�w �ً����#    0p    `677]p`��z�7�Ã�    ���    �sr��iWJ����:�   `��    pN.�0�J)��u���   �Yf�    �9����؟s~������   �Ye�    �9��}w fB)咓'O^�   0��    8��'O��  {%����p���   �Yd�    �9UUuwJi3� ��y�^����}�!    ���    ��r���QJ��ԩS�Gw    �w     ��Lt  �j8>%:   `��    �U.�0k���z׭���   ��     l�� ̜R�%�N��<�   `V�    �U� ̪juu���    ���    ���+:  ��7��[U���!    ���    ��r��Y���`put   ��3p    `KJ)�  �~�i�DG    L3w     ����}#� ��R��VVV   0��    ؒ�h��� ���z�(���   �id�    �V�� ����iGG    L#w     �$��; |�����ӣ#    ���;     [RJq� ��^�����D�    Lw     ��� �ۓ<XGG    Lw     �d4����9����Ew    Lw     �����ut �ԛ��֞   0�    ؒ3g�|#�4�� �lnn^_UՁ�   ��3p    `K���(�|=� Z����o��    �:w     �,���� �V����u���   �.3p    `;�������%�    ]e�    �v��};���]�����   �.2p    `�r�� pn����{g)%G�    t��;     [VJ1p��ya�4�EG    t��;     �a� [�����   �%�     lY��+� �!�RJ�?8:   �+�    ز�h�; l��^�}�����   �w     ��̙3�REw @��R.)��5�   ��    ز��Φ�\q�m*���i���   ��3p    `[r��  ]TJY����;    ���    �m)��yt tT/�������F�    ���;     �b� ���h��cǎ�?:   ���    خ;� ��p����J)9:   �m�    خ�  S��M�\   �6�     lK)�w �j8�4:   �M�    ؖ���Δ�(� �@�9��i���   hw     �����9�/Gw ��8��rC]׏�   hw     ������ �"O)ݴ����   �h�     l[��� ��I�~��UU�E�    D2p    `�F���; �Y�������   �H�     l�� 0���M��Zt   @w     �mcc�� &��rm�4/��    �`�    ��=z����NGw ���R޽�����   ��f�    ���KJ�O�; `�͏F�����   ���    ة/F ��{d�߿imm��!    {��    ��9��� �O�Fׯ���   ��     �H)�D7 �,(���ӧO�����[    &��    ���z��n �YQJyi]ׯ��    �4w     v��K/�RJ�dt ̊��UM��Zt   �$�    �#9�R��� 0KJ)��u���   �I1p    `�J)��n ��O)�{8>3:   `�    ر���; ���?�����   �q3p    `7� �Cz�ލǎ{ht   �8�    �c����|J�Dw ��z�ٳgo][[{`t   ���    �c�>�R�3� f�ś����رc�E�    ���;     ��G� 0�w�=�\_U�\t   �n�    �[  �����`��RJ�n   �w     v%�l� ���_   ��     �������F� @J9�W7MsYt   �N�    �+G�=UJ�bt �m���i��   ��     �Z���E7  �_.��v0k��    IDAT�4�8:   `��    ص��F7  �e_J����yVt   �v�    �k� �>��������-    [e�    �����}.�t6� �>(�|���'D�    l��;     �v���o���{t ��r�M)ݺ�����   �s1p    `,J)wD7  �����cKKKF�    �w     ��� Z��r����G����n   �7�     �E���)�� ܧ�ollܲ�����   ���    ��XXX��RʟDw  �t�h4��o|� :   �{�    06�^�� `K~������:?:   ��2p    `lJ)��n  ��y����UU�   �[�     �M���Tt �-��<~�x?:    %w     ���K/����W�; �m9t�ĉ��  �60p    `�>  l��N�8񶪪�!   ���     `�J)�E7  ;���`�#w    �     �U���� `�~e0��Rrt   0��    ����;SJ_��  v�MӬEG    ���    �I�-:  ؕW��jt   0{�    �R��; tߥ��p   �w     ��{�-�4��  v'��4�U�   ��0p    `쮼�ʯ��>� �^)�u]_�   �w     &��r[t 06����?DG    ���    ���9��  ��뚦�*:   �n�     L��ӧ?�R:� �O)�F�   �$�    0UU��9�� ���;   0I�     L҇� ��+�������   Lw     &fcc�ƔR��  &�5F�   ���    01G��rJ�� �ļ�i�߈�    ���;     �vct  09����   w     &j4��  L��;   0.�     L�E]����7�; ���#���   ���    ��C�m�o��  &��r���7�Rrt   �M�     L\)�� `������zUUޣ  �m�C    ��;}��M9绢; ��QJy����;����n   ���    �����Rʭ� ��)��t0�k}}}_t   ��     쉜�� ��;t�ԩ��:?:   �w     �ķ�����6�; �=��auu�~�!   @��    �'���ʯ��>� 콜�ύF������[   �v3p    `ϔRn�n  �<���߶�����   ���    �3����)�� �����͏�   ���    �=s���/��>� ��9���h�������   ���;     {��r}t �I���[]]}Dt   �.�     �R���ft �GG��kkk��   ���    �=u�ȑ���>� ��E���c+++��   ���    ��G  �PJ����}r8>%�   �g�    ����z�K)���  Z��9�ۚ�yZt   ��    �=w�e�}#�t[t �*+�||8>#:   �c�    @�� ��y`��#+++ώ   b�    bcc��)���; ��y@�׻��럍   ���;     !��⊿I)}(� h�AJ�4M��   `o�    ��r]t �Z�K)����   ���;     aΜ9��W�; ������>   �w     �TU��RzOt �j9���4�R)%G�    �e�    @�R��D7  �WJ9�4�۫���n   &��    �P���_H)}.� 脗�߫����   `2�    h�� ��x�`0�qyyy>:   ?w     RޕR�'� �����[�����C   ��2p     �����RJ7Gw  ������}ee���!   ���    �
���E7  �sq�������c�C   ��0p    �Μ9scJ�/�; �����h���pxqt   �{�     �BUU)��Gw  ����Ǜ�yVt   �;�     �����[RJ�� @'=��rK]�Ϗ   v��    �ָ�+N��n��  :�`J�MӼ$:   �w     Z%���� ����R�3_   l��;     �r�ԩ���2� �~�y���#�!   ���    �*UUm�7� 輜RZn�f����c   ��1p    �u677ߒREw  �WJ9�4�o?~��   ���;     �s�ȑ/�Rn��  ��+N�8qCUU�C   ��f�    @+���  L����~Ht   p��    h��/�����; ���R�'���.�   ~0w     Z)�\J)o��  �K���sss��G�    ���    ���FoK)���  ����9|ee�'�C   ��f�    @k=z�T)�]� �TzP���h]��$:   �w     Z-����R��  ��y)��6M�C   �o3p    ���8���� `j�K)on�f):   0p    �J)�F7  ӭ�rt8�������   �e�     �����SJ� L���N�8�����E�   ��2p    ��r�%���� �Lx�������   ���    �N8}��;RJ� L���Omnnޱ�����   �5�     tBUUw�R֣; ����~�G]�O�  �Yb�    @�K)� ̌G��>������   ��     t�����RJ��  fʃ���-����C   `�    �)��ՔR��  fG)�@������-   0��    ����/�?� ̜~�y���+�C   `��    �9��h9� �I9����i�ZU�\t   L#w     :gqq����g�; ��TJ�����﫪�@t   Lw     :����  ̮Rʋ��ǆ��â[   `��    �IL)}!� �i?�s�l�4��  �ia�    @'�K�y9� �y�)�|�i�gE�   �40p    ����G�'���� �̻��rK�4/�  ��3p    ��:��s^��  H),���i�WE�   @��    �i�������W�;  RJ�Rʛ�������c   ���    �Ç+�� �J)���y������   �w     :o4�VJ�k�  ��O�:��cǎ�?:   ���    ��[\\<�Rj�;  ��O�={�����GF�   @W�    0J)oL�� ���~��_�����!   ��     LW��{D���u]?7:   ���    ���; �bJ)�2�it   ���;     S�w ����9�{8�  ��2p    `��� �\�9/5MsmUU��  �{�X    `�,..�)���  ���rx0�����[   �M�    �FoJ)}5: �^2??��W_}At   ���;     Sgqq�LJ��� �s)�<{����4��[   ��    �J�O�^O)�Yt ��H)�3u]?':   ��    0���:�Rzmt �]�R��p8<   ��    �Z^x�J)�qt ���s~o]�G�C    ��;     S�СC�)���;  �!��������*o�   ��     L�����O)�At �v�R��Ͽ����-   ���    ��� �SJ���`p�p8|Xt   �w     �����GSJ�Gw  ��3r����{�����<���Tw��B% ���"�����^���"Xd!�lS��݆��H��:�s:)�ڄx�!�
F.I 	$���d���2��*�m�ꮳ�p$�tWwW�>���/x���k}�~�p8|T�   �	�     ̄�hԍ�Q� ����h�����'�  ��f�    �Lؿ��RJו�  8Kj�Z��  ��d�    ��h�Z����Kw  ���RJ���t   lw     f����G#�5�;  �AJ)]�4�k���+   [��    ���n�2"��t ���9�laa��UU=�t   l%w     f����?����  8W9�����+�8�t   lw     fή]����?/� ����ɓ�o��KJ�   �V0p    `��۷��xU� �-�Ȝ��u]c�   8W�     ̤n�{]D|�t �yPD�s0,�  �sa�    �LJ)��DD.� �E�R�n0T�C   �l�    0����sοT� `����u]_]U�\�   8S�     ̴v�}0"���  �b/]XXx����B�   8�     ̴N��)���  [-���v�}�p8|x�   �,w     f^J������  ���F�9r�1�C   `3�    �y�N�Μ��  ��666�?��t   ���;     DD�߿>"n)� �M>'��Φi^P:   N��     >e4-EĨt �6ٝs���`�C   ��    ���߿�wr�W��  �F)�t���k�=��t   �G�     �i���e9�/� ��^���������  �Og�     ����|<"^U� `<e}}���i.(   ���     ���Ǐ_,� ��"�|�����K�   @��;     |���F��(� �>��j�2�^:   �    �^�z�ߎ�kJw  쐅�h����e�C   �m�     pZ�֏F�?��  �!s)������9��1   �&w     ��N����  ;(��.o���G��U:  ��c�     �p�ر�E��;  v����ޱ�����!   �w     8���F�V�"�D� �������>|xo�   f��;     �F���p����  |����+++_U:  ��`�     �p����#��Kw  �V����i�Q:  ��g�     �PUտF�+Jw  2�s~[]�//  �t3p    �M��z7��R� �������i��9��1   L'w     8sss?�\� ����i�TU��J�   0}�    �,--�uD�X� �¾g~~�7�9�٥C   �.�     p�������?Kw  �-�>|xo�   ���;     ����ōV��҈X/� P�c���>X��J�   0�    �,t:�G���  c��ަi�Q:  ��g�     g�رc����/� 0�sο�4�+J�   0��    �,UU��s~IDl�n ��k�����*{   Ί�     �A���`J��  �"�oϞ=�����n  `��    �9Z[[�ш���  �"����ht�����n  `��    �9���_s�/��\� `�|�������ˏ.  ��0p    �-���o���/� 0f�j�n_W:  ��`�     [��ɓ?Q� `���>/�t�`0��t   ���     �����%����  c輔ҵ���*  �x3p    �-����o(� 0�RJ�򺮯��j�t   ���     ��ɓ'/���[� `L�t~~������C   ?�     ��<�/�ȥ[  ������m��ˏ(  �x1p    �m�����/� 0��n��h��+K�   0>�    `��޽{)����  c��9�[����K�   0�    `��۷���ȥ[  ���h4z[]��  �<w     �F�n�Ɯ�kKw  ����Ʀi�[�   �2p    ��׍�?. 0�R��'�~�ѣGw��  �w     �f�~�x���#b�t ������>�Y�C   �y�     �����9�å;  &ē������ὥC   �Y�     �C�?^E�o��  ���������'�  `��    ����d��~aD�Y� `B<,"��4�3K�   �3�    `---�aD��t �ٓs~k]�?T:  ��g�     ;�رcWF�M�;  &H;"�j��ʪ�l   ���     vXUU��'O�("��t �$�9�������n  `{�    @�XJ饥;  &�����o^]]���!   l=w     (���%"�P� `}�����M�|I�   ���;     �s~eD�q� �	�Ȝ��~b�   ���;     ����G��#b�t �zpD�g0\T:  ��a�     ��z�ߎ�/� 0��K)];��!   �;w     ǎ;7��  �P)�ty�4���j�t   g��     �@UU����F�?�n �T9���Ͽ}yyy�t   g��     �ā�""^^� `�=��n߸�����!   �9w     #�^��9�)� 0Ὰ�j�~�ȑǔ  ���    ��9��RJ�S� `�}��������7�  `��    `��۷����"��[  &��F�w��  `s�    `u:���_V� `
��R���`P�  ���    `L����s�GKw  L��R���뫫��+  �}3p    �1v���K#�wKw  L��.,,�����  ���    ����V���(� 0r��9??�`0xH�   >��;     ��N����Jw  L��I)ݾ�����!   ܓ�;     L�~�}J���  S�����~b�   ���;     L����}�;  �ȃ"�݃�`�t   �d�     ����F���"��[  ���RJ��W�  ��     &�����$���;  �L;��SM�\YU�-  @A�2     �0�n�M)�kJw  L���={�\?�_�  `V�    �Z[[{eD|�t ��I)=g4�X���n  �E�     0����k4-F�Z� �)�u9�[꺾�t  ��1p    �	���?�9�@� �i�RzLD�Q��J�   �w     �`�~���xm� �)�Ј�y8>�t  ��0p    �	����ʈ��t ��Z�Fo����C   f��;     L�K.��D��^���*� 0���3M�\�sN�c   ���;     L�����N)}OD��n �V9�}u]���ѣ�J�   L+w     ��n�9��;  �YJ�����n8|��g�n  �F�     0E�����  S��sss�5MsA�  �ic�     S��j�PJ�wJw  L�/�9߱�����!   ���     �L�ӹ3�����[  ���Z�[�~Z�  �ia�     S������x~Dl�n �r�kMӼ�t  �40p    �)����U� ��;�����*  0��    `�u��W��R� `����u]_SU�\�  �Ie�     S,��G�ы"�J�  ̈/,,�cyyy�t  �$2p    �)w�������O�n �9秶������K�   Lw     ������ED.� 0#���ɓ��u���C   &��;     ̈~����X.� 0C�0"޿����!   ���     fȱc�^�s���  3�A�V�݃���!   ���     fHUU�'N� "��t �9/��Ku]�H�  �qg�     3��.��V����-  3�W�u=���^  �>8�     `u:��o�Zϋ���-  3fi~~�W���_�  �qd�     3����fJ�`� ������7>|��J�   �w     �a�n�N)]]� `}���������t  �81p    �7??�����Jw  ̠����+  0.�    `�]r�%'N�8����-  3��SJ���K�   �w      .����O�n �A����h��    IDATC   J3p     ""����AD\�[  f�y)�k��yE�  ���    ��������t ��j�_�4͕9�T:  �w     �z����5�;  fU�y_�4o<z���-   ;��     �kkk����Kw  ̰����nX]]}`�  ��d�     |����{vJ�c�[  fؓ���o�/  �S�    �{u饗�����wF���-  3�q�������G�  �	�     �}ڿ��r�GĨt ���v������o(  ���    �S�������  �qj���j�晥C   ���;     pZ�n��)�kKw  ̲��rο:^R�  `��     ��Rʻv�zqD�R� `�ͥ������J�   lw     `S���ww��zvD�Q� ��"��������J�   l%w     `�:���s��[� �x�������K�   lw     �����?o�Zό��[  f]��;G��M�zp�  ��`�     ��N��RJE�F�  �kw�������G�  8W�     �Y�v�o��~�  ""��v�����G�  8�     �Y��zGRJ��;  �����������!   g��     8'kkkK)�_-� @DD<(����i�Q:  �l�     礪�QJ�{#��-  DDĞ�����KJ�   �)w     ��u:�;#�Y��-  DD�\J���`P�  8�     ����z��n��#"��t  �RJ�7MseUU6"  �Dp�      [fii�#�"���-  |R�y����/TU��t  ���     [���ݒs���ȥ[  ��������oX]]}`�  �S1p     �\�߿.�ty�  ���}��7���  �/�     ���v��="~�t  �.���SJ���G�n  �7�     ��YXXؗRzW�  ��F��-+++�/  ��     ��K.9����숸�t  ��V�u����SK�   |:w     `[UU��9�?)� �=̷Z�_�����C   ���;     ������土]� �{8/"�k���!   �     �����j���T� �{h��i�åC   �    ���t>�j��w�n ��r��������I  �b$     ���t:��9_�[  ����+~��ѣ�J�   ���     �q�~�m)�W��  �3土����W]u�|�  `��     Et�ݣ��;  �W�z�w�x�С�  f��;     PL�׻<����  ܫ�ٽ{�-��ˏ(  �w     ��.��Ҝ�[Jw  p����n��4͗�  f��;     P��������_��n �^}A����i�S�  `��     �UUu��ݻ�*� ��:?�|K]�O)  L7w     `,�۷��-� �����_�����C  ��e�     ���U��zJD�]�  ��yq�`0xY�  `:�     c���|$"��J�  p��)�����*  Lw     `��z�ߊ�ň8Q� �{�RJ��A�9��  ���;     0�z��qQDl�n �ޥ�zMӼ��ѣ�J�   ���     [�^�D�K""�n �>]������px��!  ��3p     �Z��{c����  �ҳF��o���>�t  0��    �����W#�'Kw  pJ߸��~�����  &��;     0z���9Kw  pJOX__�eyy��C  ��d�     L�^��K)]S� �S��v�}�����  &��;     01RJ��.�$"~�t  �ta�պ�i��,  Lw     `�,..n;v�qC�  N����{�����!  ��0p     &NUU�ǎ{nJ���-  ��g�ߵ�����!  �d0p     &RUU�z�ĉg��~�t  ����j�z]��-  �?w     `b<x�_v�������n ��vG�uMӼ�t  0��    ���o߾��FO����n ���9��5M�)  �/w     `�8p�/Z��S"�oJ�  pJ)��4Ms�t  0��    ����t>�j��/� ����u����lW  �{p$      S���|8����8V� ��zŞ={�XU�\�  `|�     S���0��숸�t  ��Rz��={�[]]=�t  0�    �������w�n ��RJ�Y__�ayyy�t  P��;     0�z��;#⢈8Q� ����v�}�C�\:  (��     �Z�^�)��#b�t  ��ջw��+�8�t  P��;     0պ��r��#w �I�'O���i�J�   e�     S���_�RziD�J�  pZ_�s�u8>�t  ���    ����v��DD.� ��]8�n_^:  �Y�     ����z�����  l�CSJ7���<�t  �s�    ������L)uKw  �)i�Z7��+  �w     `�t��a���Kw  �)��Rzw�4O.  l?w     `&���*"��  `S�Dį�ç�  ���;     0�z�ޫRJ˥;  8���F��ۚ�yN�  `��     3����hD\U� �Mٝs~S]�/,  lw     `���r�������-  lJ;"~��뗖  ���;     0�>5r���x]�  6����z�t  ���     �#��{��<�tm�  6%Eİi��K�   [��     �S7���^�s~K�  6'�\�u���  ��0p     �4UU������\� �M���뫪��� �	�Q     �,..n�ݻ��0r �$?4??��믿�]:  8{�      ��� `"]���}��=��t  pv�     ���������s�o)� ��]t�ر7UU��t  p��     N�K.9q�>/�� 01r�Ϟ��kUU�+�  �w     ��X\\�ػw��a� 0I�m~~�������C  ��3p     �#w ������������!  ���     l��; ��I)}�]w������[  ��3p     8F�  �'������VWWX�  85w     �3d� 0yr�߰��~�p8|P�  ��     �#w ����:���!  ��3p     8K�6rO)][� ���9��ݻ�S���n  >��;     �9X\\ܸ����� `�<>�|ˑ#GV:  �'w     �sd� 0yRJ���ظiyy��K�   ���     `� L�/m��7�Ç�  >��     `�,..n����0"�T� �M{�h4�yyy��C   w     �-UU�ɽ{�~oD��t  ����v��#G�|Q�  �u�      [lqqq���("~�t  �v�h4�yee呥C  `��     l��R�v�����*� �����Z��WVV��t  �*w     �m������(� ��]�j�n��-  ���     `}j�+�[  ش�G��{����!  0k�     v@��;�s>X� �M{hD��'w  �Y�      ;���/� L���F���� `��     �~����  l�CF�эu]Y�  ��      ;���5��K�  �)�G�MF�  ���     
��z?�s�$"F�[  ؔ�#�#G�<�t  L3w     �B����9�#�d�  6����#w  �F�      ���k�� &�C766�5U:  ���;     @a�~�����#�D�  6����敕�G� �ic�     0���䜟w�n `S�j��� `��     ��~�����s�� `R\�n�o_X:  ���;     �����h�ZO����-  �^�yoJ�}G����-  0�     �L��y_D<9">^� �M�`4�l�  ���     `�z��J)}k���K�  pz9罣����`���[  `��     ��n���)�o���,� �����Z��� ��3p     c�^����'Fğ�n ��r�{SJ79r�J�  �$2p     sKKKm��O���/� ��\����^#w  8s�      `ii�����W� �M�pcc������C  `��     L�K/��o���7E��[  ؔG�F���9��!  0)�     &����?真7�n `S�xcc㝇zp�  ��      ���߽{�����V� �M��ݻw�g8>�t  �;w     �	�o߾����#�ͥ[  ؔǏF�w,///� �qf�     0���Z߻w�E���-  l������p�UW͗ �qe�     0�7���KRJ��[  8���7�y睿ZU��J�  �82p     �p)���t.�9ץ[  ؔo�������y�C  `��     L��R��������-  l��N�8��UU͕ �qb�     0E���rJ��t  ��s~��={^_U�  |��1     ���v�ÈxaD�,� ����^0??��;  |��1     ���z��s~nD�U� �������+KG  �80p     �R�~�m)�gD�Z�  N-��ʦi���  ���     �X�۽9"��P� �S�9_Z�����  ���     �\�����������-  �֏�u}Y�  (��     `�z�?h��O����n �^=��#  �w     �������h������-  �ZJi�i�,�  ;��     `��߿�oZ�ַD�K�  pJ)����i��t  �$w     ���t>�s~rJ�]�[  8�V��皦���!  �S�     fP��?������xs�  N��s���p���!  ��     fTUU�{��(�tM�  Niw��-u]?�t  l7w     �������t^�s�K�  p�r�������<�t  l'w     ��R��~��s>X����w�_�_u�ǿ��NubW	�L�f��:��B!�$�@� �bA��P�u��Wݝ5��'��ΩN"QCX�ED.��%
�B�$0r]�Iw���@����RU�\^�������� �Nݭ�j�����D�  �(�      DDD]׋)�GĠt  w�^9�w-..�Z:  6��;      ��v���s~vD)� �z@��~ϥ�^z��!  ���     �����M)=%"�n ������;�����!  ���     ��n�����#���-  ܡ�:t菚�9�t  �w      nW]��j�Ί�/�n ��===���i�� ��`�     ��t:��n�ψ�,� �z����5M�� 0��      ܩ����mٲ�̔�GK�  p��=33sE�  8Q�      ܥ�;w~��O>+����-  ܾ��Kz���Kw  ��0p     ��رc����O���J�  p�����N�  8^�      ��io߾����ե[  �}9�^�����  p<�     8&���ku]�(缻t  �+�_����Z:  ���;      ǥ��Ŝ�K#bP� ��h眯ݷo�y�C  �X�     p��~eD<'"��n �6�Z��u�~���C  �h�     pB�������q�t  ��Ã������{P�  8�      ��n���"�1��-  �ZJ鞭V�]�_~���n ��b�     ������������-  �Ə9r�W]u�t�  �3�      ���������>*">Y� �[K)=�СCok�f�t  �w      ���ݻoh�Z�GćJ�  p�����&�J�  ��1p     `�u:���ύ�w�n �6~yyy���  ��c�     ���������'F�5�[  ���󞥥���;  ��     �a��Y�v���9�-� ������~��Jw  ��3p     `C��r]�MD쌈A�  �M+���^�wn�  �w      6EUUWD�s"�p�  n1o޷o�ϕ �w      6QUU��s>?"�U� �[�p��z�����C�  0p     `S�u���8;"�R� �[�����ޥ��{� `��     �骪�H����-  ��)�?^ZZ�V: ��e�     @u]v˖-g��>Z� �[�BJ�MM�l) �d2p     ���;w~��O>+����[  ��۶m{]�9� `��     PԎ;Vn��'E��n �_���������  `��     P\�4�WVV��R��t  �*���^����  Lw      �B�4�n�;;#bP� ���xe��b�  &��;      C���+RJGđ�-  D;���}���\�  &��;      C���1����8X� ��i�Z�����+ ��3p     `(�u��V�uN����[  �Ss�o�ꪫ�K�  0��     Z�N��[�lyDD|�t  �s�:�4͖�!  �/w      �����g>|ZD|�t  q����  `|�     0�.��s��F�;K�  L���z��|�  Ɠ�;      #��뛶o�����kJ�  �^����  �w      F����Z��ya�yo� �	׊�7���G� `��     0RRJ���&����X-� 0�No߷oߏ� `|�     0����5)�����]� `R���R���.��GJ�  0�     Y�n������WK�  L���Onٲ�M�L�n `��     0���˜�i�O�[  &UJ����W��  `��     0�>=�H)}�t �{n�׻�t  ���     ������O>���xW� �	���~�Y�#  ]�      ��;v����<1����-  *�_���]: ��d�     �Xi�f��� 缷t ����9_����t  ���     ���R�u]71��9  ��9��߿��C  -�      ����~;"��J�  L����h�fK�  F��;      c������F��K�  L�sgff�JG  0:�     {�j��*� 0ir�;{�ޯ��  `4�     0:��?�3s�]� `�ryy���  ?w      &���"�#��S  &�I���-���@�  ���;      ��뛶o�~a��wK�  L�{�������Ҷ�!  /w      &����Z]�/���1(� 0A�j���4��  �ˡ     �Ī�ꊔ�3"�;�[  &E�����ӯ(� �p2p     `�u���r�D�7K�  L��---=�t  ���     ��W���[��#SJ7�n �)�tM�����!  w      ��N������E�ߔn ��D��O- ��0p     ��ڵk�?�r�)gFĻJ�  L�S�������ʭ�C  �      �}v�ر����Ĕ�kJ�  L��n���W��  `8�     �h�f���0缷t �$H)=���wJw  P��;      ܎�R���9�jD)� 0�r�K�~����  �,w      �u]�.".��o�n s������?]: �r�     �.TU�ވ8;"�T� `����^v�e?R: �2�     �(TU��v�}Z���[  �܃N:�h� `��     �Q��������#s�(� 0�ι�^^: ��g�      �`Ϟ=�غu�c#�J�  ���---=�t  ���      �������n��s����    IDAT{K�  ���R�fyy���C  �<�      pRJ���&"^��s  �����.--m+ ��0p     �PU���9?-����-  c�gRJ�) ��0p     �T����_)� 0�.��z/- ��3p     �u��t>�n�O��,� 0�����;�t  ��      �����g>|zD|�t �:��jX\\<�t  ��      ��%�\r���ʹq�t ��w��~s�4S�C  ��      �Κ�����۟�Rze� �1t����b�  6��;      l���ٵn��҈���=  �$缳��?�t  ���      6PUUW��f#�;�[  �I��U�~���;  X_�      �����[r�gG��J�  ��Sr�oڿ��K�  �~�     `�u��v�}fD\_� `�<hmm������ ;      �$���o�ۧE�ߔn #O����S: ��a�      �h~~��9�3"��[  �E��7z����;  8q�      ��꺾iee��9�K�  ��VD����ݿt  '��      
h�f���E�Έ�� ���뚦�* ��3p     �����"�4�J�  ������Y, ��3p     �º��[rΏ�9�t ���9��^����  w      u](�|ZD�c� ��"����@�  ���;      ����O>|���`� �w����7]y�[K�  pl�     `�\r�%7����o*� 0�RJ;|��R�  ���;      ��i���v/�9�-� 0�^������  =w      B)�\�u;#b�p ��J)�jqq���;  8:�      0Ī��"��K)�o�n Q3�v���9�t  w��      �\]�oM)=:"�\� `D=tzzz_�  ;      ��N����i��-  #�%�^���  �9w      u]�ȑ#��?P� `������ݿt  w��      FȞ={��u��Ǧ��-� 0�~$���K�  p��     `�������t��s�[� `������?��Jw  p��     `��r]�MJ�yq�t �(�9�|ii���  ܖ�;      ��n�{MD\�*� 0BZ)����z?Z: �[3p     �WU�{[�֣"��[  F�}rί�9��!  �w      �N�c�������/� 0*RJ����/)� ��1p     �1�{�����N��w�n !K�~�!�#  �W�      0Fv��upee����-  #bk������SJ�  `�      c�i�ժ�^�s��t ����`pY�  �     `l�u�ύ�å[  F������#  &��;      ����^�s>?"��t ��K)�k.���+ 0��     `��u��V������t ��������rΩt ��2p     �	��t���n�)� 0��_^^���  ���      &����s�gE�;J�  ��^��KG  L"w      � u]ߴ}��#�wJ�  �����~�i���-  ���      &����ZUU;"bgDJ�  ������iJw  Lw      �PUU]�R���C�[  �Q�yW��;�t �$1p     �	��v�27�n B��x���Ҷ�!  ���      &�����G�'K�  �F�R� �Ia�      ���§[����g�[  �MJ�E�~��;  &��;      �N��SSS祔�-� 0dR��5�����t ��3p      n177ws��yV�yo� �!s�`0xM� �qg�      �JJ)�uݤ��GJ�  ��,--=�t �83p      nW�۽&�����f� �a�R��~���  ���      �Cu]���j��/� 0$�>^U: `\�      w���|��n?<��ץ[  �AJ���~�WJw  �#w      �.���1"~1"�^8 `(�/����+� 0n�     ��R��M۷oJD�v� �!p��`��  ���      8j���kUU�E�ΈX+� PRJ��^���  ���      8fUU]OK)}�t @aW,..޷t ��0p      �KUUo���#��[  
�[��~U� �qa�      �n��w�V��[  
����]\: `�      '�����v����J�  t����}KG  �:w      �������֭[וn (�n�v�wJG  �:w      `]������v�K�[  
yB��z� �Qf�      ���R��j!"vFĠt �f�9���+��g� �Qe�      ��������G�wJ�  l�=|��m  ���;      �!��zs�����f� �Mv�}��+ 0��     �S���[����-  ���j������.� 0j�     ���t>�n�ψ�O�n �D�������t ��1p      6�����Z��##⃥[  6KJi����i�;  F��;      �):��ק��Ή�7�n �$����W_}�I�C  F��;      �i���n޾}�3"�ե[  6�Ϭ��,��  �      �����]���9���K�  l����\� `�      E�u�ύ�#�[  6��-[�\Y: `�      �TU���� "�n �H9�󖖖�Q� `��      EUU�ވxLD|�t �FJ)�߿��Kw  3w      �������n��*� ������#  ���;      0���?�e˖3"�#�[  6Я///�B� �ae�      ��;w~9�|VJ�=�[  6Hk0��i�-�C  ���;      0T꺾����O���J�  l��ݶm�KJG  #w      `�4Msx�����^[� `#��~cqq�;  ���;      0�fgg�:��r�{K�  l��v��/ 0l�     ���R�u]7�3"r� ��6���[: `��      C���+"��X-� ��r������Jw  w      `$TU����S#�P� ���R�ɃΕ�  �      ���v�oo�Z�GķJ�  ��W,//ߧt �00p      FJ���@D�_)� �Nf��b� �a`�      ����>�n�O��O�n X'�����#  J3p      F����g�����-  �!��ʫ�����  %�      #k~~��G�9+">T� `����_\: �$w      `��ٳ���r�y��-  �`���ҽJG  �b�      ��;v����\J�  ���E�o��  (��      M�޾}�3s�W�n 8)��/--�l� ��     ��1;;�V���rλK�  ��vJ���  %�      c���ň���A� ����^�wa� ��f�      ����~;�tqD)� p��W^y���  ���      [�n��)��E�ͥ[  ���9���  ���      k�n��9��E���-  �*���}��ݻt �f1p      �^]��;"�,� p�fRJM� ��b�      L���>�j�Ή�K�  ���󗖖~�t �f0p      &F����v�}FD�s� �c�N)�+ ��     ��2??���"⳥[  ��c{�޹�#  6��;      0q������/FħJ�  ���il� ����      &��ݻogF��J�  �����<�t �F2p      &����9rVD|�t ���9_�4���  �(�      �D۳g�7VWWϋ��S� �(�gzz�%�#  6��;      0�v���͜�y���-  Gaϥ�^z��  ��       "꺾ijj�	��-  w��[�n�o�#  6��;      �w���ݼ���􈸮t ���9�xyy���;  ֛�;      ��i������/�9�^� �;1�s�[: `��      ����ٵ��~%"�(� pGr�����)� ���      nGJ)WU�3���K�  ܁VDx� +�       w����w��  �=9�'---�V� `��      ܅��SJ/��\� ���~�t �z1p      8
�n���xQDJ�  ��3���cJG  �w      ��TUիs�ώ���-  �/�|Y�9��  8Q�       Ǡ��k#⢈8R� ���|��{b� �e�      p���zsJ��N� ��I)�f�46a �Hs�       �n��')����; 0<�����E�#  N��;      �q�v�2��J�  |�+���R: �x�      ������D��"b�t @D<hzz��#  ���;      �	����"���8X�  "^q���v� ��a�      �����`08?"�U� �x����� �$w      �u����qvD|�t 0�RJ�W��Qd�      ������`087"n,� L��p���#  ���;      �:[XX��`08'"�V� �\9�5Mc# ��      �XXX��v�}fD|�t 0�RJ?�m�6�� #��      `����<�|nD|�t 0�^�w `�8\       6P]��s~L� |�����  8Z�       ��뿏��"⋥[ �ɓR�$�Jw  w      �MPU�'"��0r 6�C���y�#  ���;      �&1r J�9�)�  p4�      6��; PBJ�}��=�t �]1p      �dUU}bmm��a� l�V���t �]1p      (`׮]�4r 6��~���#  ;      @!F� �&KQ��  �3�       � �)��������  �#�       ��ڵ�qND|�t 0��kkk^q ���;      ���������_*� ���ү\~��?V� ���      �]�v}��j�_+� ���kkk/* p{�      �H���XJ霈��t 0�������SJw  � w      �!��v�n0�_/� ����=��֞U� ��      ������F�7J�  �)��m�Ɔ *�      �!����ќ�q�t 0�<33��  ���      `��u���`p~D��n �Oι[� ���      ������#w `#����Z: �{�      F@UU�9?9"�n ��`0�n  �w      �Q���Z��S"���- ��H)=}qq���  �       #����i�պ0����sR�����  �       #����i����X-� �������*� `�      0��~kD\k�[ ��p���駖�  0p      QUU�9"���- �XxI�   w      �VU��SJs�; ��p�����JG  ���      `�u�ݫr��; ��7~�t 0��      �@]ח����  F�E�^z�=JG  ���      `L�u�D�o��  F�)SSS�+ L.w      �1RU՞��r� `������� �d2p      3UUU�� �Ⱥ���_��� �d2p      3)�������ҵ�[ ���j�^P� �L�       c�i����w��D�u�[ �ѓs�`yy�>�; ��c�      0�fggצ����.� ��-��๥# ��c�      0����nn�ZO��?+� ����8�.� Lw      �1��tMMM=!">R� 9�����S� �,�       `nn�[SSS��?^� �V�� ��b�      0!���:΋�ϕn Fƅ������# ��a�      0Av����V�unD|�t 0����>�t 09�      &L�������"��[ ��Rz~�9��  &��;      ��v��s>?"VJ�  C��~��� �d0p      �Pu]�e��I��- �pK)=�t 0�      &X]���9?#"VK�  �+��KM��P� `��      L����(��܈�n ��o۶��� ��3p       ���SJs�; ���j�..�  �?w       ""���^�s�[� N9�s�[� o�       ܢ��&"�(� �V��~f� `��      p++++��xS� `(]\:  o�       �J�4����gGĻK�  C秖��V: _���v�������=g����"b@J���Hc��	�((iAꚲۈ���")�s~gN;��h��f�	����(%!�>!o �T�HDH-�(�
�Y���9_hл��9���z��׃O.      �G8y���d2yeDܗ� tK��w ���      ����VD\[k�lv ����D۶��; ��d�      �cj�濧��/�R��� tC)��]v��fw  ���      ��5��\k�&"�n :��  `1�      ������^�wMDlg�  ��˛��Oʎ  ��;       �d0|��z,"v�[ �t߷����� `��      p�F����Z#"��- @�� ��1p      ༌F�{j���  W��m���  ��;       �m4����dw  �.[YYyyv �X�      � ��p�� ���z7d7  ���      �RJ����7G��[ ���k677�fw  ���      �ֶ��d29��n R\���smv �8�      �(��x���,"�-� ��Rʱ� `q�      p���־���~����� `�m���� `1�      �/�������#�Lv 0S�����$; X�       ��`�R�q6� ��Z�� `1�      ������#�7�; ����m�C� ��3p      `�5M�Z��ew  3󴕕�fG  ���      ��4�#�]� �l�z�c� ��3p      �@�R����Ɉ��� ���Z��ZKv 0��      80'O�ܛL&���Og�  ��S�N=?; �o�       ��x�5�L���/e�  k:�^��  �7w       �x<��Z��� �@� ��      ���F���z7D��� �������?� �/w       ff0| "^�� ��d2yiv 0��      ���i�o��  F���� `~�      0s��p\J�'� 8/m��Pv 0��      ��RJ��ں)">�� 컧9r䧳# ��d�      @��m���������� `���k� ��d�      @�������5�֯e�  ������ `>�      �j}}����#b'� �7ϻ��;�� �w       �5M�w��#�f�  ����8� �?�       t�h4������ ��1p Λ�;       ��4͛"�=� ��xI��dG  ���      ��(��^�wSD|4� �hϸ�� �w       :e0<<�N)"��� \�g  ���      ��Y__���t���8�� \�R��; p^�      ����O�Z_�� ���Z�m�C� ��0p      ��F�ѽ�����  .�����OdG  ���      �N�F����  .؋� ��a�      @�>|����gw  ��j� �3w       :�[n���ٹ."��� ���j��pv 0�      ����_��od�  ���+++�ώ  惁;    ��)  GIDAT   scmm��_��Iv p�J)/�n  惁;       se8�EDldw  ��� �|0p      `�4M���{�; �s�¶m�� �'�`       `.mmm��ew  ��G�}nv �}�       ̥�m�u����#��- ��N�/�n  ���      ��u�m�}��r,"v�[ ��WJ1p ���;       sm8~��rkv ��j�?��  t��;       so8�="ޑ� <�g�u�]WdG  �f�      �BX]]}}��o�; ��Vk��� ���      X'O�ܻ�KNDė�[ ����  ���      X��z��R�+�|3� xT� ��2p      `���O�Zo��  ���������� ���      X8MӼ;"���  �x�� @w�      �����g�#⯳; �GxAv  �]�       ,��ǏOj��_�n ���; ��      XX��諵��#b'� �6w �1�      ��F��GK)�� ���R�n���� ���      Xx���k��� DD�%+++WgG  �d�      �R���7�R>�� D�R~<� �&w       ��`0x��r""��� ˮ���� ���      X����WG�4� �Y)��� ���      X*������� Xr?Vk-� @��      �t����Xk�@v ,��ӧO_� t��;       K�m�i��UDܟ� ���ٳWg7  �c�      �REĉ���n�e������  t��;       K�i��j�Mv ,)��G0p      `��F��E�{�; `��Z��G0p      `�M&���� X2Wmnn͎  ���      ��7��z�ޫ"b'� �H������ �[�       "��?�Z׳; `��Z���  t��;       ���h���� �eQJ1p ���;       |�~�SDܟ� ��w �{�      �wX[[�zD����� X� �w1p      ���4�}��qv ,�j��Pv ��       �(��yk)��� Xp��=zev ��       �(J)�����g� �"�L&��n  ���       �����#�DD�f� ��*��Hv ��       �8���/"ޘ� �� �6w       x���wEć�; `A�pv  ��       �ڶ��z�_���[ `єR��n  ���       ��`0��Z�k�; `��Z�m��� @7�      �9�F��R�(� L�ȑ#�gG  �`�       �a:��!"�%� I�߿2� �w       8���LD�*"v�[ `Q�Z��n  ���       �S�4���� �(j�Wf7  �`�       �̙3wFć�; `�R��n  ���       .@۶��d�x(� �U� @7�      ���_���fw ��2;  �w       �MӼ/"ޕ� s�m�^� �3p      ��4�L��gw �+Oy�S�� �3p      ��4�����#b�� �joo�� @>w       ����.��-� �U��3p �      `�lmm���� �9e� �      �~i�����_��Iv ̛R��; `�       �i4�}Dܝ� �����  ��;       �Ç�vD�Sv ���w       �w��r�N)�5��� ��j� �      �A�����9� 戁; `�       �̙3wD�ǳ; `N<mss�I� @.w       8 m۞�����- 0��?���  ��;       ��h􏥔;�; `�z���n  r�      ���ں���� �� ���      ���m{6"n���� �^����  ��;       ��p8�t���� �e���w Xr�       0#gΜySD|!� :�� ���;       �H۶߬��5� ���b� K��       fh4}����� �(w Xr�       0c{{{�F�W�; ���`��      ��mll<Mv t��; ,9w       H�4͟�R�*� :�� ���;       $����� �!�� @.w       H�4������ �Y�  r�      @��/��TD|<� :�� ���;       $:~��$"^�� �'�ZKv ���       �5Ms_D�qv t@�ԩS�fG  y�      �vwwo���;  �t:]�n  ��      @lll<Xkm�; ��`��      @G\q�o��Oew @2w Xb�       �Ǐ�L���GD�n�D� ���      �C���?\k}wv d����3p      ��9t��zDlew @�^�w$� �c�       �����R�� ��Pv  ���       :hkk�tD|&� fm:��� �<�       �Am۞-�ܚ� ����|p�%f�       5?Xk��� ��Z��; ,1w       �QD�dG ���R�� @w       ��ht)��� 0C>��3p      ����ݽ#"�� �Y����3p      �������'"ޒ� �PJ�g7  y�      `loo�.�|1� f�w Xb�       0ڶ��t:m�; ��Z�`��/)���564�    IEND�B`�PK
     ��Z$�8��  �  /   images/b96c8ad8-7845-422d-b49f-326b2968fdb8.png�PNG

   IHDR   d   �   ��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  WIDATx��]	��y�_wϹ��^i���@� 0�q���$Ħʮ�R&�`W�Ul�T%8v�rQ�6�������# � �s��fv����������jzv{v�z�;�=}���g�Ò�!C����AH�� $`h04	�B�!C����AH�� $`h04	�B�!C����AH�� $`h04	�B�!C����AH�Bv�['��G$I�E��vo����6_T{���V�Y���'��1n���]+�L�p٬��J���ˉ��!��8��{�$�}�`�ƶO�LIʁ��;W$����}�*��>��&QȂ��N�cJȮ�����ݻE	��T�RC�/CE��aǁ�%�������>�8	c���΃b�����6�mz�MB�Ν�~��"ᰴ����Ƅ�]��&��WtG���E͞Mu�BNA���
<�A�H<�����Qo�BY�r"Ρ�������S�l�&ټ�%�}�
���%�)!��9G,���(����4���A�%�U�)^��Q����$A$��Aƛ �(���nH�'1P�A&�f���^-�w��2D��H�r��T���������R��|�_R~��s|�Æ�~�	�ļ����ޒ�����R�A�� �|�.4�0�]*�%���y�P�n	�㸫q���������:tZ^]�_	i_�F��+���mߊ]G��zW���4Ř3��]]�N&��C��#�/KȀ��]����|�����--2��$��WE1~ �����W�S�ID��$v�q�*{��\n��\�O�Nw��c�ſ��BZW�>oE��-��鑝r������7|!�%�3�$��C|�Y�$BK- �u:��}���ʕ5u�i}t���۲%�ٴ)��ޝ���{��J�a��z��j�JO��|������'�&�d0�S������r��T�RB����{����Uxժh��c#�͛3��^J����ʲT���
���b�B4�o���D�MJU���x�G��>2~���V� �=�Ւ�g����Q�����	%�Z�,�y�T���n�_���$~s%$���7�?ERv�]+6l���a���d�F��A3�Fe�V��mmV�g�n�TK
T�}��cC5���p�N�_�T$�"g���8"������|H��D"_�6��E'!{�:KlF�^K_�WS���d02��TdݺX���ned�:���}e������t�C%��K����QxLfAR\�c.^�_yesߓO&ac�**%�R���hd7I4�z_-o�!c��"��ߛ�f��fRSl�&���E5�X��3:ᄈ��餡�K*f��q�y3３��ȆV�GN=5[b�J˔)F��˚����Δ\��])����k�:�5!�'gh}�x�� �J�Z[�إ�6���C;�z#��#)�����A�{HCf�ƴ�m[.z��q��54���PH����ɼ�V�y\��$w�������?�Yiy�y+������w��.�i�5B2\2>��f�ԤT�{�vmO��s��:��뇇<1�J�zc^�duTx���ʼk7�TJg?�0[dS��C}�\�m'"{K�NB
�)���#p>���F+4��5]� #[
T�Pg��~ՋH[���:��GM�pNk��~R
/�L�.�����/{]O���L�����-Pa����+2�����N�����)/2PU��a�i3��IF)l[s�Z<�o�����|p�]���R�?���v��[$�ba$�tt��C�#�ɗq��A옾L�\Bz{��O��Ԡc�?r�Y1s�|k��
��Wӧj�4C#����P-�=�x��88?U���ӺH��*#�������%�1c̤�"Bv_|�@����0�.^�|�� �!�+"�� �r��_L��|SYŀT;��;��=�C�ǂ0<�.Ӧ���|�ub� �А����ܥRo�b���ڵ�C��*	�c���e�o���v�� �i�C|��b�~����sRKT���i�ݷ�W�̔ۡa"'�5f�0G�����Ͱ��sU�����0�L��h�1F$�~�K�a�a /�ҷ|�s�L3�bED�dĩ�!uB��aK��K{��#KH���6�U/���
.(�Qpa�%���QM�	d��g#N�C��K�8�\Y���5��Ȅ��^��87|?! ʈ�_n�u8�NЀ���-H-Fc:���bdB�o*fΊ���a.]j�v��y� U��٦7���;Ꝏ�A�۬!�%����Dx��b|<BJa��Z�4侕NB�?�qc�I$�:��l<���5g�Ȏ5���R�ީԱ��,�� ��\#�!���ν�^V���Pm-EL�W���а��e�D��.�=F��U?h?]�{@:r}�uz{�U:��xN��?B���^v�0�HiRa�݅}:��?.�ukV�z��Ji)o�2@^eQ-]t��'��Yg�.H�������o|y��Ǟ!��>Rx���8l�F���3lӤ���aOB���aU�|������ad�W�xCH�+��𵌃�Y����_h=5���f�QB�ǔ;N��5�4v����]D��&RQ�
OH��Qe�U��t��`,�E�a��*�1�u���!C����AH�0�Qe�X pR��K�s�� �:jY�?�)!����dc���I������.ێR���aY	' �R3B
O֑J5oO���1�ԙ�f����C#PA�n�D�۩�܄�Dǽ�ˠ&��%�m[�}}��l�L�Gc-������l����Pwq�[<���"!E7,A���>��DQ"�@��ߏ�#�4�f��Hd�nlJȮlv��\nJp(_	�im��ӱ4�c,I(��!f���ؓ�N�B�J�!4���t.g���(�Q*G2Bؖ��R�;��d2_%��<>d�d�*�uJ����we2��NQ�q�k�C���R2��m����kB��ТG�m2�t)ݶۑN�q�~�W�-!$���6c
\�R2z��n�d��.	)������香,%1Fd$Æ�WOduI+�%�
�:�[<o" l�'D2���]�U��a�/�T̆W��rM�XF��)Ґ�O@FF��"YW���y��7�0R$A�1P�Ok��T2
�B��"�4ா�yd4'A��e�j�� �d̂[�b�}�o�H��Օ���w2����rF��v��{�߷d�h�d�&�>M��"�L�����	D�'!J:�� �1E�\�e%X�/�w�v���}!�G?�x Cl��q�i��6��5K�����@��d�6߳��7G$߻s�ŬYR+TC�w��9M|�4��3�PSV2v�vt��D}VSZ�FSR�8��s28�c���|���?_q{�Q]E:�2�mU|�9�P�ɲ2��~)BBe:l�j�0r(�5@��
�]�#`��pJz.ǽ&��TZ�KtG�UB���dG[�,ڶM������Qԫ�"�a+>�(�Z�;)O��U�a���ǆ����ʓ��C3�����M�c�}��Bэ����aW��Ve7gU���$���<><�t4�����U*��1o�,�q���	A �J����+)��@�5*����cuuɶի�ͧ�GK�rorr@�_$�}���$����Y�>�[!�7���'� ��A��Ⱥ��{���o�|]O��M�*'�D��&(WJ��ڣ�U_uu}���Um�^��*'�Kw��':<�58�g=LE�\�r��i.��	Q�W�Ji���T^;�֟o�켣�si�0�le��u0h������C滴^�>{�2��-~\�2B�Ov�A��y3�q.-��l?�8i}睪.3�8uoe��dC���(���ž���ޫ��②�Ǵz]�#���G��p	؏?��#R0�@��T@�P��J\�S�Mw�ʮ�Ď<��:4�cX��L3e2���-w���ގ��ի��>�{�p8�P�X�,��ϗ�M��T��Z�*&�0dl惮|�)����ⱅ����}>�^B��r.����♧#�@W���;�._	���SY՜�T�K�)��hѓ5.�#�+�m�؝{d�C�3KE*z�1q�8�%��M�$ħA�#|��%������I��z����Qv��i����(NgǛ�f-�-{��-����n<V*!�F��LB�\���dj�/j&��И����TW>�Ri�J��[["���v�K$� �,+$A딻3B�+螞��9s���klG")+��wɈV�ՠ�,.o.�
��ް�ǹ���W]�-��ch�Ɛ�����������G�V���Jq�/'�}{ЂpAU��C#���b�J���q,ٺ��ˎ�D�\��kM5%ׯ��#�H��d2"P�e;���K����bc=�G�Ɂ3YK���*�=��f���ZN�:. pquWW|���C�%�[Ϙ���+��z�s%�ٳ����t4�p�iF݅�Msb�U�;;+%��=�ܔO����,/L��۶I���t��sU�Qy#��Pȩ[R�X�3ཽC�J�[;�Я��v<�z7�ľY�u��@%s�{���fx+�^pW<�^x��:����h4',���P*r9*jH~H2JSGJ���ӝ��Z} ��܆��|�9��k�tv��%�(s�\��I�84�P�W~����
A��zS��+'���1��G�tp �O=�G��r�����	�s�'���w���l�K煙�������m�h�����V��[�TQ7q��ʲޔ�4T�}��:y>�����˹gΔ�9���O��/J�C��Hd�:eΙ��}Sg2�=�P�>,���ľ���5eE����2�{fx�ᰄ.��[��|�omܲ�r�*�;==hԅ{����F��
����X˖I��gtv�F��l��O��I')�ǚ�%�0�Y���D3}$�ݻ��G��ߗxC�\H��2��@�(���Q��3�5L�ȢE^�D,�.��1�a�v.����E~/�_����cP�>��-F%����T�>{��<�H���r�H���O=��d^]�׬Q��+�$�[)��V	�8г�={$��.9�*'��$*_q�K�?���c�!���,\ۂ}����5�g�q���u�ђۼYl%���O���8�*����&x?1<!\e��s��������v�a'HK��3\2/��s��.�����Th�
��9�[I&$�%
�r�i���%w������%N2)*�P�"0^��Q�{s�k��3��]L���Q�K��S)�}�d7m�܇z��^����%�8�
H�\Ɯ���7F�ituݮc1z!����W8��ST\��4X���}Cj葙l�G�E(���*�@0��/�KIq��t:��b�a�Mr2�5w��Y�\?��4�6?��h����	�b�H�O;������3� a#��)=.��lh�^ɴ�I+Tp-0,!� �;P��ԩl����@d�)�h[4'�	���O9ER�>*YcC��h�i�db�L�0d �w�L�+(7��!X��9�]R�1��Sl�+�TI$���0\Ca��]ǵ���c'����n�y�m1F��EБ$EC%DW���45m���	Z�l��\����F�+|�;w�����$Ā��e�Q$?w�T0������W��C�*��j���q?�	_ ��>ށJ��{�
T�V��N�0�.�JT�e����R��_/�����~&�x�}��3�`�K�[H<�+�m�yr(e
�J�9��y,��<��*�X��	 !�҆ћ+\�6�;Ј��Q�3��MM����4��F�
)�5*v{[�2v_p��W�����oy����9�替�}+Z�Q]���HR~�_��������b�6z���@���'W��}Ar[a���C�?�쀻C�񩫯v��ޙݲ�0�߅��bU]a�*u�Q�`�+�ȝ*�N�������G��fF.z�U�=�_.�W]%]���Ad͚�R�>�� ����绪C��-҃���.H�Ǌj0o���	��GF�{�a��)v���}�=9��|�kσ��a��G}��8��D�ZG01jP2�cY�,��A����n@�`�^����hP�P�ּ��
�g�q�L>�������^W��s����.�t��b�7�5+г3����4��=�����9�<r��ٳ{I��d�t�׭����^���\��K"(;@�m0�+�9eL3��c����e&�e���`����|���~��s��{ͭ��w���Ҿl��B����Ά��8���k�˝��ƾ66���������@ʝW\!6*�5�TW��}p��2��N�f�$h6t�Z���#ɤX�ؒm�R��Ê7*�DEK
tϚ% �c�B9�����>��x�p*er�]w�)7�t�H�Ѣ�kU>�0�=T��t�¶�X�V&�%��+M *��-K7m���A3�Bw:���¼��$�ױ���m�ҥk�S�HAhAe��I���K�k3����t��pg#��A G�~`�<Wu�z�y�����<f���)&K�q��/���~�k�WA��z�%��u_��k]yʫ���6괋Ҹ�?/HP���n�q=��w�H�Qx^�w2�cy�������-?�Bc�	)ڄ���9����%I�dF����AH�� $`h04	�B�!C����AH�� $`h04	�B��J��w���c
��Y�yLVB�B9��!H��;!I9<Pe݋�VطW�CJ�RM��(�+��P�R�.Gp e�a��rp���,�t=ޤ�;!\��(�Tq�kA��Z�/X3���;!�O�:B��W8�Z�٦LB~+�DL��*�CR�F�3��x�R����Xa�u���NKR�G��;+�X�R����Y�����Z��?(_Fy�_�%)uMH��7��A9ՇSӞ�G�ʏ��CO��o�Z��	)���x*���1G��,@�.�`�Rki�{BJ�������Y>]�;(��H֒��'�(!���R�GQ���U�o�ˬ�|U�!�u�]5Q_����P.����עp��kě8�&�LB�R^D9W<R�|�=/NAx-?���JL(B�R�D9�7�%��_��?�&?�mO&!D	)���<�r�O���c�򃟤LHB�R:ĳ)�)����*����k�B�������iD����qʧ�3	��	MQB
�������闣�&�
�EJ&<!+����<���t��T��q��_�����&!�7���XZ~&��s��['/�{���LB
(Qa�7�ʏ�<-�5����Z�5�!JH���D7߫�|�O���*oM&k��RR��r��#����� �:���7(�P>u��;ʏ{�Ԅ��+��ʓ��{�Ԣ�V�*i���>��u~�    IEND�B`�PK
     ��Z=�W2�@ �@ /   images/14f4e0bc-85be-4a63-979f-9a3c78ebf9d5.png�PNG

   IHDR    [   ��3�   	pHYs  �  ��+  ��IDATx�̽Y�l˕�b��Psՙ�Dށ�l� �lv�a[-K-��eˆ�b��6��`����n0l@6?�C�ղ��9�&yyɾ��Ԝs����V��]���F�� OUee��b��[Sd�G|zyyu�}�<y.�g.��J� �o��|魷eggO6E!eU���8'��R���"I��=�,J��o����x]U���J��xVߗ�ex����k���R?��w�U���|x|d��׉����������?��������^-$OZ"�0�k�z����ch�CǠcYo��y9������v��1j���J)q�|F�E2}�u+I�;��cO������޾a�R���~���x�p�����>�Eo����~r���D`�0-X���5K�F�fc��%�U��pa���T��u���!�6�Y���>U�y�W��c�����5)�_��s>}�O�A�Y�EǠr�׫O�H����O,*ʑ�����]��De��$�&U�їٵ��ki�Ey�6��^�� �����C�
�ǂr�Cl��jez}�����W��z�\_�U�1ŉ���i�󪲐B_�f-�::zo�h���|-�Fe$�e�=���u�ת�o��_�7����]l6|�[-I�:'��LN�m�v�����~K?[d�*e��YWz�����]�nG�����E��ɤ���b1�����t~�\%�M.�~O�^[��u�������R*�|���/Vs]����=}t���>s}~��a�qa]�e}g8�^���]��Օ�o[?s �~_��\��]���!;�M�?.��]��k���#��k�Z�V�mw��鮥l�:d]�5�$]s�F������ߗ;w����X���έ���G�I9/������c^��5���h���+��d�k�}�;��{�����T�[��X�M��u;��,�c�jK�9����k:z��b)�j����^;չW����F2��?��l)�������۬��m��A����[�Z���g�;}��B�W�B�;*�mY/!k*���N�s�Q��	�ݖN���^�Z��{��1�k�>�j[�j8�QUz�X�L�t:��\ ���2�!�2i;PP�`��*����S�k���Awy���*h'��D7b=K��o�n�,Mj}
}�B��c�r�{�V�׬T~
ݗ��^�K��$�sA��ԩQ�ySSb
_�}�O?�*�[���	����`N��J>�=]��A���q��2��p��rOQ�u��e��7a���̙������z��x�,��>��zM��іƱ����l>.����6*y��5�U7���Ma����5�����#�k�[륎e��ƽ��8��,��/������{�,�&k�:.����ƨ�ƞR���N��I�IV9Uy�L�nG%U7eO6j���B�?+���>6�#/��C���6���/��������3��l̓ q�'����?`#>�E3���`n��<Q�k����6�gx��bX��'Y�Qx{K���s��0�(���+��+��{���o�ϙ��埼xs;��vƹ����Ϩr�}��D�>�;�q�7�~T����_�� �����������Od��OD��X�����۹�����|���f������������ο���;�7�+{���gG�'���B͂����\��Nd�F w��	���nz����Kh<�ed�@^�����w(=�V�a@5��oBM�^�}3b�2	B� �:����=U&j,}Y���mp�n	���*CUpI�X��=n##�y���+�Hc��GM�3Q"5٢0�vCcjJ���a4PUe���FB�.q�g��#�qP�X(�@6��`�����)� ����h߫@rI��=(��"�F5)�mb� �Yb�2̋��'��|�i�T7��-�K�`�	S�"�"~��@t�@��^i�r�I���}=.)�5�'���.5��I"��m6v��8��H���O�>���P˥��E����Ś�t
�*��f �
	�������L�pb�uϹĘv
�r��U� Ҕ|*M�h9���Q����p,��.A�|:�Uq#y����3�m���J[?v�k�����T
xW:. 쎒�T��c���$d���FIN�,9�%^���5�1��S��﹙**���G�fs	<ֈ�^���ݗIJ����s����0�9tI(�� 0p(@W���P�G�� : 񎒁^�G�7[̨Gzz�^W�b[	�x$��ޓ��#�(	�$42 �k]��lJy)r�\�~�X*� @��8ǃ�<�Tfz��{:�C]c�D�U�m$
 |���b5���@:: <&%~}�V��l1��tv�}i+!���Q��k��ʌ��ɂ��S��U��Q���A�DCn W�W�j��HI�P�%�Ìs��(�ֿ-�.����f �m���\����:d
P� ��r����aQ`m@�@�u�2�\�]����WB�9[�P���ެW9��y���=��b=�Zt�wt�2Y�g�z��@�Ľ� ќT%ǅ��s_�t�c��!�W��e���ls<Щ���?�['ц����c�$4A/�@:\�3s�T��t�4t�8#ep.���U�'±��1�-	�*	��L��N~~R����(l�5ȱ^k���_A�\���c��g�3���\�P	���� ��şPN+:� s-ߖ��}��̂�l C'vun7�5�F�`���n�|�XD�jx��E��q�4�D�K�Sʱf)IGY?Wa�ws݃��:A�U����; �Q�;ld��������J�	��Y�s����`���d�p��<���H�>^�jHx�mq0m�݋a*#���@>0�I4Ppj�I�O�c|U�.Ա�8 �zR+>��}�e�@A֑����@�	��z��q�]�[,$b}�2�l|Ƭ`�{CUc�-&��Y���y�
�?K����@�����D$R�2�x�% ���/���_���$!�g"œ?���_����j�DV��ˤ1Hx�W�ߡ��Y���_�����{�[��ֻ�}���z�Խ�z�7ޚ�������7�7�+{���'�n���b�� ��M��f��ȅy{�K�p�e[s���ӫa ���Ge�E
���2P3m	�[ұo�<~�cA�m�F�N�h^U�Z���%�"��ڌ�Z6��΀^�f����SɖQ�o�O`��H��N"�c=mBrd�^	Fs?�x+ܜ��+l��.�·�ʖ�S����vU�������S��z���-�P����a�0)�:.��J̉A�<M>�1З�U�T�MS%f|�M�U璆�Ai�t�m$�E��g/	*Ŕ���TQbBƐs��Sj�V����I�"��s��4ڜ�)����E��M���B2��f�[��*�(�cc��7wPTau��N�>��\
 Z0<�
��V[Z�.�Fe]�0�\��Xv v��`����*���&9I$���HDapaߐ�;�� J�#t, F�;oX	J:�f<0H�6�
��4=ͪ>]��篤w�E��C_�nhuF$PL-��(���F������d�	Cip���Ag�U3�����(��\��ɜ�˻>���%�}!C�ϋ���e�=�9�H��{���N
�,�2[.� "���`��"�T��L����OH�m�F$'�ڎt�M�����? �W�W�/n�c�[:zKw��e���W �ʣEW@�JL+%OC]��^�<ș��� '�9�J�#x�U�z�-F�Z$A+�]I\O	H�jC���e(%B ��W$�]}]�����U9�|�A[	F�{�T; ��e4����V��&��*ɀ�$����R�����e�R���ӵH�j���B箭sOIYK�t\m�˖��=H��У�~�6�AX'J��/�u������17�xg����:�IJ@�q�r.+Y����uП��$��`/'����%I&NZ��	 ^�Iݨ�A� s������JI�l�!
����,�`�,u]��6ɿ���/C�B�l�X���G�%�#�O�S͉=�>5s�҉��5q�ԢM�?%6KF�B�?#�QrD�+!����SE�*W*��8&]��<B���M�'tD�`��:z���I�S�����'v=F��t-2��!�63�\o���e�dd���"�}�	)͗f��1qkO�l2�3�Q����G�2@W$!0�����e�c�*��T�p��(HI�(�&H䕹�ŵ+����H��F�5�rf�8D2Ӡ1��k'�.�I��4�0ͫ詊�]��b$Į��l!֐�碃�.� !Q`\�6��@D+6��pHɇq{ҧy�5i~Mz��_Hq�c)����?�\��v�4ٿ{o5�?|y��Oܹs|���6������/�x㍷F��;�;;�_��W���_��?x������q���W��[��2���g��/����������7�+��g�W���$k�C�¸ÓO�8����&Ơ�xں������.�[��\�y0�^����%����B�Q�]x�	R6�m����(�.���0��lA%v=�Q� ����H>�w�r���W5��U��l,��a՛�����H\��Z�\_;z5�=|��y[$���e�8j<ˌ�ޅ�.A�|���{�u��
)t�Q���KL�r1��!
xe~Mo��T��\���b�Q�*�@c8>��pP�4�Z3�^�����
��W{���r��|;3����b��2�6�^���_;W��b���)"_�����04&H'aL=�@hЫ` �xh�,
�k%I��  & sR� :�� -���J��]È"�o_�!Wи�\ ���W�H+A���s��������(-zG�[�@�ʭ(�8H�6S�Kr2�� �Ԍ^�v2�)bi0t�r��0�����eAɗ6>�{G��
Q�f���9�~�ǃ�# K�}x���iU5~G�eY�������F+6/'^.&+���;k��KY�3)л�t�&�?�Uo�i����:Kv�\����R��RY���ֿ�X��bV�z��][=��إ��՜{��t�*��(x��
�3��#e.�b!�������ޫ ���k��.�� &��\�d��p�v�=��D�C�f�����9�r%c}�2�xD!a�B�2�9��y���J��,R!]�h�E�q��éc��@����gJ@n���isp,-�K~n�t/#}Rd������n�C���VPy)���sL ����!�.���n��I�H	��{':��1El_��l6�*�ۗ�p��	������k��=�(P�ӥ<.U��3]
�~�����r��2�/ ���l:���|]�]����v���Ō���ku��M������>u��Մ��<W0�uFza�Zl��Ǳ���x,������"SH�l��Q���[����s�D��IU1e���@����)� �H)��=#u���ߓ�v���U;�9:�)䵧O��4��z���]�ף#�d���ѐ.}�A�ꠖ�����:$S����ǩs��%�T' b�ZʳgT��R_X�aWF�� mm���5S�֌vl�>#"��E+�N�΄nԵ%"X��,��l�1�*I��11�UCf�!�:����vbiƈx �6����(�U�����"�*�G�Ĉ����`�@ ��a�t�pt� �k� V��n�O,�l��.��%R���ĹJ�3mQU5�aӓ��0;�AU��!;�
�V�kh!��6��[����{�s�K���K�������׾�K����|;���\^?����ܻw���}���zz���z������8z��@uA7�H�>���� D����}�޽�Ϟ={,���O��=|��^�R��F7y���
��M�P��z@i0�W�[C�j=H.�#z�ొ9�[b"����2��s���/��zK	B� 0Z���Y�2�v�<�3q�T����	�ka��� ����&c�8��ћ쾎�l�F��ͫ4o�����B�L��깱�^3��*lT&ʔ=��!x�Ґ�X���#{o��\̫lއ�Z��r]|��w�-x��4F�*wӒ�M���	A���S�جE����2��4(�Ȫb�Ӗp��m4�o�I=������ؼ�.��P[��.�AC�$�����'\�ٺ�Na�\��gk0`L��#�� l4��3H^���NB�o�e��7�c�W�@ص��Ҝ���,�| (P�W��E^K��2R��{J>F��L��T���>�c.�T`�L))�M���j>�2�:X^�0jDK^B%k ��&o` �[�-/dYP�1q�r&Q�bX��h��v �A+�`!E�$x;�0��,$%A`�tQ�>K�s"��Co L@N�*�;� �K�+��#e���,�4� "SD���|���F�����>Q0�;�:9���\���i�u읾>ZJz�֧����e���N���6ט��R�_�VEf~FZ*Qj���B2r�=�8��P�Xl%D�5�{q��Y!�~�G���L"j��v�9��K��R� bX�QΩ�����g�S��� S@�}5!X���� �I�9I�qG����s}O�z�'xb!����g�����o��ݱ���꼵H�p���@=^�]�3x(�A}�D�<҈����2�[�o���ы%�wp��C�V�svv5#I��Δ�����*��Dw�D����q�B��TI�D��H����B�ۮ�8��͊�� �I��*s���\]��}+1]mH�0����Y�y�׾����Q�T��S�on��?J$��=���u�PW��)��5"4J\1� 5�N�)���Ŋ��u���v8�󥒳�$ |����Be��`�U���]�V�@�t�=����zkM�Z��r	�1�u4M��n��>�L�T��ZNF^�:n�rڡ�'�,u.�+@8�c}*B-*����tLƴݰ����2�d�e�0NG]���sm�+�Z8�#�|�P��]4��ӓ.H�j�
Ia:E��0�T*2�GE����.ߔ���i���e���G�w�C|l���UO3J�i�������*Қ\��@W�x@g�`(�^7e��@M��$#p�\�nX}PL�a�p�J�&��y�����tk]���5�G����F[����x�[\X�;��G� ��kܨo`#���W�n׋M�e�X$�%�P����|��4��W=r|r ��;_~�ͽD�+Y/�󁒌7�x�M���@XS؉�*���2*6F>��}��7���O���w���g����G�����R~�_�*�����^hb�5��A�)H�|>���
��kH���Υ'��n���F�a'A��Y4o�H]PN�B$���s�(���5Y�-$��9���{���u�|�;�X��T�D\ S�6w�����-ш9�_\5f02&���WĢ�,�qi�q6.�����{%َ�
N�kVA�0T��֛%�)�H�ll��6>3bI�pH�A�� 0,�e��i3�!C^v�k�c-�S����k] ��"��b�c�F�zqi-6�d�}��ӧ����~N�0����Hm|�E���I}�d���+�$�m��2<b���m�s�UJ	b�3�c��S�0[�@J��3Gu�P�����8az%��΀��s5nn��iC���[��*���S��b� {�	)}��g4��yR\�R��"�3�<���m�uR�2�$��a c�:kY�*#6�!uZ\�OKL(�f\m�riE����` ����aEpj���"��Vg
�
�u�*�I�	�*�f�-fV��m) B�����@�CBPVy�.k'��כ#ǐ��3�}U!�;�#��`�0�V�/mF��s�Z�$6�>XTiI��'�(�M��L�� ��D]S�	5YUL{؊�Gt-�擎Vg2�Z?������gz\e �Q��ր�F�];�m.]��A���:e�' �����%��0�W�D��7��{
��h�e��J磚%�h����SOV%���56 uh� o􄲏l%i�e�(��٩���7�����c֮���|.��jS�����յ��<�;w�ʍ~jPN_����S���Q��R�K��O��^\\�l2#��� ���� Ur�d@}�6���$d:� vv��ם*�j�^>9:���_�O�ɇ�L�<~*G��l������w�Qb4��l��1����\�_���F�߻/{z}�s}k���CB�'�sP��
7�yy~&W��)D�Pos=Yp�ZYGm�H�0��7�,]:@t��b"�f�{K��T�������a�!z`�+����F]];#>�:A��rB��j5�©�y�����l�g��C#@h| �,�NX��Z B�_����@�m�[Y����2B���&�u�����Fje2��|-���^BTQIdξ	s���sX����#VGk�%�1M�����>�h�E�����6�1����de��hm:����p�՘�+rs8Db���44*�]��E�5O o"ٲT<*�2`L^�=�{�����	�D��j[#I|6:5>�u��3:�%��l�bT�	2�Pa�/µ���[�SG_
�ӽ���� *>U2^()������:�����;G���'���`���^G���F!{����+洬�-9::>������z�����Ϟ=���~���5�SP27�<��a��L(�SUP��l�V�f�&��ʃ��W���y�k�p�w(=����͏�n'e(�RP<�t�P�l5'%��m��!O�*���W�(ֹ�����;�ˋ'��T��Y��*��4A+�����e+�M�� ?ַ�<K_��Uv!/�V7�`��)FV�mE����J�Zt�u���5������_WK��Y�v� EM�qe^��כ������X!] ݚz�&×�o���%R�9_L�1�R����J>| !��V�'lfP��&[O�K�"��m�I���|T,U�<$x��(c!����6��s$���!�	jc="��YfX$�-":SRH�`-HHI�Ji
k�/�b%�g��9ƎJ���w(��%���]Md��灾OIHG	ɦZ2}�����"ӨpˑW"��9>��,oPڧ,�4Ȇժ��ۮd�A�c7���Y����n,��h!�NOVx_0v�$8���i�ع!
Q2z�*���O�Mx�*ԍ������;+���Z0�x}\И�.�-UG߻��*������j7������M)���b#L�A�&�|�=�23��^;i�d��X�PŚ��60���i:ע�7b�ü�4l� �Up��o�.D�*�<oLh���
~KE^Y^ѩ�Cj'�����7F��/ j��~�ggF�$Tr�}�u�IB���m���8�d;	��d�@MC.�Y�D't�!m�kĲz�E����6rr�P��ɽ����P�]����v�G���X>���)@�2 �\�'O^\x�_^��ˉ��K���U{9!�X�HǉFh. p�V����B$d:�����ޮ~�>�%/V�ڣ)N �w�R��� ��*H��Og4�<�����k��3<P���0�w�&_U��X-����H�~�˔��K%CәELt]м ?o��ji5e��/t<� ��� I綟���^&J���o�������/��w~���aD7�K%y/�������a7ө�+)�h+9oơ�H�z6t�@c Y���"��y[Y��|E�hT�9Eݐ���Q���l�g���b4�@�"4��������2���5:��!%��B�}W�Ar���TV(_���ںF3�O� [��}�܄��*���N
XŁ���s���4���>�[4���е��f�!�Q vV�����"��,���E*l�}�Ɣ-��	"�*{�t�r��lT�t��"J\����!��3][��bϖL������`��D�c�1N��x���TT�5	�d�4�C��9`b ���k�O�a
gMj\ p�FVK��#S$a�+��p�2�D��}-'G�r�ޡ��y<*�=�宎&5�B�(vҋ�4�Ps�okeAX�ܹw�w�������G?|����~=�_�W����߄�9�ƢQx��M��m��ww���ݶ�jUm=3��R\w:��cf��k+�K���%��wTy��;7zIZ�yx�h�@�����Ghu5�3t��.���t�q�c��uh�~��t�t�tkPZ�ná��um�H�aݦ	�k�o�EyG�x�Q��E@|�BɊx+V�Q� �c�Bc��	e� WHeѦ���=��y�Hg@abhk�@��Ʈ�*�U��j�f77
X��X��"���E� #jD��>�HekwЕU�nA���+�^��-ז��a~\�\Ü��7�_ �%&��E�㒘ץ�l$�,tc�n	J�{Y��k��&��A|�y<���Ђ޼<Ie�y��LI^���@sW	6�!�'V
&�J��/ksW��:�'{9�����5�LINr>[Y��J�॰��N��)�#`(��ʯgL�`;Z1#"�ei,�'I�=m�����#L~�7���9MP��T��$O�����f}I��Cbk�z?��'i�'��E�^�6������UO���2�`��۝���ْ-����a{E.{h��]D�_ȳy�lh�T�\n�<� ���u��f��:]P]Y}�J��nk B��ӈv��{��j�!Z�%F����V=�B�$v����Y�w$/Ya��Cj�D��b�XB�-:�U�'3:s��T��Im�V�Ҁ�%Fj��+k���|����bQo��'���kK�@TB���C%��}�Gm�`~]2">��U��䎼�ޗ����'���Hfx�L�y��|��gL�z��\]^0���h���7Rvvw�i^�]��O��.�uς \^\���^���[6Wh֒�S�Pz�!���nD���)���*Y@f�qk�NB��T��Z��B����Z��f��x���;C��R���aggL ��U/O���"ꂴ���/��>�ÐQ��lF�=��cJ���5ea�gD>ؖ���k��m�@P]�ny��[�֛9;�f6�ѽ{��HD*�|1#)��=b�n~=��/�><���>� 爞#�V̀��C��)���3)O[�;�;�B�&Ss�����R�0� vП��=/�$OH���CKkD�P���}�y.֘Ŝ���1���e^z�siS��A�_O���4�o��[(&l%��:Z��C]�E���
���B4�3�H�uM�ۛ�#nr�9`����p��9�ކ��@��ӷ�e��&83�B�e�"��2�_c��9E��[�+OJ;N:��4�hd�e]9�2
�2�"�eL����1���z��C��������ZZ#�*�q5Ҽ�:�*��E @=m]\��L�^Z���ҡABl�J|�u8����f�딲���c����s��-����a-�n���Ƀ'������:1��1�ÍT��>|�o���!��A�:������������;���_(�P�����^�y�E,.B����fQX h	�Hm�mt�K�M#�С+
½WWW���\��e~hH��렼���:�=���!�����:��0�����n��6�0J8W!M̸(���z��Q��f*���{}��.������W��o��ƨAț�<M���=��ߛ�ߒ�-��h�����_!:<#qh�{ؾ�qU�}�v�V8˺v��l�@:F]�4A�R�.O���@[��6��>�h��x�����yK%�9��+�Ǝv��Zj����9��ʖ��7���I�^Y�Jn�Ȉ��v�l��ݖ�[<c�Da.#y:U�g~T |�1�H��-�� �
k�ܕ1zU8���G��7JW�|r-/_>W���2H�Dx� �`F ���S��z�����K5�s���Z=����K�x��=00��R(Qyp���=��^^���GvbD�A��6Şų.��u1���V�ѫ�Hǉu��~ABĳd�hA<�ѫce{��]�sq�mM���]����F�1;��T�*�4�8���C�w2/�]�k�@�
 d��j���	SŌ+�~ۭ�i!Y+Dn==�9<�:�i7%`C;Xt�j�(�{�bQ�SR��`��Vu����a<:Vݗ1�`*���гn�0D2�=#>̧�����gWX�����/܌0�\!]+Ѡ�]�t�hm[���*�1��n�Y����L\�6�8���]
���@����tى	F�S��B���y[�,�__^)`���oޗ�ߺ/�����:y�����L~��3	��.g����#�ɐ҅sjP��|�V�H�C�H�1�7Խutr�zq�v��pCV�s����ܽ�H	��R8R-���W�9���Qt�m���v7)�,Uݏ�����W�M�/��������>�L{1�b5��c�>H�Z,��Y8�iY�9S]��ctG���'3Nūb� u,G2V���d9�}��҉�V���5	,>so��1���d����\+!����:H��R���\�`X�g`���D�`c@�z�����`���}ꕫ]�5E�Eu��ѱF�4D�A ��^��\I��J�����ZW!}�D]�R��%eQD?,3ĜoI���������*�fl�^g��0���@֑������F����Vӊy@ګ����(�m�١^E=�
2��Mhzbz���E,���	�Ai��)�tj�T�Y�B��Ǿ���]��#�ET?��!���p��Kf�|�y�HVf�jЛ��{BFm��podV�kON�ȏ�58bJdԬyĆ�,
w�ALG/C�>��$��9��$L��χ��h��ІF�
��5*�w�3�rJ6=p�&Qؘ#�zl�B������ߨ{�U�(��a�%w�Ȟ�� U��!�X��"'��t��zL��Y��(���u�ޚN@O��^�T�=�����?��������?����"HH��G?����+b����O�_���p�֝a�t��L��P��ʚ��Z�)�L&�6��u-�B����������8������Vi��V����+�����Cc#������Ba]E���n��2"Q{d������[X%z4_)_$'���hF?$�S�Hl����u���U� 8��T��@HDj���a�L��/�'U��Ʀ�ਯd�r�����KY�AY�R�On�Z[ t.�>Wx��1$�X�e��Hr�JG�h��9Q��U��{��*9��������LfK5<+��CyO��oΥ�e�{�2��k���^G���X�����]��5	�
���M"���m�f�$�
a�·�X%��;J��T�����[��5y����gS��}�Z����xHލ������v���9�� ���Gw�+5�Wru=e4�X�� ��z�b��f"/?�Y(�����������j�z]6	 #k06!�=�Ѳ�Q+��-EXW���s��-���i��*���A�}�~�(�����jٯ�0a��A!�	��E�s����?��F�U�Q�V
�*����1��P��n� �}�7i������l�*���%S9�m�W;{�Ǻ�#�Jzf];� ǹ��LUK�b�D
ƨ�*�(e6]��dB�}���3�W� ���Z��E�M�-�Ģ�{��c�(��N��$FVvC�Ix,�����ZG=�Lf�S+��8
K� c'<v������ ��a�� rL����.��\} -t�YJ�X�T�!��d�1pB��\6��\߬YSpr�'�Wߓ��c���ũ���?�O?��Nf�Bb�\_�lZ>[�v ��������D�"% � ��drM0X��c�	 ����SQ� Ђ�U��:%������hG��l��*��"�KY������t-�7������ÿ��-XP�����0�V��`��(���w[hB��9�S%m<��LX��bw�[$m�ob�FAXP����Y�Mr[��Zz�;����[J���駟ȹ�jj�.�HD� !:�ي8��Q� ����R���[]EKv�v���P�:�g��Hp��-��|xR%WB���Z�=��- �"�YGIC�U�o]R�)/x/[��Ό-�g�qn@z@b@�1=��D���ۋ��a p��V1����t�B���j[[L�M�� �)6�r�"�а�[c��tJ�E�{[�.S��س���NA�4��:���X�)�Xk���˥Lve��V�Ķb��#��_)�Z}�C���Y1��ڹ�8�N%��ln-�~D���V�t)C�Iў�i��kYE�m�l@-)�6t>S�LNC&�҅�� �����q�y-1"��Kg��2Fű/6$���� 3#͎ie�}�@Up&���g�5�ܘ���s�6xr})O�>ֱ���Il���pε�\�3#�K8�+�TU�p8�)�h���	e	�]����������js}q}����������l��[�-�b��:�xqΟ���2��;K�����҅V�6��G�<�1����#�����(>�b��iE�VB�Q���UHn�IE�PxP�{{�2]܄V�B�I,Ff^����-r���(����� ���A�X�� No���5u>z����ed'�G�\��淢��'u��ќc�J�HR����Ў������3SVS9?;���b>�
y��'_�s��C������������R�ē�$j�ת0���,&s��`�'��H�F]ݩ`$'m�o�@�z���c��#"q�|X�X[�g�54׼����$����j�f�]9R����0\�bz+�m��;�î���C��ۯɃ�]%y}y���p�����(؀�F�6q6R:�ǌ�LIN����z�������0ͳСi��D��G?�H>;�L�>����I���D�/-������f�K##�>ʼ�jBf]��i>�]�5%��,6�lc:R�l�����l+���d%x�XC�Z
g���x�(1�-B�"~�Y�����t�%�v�
����-3o����;��2�"q�a�l9�Fu����ZA�%�0��&vZH�I��h���|U���ur6m�'~�3}��.�]�'����������P.�/y�2�R%x� ���. ����t�E~0U!43Hc{�>H�'Љ5���A��[-5!4�n(F��}bs�J֨X$i1�p�����j��2DDpP&A��4�y�`�h��Hv��K���nǶ�H����%��>r�{,�_�W�B
nG�ߕ�^�w���W_�/}�Ӌ��>��}�/d�/�]�syx�R���Ɗ�qf�ݱ�Q@����c^@�&h�ކ�L���Q01����ؠ�n�

Lp@�t6��v�a6�0M�� ��Ëӗ2U0>�i��<Xm��ZT��;�77�ymy��G�tv�D��s֩<%��S�d�ΐ l �X�"D���R�rZ�ҭT� ���hް�YBF�,�a]M�����M` ����p�P��4���ݓ��=�����*����fr�ή<zxL�%jR�D��l�����ۛ���:ȯ���B1����U[�@��*��r`��T���R��!(+;ׂض��<��iuz�wH7d
�VU���`�Sk�Lo�7�oQq+L	�S/��`��`"
���K�;P��b��x���$��H�a�o�;����H��.���:)�%#�v��p�!����#FҐ}�C�
��ګ5OmG�+k[$N��ʼ��,���՞tP���1R�	��b�PۄZ��rE�9Ǟ�#���!��j2���<��Gc��G�(䵕 z�'0��I�]�E)v��RXM���.��~q��z��XG��:���c\8�	m�q p��m�����b��3}&账�	��n%L�j1u-�H]���Z�ާ�zk5�=�T-������lB��?Խ�D��?�TO�yK��BD��� �����(;kϛ3I�|²�J:3xH�V;u���}����o}�[��?��?�_�W��gRl�K�>�}��xÈ�4��=�(q�}[H�/�5EQ?����o<H��$��.��I��w��N�>0���kEKYH9J�m�2� ��-���Q�hT�����Hu�l=n=���_��y�# ���m��~O|K��_��Q�@:�P�+U��x���6��.}@D���g�X��}����(S}��so�����o�/���B&j��l�]D�D���t��['��	��p<	m�م���/�)qx��b=���U���� j���LuU�=����\<}=�Q���k��W����z
c#]�%,qɚ��j����o<��"]��.��[x�@D�V�=�i�8d�����Z/���\..�����ٗ�h$�7K��
p&�v�x~�
[�Rg$�C5�
��'�$�wv�<sg� %Fa�ӗ��=����P>��'�ӟ�T�<y"���T�� f�Ս��z�[kʌ��Y8���L�ltjsU�(�-)tu�*>i'�F2Q�{�k���P�m[��x�5���eM2�!^��	����������L�W�փ#��_��ܽ_6�7&
�
vvzc�/�t@@#:\�`,���}vv)?����O���9Sݤ��;R���w����,�er�Dq�X�P�F�:E�:g����Z�u�*���"2��������"�����ԧșFM���'u;u�;���B�M<Ke�i�r�=�SC�M�1_/8z���Ӗ�v�I�?��j����l�)�	�輈����[��T���ʻo�\�n�̋F�_�TD�X��ɬ���\fW�JV�r��k����Pu��\���3�m��<�:&8������?xxO���U������h8༣fc��ZmM�{r��j�c3��d�:)� �[�~�Β�������^�  p�
�.oT��^�i���wG�CDLV�cI��;��yө����~�q:'%Gq��l���K|&��X7t��QN���p��̧s�>>�g-^suv*'�(�?�~Ga���+��جPT��Q�'{$��Օ�SS4�'gr����'wNd:�>�(����{w�5]���=y��M�j0ntn�����}*O�V��JFCD��9��й�2��&+%�V2rqq�
���p����"��3��8Ǣz�~��m'���	<m��2��3��l�`D!<֫�y7~]v�u��c}�5����,|�(��Jd� ��*#�[���iOh� }�\�nbQ���i�+�G^ъ6t�ڗ�+
O�V����ڌY�H)�N�Y&���q�#��뺻�5E�>棓1B�� |G��IGnY0Hwp>�2���t��	������"�p4�h�@ڲ�\��}HAk��E��*�K_h P��Θ���px��7�\�Yb ��{����0W7)`����j�`:�)6_�@�����T��������R�g����r�w�cV��_�I��QP'�bwu5���j�N����υ�#�������@�@���P/���;��yDhYS��*鰴�#���it�&w��֫�|!��/�/tB�T1���Y݅
9�Y8�����R�Y��C!*IE0J,�X�U�\����Շ�5[�Zx���\�ϊ����3���W=3�Y��ǡS�0x�:}�EN����Xπ/��e�Ō冫��.oy����M��,.��(1O�k\��h���o1n<t.F=�a6r��*�!��ɠ����^8S� ��_U@=��G{c�s���h%S5�/�� �!��R`�*��K��F�͂�d��.�m�.��*#Y<�
���ҿ5g.xT�js�Fo	 u�F�Z��������tCw�z������m3��z�H­��ùp��<5h��}~\�Z��k�������D������4^�ف�|�D���=zkvr��|�Ͽ/�gߕ���g�ף��"O���P�+�	(��H���͑�Z�s��A���s���~ ?�������s~�A�������v���B�Z$�A�xP��}��	���*�c��ǿa�~��u4u�z��=ȴQ貱Lv�'"OB�Je`R����a�=
PW�P�B������U���_�e991���K%�];�Z�}��yR4<��.�{�H�y~z!c��
 ������5�V��+��;H�0ԫ�\�n�۝*!�P?�H���p2|����� �^�<�3�Z���U.�XbZ��u.�E���R��`�����O��sZ�oSY�������b[1b��1ޅּR
ڀ'�q�њ�A���;�v C�RV���F�=�T9����w�W�K��PuN��/�����@�\p�v$�ϝ�_����j�ϔXO��2���H wO�=��xO��x���W� ?�;w�e8P��� B�*�6b^h�-R�a�Ā"�H�8`+%�H�[��rw� [-R���������;�W��:����
��Y���|BOyKep�Ȅ�������*ۢvڶ�,�qDc g����K����{@�PO��q�B��*���h�j*�E�t4Rw�.a!���v�)��7�Î(@�?⚣хK�;|�6�Է��ȆX3��S���#֣aw��_|O~�Ï�g?�D?y!W�8ɦ�ؘ�d���g2�z�8�uuun�fWr�K�Y��<�]�E�J���x��2�\�.<�����hk��a�hn�X�{�2/�Ug�$h��,,X��E�5�젂��G�Mz����t4����*'h<�Q�0�XԣR=����*S�hl^���3�<�ǚ5M���V#�Mm�#��(��f�s��\��i� �� 9�%�/,r��킣�iw��`l J��6�}h������X���jz�x!�yC�c����֒�bC���np�%��s�Z�����8��>� 4��[������$8�A�W79[��Jܠ� �*�GGG4Wp8-=Fc���YΔx�����qW��eoؒa'�9�2�M6�4�U5��O�R�P��:?c�����	+��P�=�� �B'��ܑ��~���M�t�wN�2M2:�������}Eb����ݖꈩ|��g��G?�����lJq||����;������G�u����<8���{<�^䁳+
���Z2�
>|3�l��~<�46��.6-H� ��TJL"P�0#.6���ANy�N����f�7tk�o�ׅ0a\�V�U�)�N��0:R��_���T���I$$A�V�j�/�A@�+�p8�V�5^]{Ҹn$��[C	Q���������0*F�T[K_A�Ѿ�}5кDS�/>���<}��jA��t鹴����@�
:+�����=��3���dy(�<x&AL�v��H�>N����2�����ށ��VO�h�Fk��پ��=I���y���ȇ�Cu=��S���iF-bJ�+kxk�j����O6��ϳs*��*�>�^� 8�,-�,�����}�
�����?����Y��\r�7��He�WcأBF^(�ɞ
t��-^�\S����1QE~�$��������G)���B�l��4�P�V8gm����,�v"�Zn!oQ��A�c6`���B��Wd5n�$N���)S���������'x�v;�"�4����p����SG�"��wz������)9� �1� o��4�騡Q"�:s2���!ju|�/�?<���{�'*ߗ��9���wx��mz��J��a;��j��x�}Q�RGY�.�u�1}���5�xR�ҍu3A�lɅ�5��>���a�l#����f~��
�%�_��d�N�B��k��t��ֺ�9�Ä�Ύj��0�O&�qz<tCY-t˫�ꨬ��+������8�CK�@��bIc݅�Xu�r���kJ��y9;;�sz/E1�\�ڮun��6=�(�(0>���}�]�w�.��h�M�рx���辻�v
�����k���z��:�a⊐����-sztc�[�����]�ĥ�;��g%I픃=e�Uj�݈ � 0��b�s]��ag�kS%Q ���\�#
��|>Ri�Gc�~���dj6��V�He�P�q�S�qƐ^_����k�Һ���f���+_�y腮�G���yR���VSbi���:�����1����<~|(Ϟ���ٍ~�5���0dp\�����<s�+̗�R�*�$�ۺm�J�vu�vzc�F�tO_��v�<���c�%���C��7���
�Ƀzg,X޹�=e���R�R�I�ɰڈ�������1��'E&���\�KPwF��B�oO	
�w�*���L����6���g!�!f0,U,@FS�@��t���<tMM����{�{����*Ck���d���ޞT�F��m����r5��A��ֹ �p�t�DH���D��y�~_�|=cT
�0���L���<�,c���<�(��T�k�4F�����pօ�DG_7U�ȨH�>@�.//��@�ɣ2�����<b^����L:���?ܗ�^?�/=:��a���B�M�"����b�#3Xǁ�+���lT�ˌ���.����
�u� B����ziHf�yH��v�#��� d&�76*A����Sy��m�b�b�����������������ދ/���+[�f^Y��뫉��wnE-�AYAKe�W�kCr��q,�x,l�B?e�����	3cDY�7��@$�i�/O!X�a8:���؞��Y> 
��.�]f,���&�Y9�}`N�rdMR@jovs�^e%�������ⶑ�۠J�=�H���=b�H=Y�~��>�j �\�������;�ɝ�}2��ՙ��>��gOU�]I�.�y����ktP x�������#ꁴ�x�����.�|�V�ٳ��2o+��!�E�<�Y��[�G'�2c�	;�h��D�j�v����}Ĺ_ 1a-D]�����"ȍ��o?!��[-�����i���?!�Gy�;�����$�jtqx`_-��|3��,�ܶZC��Nى&�Xx$�ю�/�j$F2�Hv�|��tN�%�z���Z�b�y��A��8<�����e��sz;#±�q�y��|p��2��g�Y����:�u�ĬI��h�kpL[-lI_�c����3�	"2V`m��a���w�"y��Y�����?�L��@��\B�Mv;=�`Ee~�#S��Kr#r���d<i{�`,��_�~��`�+���_ɋs���`9���PM߈Ӆ�U�~��(����@�B��:?CBC�2�W����:�E"^��J��{[q-w�aOo�x���.����IY��I:Vc�[q5�+�{PR��S��d��Ct`�q8���ֳ�\+�l?8�A���ഡ. j��1C��+U�M�����޿ǟ��gX!�b4������U�_�u�?�g9fD�㱌t�x�"�(O���A`����s�RV�F��~8w�'��Z���Ν�@њ��M�ΰS�	�Íy�{\C��#M̺�W���È�a5�m���� Н��{ܗ�p�>���!��
 L�	�H�.��%�����9M�Α�^���BN�w��߷�X4�������W<�;!PX�	2�}7k�=m>҃0Gmt>-k�^e�C��w;:�]9}x,��N#'��ijS�ES��#%uG'ǲ�����k
�R���T87,EK�]9<��s��oXggi�	��P،h�(��#��Z�8rrsÎT|�<m`�hC�a���L�����j�K�~LBJ��CX����9���;o�[��㞐�D!9�zR�N�f�_O���R^�"Up)��v"�J�ݽ��ە� �p�h7�&h}�o�}��s����)�4��Q[���]�K����z��6 ��@�n��_N�N]_*Y��fJ��*tyt�V���� ���u���`w��Ԧ-�]���	A7�*�}����u��C�HH�Xc��fgzC���%8�ɭ�D�����8>�O`ϖ�D�f*�v.�w���=����%�=4$)���i��L����=%"�
��C/�9h�s@ʱ]t�=�õ�N�e��.��U�u`8p& �[-RB���C�yO�qq�L>�qKm�.�U���G���������7��������������?��?��#�k����=y��`8�''�̿��ݣAh�X��W��Q\�D#p�ei�yX`tI�� ������!��D^@����յ
NV�����	r���P����pº�+Rr,<��[J+����g.O���]j\�����J���򊗺�h ����x��?E��"�%�*3�!<�\����w��/~m_{K���l��/�-�R�հ�5#/�~*7��^����#�{o_(���#y��7T��eN���.s�c*|@r��
~�P �0O?��?�T��Ǭ-���������N�E��R�*������	����Kv2+,�4	�!5�,���;x."�2"f �>��(�e��aA5/$�M�ZW��n��dK�\\� ��e�eg���h�~*V��zz�CU�(ޔַ��F��"�Vԙ9zkp^�+9ZUOs떥 �?��Ss�k���d���15�l��%�����0�_�\���5�Ҝg���gM�#yv�%.�F^�p��	�=����0�3Wn�mc_�o ��S����j+�5��5�|'���:k	#,��C�]�=C�5���!��1��G?���0;F�Lp��h�������6�eR��#���J��������]vw���_z��y+5����bκ�g5��Ũ���Q����Vqw��Jn}���^!���L%	�QSoW���k��ژ*�������I��e�#Ύb!����	-���:An8���H����\W�fR���JLfkŔ�L�k7ʘ��B-`fi_l��<{}R�������م<{��6��6r��P�.�{�7^'���������XM�5RS�� F��U��.���ЛϥaÁ��Wt�txcRKtTH�yr�����ܦ�mI�_�$i���^�i��Lǐ"�nt#>�-�[)��&9v�����U� �)K�SaKJ��eZ �ؒ���ޱ��uƶ���)B��cw[iлS� �H�t�A�p�jv<R����H����쪵p,w��ˮ�b��`Bp�s}3��ɔ��JO���ե|��s���B.Wv�"R�vwU�dlb3�.8^�c�9���(�j�7�o��hV��Ս<}�T��3����C�Q�,�5���Ǜ� ��,��2�֕:0qu-$���;Ǉr��<|x$��ٕ�'�� �h�멳#�u����{�>�9��]U���@���?�7���CZYʚ�Ng�������?�r��ť���P�t��?���U��
��L�+�jU�͍�����/���M��6�J`��do��v����\��J�k�0��݃�*�������()z��JI�x�6U�.]���#�옥�d����m--����ItT����kzT*FY���q'2�Vu#�%x�\籫�x׳��e���w8��TF������RIhV@�$tf�V��n"e�~S݇�ǘ�����k�+��ΈQ荜4�T�8W/�ߨm����R�x�"�I���������������o|��߄�`5}8i��14L��F��BްPA��qS-�>��ک����	ʪ�tc�6B�ؒ�	QP�T����E5,״��4�Bu;Aנ��I�l�[�D��աTaC�Y�ԇ�����|����ID�_�*��d�?n=����H�B)"���~{�[Ci����%�j�n�\�=ac|}����XݎS�|.��3�ɎT����򕯼�����ܻ{��<�2�CJNEBR� ��!ġT�[��"8��+�������@����G�L?~�|JK!hDh�[���21�=b��Ju��!�/dU�g�����p�{0x}����'m3�^�_�3}L�"!�cS�$]���~7W�A���}3�%����=��/q`��gN��U@���5�^��=���T��Z�.��r#g�ܻ�Q�]�&�胱yq�1�g!���}_x��S�%��R�����m0�WwBS��{����>�_xw�X7^��*��7Ί\�^� �5�ے(�=I��-�Ym3�Ee3��Adk�sts9Up0�ga�zaQ��0��]��\&
p盅Ȼ����\r%�w�.V����k���G���-z�aԿ��O���a[!�<���9"vnEU��6� ���[_���i:V��D�����Z�HS��D����o�j��訤M>�=\8���@��am���{J;���ue)���oP�����L����-�`H�AxT��'3���g�z��dz���o�����Ηy���ё��^XN���G*V+�8
Z�QFs�9%�e]lv�c�P9_���<��e0��ԝh�"˓�kN��b����aj;�^����Ǩ�+��3XK�>�58�ut�@�@t]]�X��k�8Dy
���[fu+��]s�������%��5[(�5�\R2���sU�;m��#��0�wQ�iب��wQ/��������fS��ק̨�wgOVҒ��O���c��v�@@�ϘXZD5L�Fw�=������x�N_u����,/���[�b������n�@�藄ŵ����k������C��y��ϥ|�'�{*���;�d���;��'�\f�D�r��u�v����#e��_~(�=���.�(�Cq����k�����N��DV���Gr��P~���������̂��l��������FN�g�/o��dI�\���x:����-��Lc�.��/4m�*�k4�~��0.0���ZT��J�^>qy�q�7"���K6�-;��q������"�'c98��N��d�y�����(��˗��Ł�O�}�qc[�}C�y�M�N��:�`}uh^�Y�9���D�G�����I�+�~n���&�1�N,��9�E���S*��`�L��<;=4��	��C0<���VX���
�GU�<)�Ś3���5�u����=#U�<5�3�9�l�vGo��^^Po�{K�}��x�`���'Z��G?��'�7����ۇ<�J~���W��'��`����\���c#��E�%�M�D�:q�#uֵ:d ��v�,�@�8�a�Q�7��q���){ބF66��cA'�dz�46-�y����80�H)"�3�V�#��オ�B4��͹����
��*�aغ�Fh�KC?z'�{�=���NQ�z��hދ�_Q#�3X��ѽ�GY�do�1!Wm�������G�+����X__e�-`mXZ�k����i�������ZN�T��)�{�Np`6���}�|��g���S9�?fʝp��\���Ag�,y��B��J�VHՍd�pƟ�"�������E�^%
��	�3�}Tb��&y@��DL��UE�unp��N;�3B\��j7�j|���̏���G~���Fb�I��i�ε[r'(��M�9,lk��$���@���k��f  h��6��`_�^��`C1,R��qtt&�)���V�/Ϛ��n�C���"1�"�'8:�:���p���^�[����5n�M�<Qh�R7��~�=!.�5�=�{G����� �%d?5���æ���(�K�E�eǋ0~����8<��o����[a��rg{C~t�����eo�PN�jt.�jf�Ũ(kh3g����jr�"$���N�߮r<.��e��&�!�9���V��HuGq��.2%�5�16���I�ъ�@��sQ6����e?e֎��xd�9�<����y���<{�P�����$8���[o����v�7w����á��D��Aw ���4bZ��f�G�1Q�ś,1c^���ݮ�Tz�0v�� +�UŬ]t��W���>�{Ik�ד�t�����b�M��}_���>��N�<g����j/}f���e��q��4Wws�^�c��{���ʕB�R�Ǟ4�����Q,�H��T!Ȭ�AK�Y�MA��ƹv2/2>��6kکsL��p����dA���e4o1b?�,�Q�ƞ�f�t����x����F�ȣ�#ۀ&/a}����Da���9DeT$�)�>t��Oh�*wF�
Jjd��ܠN	��ȗ�E�G�^I�/���[[��#3F�i��+��#�`�8�U�ũ��e��+��}WV�����0<�
���N�c��9�{AF��Y.�'����dw��Ίl�A7�f�u?`0-�sy�d_���rp��4�n*o߿!�7���[����0��Y�3G��3�my����Gw�����y�L\%W	N�D랰�����~RkT]m�4�Q��E-p��f�Y����2��2�#�%j��5��@1����Yo8Յ�D���Z�Yk���.fZK���iE8���b�*/��ɬ�H�Q4{�x��F&�iT �
���~���w����qX]][�������o���cp>����<Z�R��D���&Vu�ӂ5�H�e�,�oT�Df*0_`�aC��.x�K������M�Y'cQ*�.���5�V�fT����}{[ej\E��5̜R�"��L*��+���8K�#��WU����oԝ5�U<Ot<J�꩓3R�6�\�۹¸P��0d��(��(�*���0��q}C�������"���M�V��4��n���w�w��)�)���~@h�����lmn�d]���gŗr|<��.����1:=���:�77V���|4�yY{`o�+o}��2v����"��S�[���P�s��K�^���?Hzv/�Y�3Y$��A�	���r�k&?e��B0�L�%a.�r���H�V�Xx��'��ߖw޹/����X��5�oSЂ��d`��>�Q[E���)��yY�X�P|���|������w�LȆ|���2���2V��v?ܭ�M�N�W��^j���5�X�x��k�B��]e��ٰy���aʒ '���:[�:ͱ˺��4�x��m@ޔ;ש�Y,Ʋ��%[ׯ�6w��T=9������Ͽ`�
�:�������p��,������wߔ��޹<y�'��X�OjH5�Z�����0_(�Ι,�Ϟ`hR,4��t\�ԯ��&m�z0%��~���ޱf�qn� ������l��.��N�Ǽ��hN�0 ����*�|r0d�~�@N�v��q"�Q~;Ȳ��o���v�+k$S�#�{�Xϱ�}�r�UŦ�i����8p�(9���
2�!���k�BuD��ni�h�x_ԆX�22���L�y��Zݹ���I��龓���-�,ǽ૵@��(w�Yi��Ԏ�������n�Yz��򬻨t���\P��c?�`/,�2MiX�����%KR���r?#��q���ϗ�	�Z�w�'��Q���{
�O9���@�O�o�N����De
�����:q`G4�s:89��A���AP�Y��D���ӂ�q��{T��h�����G��.�9��$8J=���N>x{+���fd�`Mex~~N��QV=0Va_�ܕG_e��My{kM֯w��s��J1&5���q�ЉPiGY���n�+�w{S����C���~
wq�Nő��>c5������>�ѻ���ߑ�;���;���y�셜��=���ޞ<|�@ֶ�r��2��d{{���BAí椢
����d{w���;�`��~�j3a�a�ú*|O����		-�����>�Sgfe��t��"����P�C��O�Ԝ}�T�eV�k�w{a��T�PJČ&��E�!8�Rx��aM�T	Zy�='euue������۷�_������+?��BS%�q����Yܵ��K��oi�?����A�77�Q�3�"8tc�=?��I�o�3���y �#�xܕ1�*%l��Tlc�a�A[Sl��).�b��F�i��-�ᘙ`4�� MA[�������8^(�uK�V{!�j_�Bq��ě��l����|Շ ��[=�e�u�S�ظ��!?��]������x��ܻw�LJ�
#�"�1�𺧋�;M�G̱�P���۷	����;7n���w��X=z��)1���|:���36W��ਆ��`Ͷ9����)
�f�U�@r��5*Z�jUb^�|��P-�L��ԣ{��,���T���tꬡ�eץ�0P��r���1�e�S�#0�L�'�rtr$�k}f�Px�]�Q��������w˚�2c�G���%Ǡ�<}�0��t�+d����b�NG����Sy�䛠p�0����f3쫱G^�ɑ�3��I^_2Jj����W�ڇ����ې��q�.�P<�\��˪w+��'۝p �	��:M,�5@>XpoG����7a�ACŻi�L6��$�?�����O���o��/>&�d��,��sY�蛧ҟ��z/��~�pś׶d'8�/�ĵ��O,\A�]�+����Ph�eC���Y�5�����ׯЫ��\�	��$Sj�e�
�������O�4Mgd�++Y�@I0r�[���Y�� 6���V;��;��~!������3���țoݓ����C4C#����Jc�ў'Qe�^�`6ʀj�*���2�efD�Z4nYl�c*�_r��b��Ȣ�s�����ln����R���h�����W��R��)H�B&�֫�^_�D���(:�.�ϸ������֭\�eV��l���E�mx�vF��F�X��NBZf��$&@[� ��CrRڲ��|���FCG�5�~��2�!#���o|.36�k���D���e�����D���u�Ψ�Ї!�<���m�h:��� Wc���4R�80=�_��9>
�z~x�y[L31�{<�YѲmޖ��$���&�*���ZKN���-Z�ϳ�|tِ�N��b�Z�,�j� e{��$��Pn�X�}xG��:�N��4<�dt!g'������`/�c���g�	�/�z���{r#8;�n����ƍ������b)迡�ؓ��8费l=���*�gcy���<~�(ȁs���r��^Қ����`m�[Hc�8I�9J�� ��@�A�N��zi��tC�)��	Y�
k�����A��y��HYG���%)+�A^���H��#���S��2`��a�k}&�H���o�Mu��_J��,l��p����7g�P~ࣅ��:k���7� ��N���`C9uFȜ!�mwt����z8G�*�#��Bc
*��Q߁�	`W�����j{��m���}ff1�&ll�E^F��9E���F�������.1��)�_��/i�W>^[�)lF�|�K�F�)yu��juœ�}e�����: ����
����zW�������_�T��ڑ��x0:X�c�G�Pʗ��/�w���t���;'0�����s8/�B�_��p��?�f�Nd��"�%t�xM%/�U�]ެF�=&+l#�P��7G6�D0@��hU�U�����5 �:�<7�ޙ�;�Qʵ3w��),����|<���� �H�)(Z�-E{||L�&[.��=���څ����q��P�v���_[놱�A�uq>b�gD`H7�N��|����پ-���A!/���4���d2>��D&LWs�-�j��:sҫ�ߤw�@��)Q��U�����}�\�+�:8u�?�|�6vA� �+�ĕ��lo������S�Q���O�q,wI��b?`�σ"^^�H���p���?|y(ߌ��ɝMyy���Knݺ&7o�����D��u%�`>H
k���S�2R�[���5C���H�\����}/�y$�v�2�{��3�Ι5�WrQ��Pr��;y�XÙ�����V���H���3��?���ꗿ������Z�.���8/.�q�5":9�Z�Y���S1��7�z�wy�1�hc��t���.�`�,%�Gٝ�5eRɲ�͍fub#V��rƲ��s"��siO����Q�Hu`�˒T�^f}u%+М��[2��9���i�][�WC�EK�Q1����Qݧ���q[$���T�)�^@K��P�����$�-�I�9M�7�Y�p���ss:�T1Ͻ��d�0�Iٖ���&�ȴC�)]�PN볋1�kT��Ђ��ֹv�ؒ@�R�ʕ�>��Y/����Gv_sR��i�N�f���["�np0��1���)tK'薾w�
�O?ߐ�l��ҎL��2���6
��{05�Â�>:~�1�T��t��F�>N�F^�e����s|Y��%�/@���z�%�5ws�:޺�#oݾ!��͍�\���ݻ���dҽ��˳'O��������"����|W��c6�����,h�N�#��J�U���ߵ �܉�z�9������Y:�c9z�t�r{��$��C��D&���V��G��~ƙ-mo�EVW��TI{[	�4��}SQ��l��$�6�ã�`s�{{�:�M�J���w�omoo�����Gk1�~0������|��O�bռ�,*����L2�.yV�j��Khu%��R��,:u���b��]=:�Q7'30���P��h��!ZC#(���U�n�4���z���y/�=Y����B���I��#��i�L����Q{�a4���!��Fg{iY�7փ0X����)?��˻�ň<k�Y(]� �j��HV���1����@��r��7A���EJY0��f6�����̓'�_&�A�L��_Zc�'	��G$S�C�Un1��?�`���x�G�r9Ia��~}m�"]o|W;�."h3M���˂]n�Jy	
ϥ��M�AI�5>��<3PX��@��h��Ɉ�ҋ�M��!?<��������~��-5�no���W(�r�.\]��R��O
%4�vm��Ǔ�4��ݚgd�����������?�����U���k��ڨ�Rˤ$��fXņ���Q������M5���)�J��Xc�ڳ����͠`_��yyu���# H0�zc�WZr}gS?>b��^	ktUfgO���d��s:���X���0��Avv2HA5����E �j�a+FGc��<�C\߷���	�|��}r�sY�G����� �y���UH��&U�K9��<8/��ȓ�ʯ�k��_�R~��_˛o�g9����7	C<�zsk[{e�4��Q�& �W#�`a����z� Xn�=Q���s¤�(�*0:;�.u���dh�ue�V�0�Rx+��	d 
�\R/����%�)fdF��2��9���ҲdTfHuh��]l��P��>��n�/�pW�E�dk�Y�׸�k�l|��m�٤�X��$75/I]j6Fak��(B����T3�F/LB	`k�MA�,�p
\pBvLA{ ��BƗy��@��1b�$�2#8dc�RW"�b0���#8���=�$`	{}>�	L�@��˲��s�|�K�k_��A�_5�=�b�
�[�u^=M"gǳ����9֬-u֤��88� l�"���oK��9�� ��G�֥li �k����Y�?������k��h
�g<n�����'
�C
�!��7�esu��]���~);ח��{���l,G�GrvqB����p�a��� IJ�j2�;�T��Fs暈iH���oU0��W�\�e��ь�*�d��S���,zF-�6R�h�!�Wh��E�<k��q��z�sk��'��:�?�#��f�
�b�JQ��{g�������Blp桻A�y�������~���?��?��\W���hA��׾0� K����iS����d�,��.9ٹE��]8pfaC��� �Y�`�[�#_52�KGS3�����i��]Ί����oq�96:����<�u#Rj�Ԯ�%
�;���Yf��۽^�盫��P����+>��/�a��C��R1�k�ݸ�K�]~��{�ט �c����#��w����sc�rt�P���bT�rB������۽� �A0� ��y�����?�ׂ"��u���9�Q̅�.p�;4{��Dfze�Q Z���&�xN���7�	��f�Y|]9DǤ9���0�¤n��s���8.-��)�Ð�x��yp@�Q�ʂ��Z�et>?a�x�#�.�C���a3�{F������/5[��60�tI���34'��V�>=d
v�P�Ie��ݻ
[$fy����D�Ime��*�k��A�j��W߼z�\N��t��Ai�z�}2�f�ڙ7���XOvxx�L�d2����f
�4�(z�Q��D�6�.�����lL� �w
�׳Sm��0��I�\7(�1�D�ZF$Qn�uv��+>��L�W^�9�������g�3�����T���2�F�L-�t$8I�Ow������b$O�=�Ǐ����Cy��K�ͯ~#�<��8�<싋�X�,0�=3���:�Y��P
9UX3����)D˅D,-�ABUQ'����@�I�&-&���O��G:r�8%�לE�jX�X���`��wD0�5����=��w�.��x���mueU������r��T�g̴�m��㰟I$�i�y֓¸�|<?�o1���v5�_(z z��0t�6 F��N��ճ�!Ң����z��:(�Qw��[u8���v����@@ɬ{l���{M*�\T�Aa��~ClS�g�X��.���`�M�W�A.�o���m9>����.��\� � 2�kۓ�	��b��� �QfЌ>/)Ӂ�3���wW�榯���{�D�#W:X-�	F8:}w�p�T��9��m)�oy	=q@�����<���^��������ځ$d1�����@�a+�@*�
���=�L����t�~���j��&H\ ��w�ݒ͕�l���"؀�\�\������}��)�2
�wxz.��������Gq�,�����6�+��b�P$f�b�fW�J�8��>�DWJ����-nI�^۵e1
k�����S4<�H7��������t��Xg��[a�H{��|Č'�h��r�f�wӠ͆^(���T�.�0Me��P��ĢEv64ΉDa��5ȗŏ��?���ޖ���т �����BJ�0��A����p<�v��T�82K�h�E#��(,�>�m�'CO�A�^c�"F�i+yd<0�X`��@]�5��H?�bD��{�_7j`�&�K��(Gsn��P�p�R)�
�p���S��W��S�UT>�W�����@"�Ht@ ��\;�͝y������oH�'f�|t8�Z�d�;O9	�(I`VE�WC>}�n���y�x��IPg2?q��Y^P��Ձ�@+���_�a$��(�����N#Y$>�_4�_�wt>���5o8"�p��Z��#�0�\�	fp��ߘ�^G��3Ԟ���P����e'�E�B(���x�(�6���22WgmFcC���5�M�|�ŗ�駟�o�;��Jp�n�l���5y�������"��{�4�Q$Bc��cA~t༕*]���ו���_��)���|A⚬��*����s�z����A�T�G{r��-��g02˹��\���W@W=+�<Wk�#�==vOv4�Ά�a��K�������򋮼-ݙQ���`�)����q��x)�����G��r�$k��U�5`�j��kͅ[��v?8�/_���ٙ<����+U��rO�ΏE�K�5�>�:�)� �L�-���f�g�9ur&O��`A;�0��`���=:x#HGD;R�n[����;�0��a�C�B���l��[R��Z]{t`����ʸ����L%�P�@�2n��zHPh♵��AE:Z�d�1�n�p@��K�����h�g�gā�k�(��lmm90���}6]��[����9aY|-�/��;X,ѿ�Q+o%�`:���n9ͬh��lH�7�-���Dtk�R30h��`n0&�@��tt.S4��{�a���3���Pr�\�Y����0�SY�l��r[.�%^�(O�L�e�X� g�<��n&�
R�f��)�[��5�U��B�7b�{=���I ����9	���2��D���i��tA�3SV(�f�0����{dN�9Lǒ�d����[z���Yrd�[^������$lֶK��!2�v��$�-�N��%f�Zpd�\�������ݷ��X߈DK�@޹�.Ƿ�roﺼ����ݾ��}	�	�hS��7�U�y��H����"�D�P1����\��f>�L#���#��9�����g�(^ޤ�H���
:�k��U$Z`-to�*ǅ�F����Θ;�&�N��:��0S�2�G��>`q��U�4A6�vvn�1�|��SyN	!��6(n
��h�$;�b�!"@|�c=Hf��-�	�X�6�n�X� Ƣ�
N�u<{D �9�n��nX�zD5���>���}Lٱ��)V8Jx��v!%�4������GC�M�l^W����W8�ô��2��)˴D!y_����}��q�[�4O���׷����k,6G!w�ԨBt-3<bReY�R��t�z��R�U��qe�6��<�C�Ν��޻������QPl{2A�r>�O��-�ts�+�D��������H��������]×L�_�b.9�U������o��xx!Axͧ�ރ��_�2A�n�E��/DO���/�	8�qS���t��`�#��V3f;�CO�6/s��|��!��q�}#�?�������̓o�G~��uy����'l�u��%a��Uc[�p�G#�Qrqn}mh*��X�i�|s����w��}}�&������[�mw��E�T�_�CL;��뼳�ݽ.(ZgZ�;�������`mj�< ����`�a�sz�e)����&�щL�6����ږ�]��^}��9�c|��w��٫�T�_�1_���:*I7~�_z�)Zm2j2��z*��O�œG�d�[�����E0P��B��c���Xh�`��;d��&d&�MG���s���(�}�epj�H؀n�X�c]+`�a!3��X���e"�����k��aF��w��ă �[�����аV��p}A�"������<0��"d(�N䪗��`]o���0F����;��$�������i�Av�^�,@W�	jw�C�H��^
N�+gg�t<4��Y8���2
4�h�:<;�|`�@e��{��RA������{��������̠3=��������T3R+K+t�0'�'\R˫�ҁ����vj�����<8Up��>,�d����"��r�¢7e������m$�J�nAM�eTC>�tn��Xw�Fb���x%J�S=����� : Mf�20��������Oek��9�ݳ�'s����r��]Ƭ�}�;��Ƭ��2 3Nq���=l�1FX�
���-Y	�V �X��y�mP^oǲKH�d3�n�-ks�-;�7���m��|S�?�6��1a���}�S8�O���Pt� %�'I�]6S]�%�o��ɬp�V��`�4���`}e�'~sY{�`V3c|K�ZA����,A�{�(u�dYd�T�&��@#Af�'j�'J$^/��]й��2�� �Ap�	m��&-��������n߽{�֓'O��t�H{�4r����v8/�e�냶��N�1�+��\V�+
]dG���`�z�fr":�Ll����9�l�[J���h�(�S��h�A�P�}N-�D��S�L3&��k͐t.SC`6����	��0/81^�����*j0v?M��#z"�\��5CX�s,�vJ�aS�L�om���Y'X�]x
D4��i�D��Ն$^&�d*6Ed�P�GH�\h�0���s_��/&Ϟ���yXK�Pj�[� ��)â�ke�הw��]�ѥ����9z'���R�?}�
_�U��y�	����GH)�E9+�� `f��ҀS����{s�B
(���R�6hu�k�;�ǋ��|��?a��
5�˽�}y��������0�"�[�����zܓ-�"�e8]����1kk���%�o���o76�忛�vRS��%n: ���m֊Y5)�k��������1���������@��7�ړ�E�қrz<y�V1����{89E���e��8g�3P��bfk�+~9�G�z�K���c���D�Tݟ�����q'�p�e�Kv�\�Nb���k&F�`F ��m0�'anԑ�Q�vGͦ+tYQ�=��0��� %�����y���|��g�_����W_~Cx$�3j&}r�!�>BS��M�w�b氯�(৕+]/� 0�����|���;}�`T�7�W��F�g#��zS@�BG�'���� �/����}:%0�!;u�a�oR���b6aP1y�����pGP~=��*m=�+ � ��A9X��@ˍL������#�#oi 1)i�0S1ss���g�{+�	���^w��?ٴ6�:�"0qg��6:���?`Ĺ$T|�����CP���&�(�������{عq�rm)�d!�cey+���=6tM�l<<b�k��-�[`���YL��tNEC8��p��$��NrluQ48#�jdBI>�� ���ԷQ�M��e�A��܂58��t�(:#�! ������@޻Sn쬳9�����̃��"�on��W�|�Ă,����J�&z�L{��������t��p���
e%��<{��w��#�w/�g�E�ga~��	{I{��:�IV��}y]�>_���<8���s�5̀�X��B�7 3�n8Z��`��%Ic�K%]��FS1�0��zs��Eƞ#�ޡ^2�V�Kn=A2�Q=0���d�.�jR���f�,c��eiB�������w}�����1J
��FD=g��gEp��y��g����u��!�O������O~����_���S~�;L_�ۣ7�ߠ'O&�X��C��"�9��,�*)x�Tt�*�T���Dvi�I�d���?��!�=�l�1�ʺ���H�f
87:�*���9�w.�v%��;�&
����{�\d��K!��*�Pa2]�J�1z��I���"�΀5��Ks��a?�~�:5\͈��&�>�#݊����%#��Z4�h}uY6֖dk}�x[8y�1:��������6.�$��oD�����u�����
blp����{��7��%��4���Xѣ�q6��)���͆�Q�a���Zi*��ו�x�B�sQh�MJ�@,�d�>���˂T�!��H���0$@;��}X�ax}�ױo2ץ"G����39>:���C�G�`�1�L��/eoo��v��m�-��(v����b[j>x�5�`|���}����������O�s.�u�U����K��O�hl700R������T(������3ψzh]ߺ+��֯�){��F��A���k�K�����~cS�8"Eh!4)�)U�B^]r���q�r�J	�nM���5�l�+���_��o���L|�ì�-��b}A�����(�f������3k2��!�|tt���y�-+$G��ӡ��/�k����A���AK�į˴��XZZ6�ゆ�jD;��&����|\��
�� ���?<G��dB6I�+8���ẇ�#�^�G�|��Kh.��.������� Ԋ���O��µ�%�/��u�B�$2����(t,�K����Ny�x�� [�.��9}��}�[0��>z=͠F����|�9�b?1���g�
Y�P		+4+�1��A�$�0-7�ᾰG�hb�-;��?��Bp���>��@f�ןLp�p=�1��C)A+��Ko�D96�����
���/��
r�-K��9D_,V�*���:dHum*�@�9'��p��\��H���ގ��;|�}�5zv��>2�jE�̼����f̍U,\�����5���g��o�ɹ��!#T}����߹gu p�f�O� dX�gh�$
\��1??;�q;	��N�ƅ:"B�fC�G��oߑ���:ϟ��YX��n��F��A�ws�\�������ٔ��a���!�}�!�\�J�D�<3dT)�QS�0fj6�K��׋����=����:3�:�-�)~%�1��Ca��3�Ŧ�*��0? ��r�p�K�1V!h'�S^0�Q���^[_[�-��I �s��5$-Ƥ��8Nw�]����AԤ���΍n���!�8Z���ɶ�
�L�`��Z�Ԯb��aZLłr�e�.ʐ�V�0��K��E@�ȃ��C¨����4���c6��3�̈��{[�a�9�-��/>��u�u,z��G4�t�0l.A�F��.e1^w�j�'�U󠤑�Eԋ��!Ć��Y��Rֻ b]7Y�P\�5lb2��Aū�����Z1���b��R/(���<bOC�����K���\sC%��;͡��*žJx�=��r_�x�������O��q:r�9[(T��l��X�^f�16#ri�kϝ�8E/b%y���&ϒce����z��2�c2��Y�<������X�N/2RTpO�>� Xܷ��#��K�4`�S:�A����<�������<�ܰ�9���ޒur�eye�?p<`����8��䅥�*C3
[_�h��Vak��q5�\t'Eܟ�o/��gK��Cm^����fԬ�Pn�z��.���(X3�Fi�W�<(����6���,�O!�*L��1P�ZP$�q�O�$w��G�Q����Ԑ�ȣ��ٕ��=�ֽ�4�����\Wdx+�)��~���NiW��?���e�À�S�(�ۢ��mw��8�s��ia02�� ���pt�U19D ����L~��7���}"���o��/�F������x��U���Z`�\̈
��0�C��{-x���9L�<�<�Й-�F��H䢬~��E��8�����e%rf^� 燬$�����{hK��j��1ӂf��w�.Y#�yrȩ���Y�0���ǌ��IA�^O(�`����Dy� ņS�+�ǆ~�9in1'�7��AG)��C�ZE= !�h�Bƴ��vվDS`�as�����p�])\�dX�Yc6d�[��F@�P�
�#�J;ڦ�S��?V��0��jc����Q����
�C;�H{QXQ�ѵG:Ug�H�(�1/�"4�Aj���<�k6OӮ��	�BJ�]Т~���@��̄� [���&˽����Y�]2�@�G.�ol��
�x��eAR����a/��lT�ǣ <.�e@�&��)�*Z�V��d^��+���oʵ�rzx,_~���x"�w#��*[}�B	�;м�֭5���)�w�d���$_X�?OK�B�@����[L/��8��ᕎ��-m�Zg�P7��Z1.�c/L 3נk�'̪~u���։�Eq8~��k��Rf`!ˎ@����gP�<YY�)c�ߗ���z��A�`N���LY y�����1�����_~!?��j�ae!�|�(�Fd:T���1*H�8�� j��<,����dF�+�A�� R��+������G�5f=�����`ڐi&S��zUx+��Z���)b�[�-]���}N/8�w��U�7uV�+���@�Hu�,{T�Y¢q>)��y�W�Ol����.�s8�~�Ez�����В�|�u(V2��l�Z��Ü��hR�W��@���6\���61�ͨx����m��L��%�E��R�����)o��ُo�}��1�����v��LI����XXM�z��K��QLC4��|���*#-���s�[Iaԟپ鵶��si1�Υ�ӄ�b��ܩ��ڀ��������͠D�,(��x��})�~�mP$+am_'Lnum��m	Q�3�-�}*��xH�6�v8�Xd]�5�nn_�3#����ꈖj�a�2_��a�X�P;g��7X\��y�y�����F�eW�/�{�U�\�'��X|4r]¤〳���s���/(�n��	�{��:�lʊ���"��㰿�� r��q%�Q��exq*�~&à��Vd6��ÂE�.Y$�jܪ'iF��u�}o��Թd�h.Ԩ�j'�R�|�dߑºr�\=�x�1���kr!16��Ei��g :g����~�x���<�%!r�7y7��YX��Ů�����/���uX��yHg�"�T�6�FU�3�`FY�Jw�t���¹@'uF�M�ĢRw�3�֢�Yx��o�U�-,:�#���`�:���`�"8�����9�Qt���"i��(ůQқ������$h��LY����z�̵�E۲�YwŢ������x��'�8m�
=WQ��WJY�SA6�@=��N/��p��Յ��8S�u7@;�a#�#�M�it��CP��l����ǥks f̆�]L���E%�PF#8�v`�R�ޒ�qGj��x��-3��&�M������+��'�B���3e)��8� �O���lb����F��Z��B�N�i�B�,-�s�:�`8-�=���Ԧ���ކ�`X�1)��'����g�E���_X�n��Y�«�S������7�o?���cy���ܾ{O�6�=�%�I��u�ƺ<��%wv��W�zx1>�� ���A``��GLz��%�qU��I��OT,���7���'{%�P+2&�=��ұ�ht�lȌ,r�8�(�oe=�l2�((����Ŏf#�3��Pߊ�!��+OLg�Wep~��3�'�Bl�6+���b��� �F�L@�{���i������Z_��������S0
��<�"\<m�ֆ�¢L��PE��q0S2Sj^l0,,P����1[&�V��,Z��30���4�l
Ϯ�޺Hg���ʴ���NKk����i�2�W$���Ҫz����>�|�����7���z=z�ӏʺ*����+Gf�~���+�
-��|T�i*��(�M.h "2����i����l�\N4�4�_*��g\#2��oXZ@��]y��{r�7�p�-G���b�c@�W΃Ԇ�밣��$uu��W��hN�T�bfJ�GY9���N����'C�Nd���T��F�XSƼ�("��~+�07g:�`"�̩P����p_���k�{�F>m�v}�{
u[��{��kS�Ö~�|�cF,5b[����a+�6�\YYeA5�?1����HLf�6g�?sq�2.���jkBߪ�A��Ң����5����IT�
K���v�NlF�
���w���͍u�~}���Ҁ�P�2���;��Q�z�4. �Z��;P��d{kM��iE�?����ʠ�e��;��i�0�(�Q�ֳ���ҭ����I&��|}�]5�0MEm�Uu_"Z�t���h�e�P��y�IZ]]Fʪll\�1˒���a A
ԃ#��{�:�O?�\~��O�7��X^>��~�}�(*zK�¹�VA�޶&�e��$�Ь�q�PYo7����K"��$ə1�Q
�&�z���"fQc�x�� # �8�WvHRo�jt�\��*�#��v�N�/�Y*AF����s��4N�"6\�m���Tu\����Q�#�(�"����K�9���ե��]��XPÞי�1[�D���]����#6I,�u̻�ܘ���uo��3�jC�p�D�:�m:_%)�v�oeE��d�k�QE]LD4c�y,6.1�Im���)|rtI  �4���h,�U�I ��\� ��C�<|�08�Oeo�s���m/�4?���7���]:�.+8��t����N>�e7؇��j�w��hν	ĉBg�4hi�
�S�E؎3������}���w��P<}*Ӌ�|��ײ��C������h B(��Ƚ�;�ͣ5y����0�a���0�H�wB�JB�0�FCܐ?:^������Z��Rt��Cb3N����4������
��ح7�!B�]$��� ��sf��[�P�Ʉ���E`��,9Mh�����`F�wvEɴ9flm�vvA�>�z��
�1�n=ٛ#��_��_|�����h�dB�`SA��e��Դ7)�b��	�����i��R���Ū/�\��lI�S�}�����n�rN6&���W�n�<-,5�-�:��ȉW����#R�/��p��,����,�	�QFOՈ�Sx�I�u�E~+#ӻ(��"~ĩr�ڕէ,�I[+)�&I��m�*��^�47R���B�r���5��`�ٝ�[|�i+�j��2�����=�#AZ�'�G$�c�t�s
�767dk{K����0:ku�
�Č��v^s�l��������~�tJ���ߵHV2�l�G��]z|�[jz]�б�w�y���|��������>�ٓ��0u�/F8J��Ě><8����4�
|9��������0!v��a�ږ��p"ӌ�g����������=�QXB�)�Y����.E�/-�+�j��2�k
#f��O=�6Ǜ�lvD���`[��<<g�Ө899%,�����T�hF���	�������y�o�!���O�0��������Ѥ��׃�s�e=�}����]�V[����һ����o��n� _����s��t%���{��@=���Y_9W?S�Su��9�PC���\���[d�;d��[����P�a|O��H��l(���O��g��{@��n��vU��\{{ �ӲL��
Ec���  �j|�7:���O���3��T��S��ēTWe]K�<�^7�����!<�J�D)Kj[I��F۩�5g��qR�R��y�_ḁ9͘��Nϳ	�ם-�̩¬ud���� 6���%�T]��5�s/�ꛎ
?���љRy�E�z���ɒ[d�N�@�bYW��E��o1-�)���l���W0��LH'0�]��BJa�N��N�.���:��(ҨOt�?����ԵF$�]Y����"8���_Ldi���%ϓ�cy��\���'�٧߆��(����fr�ލ�/�dekY��W�t9l.�ςwN Ϗ{`�È��!<3L�hjp^����{^޽��l��zi$��|qp��I+|�����͛��ñ��ɋp��oߓ/<�a���l$k��T�m�~��\4�D�m��*�jo:=��y.F;A�_�jv:O{�d��l��>E�k.�s��RV6�XA�(��̒�-�AA@d2�i�.�v�KH�`����^|&�n�뺋�j�؀z~mmU���k&��O��w��%e6ʿ���z� ����Qg{D}��G�������`QnA��Q��E3$q@YC2C��L�	)���(��\��Z�#:U*V0֑�f��k��B�&h#ŝvn-��%�#DΑj��M�����͘����?&�R���P�����"�ޢ��-&����F#�ti߯|����cO
Qa[0 j@�|r2���w*�X#b�R��@!3�%�L��/x��T�8�+àr<LQ���j���h�M̺�7��ƢnD�� �>߾�E֕��Uy�wDJM���0L�{��.��F�M�]d�l���K���B�3�r�̡qƸ#���`��~���B#��r��~���u�g~"�݅��a�v%�!{y��ԷP�P,�|�+K�`�Z�� g�n2>�qp�f�!�����g�UE�9D��ܿm��`�:�1;d�m)"a����d���5粙qx���G����o�����9j��뗶b�&`���S>�kg�!^2��B� ���zA�8��U`�ʴ1!�$��#3��/��CC��p��G�Q{ȍ�xyP/ϴ�k����w�QsD�K����(��C���Ԋ7S�x���B}�|z�q��F��_RY���}��p�lc�3�v[*����i ��0�X4#{�����]p<~������\�ᇉ�=E⒬!��Yp�^�R���g���N��i�!
H�HG����yl}'��6.���̄���<��i��R����>�s��e'Ču<�6��+3K.J��?C�	����[�2B/� ��!��ߡ�(��<�`f��戱����IuJ[�����Nҳ�Sr!�Zӑ:Y�>i�����嬶.k���!�fiG?d*a��}v	�l�P�t�l�����>9����5�<�+���h[H-�U�$��h@����.����.Y����)��!����BΆ����npD�2�#�ǎ��`��7k2�؜����04W�dy�HzIZ�Ǡ��Yǜ�R���1���ڔY�v?������G$���Ќ�w<�?�k��;o23�������q�G��W�<=	�x{��N��<�"6�e<�K|���VM�Tv�kȲ�^
���b�Y2�C�F����#�ֶ�\d��'���p�T���6[P�����%֖Awg֤��*�E�T�0��`�,BvN�C�d�Z��"d
�Qc���Q�(e��.�<��ۯ��׿���=p�O2���i ��`�@A
�r�V��^O�]��ȀR���ln���C,
R����b��R`o'�b�����L�N1�	7i�E�D���B)~�'���N�-������z˃��A02]����%�`XÓ&x�2y��*L����^��Q������D�C�m��=ϛ�����;F�*�c�L�S����J�[���oZ�R�M#ςp��䓏?��~�����]�X]Qc�Õ��̌�
�n&�z��?�vN4~�����*5n�u8X^����`��/�Yh9�sRL�n��u�z�kQ����MAb�*B�rR�)�*�@����k�DRQC���R��<����x�a\�F��,"�D�a�n�������l�\#�.
�a���� 	�	2{�cb��b�}F,4;<<�����a���M����+M��g�\���&l6�B}H����.�65�G��*G������.���Qm��N�Z�5�"�!W�Ci/��~���ix0� �HhI��Y�);a�؟h*���@���dO.*݇.[0�N��2��#;�%���k�T�#p��wA"�sȳ�RV:Ut���%X���pD�52}J�i�J1�����J�jB����|-���צP�Fd|��2F�k/K}EDyh�Qh ����`163F��7�p��?��M�p�O�<e�G�	ĐA4��-B�Rc/�)�%h�4�]��m[�I�Y�T�ĤX��Z�U�Q�	�Ojtc<j��l$`�*����i�זA�؍]��ަ���>\eK�u�j����yt;f� ƾ6�q�|�9% �ps�Y�2����GiNR�=&����V�e	xK;u�ँ�-��T$	˱�%�kd~�Fg�X���&!j�%���YfR���,{��M����
J]��&��T;=�3G0U�����n�5�´2@���lg���~�lB�M\ c����Q�{�Ŝ��^H?���1��Q�:�f0�x�1 ",�u�C������_�����	��GVV{��ڗ>xO޺��r����d�HΧ�������(��C�⫧r�Ύlm.cٳ�z�ܻ}S�_<�^��y��5�=Y�N� p�L�m�@+��?�-����2�n���{5��5��M9�f0#˺d���P�WX�eR�k;Cq����5�˧Z� �2W @�0��v��h�k��:� ����."1��ߠ�n[YYa�����������#�G��p4�Ů�a�F����]�͢�caXEDdM������C1�����!��+��kY�Egi>pcpT?(��'�'�o��9�I��P;�^�9�MVfsq0�V�H׆�}ɗ6��q^N�p�f��(ւч4�GZ����_h�P|J^x�X�9��(�c�L8�Q��K�UQ�JIէ��~��y�>� �ף�R�^����oW)L��J��Α�x��ԓ;�׉��1���4���dХ�˟xԿZw�|���a�5���j��������*� �aQ*�.)�d��K+��o;U�zAyƴ=���!-�HQ���b�1^��8!Y6�"9JA���ط{%m<��ب#�`!���N���zX�+
{`�+�eļ���}9����n�>z��b�;�ꋦk���@[��*� !ĘB����iP� ���3JH�#Wc41¦�P,27h[24�G��l���������+����+a^Z�{��/nwfQ��	06�U�x�l��/>���ٟ�RѨeRy+{�X��rN��t��X����'s%M�sq�%#�(4�rY�?���	р��ӝ4��Վ�3��u\5�Q���×Ne�IJL��Mr4�b�Z������m�}s�It@4��DB��j��Ui��p�[��M�ʩ��Y��z��%Y	ju G ��{at·Lw7��.��bQ�i?�"����k�ч��(k^Y��)'���ury��k���L�EQ�sP{��Ʋ�=��
�3�d��N�qV�f\��Wy[��H�:���uݜ��͢3��J�ؕ��h8�)�1K��5㺾:�ߛ*VkʹT�c��!�|���a�'�z����*���R��s�*Έw����~E��8�-�+�)����Lލ��8�)k���x'䁤ߥ��(:td��hL;����������L��1{������g����m�NhߍQ4[���Nw��QX?�t�A�n�O�����=�������b2��/���52��*�[��z�~p>�{O�6����P��<����2�����h��~=�/�x*o߻'׶�esk�U��6��lnH��p3�[�A�X��wv�,����i�?���1����lmm���;��E3"��?Qkvz:RFD>@PT�ƨ�٣�H��g�K|�3iI
M�c�2g��(Y��;<ؓ��e��;��� @a�+���X�$5DG�+��E������O�(�NG��W��Uü�A@D����U�2kF�Ap����
�І�l����aZ�ɭ	�XmG�ia��48�i[`��(?��0�0�fs�Q�� *�E�8Oԋ0Kܦ��U�x�Qx{$�A'�j'��d��.��w�7�C`�"�WG�@V>��� u�)V(m����!��dʄ��i�E+�L�����v��oJ7咝4�P��������Hơ�Ӳ�'��h.�~�T<x,׷���[7Po��m��y0�(W��ؘ��(�kn��w��u}h��H�g��3��]/d:�ڈJ�����ǧ��u��U'.fDzi�������]�ef�����ٺ����qǺ�ւ�^v���ba��$Tȃ���`��5���6S�`�@dͲ��rsgGv��E7����"�Nx��9�H͂�r:-$��ZZ@�g�������,-����#C�4��^�4�ke������3�ݤ��J��5��#��ֿ�h�7i�F�SD���E����a?$��7�A�����g'#���8#ų��V�Z�vr|���D��=��vN(#�Ff����T���UV�B�Dn�ٲG�f����k���H�x ���t1��(��hp3�2o/�"�k�4���o�L,������:<�#9��]4R�E36�4@w g�ZB�X�+.��)�A ����s�6B�s[����jQxwI0�}ef������F`������K[��1�1��n���L��w{�z�#��j�W���Þ��urB��=H�$EƟ��j��ulH�x0��U{�����̒<��h��־�V�	���Kf��];j.6��z'�!'��R�Q%=P]'}+���ڿ���	��2�Yj���z��@F�Un;�|�����#����1�"�B�I����ZO�E&Z�Y��N��|!�A.��Yޢº��z���.����2>�=��%������ �:h0��A������n�A�,�	��h�>���	�EW�.)J�)I�6��%�x��G/���r8^/_�˃�g��g_���l')8>�6��Wz���ܑ��i�{K4�E�_������hK$���U{�Z��؞}Ł������;�.�Af�n��T2��,w��*�F�Jiw�{�m��QtbH�f�*�����y�x���:/_�O
 s@� �[��eސ4�!-��c����!�A�VX���󓕵��w?��ï>��3�����ܳy��u:�v�&��˅ ^]���hJ��Ku���Z#�c�N&
��v�BG��L�R�Դ��E���V�u4��+9��
Dzr.&(�6�v����ģ�X=x�Eq6YO��"ok��[&�q���H���8�[t����X:�6�F�!7ZK��R�����lQ�"�	�R��e��2gX�J������qQ;�)�G*�!F���i�Ef�m�K��~[
��y���酼x�'�|�@~��{Re!%�ϒӔ6��#1M���\���o����0����L�¢�8�F�h�����i8cu��������P�I�1���i ��X$��Xs��e��s>2�����xs>�����1�� j{6��c�O�uz�T�μ=d&,�G3OW�λ���"�������6�}M��LY������w­�������vA�f�h,�| ��gH�7���w�B�d�h`�Dv�
��R�2�_t¾�٬M�����{+����~��sՉ����(��5"��Nq���.=��p6�k�r��/���Ύ��ap�WCF�����@�u]f��G/���d}8�.�s5�>�_�}D�]�a����@E�2���b���W�y��p�РJ��<�O(8�<jU�RC3ӧ���@�:C���[e#������z����[��n�^Df!���H��4j�@5��R��L��|Q��[5��90���T�R6�u4؉��e	�#���y^X���4Ǡ����y���z��.P��M����{u�V��T�7];���������C�t��{�rV�5|:�͇�Ke�ٜ�
VI� ���A��gW��}D�����x��������Jte�
�im\��*P֤���8.9�x��m�X�0*_]�k�'4F���W�f���*�Us�����ɷ��%�*Q�a���hx!�#�}�����ݥ������Jp2�H1�R~&�^�z`>UR��f~p�hX��}x^8F��9<��f�-/�B�%�G��1���#���_��0�yz8�{'���^���aj��͹o�=ݗG�>��Oޖ��eYN���ܗΝ9_Hy;�oB'H�"#Fc�m���������fN��g�k�2H~�ݒa�'{���m+���W��̖�i��'غP=�+�6��,�%�I�A�nwLJ_�p8m�k��ZN����iK�L[о�����ٍc��9iYfY�Z��${?���~�����˿�тAz:�b�3�����r�㽣�c�����.
V�C	��@���I�C�U��� ddA�{@���`"��ެ	��H�W)#x�-+x-"��.� ¿1�0���@W	^�Ea��a�	��`�-�n��[��-7n��Y���]���ǄYMP����
���� .�&��Φܼ�!K�u�b왶,��p}���|��cְxǥ���J�_�B��g�dm�1��3��TD�����%+�e`bm��^�Mۤ�ݴE�]�:+a��,������M?����33�9<5a�p@*%�
�_�i�\��Iqh�}T D0��:��/
��NσR�ظ�d (�	�$׳t�҄���K�DEa�
-��a��ɠ�7磌�P
g��̊a|�H+Yt��y�0�9�Z�#K�=m\�(u��#s��08�]��@
 T�`����Yؗ't����'�����?�\�:\���)���	��BD��',^�I�Kee�ⶹ�c�76Ī]���%�z���ɐ���P��W�y�*�)FH�լ��nZ�݂ΑE~�.,8�U��g\3`y�}�B����'tЙwK��L�#�w���v1��<��hȨ^�s��C�}A"Ud�kPQa1��@-vf~H��Μ�8�^f#��m�I��lL�7볻T��ط@�A3Ǩⵑ����(��#�c�?yXhL��Z1Cj��V�����@�@t�&[e���2cY'ES0آX�Ep:`��y��[�,��=�4��v'�L��Lb�m}�E��8�;*��"�w�Vjxt��+�cf�4���09k�0�]��d���`*�U�/q����/�LG�ܯ=SC/U�����;��;J�z�[��D�Z5�K��: �~H��"�y4��T^������|���
/�Nr
�2���y
�@&�(�
E9,�k{>�>�Z\�g,�|�[9<�nd8)��ߣk��Q�&���ɴ���vxG���%i�������`����a���z}mkE��aW�A��xi�)e�U����V��ó������UYZY��҉�]�y�[��y9溄�������vp$�&%�j?~�+�^�l�i����}�n�/^���o���Dn��k�d�	d\�~?�m�9�}�5���� [ru#wϫKE��i�5~���*�\�@s���%]���Y�q'c�%��%�K����vn{IdPa���8�l Ԍ]�*?���$"��.>~�D^��e���> �
��t:�֊وq-���Ac­�m���+;t��Zp�VWV�7����={)�G��Pvy�l���3��x��?~-���:��(ZbI.ƧA/XP��>`���x�hR+�+��\5z�{�A`̢H�:�� J[������r�׎�ڢ��`@K�����P�.�y�3��/������o�c��mb��~��`ȭɓg����������<
F�r�lp��&���ȭ��򳟾'o�ySn�l�Jo��ݦa\VW:�O
�ç�7�R>��apj� ��,"^6U�	![�Le'5P�4�R���XQ�}T`��,L�����
K-���F��H܎�����Sn��X�����P���K�q}����=�$Ɏ+Q�H�3KW����$�����5{_�/�l����`f�Gu�(�Z�x~��Y��4"��.��ƽ~��?�ࣥ�Y��A�l�m��i���!?������Xsa4 �>�Ң�	�#�����qá*��j,] )(흰��u�@���%{�s�jm|�?d��f�e;�0��)�$�jX2
�,��K.�X� ��W�gʜk���F�����ud�@�§�y8�G:���"�eJ���r�Z�]5��s# �¨甌�p���=���]�uY��N��pD���ݳ�M�y����p�����O���}:�k�ݛ�ȥ������\���)y�X��(=]~�� 
��&M~T�U�>���C����vMί�K��'��m���Y����1Vo�#����2]m�,#��eSKl���2�8?��@I]�N8)��H ��9u_����u$V���R���bf��)/�D�d�*����\#�h�g�%��:~�=P�t������ƹ.�H ���J�����;IPrp�Q��=�S,����*@�C�@;ښ�*����zMY����Ș�v&���w�Gq��f��B�N�	h@
@#~.��X��:�]	�$Gn��ި�7�t�;��$Os��_mR�/�r����r��s�s���l%�U"i��I-ha�]�F�z"�-������z�TYJ&�}q���������Z���q�$����m��=���~ ����@��X�\Q�]������X<-;�N�����y}�h�T�
��@�\gZx.n|)��k2��cyxڒ�~���{�@r�:q��TB�����~&C��ҽ��Ϩ`���d�'���A`���Y���i�j�28�I�?���D� a��������X��I#Bd=N"'�^���R&��<yz%ەmpm ,��Gq]jIK.n��գo��w����%Xd*M����'(����	�bPҐ�]��;���_|� ���T��E�,~���
��~�VA�#1��Z�dv]f�Jg�>k�\�:��&�����h��]س�S�C�!���R�>}����u�����@��.�Nv�7/9�F���z�N��9;�d<�����9nRh�*��)�2}S�n���ֹ�������J�.���%(Gr�+5D�ײXN���7h�A�n�.�I��T�&oi��q���']+�C	i����z�X��nv%*�|��rq1$���,���t��(ٯ��Q��H@�i�FU�?��<�H^�[o��`�5"�~����\��H�H�<�և�T�ߖ�~��^��?x]���ޗ��8V��U;��Z]�{=uB }�����==�==�'�������V�(^gZ�� A���sc��S�;0�V���ZZoU6?�4/��MɃ.��ViF'r+c��8�b$$D�J�˚�x\)���?��{'�?�K]�G�Xt'�i(�Vv�aN6��<:�mv�]C��. ɢT�� .a�$�K�)�'��d���M<��
w *��/��p�G/a��)O���1E'^;�r�S��u�͓�QVR+&�<7	��y�=k-V�Q�k���@
X�[�L��$�:z�*�0��֮H|1�R����J������Rٓ��t+/����`�+F�����!y�����0I�%�B�9�0�Ad�nЋ�3}��f��j��y�en�Y[�9��d�B.�O=��\F�	��~�`Q�k��L:hmV�N�h&��.��Wޔ۫鵚��D�f��7����y۴A�	E 	�gm�!�)o\7"�p����ڹ5�M�	Ƥ����6��g�VɟA1
7|��v��y�,��z�D��M�}ň��2�L��$4K��6ƭ��������h�A�ϹQ�1j�<�+m|(��99����z�5��#��ϳM�@$��R��$3]Cs��n�[���V	0�����׹�EGeu�bȱ�l֘�٤��OF�k��
Ϙ�����_x����LHKs�کy[T.��:�W�cM��*��Z��]K^�jK��GP�ۣ�7NO�l���M�e{��GI�¹�@�]`���� wȝ��(a?����q�������WF�*Ԟ}6w7�� ;l�")�.�<�F ;C~����?���G�EO\� Z�8��;]�V٨������g,�,�(���;���<�H�ߤ����ޢ��܏ BRx�#'���Y�=�uo���@�uf��_u�k2�y����g2[MtM�W����������B&cN�'US���ڀV�-5&�vC�z)�~S^�T�z�U���m��̖���E�a��ҥ��g����ɅD�K�
��"�Xk��t(����嵷N�_�'����Rn�?��D� OG^�u�Y���٭܌V�������;����Js�)�&<<N)�Ƅ_#��� :,lu��24�;1E�T�RyYaֵV/��=:�������F��������\���=����8��@������q�}�c�k�����L.o3�L�����{?�g��������*S�\��!��ѳ�B*��l�Ȉ�5t�l��4d�h�ᠡ�%-��%j�We����� j��F�XL�T!R�&4"+y�{�����:����|���z��2.�a��:�urb#n����kɃ���������O�I���E����7_e!�l2�A�ʃ{}���}�D�d>�Շy+�����D~�7���/����'�@��Z��̞ot#nI�՗W_Qg1<���9�~���F6�9
u�c�댎�gE��U`��� �Q��DNj�E���R��EO��e�w�JLF+}Wn���r?�����eqe�E�n���F���{"��U&���ٙ6Lrex�q�R�����o$�ND,��m2��9�7��Rnn��8m�c�c�N~��\�c�,
��v�J~��0DZ��sd�'�K�9 Y�$p҆%��2H\{�'j�alSס6��
�n1��z�XL)��C�X���4tM.8o ��9��.8��1{����F<O���Ź55�5*D�cC��-%�龼��kh�^d��'S�0,z�(�����#�~콋�? O�):�c�<�¦�9C��{�����w�R�hk�cq#��v�|1���!�#��B��i��	��e���?�ǎ��ֆ:��"�KF��=~���hͫ����mu�����3�0b������'{�W�9�U�7�����d9�g��J��,s�9�wd�%�N�6��8hPnV)�Bny���>v��"BTI�ó]�Vu�5i�fXS����٨���t���ݺ4�3M,����
�u�+��9��gP����M$��F�����_��B��J��λ%�%A�bm�&���A�0���ٟ2
3+<X��c���?�G�~�{N�uwO�	��s�+�_����$% /v���*e4)D#�)�Y@����Ey/����^�B���9fS�T8F�%b3��LZ@��cy𞭄̏M�(����.�,tv�֔�N��aL	.Ɏ�)`���1�֦���/(�f���Z﨨�̿�օM����1�q�q����;�)A'莠w�D�@;5�y�a`�ī#����E����d���wG� 37`t ��R�U	mӪ\Wrq���d�C.Z�v{�Ǉ�lJ�s �>LZ�����/~���;M9{>���t��;%Y���� B)�ȼ^���o��P���ߨ��S��j(��F]נ�c���}v5�o�1�o��
ݶ�����\c'�T��$��WgC������#)��US�r��N�O���+r1K���S]�����ܙ"/ {��i��FF��=����F��\�A���.5;cfb-�a�BT�Lm�@>7I���zE�^�A,8�z�z�~9�oonY?xrr*�"?���1i����
�]��Ay�v�Xƌ�+`+\c���>����*eT�K,�W\��n"kE�H�Z�M��5�\i�ͩg��Z4���+���)S7�.��R��5~��D}����tpʌ(G�|l�ciwK���9�-:��5��g_|&��&��[2�?�`-�#],�ִB�"8��//F��w��ݣgr~v!��R����n�Uy��@�>hE���2��C{~!��7rrЖ�}E~�ʫ��s�*`���>
��^�T��P���9Vԓw�;����.n�O�Q��O.��P1��@ò�D�@'BE���Bf�굒S��蘂UOߥ���m����C�{6Z�9�A��hR ޹��ktZ�v�����O���$~��7��cU����Bs�Qv�sD��hP핋:�Y����l�މzMy8��h�����3:^PZʀ��4u�%��]�7�" p��ȊR3��`:0��
�Sw�{�&�G؄Qn�/�fP�L�tFc2��_��N���\B蚎e�ѐ�lB>�|1�32�1�E%����*bd��f�-����g�N�ݟ�˅���� %55�0���p��)�֥��A
�QO<�,�a�eQ9g�w�V8��ʞ��-���1���;�{���G],��|�3#��.�L.t6
W����fd���F8Y����D� �P�QSC���5��h�\�����7�������<��j�g���A�-���<ԍ� ID����w�W����WuM��^���`h�J(�0�(��8�Cnt"�����W��6��`g<�����EM��H#��3��B���j�g�@ ��Bb '�{�������5YK��N
�Rͨ�е r�yN�Ѯ��v��w���:AC�@��l2Yv�f���T7��@d�	2':'�Z��z�0'�Bd�*)���WSu<�S ҡx_��*�\����v����6\�l2t�aN f(u�k��_h��cl"�&Y��K��2Ji6�s0��"�<5{���l��'���1��Ǡ�����(:����"����o�,��� ���)�d�)�[��~��]}w&���s)<�,��7�����ى�I�����ϼ2p-&1�%F/%4���)����P(\�M�0���/���#��s�҂a��2;�Aa3 @GG�k�+?��������&3���X�&
>�������=F���|�����[�h|����r��˚��t$�j&(y�?�I�ݑ��*_?z.O���x�T�Ԓ�,�G�.e~;��'ϥM�u����h����\���\t�Ra�j��~�2Sd�*s�_������og����[�U��κ��~L6�	HOZ.��
g���i�~zy��Ȁ���CN���3�*2B]�V.����X���;��S��E��̌��/rqv1�Zs��'e�`4��N�+�t��'w�����C��k@��o�U8	�L�� �~�!
8F�׺/Xgv���9����d2��0�I�_e�|�[����ژ�� �Ie�\uP�Ln0��Y��Y��Y[�d�π�2���1�$K1iZ�
Mі,���5*ia��k�3 �f]:�6�|htx~~�(Mp�l|YX�"lt�W*
J�����X���������?��y���n�U��F�[y����ǯ���=y��#���,�I���W9:���~O�x�T|[N�����X>��������|�ct�ȍ��V^yp$|���)����r5ܗ7����wt1q��C�~����X*��N�P֐�d��d,��" g}h����vSca���d$�E8x� "�dI&���)7T�G�BP:mP��������~BU�V�KA��>z���4�j�[xEs�\�A|;+D�Ӵ��#A��,��8��� ��(!<R 	:����|Mʊ��`���E�찁kHe!�bTI\��LOLP,NV�qwm^]�S�����p����y�a��|���viUȕ���ٰ@���[-�t^e�_�M��^���^��-�;8��"����$�JT�@_�����%ޏh�%xs��~��M�<��w�޸o {6�s��;�An����[�K�s�$>���T�c�� j���C昑~h�;ƴ3�'p`��~(��|R\��gh�Xq���㳡����4lX�4D.N��equ�q\NƲ�O�h�+�P:z�WS��'3:ѓ�%AߓǷ�-TU;v�iHU��a�,�%y�[e&���c�ʁ�~]7�Z((K�FI�D��)�v9i�<T?���	�ci���F�ME�j��k�j�;�����fOm(D�+RNkz=��k��Վ� q]���x���ַ���s��sU�D�2�  �uJ�z@vP+��x��C����ԏ��d��pN��g
�/F����a�
������7jAG�z u8���e	��D��B07G.\6�<̵������a���9�Gਔ�;���fS<�(�N���pP8������K��!���$�A�9թ,y[T�����������vP�,J%G���!qb����Md�@��G^��;��ʲ+����;�󸅠Xv�/�w�E1��WM�e �_����kՏ�y6���:��>ӝ���	%��ӊ�z�G��}�Tv��;���h�� ������zaD��,l\�?�KE����c���J��i�z�U�Y��h"�'���܊<�V},Q�a�3�!Txo�;P��G���lI��ze-���V��XDs�����S�l��D���e��-ӐŮ�)��� u,�*��"(�ٟ��->���֋������ZkJ��/�΁|���z�[:ц7\v.��)̋�ؤ(�}겗�&U�����[��(({�6�J�Ẃ3�k7	b��y�ιX�Z���9`Պ����}����T�Ŝc��n��2��R���]�i֔�Ob5hn>!��+�Znn��B�l�̊���?{����j5�A�>$���JE�褬� 
��&��Өw�I�#S���*��dک2U����zd�F1���Q[�Hk��.�1|��WA��?���zn{�C�>Wǽ1�Zc���|������w�`�݅�[|��B}���w�u]=���AE�"r_~�XN����Cҵ��h�:��-E�U��ф��.�WWO�o>�?��c9;�d�Rэ�%
fP�����ۖ�����rrҕ�ݜk]�	���P����hj#���h8��4�ԔX�-}�:]e(jg�h	��cLHL��|IG|��� l�)��Q&���&|�B	��ʒ�i�X���\��)8�Q��o΄��ݩ���kz_=��yg��y�Yu�5�h i����t^m�H�/Prm3B*�!z{~~#�|�|�o��7������U>��/.ĩgٯS'5ho)v������]r#S,V��6�3�A�ɢ�C��(��d0��X�S\'
��x�un��i��H��Ѿ��o�30uShS��N�����>�]�^ժM��#O��i��d����Wbk��:u|OlR�-�r���m���+����y��I����0��w�l%��+�����uF�	����@-���&�꛴��	2���|n���Vs�\����-67u��0ˢ�"��X"���o.�R�pO׻:���x�(8��׬��f�ϯ���L���
u��M�yc���k5i,��TS�-����K��D?��y�nפ� ��N�ت
����%��Z�-���0�ӾV�K�A�y��f�M B�p}�5�ꥭ�[ �7!k���Υe��-/�����
�j�!BRA�2��7@�j���S�����q��qk6tުMP�;M�k���Le�_�Ù��W2^-(ڑ0��4 ��5�e-TI=�F^}�P�/.,�'�6��i��76o�ܼ���AV�Yr
V���!�H��������nq
P�s&������;cw�O�עY��lO��|�`����p.x1u���3�|8@'��Gmߟ�Y���Pv�2�IH�	�.�rF�	����	*��~(�� �<�}e�]���A���M�O ���x�?�[��z:���S'��z�E��.����l���=�3v�|��3;a�)d�l\��}�?� �f�k!^Ӂe��[�7Uf8oo�r}���<��O)�rq�Z\�xa���['x��su��[��;aC�jf��\_NԟB�Bm����r����i*� U���i��j  66n|�vZ�S�6���F�u)���T!��]��8�����N�jY�����(����G���l��sa_�����&bF{o�]biB&�/U��r�I��B�c͠`պ�W�޴wp�~p˾�M��Im`��3�ɭ�"�K�{�Z������' �����QY?n�2GGK�Z��_e*��2Rg�T���	���ac�թ�V�9�@��)l��xI7�Ɋu ���:���8&�U`(k�ԑ.հUs���$��.ՙE�-,�F����C�,OҚnt���פ� *߁�dP���C���مnȊܫ�W[�" �|u{+��?�O��R^ycO^�w����k���s]�kb�F�̮��-���ht��p.�NO�J��gOG��]���c�P��Y%Ɖ��G×�%�Rt��̬�>�:��魌�[��,�a��#��@>NߣsA��k��l(7�e2�q#v=@���l�h�����,�`���L7d�� ĥ��rJ=����E�Q�D�w�V��j��:�Z��|/һ �����S�����F�%�M��o�������������˖�����\���W��~"_~�L&3u���q�%(��1����Wf6ߊ�O�q�.��<e,t1/�,���yZ�N��ݣ�*ľX[��?�x���
K���A���v�P��jp��YDP��s��]y��Wt-Y�<��t�ip�@�z�lx8�j�{ai!^m�*A.$�:�9�s��{M=�L�Ĝ�U�8n�sNv�I���K�s?�i�t�/�DP��D�y6�|��C�1jW�ѓ�D�àdϝR �=�
;��#��s`�_XOu�c]W�b x ����r�f�dO@�@N���^��Pm�]�!a\�I� f�5��Nu�VJ�V�(�8��t&W��d�F�'j��=)��з�d�ᒢWQ�Mdv�k|{#Wg	V�����ה�î���;��w���z�k���d��Hץ�d��BY�LS��zt�Q��Ԩ�RQк_��t�P�X4��:'�T���@�ծ��f�(B�F� S�^1S����H�]�~�#ǽ�vKr:���EE~x�ȳ�B��L8O�ԭ�� %���Ր�iG�����!�?�A�0�vg՝Ix�_��m�(�[��7��0��fKn)����Q�2���i�?w#�/[xx������0�}^H�F���߹���z*�8D�)�̴9�pb�GS�+�)�y:���� ���� $�흘m�]ͯ�ԭC�1�@�q��.{�A���;���X�(g�|>�ۯ@rz[~ovK a[�h�xDk�?O�$�U��$F,10kʔ(�c� L�Q���ԙrz�3\��U�[T`P���p���ڀ����f��۰�0�a�	��N��ս�bY?C�����S�#'�2�t� sP����>���X��T`3!�n\�*�VU	�o(u8�ׅ͟��&�yݗnq=&�_)��F�w��%y:���&�?��w�M(/۟
bޗ�w�56�d���q��-�Ǩm�HE�y���5Ѷ�	�$q�����H\��(�G��5��2A�`�������!�&ŁI�=�8ZWa,l�ք��Ȝ����v"��W����O�u����]\\@�*��ҫCRf����l�x�d4���WO��_�MIH3Le^�Z7V� K����9��<k�����H~8{.g�Al���ylr�@�B.7���=V���`Eg�Ρ�Չ�F��b71R�	;��y�s���XG1�"}Uc|�rE���,�:	խ��O!a:�(�ԁ�A�?>��l"Ǳ9x�V�Y	��u;� �.�2ռ(�tɍF3�G�|�H���<��x���nF2��r2c��b�Z���&� D�#�6�6���{*h��Fp�	1ZJJ=��*��A5��Uu:�0��ݩ��<Q�? d�1�S�()��'�F�b3HH�s���Ͼ����Թ}��#9:��mR��e��φ������:���ِ�
f�C+�7��f"���\���� P���'�˳g�������8�Q���bH�{��6�4�6�	\�FhQ-'%EρŃN+�qdwO,l���8˾K2��q\F������E�@0T۬�Cx��t|4Vz>�>��m05�2<K�uZ�P@�[�挺�(�Q �Ϟ2�ؽ����]q<����q|x$_�������([�#�F�4� ����͎�
�bG ?�^5̻�f|׽�Q]s^\J�_��ZG�@͛��]�ސ9&���D�5�j=�qLXɮ��l���5�v�(�.G!%����6'S��m��^���`%�$��X�[}���a�:2&ӫ��Z�,XȲ��~�#����^R�E��UIme�$'�
D����$Q�1���x~Ms�t_��tO��]mJS���ds��H�V�Y��F��92�j3���}9��y0�yՃ|zG7�Z��0D����Z�nUԎ��Tr]��� t�sS�Р��۪�rUc��x����,l��d��^�
 O]�}ypܗW�r�!�?��u�{~3�z�����nunE�i4X���g����%+N:��tT~��q<����ۭ+Xwc��Sa�Y����)����û���N%�Y�r�IN����C��g<x�\8!-D�}�w[�7�J������m�����;6G�-+�پ�Z\F&��(r���u��(G��(�N6ge����(u*/ˀ��k�~Ѝi6F�=+�lD$�#
�)�-�{2a�xa��JYq0 LÂ��Yz����.����na�y�0�%�u$�9�b�cИ�D樵���킟�=�N �g�z*H��2!	��D&�\�� � О!�����q��R{��H��~
���=k'�H�V���N���!cc���1R�k��Y��*�A��_�<Wʓ'����N�/K�i�~��;c)w���@�[��s��rY7����\_-�o-�y��(�O���$t*�����1��"c�� �F�bh�_���@��N�ϔ`W�H&���n�8���i�EC�㖄TR��[oԃz��{�7��կ~�w_��w�W|���nKG�f�[�{��Մ�
T����{9:nY�tm�)Պ�%@Gqր0k���[�+M��������_ؐo2Yp�'�d100���q����Q���P�u Ɋ�QZtΗ3F&-g�a��ԦzP�T5-y8�0�p��,(0��W���Zm����I����%�����ݓӓsA��ZmQ����YB��o'c]]1jz���܎�	�x_zSu�A����L_��:�"��gCZZ�"ז:�0�[ug,&�2�f6����w�*�櫩S��k�:\�\� :���=.Hȭ����b�eC0V���Զ�.��	���<��	��l1�_G�	���5����\�y Xp�#�1�S�mq;o꺸ÙW�˫�|��7���_���Oˣ����v�l
�S6\+�E�L�fw�(��ԑ�c�7�^Cׁ���Q��b3+8�_���9�o	�A}Ľ]��v���ꦵ�s�1�� 6���kI:�==o�ﹾ�t�L����Nd�����ce�#���@�LFd<�f�����b�ud<�+d8�t ��� r s���F�A��C�)�.m��篦�;6o�`��[�p������L�m��x@lN�Iy�Y�$�"��3 Eɐ�m���w���j�`�I�е��~4���@dY�  ���u�]Ǭ�*��`����q��ج�u��2A���&h���Ѐ/P�>(�r���Fm�bҷ��7��g��/Y�W��+�����԰I,����Z�������c��eE�g���(��:���L�Z*�T��X.�,G��S��p����iP?nT���&�Mr;��l����'�\��F�5ٺ��U/�N�:r�d ���������J�	��(��?g2�*�Q�߆jJ[�N���I�!ޤt���^-&ll�}�Z�=�4ZRk �&�n�����bR����E��K�k<�X�mU����h��{���oXV�'q��4�"Fvn��B݇���
4ހ`�n��
����<wtw��;���W�c�W��7�����YY5�M���q���Ѣ�ϻ߇���z�:(/0���'62/yn�M:�ε
x���\*;yvq5(4�N:4q��Љ>���4�[�2
o�x��h��u�}�4Pٵ�/���l
Ir�qc&�_N�Y�K���(�f��Z/p7A~��%���l�Ɍ�K�+(д\�*��3`c�!\#��󼮩a�V���^�r>9�ςig�����KQ��}/ u ��<Y-�@�I*�O��,e�G4���� ��HڝxJ}�v�b�	L!N}Pn�k�H֭>��w&�f�g�C\/�+?Dܤ�*s|Kb�I�J�`~���6w��R'Y#4��OH�����R);���:���)�Y��Z�2���w�����y��T�1*�=_7̤b�!�ԶMY��Z�k������/~��/���o���}��Ͽ������ra1�б�ҋ^<�𘎎�(�vttDN4(Pw�ϡ�Eז�nn�u��J�m5n��<��R�T���	��e2[�C��+���!vu
�2q"�x(F�6l�g�����\HY�����G/H����$��Ao�@Vۈ��j.)���z]�(��\G�Ӊ��L�s.��:�M�$�tt�����F=ѿ�Y��(�l:�h����-iH�Q���4d7Vk>�n���Ap�f��u���ׁ1G]>�64ڰ�*a*�.A��NƖ�#dXb�졂��X�o���H��(nǸ@0 �l��w�U���!2[�3�c!J�"�$v!�̍E��W
����k��W_���݇�_�B>���e�
X�[�@SX���jat��թ9ա�֤&
J��v,R���w���/���׹��c8�3�4�P��zRT��hW"��� ���tsjQ;n�iꊞ��!�m�|���Y����ܹ8gj;Rn�R�SB���ڮ���Z���Rr�-�'�=���p��ɍ��7�զ���kH�Z��*��YNu���f�(��[�H��l�XX����Y,"���L�����:����@v1�p�r7Y7W3���?�L�k'��I���5�vs(�.��6�i��Μ��2i��5u]�G:�B��R{�ߪ����S9R�	��Z��|�k~�5�z�$)KW�sV[���������Z��f9S��"�
�ձ��ѹ_+뛑��ao��\3;OT\��G^��G!�t8�N�+��F���l���K1ҡU��Z��=�sȑ���P��7�Z-%}����4��� ,��t<��'������K�� ��Vkb�!3v=�P�B+]I9���^�peqݎ�[SA�jV���)�����H�RU��m4Y���$,�@�^ �NGsY�kT��4:�����������U[�9��[v���=9������EZ����2��b8�L�J�7�}~#}�ۃzD�XO����uI6��|��sJ� ����9���^6e �V����Xq��+��  ��IDAT�B�0�.>�k��6�X��y����!�.��/?rQ����b6&#$�b��'
ߐ�xyǿ�`�ѭH\���6y#c�P�]���j'҂�h��ݎ��8�g}-�O����/^R~)�^��2��\~ ��q	 錰K@�ղ��:p��2���KN��K����l^���W!E�Q�H6��NS������ ��;@�ß��=e1P` *�؁��E�C�	���_+<Fh?'\�]+n�-�b3�R׏6yo*>Vr�F��=/>�LL��P����/��\�׮Ϙ������Q��������u�7��ʠ!,����2�V�ì������M��E�m=Fzp��Ă������`j�q����ͣ�+�
���~_��T���?����#��ҫ��M���#J�4c�@^����nU����r�iVd��E` Ҏ�*%��c�+\ތԁ���vfM��-����[�b.�hcr��&e��>�~o_n�n,�H�"�$(`�,L3:H�e)����	�QE��MẄ�­��|���Y	8�C�����9ď��V���D�~�Q���N*��Ldr{C'�N��l��@�8!!�*Z�5&Z��Z,f򬐃_c�Wk���а� ��jRE�'�a�_�6�R��Y��"d�!ي�H�)�z�R� %MW�T�{���{Pbu<����t6sE�T��8����o���B�����߾�������7ȫ�ݗZ�d�mĮ�ݨڂ?6��#�=_�1����P?~"OΞ˗_}#�<�Q�Q�1[��e��:#]K�K"�A��G�ck앛l�G��C�s^������s����{�9�!��J�Ԁ�)�/bO���t��O��&/��[���t�qȒ���+M��`�Ս���(7�c�ڷ�s�X�X�(GA9�*�p\__�hd�7�!쏀�y�z�PX�t����u.fP"M�<N����㌧�.��č��XR=t��_�8@8 �
8)�d�7f�T��' �����Y�zߝ���J�����:��)u���ꍠ�(�M��:�[]�㊮o]s4�Py�Rj4�4�5�D]M$5�#{���u�골�)����_y�Y�@�P7�+�}�~%�D���>�L��0��4�z���Ƥ�2R�L��ư���nUJ��T:mY�I�N�6<|48��"¦kv8������^Oʭ:m�`�rC���/}yT�Q�NL�1$�K<H �R�R��[ʥ�� ^��`���s!��$hj��ظn����P�V Ӑ�-��"����5�\ؚ��K{�DTur|oO���k	�H�͒LtY�vM�U`3�W��H=�\��؎䰕�j�^+�����$NI�Ȋs��;���c�'� �`��-촩��8�7���K{y
Tf���w���[��A���Y����������Ř}!;0������
�)���RP��pO���a���ϖav3y�9����e}3�����e�s��[�����_�/ ���lk)� �f�n�9�ق2�(,$�^�Q򀖓
6�@!+(L���(-\K�߽ϗ���:ɔ�?�	�6���l_�{�p�q�)O#�u���0?w`����+�����X� [�A�<i�b�B)��T��"u
��N�Ҹ�Wa���:~�w t�f��>X��`���k�GQ�a���''=�������}H�l-k��]V3�������Y�EP��4Z����h�����9����r}u����ѭ�'>8\�������_|���_}���������Bߏ�un�#"/m�N��2�|�ݙ��s��'ҋ���k2Rz�Ƈ:S����:��u�򕂈�ۉ|��R�_��f�ٖP��r�FkNVd�*3�Ņ�:A��FW��v����Í(}���|�U�L��'��r��9�T�����&9_/(kF���������/��H���y��9��?��3���f�x8sB�fV�����hć	�6��x!�@�F�6/D���9e}A�j��&7�Mx[4�麍m|!հ�4����f���v��nl}Uj�5f��E�΢uk:�p"�=�R��K�C���WKP��l�~��;9��=օ��c:��f�`Ti26� ��k�2������<�"��~_��u��:&Xj��k-�ۛ��ĭf:ؗ����<����K�(:_�����Wg�a�cbp;�CF5H3㚱x}�:-�bQ�7�����̅�^��K��Ǳ3�p���iC�9��3�b�m��ci�<.�o�����]�Y8l���
�L�/<_d��C������� :��38�hX�^���}!GG'���*MP��ͦT�Q�3,���b1#���6_1'~�:�Gá���/[*_�(�[oԜ��fI��E�b3�]<׌1�:������M%$q��9o�ϊ+��g
u���a=��-��(#U�b���(`H��:ˉ:�-99���{������9���j��FD��d�3&
֪z1m�W�g��Q��ZrTX�㽜^�XH�%��tu�t���J
 Rg*l�X���Fz_{z��t̡���n�H[]w�ڙ�����"m�c�����V惞,թ��AX��TҖ@m��<u����㵜U��WESF�P,6E�,��AU���K4񂃭�-[��4��w+
�ҭj����1jU����Q�\���E��5�{�&鹍l��iK�j�!�=;�!�i(���J�`OuN!�����|��y.�R����Ѿ^WM-N������FS�����C�QP�gS�B+��3y�/�l��h1��N�Z�:����y|�Fn�Et1��(A����lHFG\��ζs�SG��2���X��y�RmCPx�/Bw��4��{�X�;kٹ��,e
`��B�UmR쀎�X�!6^w| ������
^�t��qb+��XN�"��[t�v�<r]��x��J�����K���!^����W�g����Kv�� j,��`���}�lo�='LSJl��d~��r�{�j^2Nw��/�I�U%�=����9u�0��$u���y MM��S�$�J= ,(w�W�@�ߧ�D<�l'��=�|��GοlU�lxZ|~/]R��#u����v^�K[��A����X+]��4��?�N8G�9N}ѷ�􋍵��J>�(yv��0�o[R�����B��s�8��M���ڥ�e �W`G�ǁ/?�����d�F���?��g�}�s�_�UfR�͕,$ڢ�B�}�����:*7�n����]���1�b�YI�זz��D8�P<A1�t���|�Vg��&m��c(�<��N7�8TB�*���HH�m�9<80x꠩���Fz[�l��-���
�P�zr#��J�oo�,�E��bx}#�O��s����q����q t������:�
D��,��\���� �	��(T+�~4���i�27�Y�-�x81CCƈ<��\�m��K�W���l� �f�H6�[R��b|{%�䒙D�HꊂQ+��8鴏���W�eL` Z�r>gݝW��r���cu�n���B���;���3��Nƾ:� ���R�p��t�ԹE��vxKz�r*�:	x�:O���!.�Rkn�X{P4�÷c���B"���(*D�=��d�P��x2��G���NS���Ŕ'5{�6�Jى �d|Qa-E�F���)�MIeY-��� �Be8P�t\O�ݓ��+}O�)��zė��3��{�S�H��c��Γ�g�S���Ϟ3�
i.J�l(�ybYS���Ħ�� ��X�ͤ��>6fT� =��<��k?���hp`ˡ��L]�F�zE�� [�ڗd�PG�)����*@G�nM�(��"�Ǧ�F� Y���b�u]����XQ;S/���$�4Bd�7l�UAFN��i���S{@�U�
"�	:v��s�T������_&�lo��ǟ����z�'�G�D�`-d�B�0<���v�vuzT��hK	Y�J]ک� GG��� s
�,�k�_h4ٖ��s�?���<B�Lp�aPQ����ASN߼'�.��v+o�oxf G�g	Y��ҹ�=�,=	�u6m��js�t����}>��^Md�'F����D��M�����}�{kv}������L�u����U��#�٭�nf\k�j*�'-�߯��͘=K֛��Kݳ�
�6}�(�/�lZ��۸�@h�RP�_˩9ge����S����N������f�l��ݬ���t��}/�'�:O��9�KALZ��d �=/��f@�r��M�ZO��_��#\��Qub�gek��s�~���R�^��������`�eZ��������@��+�~��n��=P׃��w�~^Mh?� �T���>��"���N#���L<�zG��;�AO����e�rH����X��}6B�-��� \Rع�B�\�ǦL*�������������K y&%���-n'�6�Y#w�=w��n�U ���KD������KJ��a�h��ӭ�������U?��&�c�q�^�� >�J��'��ο0Zd)��:�N��&V'Bb1N���>����P|�Á��3��c{�]V������׿���?��/�����E��_�*��,�^O6DeL+"�4H}�.�i�Po�c�E�8�$��j�tI��[ȇ�������Y���`-,�ѭ�$�r��hd���lXo� ���]|�`˾h���d�C@C�������奞w�q!��m�/ M�Z���QO7���������O?��?�B�=y��3�7�wp�A��sl��*����m	 �Y3sDŐĊ+�u���@�%C�֨qk ĥ��E�`�B'�&����%��+S��`�^@��Y�Z���^���t1\�\ �"��0:�:"����chE����������6#�pZP�f{�&�k����s�>��bS�j�p�����6|�����ED�q,� �P���OY$��J�7�dNp��P�ʕ��GP0�i���1�+�k��ҋ�*�MQfC�!~�\aG��9� �H��F&���ߧ�3���`�$24.n����Q�6�Ha�ZSJd*p��t�s/W~�7�Nu]�����Q���o c��?��Φ.@��Q�l~���b17 �&�j�R�+����c����^(A�f�E�%6Tn#r1�1�\b��mRT�1ǎ�	�RVWTF�;�� 	��j9 [��-�=��]�;�j�6ֵ��oRR5a�r�k� �ԗ�AK��&n(Ѹ	�ojWS6?�&r~����^/6F�!�[K(90+���j�z�jb�O
PJ\�f[:=�Y	��!����陎�H��D�{y���t�Ri��f��ڢ���f[��c�WB�A�BA�2�����Ҝפa~4������jK�R�{rz|Č
�q���d��sP:�T�M��+�����I���r_���S�^%�J~���2���}��-�^�:��\�>�F'T��6v��Lj�����T���z�gC���<{~!��ci��xu������]ͮ���ﾌ4��NO�w�g'����lA��ז- �;��.,! U=��^ӠW����rv� �܁�R.2�M��|CVĜ9]��z�b$d�Ô�"�-2��X��>g�h�[�<���8�%��X�<ʛ���5�|�"�D-��L��]t�ih^�
ldsLQ�$t��y��{�6�2@��Ў�g�d1S�]-,�u�����_gt��A^>�iqc�ޓ��ׄ���kG�8�ہώ;�Y��`TVR�}k��3$�0
��l�"�y�<|���$qe���/Ԍ˴{����6w�/�U����*��~|w���k��ǝ��"��{�<��%L��ј9YŞf��l=�����cv�� ��S*�ݷ��] �K��݂�X%�!�}w�����l��hAqA|��V+e�Rh�\�{��0M�5Qƽ�G;	u��'4��^��]��á�Os�|�7;B��_�@�(���U��a%�L"uR�����o�ۏ�Y��g�����eʵ�kl$ȁ�*� P��g�PCNs��n��
/�$B��HL�qCc�F50��,$:Q�/p�t�^�u�W�d��|DC���9E۹>4@�1k]�1��LϩN�n��ۡ\\��tO)m�p��5JDAv9Q繥^[�5(�������|�/�w���3���V'`�N@�I�֥�����T�B��J�PH��Y�g�7aD$+6����8��Q�z((��8��n��֖m��g*D��6�Պ����w`	8�33�(�����WGz�.�DD���@12&󈔇[�;��������U]7b��#Y��:G�V [�K��;DQ�Ι�d�_k\j|��|��� k�l��ށT؁Ӵ2P��LYWȝ�솝p�i���/y���7~ި�Y�s/��^�Q�\1�?�L
�� Įt�YTО��eYw`�Bǥ���.JS"�G�+�3cκ�3��Q�˹o��w;m���a6�<H���R�,(Z��O�
�
�i���R���ٓ�hh]�Q;�Ƅ�e0�y��
ѱf ˋ�$��DU��x/2A�e�'�&^�w�/J��+�� z^s��h����,�BT��J�9;h���lV�hЕ����Ŗ�I/#S�:�1�.(�]R���\!��*�ؓ�~W���/�u]"]��~:~
B@�u�K��Y/��[��,���z�r�!:�G�L� �Ѵ57�	+���i��k��I��!G9Q��ne��d-�R�n��S��'r�Ϋ�󏎥�Z�[�@��]���ߖj ��\�j�F�Υ��TWp_K#n�y����5�#Q�@�X����=K�����Ƴ�ʷ�� �}�X�_�-�����s�Z�O߻a�r)��^k@M�K�"탎ږT��D��'r��k9r&�WsƃR�u��ogS}�Ͳ�[[Z���ƀ��ZC��-��Hn� ��T�
�/n��h<�A�e�"<l��F���v>�����w?�:���RQ;�:XJ{r+�Řs+��j˛�4�� ����?8��ko<����ɗ��Cy|9�5�Xw��4���"�6
���V��9�K������㓋.�j_Ip�D�����w�J�#��D�����3�q'y�V0�M�qփ�؜{[9ŮF���)�@�ˠ��2'��"mkr�v��=-w�_|�t�
��?�1*F�]�=�|�ܡ��ޭL�삽-��Z�mX��]Q
���If��"�Ø/��wLG=����Tp��^���V���d�_�Q��3o�7R��������vW�goe���t�י�OU�0���e�Q�+t@1
bqN�x�{�O��^�[�4z��p��[�h�\2|D�_��߼%)��l��j#0��~06�b��}$��q�8Y�X��P��Č���[fo��6\����򜥒UJY`Ԟ�=kv����ד��1}OTWo�:ja�^��������?�����/���e"-`���l��1f��u�ӌ� 8�P�\��P<��~�U�[ivGݰ�@ 3uL�l ��&�V��:��F1�0��X�K�3П:u�$N���-I�y��ci�J�׊z
8�%4���p�+�n�Һh����e}3���H�R��5ku>�LJ0�T������M
N���Į�6Ȥ����9K�{g�:�l������:&,�s��2t��M{p��,t�p��?���Xc�tZ�}�  i���OE��25p�с}�? �
}@�����ҽ-�,�F�Od�ﳫ:
�G�?�?���y�y�Ծ��Q0Y=�	�N���a� ��h"�N�hp��*!�F����hn�?��EZ���:��h-�%�ǜ�e`2w^���@B�6�����]�ʅN.23�� �P�0p�;hB[�6ufBl�����z��g���7����:��f�s5W��1)Gs*��I�eܰ�D�U7�^�®�8���su�'�r0����R���LHj��4����JƠ�Y�JH~�)o���Bc�\'�^�bZ����\*��X�`��j��u� Ĳ �v%�h)�A��4�Ȟ������� /�����?]��<��v	=-�ȁ�=���KR��7�t�N�D�]���:�豱Q�6E�������"Y-R
6p+�q�r�먱Ld��g4����;:�*)��'r���L�גV�r�����"��ޒ����m)'��u:56Bm���T���o���od=�8��ʢ&�Չ47+W�]�	��r0���~M��Uj��JǺ~FjN�RI!�=��5c�}'�q�gБ*�cK������4'��+��`_?w���v!��~��X��;���l�@��}�%h�u�L�ׯ�+�u~��
|"9�2���:[z������ڇ�T�]iK�E�g��g_�F�S[�G}�]���
���^]<�g�W�֛o�`��jr�%����F�8Թy�6�R�]^S�d��i����X�!�����<�L0z=��Z����B�{�ZS5O*6�K�
$�;�m����_�8�w���(�es%��Dn���aL'�Y/��n?G`-�6B �=t*'�[)�n?��<���%߯��}9@��\Dn�S|	䧀D�k�������Պ��D$+���}���@�şH�,��i�1z����52�lPGݘ�fI[�q��Y���;'v�%}a>yj�N�ls!w	o�s+�;���/f�����䙸�\����E`��}���{��τ��d���>�+L�ݯ̭ȁ���3l�z���N[�̊:��r!cu�/�o��<�HL�Yep�=8�-K�1Ɉ������3C�W�
��8�oS���aG�بP5ւ�;
s��KLQ�̶������M��q# �U��k}������_����dr+�E�rZ*z�咩z�l"��H�E�H�;)�o �8ǉ���M����.ƈ��N3�nt!h�J��D,���KՖ��}�QY7����<|�?�{�p���|�l��p+e=�ZFa$"��r]�MB��x}��:�9֯Z3�����3�A��gtb��w�� ���Ђ�BZ���'�n�Sp��:K��ٽf��6���5���D���,wK�Tf�^�#2�R*ن 0��P��9��.��q��n��Ԉ � C���t6WGnf�s���~�����J./��_�ׯ{NeO������-e^�dƦcb]U)%���	�,A��SW[[F�wTf2uiV	��	�g⋶���"�(�uf,����%~z�q��6�ۢُT��F�PZ 20��ٙ�*K��@.u N��D��"�N
���9aL�(�W�$�&A6���L^{xJ��<1��{2�Иlg�a�
s��ׅ.�'�*@�px#�׉>�:�ul���+�b�"����oZ�`������F�P4õƮ.�ڽ�W%�0t���j�rX%O(���@�AU��M����n�zr�����+𨳿���r�u+���j.��k���2�`�*���@�
��ԉD� ����|�JH�ȫ���U�v��6 x!�0UǷ�c�ڥ^W���xԥ�Æ��]���6�_D�V����[u�g��[o���ߐ=���Vs��k%iM�RS��h3c�l�RG�oєp�R���(��{)�uS��U�^���>�E5u+ݎ�2��c��
��VM&���
,G�]&-:И�U�XTbYͯ����\
b+��D=���V��뺣�����Um���@��n����Le��K�j�,AM��r���vp-�O�e~y+���(݃��)]��:�~��v볘QZ���g���s�1�}:����屮���M�\�=}]�z�:/�눀�>�{ǩ:j��_IM���%觠��1����2��|,&!l}LV۔����,�v�AY4\�h�h�]|$�+��?�$��Y���fǱ�[��L=:�=ž�0�L&��c�Ր9��^8�; "v�0�;F{*��e���~$�SL��;�r��;�,�J�܊���_w�� w�9&������[�zQ�6p�T�4�`4���wx��� ό�*%�OȌ�w�}���=�/|�s۩��(�����������x��^g�����4̿/�[x��+�
�E�Wo�b=@|���^���v��;��,�\mTY��V�h,�f,։<;Ru:������q���k�c� r���0
�W]��V�
��%;�#0�@�Z�Z���}����0��c@�Z�.m5j�[�,oXoY��9��ٓ�z�CfK������޻���o�����O?�����_����R4*I]�ĥ�#��mq�$_H#]2����R,���Eޚ:X'�=��_�����^���z�$�����͏���ݮ�;�J�{ù:&%�r�Ù������ǿ�=�L�d���z}[k��k��1�{�q��miU� ��D�ӳoe��B��Vj���i z
����7[J�.�L��0[��s�	�RɊ�Lz�7g�I���}\<S�NS�I$���k��һ[lg�>+��m3�]�����$���{#���ZV��
��u����v$��ͷ�Z��s:���39<>Q�җV�!��>#��i��*
�H,KW�g�q@A��@��͚/y���o�Nm��esfma*{�e���1k2h
��
�q��<h�@�m�!�=B��O�2�s�5�R�Σ���F�ur|NGJ+��T��ì���*�I)�O,�Vp 1��d�F�=P2�s�%�y��� P��}���3�����\ݨs�S�yzrB�4Di QH�l�֖�.��E���{)n����9��0��r]��r`�P���
T���!���Dù � ���@]ց�?�C�
�:�*7i<���nf:7o���c�|z�L2� '�z�z�^S�v��T��Vu���\-���obc�!ձ I׮:�H�7�M�ve���@�,=��H#l�f�%�ެ���}�T��Kd�	��#t�l���H�����M��JW�_��s���:"k&R�J�̩����
(ӑ�D*i��p���W��B6G���V��ڷ9A2F+�k󙂱�F�
��,����٨m�v�H�D���@i������͞$9��0�#�;+��nt7f ��ʴF3�Q�2ʌԛ��M��t��A�Z�h2�=DR\�`g�3�c� }�]y��q���YU���r&Q�Y�q|�����y����Z(�w$RB�u��sI[;<�K���>��0�h ��?���lD��tͭ���vY��wzt�����3��_��W����!�wv���&��n���ө����.Gtu��.X����\T�m�=xH�?�WO����.�3;!�贛�� �|P�T��v��=�˦:��'O��)���Ƴ9*���y*���b%We��9a�� ���6�ro{�o�Q��7�7ĕ��{���3���dFn�T�"ĸf͑Fg����L��x/6Ԟ��D�$IZs��Ue(<wQ����#%�_��Ԍ62�|�9r�+M3J,��`m���0�	�n�6���~�q_IN��	'8-]��'y�J	�^�1}`�^�;V4��165p>Y�(Ӥ��ݍ�L�Fj���#�99������7�.t�{�J�ʟ�M $��]ǹ�Q�Y����h��3Gm�le��Y�����{��۴=u�7�k"U�,�����A�����,n�.�,�_зߜJ�&���%:�� ���V��W��:{9�N� lf� �I�C�lW`l6+��jH�'�]"QLdAA���X��&H�Y5H��&�^��P��	Q/T��(KMoEHu�4P�'�������>������g�}�W�������_�C!�(������B�/�$�, �P��I���汓-�$�{�Ӫ�;��I�{?ا���؏Fc���D���
���=�=6DPh�^!^������Ƅ����O�"�:+�+��0d�ӕ����3V:���_�bQ�^���y�HMB�c��1F�H_M�����:�����MCZrDb�޴�t{%�y��et"�:�f߲B8ή���i��o�7uͱ�g�L�H��gk�E�(�g�[]p5ꌛ����6�o���2kF���]K�xm�&�� R/��VJ�@���0��`���t�Wm�f ��R�ex����SP�*�Ď�k�}�-�K��_:����N���1 ��Rm�
���+���/@]�V����g/N��`N4�1N�ˉ5B&P�\�1^4Oj��ْ4?D�н�V`�0Jݟ�6��)I�^5KA)�%�4^�x���J�k������kI#[ʸ�\��6�0֘}�d0�M��`��5����$~��4*-*���t�ih��+*h6�]c5���C?�r�C;]��uh��q��G
�]�-jV�����W��W1�!�ED?X~ԫ%I���x�7[���R��_x�F����s��?��V-�����Q�[��G��'�Z��K�����I�?��>�,D�x��	�
%.���geWѕ��Ja���zpǠ�)D0�s2@JFT�-?o���VPØz�"y|_�F��٘���,�x=Lgg�5&��~E�0�oh!�O!�RQ��P3c؋+RH��lҺ<oH�
��D�%����c�wYn_]^P�wE��}jn7�8]����ף��m:�_��r@�ހf�C
�(��.5��z�ڠv����Ђ����O���M��5X>��P�윆�_ӫɷT��?`P��Q�n�$Rr1�`�Ⱥ�Z+���1��}���r�ϸn�{g���p��KIΪ8YK�T��%�5N�m��=aX��*ѷM5�m���i�ۯ,��Z���ن{6�)1�C�g��Yݐօ�9���aS���Q �I�6 &A!m��v*O���(�Ƴ9�Fmޘ����E�(Ɍ�T�P6�w��7��&ȸ��շ*��� ��+ɮ�[1JM��g�P�LXX���X�b��_�܀=����L9`������buw���H#7A�c'�n �F b q����,8r����;ֶ��^z?n�����1W;���7�;�8�p���C��tz�,@�P�l�G_��ix��l�V��L�5�^��r��ZI.��Ǐ���m�=���W#:�����!�k��JT[�zc��hU��x�~�~D��^��}�z�Gh 3O�@�޽#::>d���:cW����hV���ဟ%�?��@pm���ھ��G�����G������?���ӟ�ɟ����?|�]���$G[�#ŖH� ��[$o5ݬ�N�<sa0R�.~6�-{�lTyPI�(���-�`�A(^�����m!�f��ti�wL�|���|�W�NY�%t�꒕��~�P��_L�tq�T���5O�+1
��*_�)��"�`E⽎$E���Ю�tو�ɵ��*�¾>ޤ����e���3^z��̿e�M�)U2�gF��"E�4���}��wi4'ࣦ���jZ��j4���E�ł���4��ĭ���5�Cr=�ǝ�]�ַy� ���:�Q��8��y��(�y�j��I7x^����A7|1ya���l��I��s�k ��X)r�T� T�s�D�]�]���5�&4w��
XS�#�v���1>DY�*$$��
z1�;�����y�zT,VĀ�wO�д&W	�����x4Ԏ��w�_-W�tP,�Si(7���y�Z����X��h� �~}?c��*��$������-`kJ��Kxߡ����%�J	��u:�ۢcH;�6�u6�}*��u���̓�6N_����X��L��A��w�� [��6Da�a#�ڬP�^$�BT���p�Z�&��u��mjtvyMPc����Z�u�xE��c֣ɋ)-���Bdd8�P7ɇh��!A�������D�����k'�} ���o|Pw�E#b6�}��'Ŋ1�/��"}��xMTP��:9��veAe�}N	� �RG�1�B�����Zd-HЛ���Zꏰ�@��s~��L��F�20�|H�� �X@U�ؐG�������Ԅ���H��;=j]ti�z!d"n!"�+��@*<Ui���h9�tpA�/���<W@���b��pH��L}^;�^[�m*Q�Ae$���z���`�1�Q#�"ux�_����%+z�{��U���'�*X(0���L��9�a�&�`�Ψ�[_V��>�G=nmse�FU�E��lJ�u�І�p��7M�e����Y7tу���`%O��x{��aQ>ڑy��l$fe���ڐ�6����o�vֲt�8��h$i����h�������O�q`�@���4���DR��9����}�[U�a�n?}ח�{�wLw�����������m�N��9�InN3���Ev���CVU��Ω��@\Z�������ȳ ��J3}2g�n�X�T��=��X,��y�"D�Y�U�5�<����]::ڡ^w��n�:��z,2Y��b9��ӧF��hD=�����ѻ�ls�ř�n7D={�Lz��~}��c)K=��>~������-�ԁ��e�3��e��.�Nh2��3DƱ��6�������o��o�槟~��st��5^>��K�F��o�hB���u
B*lD^J2�؂�tqH��l�$e)�T�@���/O�O����)+���#�����O�X��Ѵ��4>dewy5�����?���p����>�+ܓj�O�b:���)]\\��2�0�DqϨ�@^��A(���4b�S᪷��=���SO��1��7_6_�v�onQ'��U��7c0��}�g��z&]I�S��!Y��C7�Ob(�Z��x�Q+"���Gn���7j��7<�h�8\�`<���6
�%=��E6���"��5�;P�Y����3d!j�n~�l 2`K9A`�n�8N.%�1�ڬ`*B����Ӕ��Ӯ��ո6��B�u=6��Ώi�$\�R�#���ɑ��@sO�#��q�,�R:��>!�$`p�ַ�/_����Ԝ@�G�K���ABA���p�C�1� V$���1��`��� W@j
�@%=��i,�[{~HGqS\7�<�ဗ�O�����$J(���H��:�����������Ƙ�%D)\���������������>��l1�TK���(Iz���qB#�߫Y�r�o(�����<Fu�ݐ�:������L�'�����&?إ��.���=~��f����B9b���6)��"�L� ��r��	���*�Hb�A##_�ɠ� }MYA���1��x!`3��wM0, ��j�y��zk�GDJPDRP�OF'���� wX* B-�c��B_�(R���R�N�х4NYQ�.X��R��Z�k��*��O3WY���������x(T�6��&yu�Z@�v��,G�`�*�| 9��������x��k��q[�[,_�b2��ׯ���K�^[����6���@f|k��<��{ThoS�����	����
�zmtX��� ��q�V``�����\�	c��^GzIE��6��h�D��=�����ƮuJ�*�M�83���y�#�K��3#:mc@Je����E96���
�ȹ;X�D��^
hS��N��o��������AF�sn�C��q͛�)�Xjs'���M(C�Vp=�ہ<�CZ"��g���$���ݯ�<�nĉS��59������@w=��욷�P1vE:�N�iR��1�������oy4�?<I��vA��̿s���o��w�+v����w���ki�E�;Yi�tC)U Y�'�l���HQ�GN��!��n=����bB�y ��ݭ�Z�Dq�ރ.��=�ewY������<m0�"�~B�NK�;�ۧl{U%U�񮮮��xtt$6���֦!�'�����B�Z������+�ؕYTզ�㺾�?x�w>��w>�����o|���k�����$h�aq8�Pj]e�BH��ǚ�/�1����tMЀ5����Ҟ����@] K�l���c	���Ǝ�J��Q�0d������g4΅��ӳWl���_|Aϟ��W/�K?$:3�h���r�~��lش�|�ŗR�=��%mB�&T�qf�g�$��Qo;NnF:��J7_����Ƶ��(1�b�)�� �,H���R��`�xv�$�[�]bM%jX�^aa�@Ét5(��Q��^*R���N��}�	AaӂA�|Z�Nw��^���K�h�`p�OJ;ks�o���8m*��n6��;�-�q��J�,Mǲ
"ﹱ���dE�dٯ�8{�62�*�������&E�xL6=9�6�������*h�,�%C�$<W�Rz[��K��Go��
�y�V�͂-B��p��Q�{��54»�&�M4�u�ʾ�1O�73��I
R���8B�|d��P|�h���K��i����qK"c�NWk��5��E�9m3h��ۥ$\��ئ���"5)JF������.h4Ҁ�s>�R�,'lDu{e��xV��kZ��٭�w�1ʀ�,W�*�[Po��ٞG�Ge�_��ho�S�1��?�u���I�'�)���D%�'�A>���D�%�a�Q0a��o3^��2���A�F��x.��J�њ�	��r6����e
��)!�Z(�Mm��7�A#(I	�~���g4D?o�?I�J2AMAU��}��1Q�Xi��"���z��Dp�W*�����`<DC��lH����<��+bi� ��J��UU�2�x.��Tv�T`P 2�Af�����)˘`8�Ր��)͏�L�T����t���M�k���1��wG���5G+�E���y�c��O���'zmV����v�T�Wh�s�x��u�L�}���L�#I�B��P��/�8ɼ��̶��F�ү�pn��L�e��F]�ϴiP���;o_:&-�5:��j������T����P0�����F�7���g��}#�l>߆�~�`Y��ey��ϼos���F�����<\�ٓ�j�
�" ^l���wrױv����4-�iݱ�����|u���=^�w�%9�?��s7���_�@�^Λ/u�v�ND�1��6l��_6p�I��,:��7����9H��bs���7g�ה���k�3�ц��ey(���B�&�4�~�R#Q��N�����O�R��h��,K�.�?�U�ħR�i�_�d�-��_�r_Ƞh��DvjOac�����_����B�p��Z�Ӫ�&�7N�ŋW�m��C*�%��f̓�+����O>�x6���V�?��/_�|yB���t����s������`6 l�����d�Z����HV'Oy��]��J4_F����^���
ep@bVZ�%����څ4�׊r�1ؘFs�)R(�i���
���bD�oN�o����'Կ�E.�
#-nE�������{����/�Q�ˉ�$�U��krfsO�)8�T��~��h��� �o�5̧Ki�v���l�)AkS�O��?fb#fs��2d�e�e<�Ƅ�xW���ה!�A��j5a�i�?�Fǔ^�G�x �`"�҈&�`�ZˆJ�+��3jD2oF&��۠LR&�2�a=ҵNƜ���(�HV'��M4͖�4
�#r���޳���S��mek�����MI.��*$Q#��G�Bw�E���x��-{·h�!�Aw;m����
I�b��KG<`�@���H�ZU��P�D�b�^�e�����k��G���!͊�gt�+幱"d^"��BG�{���1=:8�-�m~�y�,S<>ϔM0a!�>�.%�j��U��m�Ӑz���]�d��a��'��4[�XL��T#��W��.S��Rg�M�[ju�hc������Ɉ���o���m�ऽU`c�AB}��	�?�4�e�k������_%^J��óH7ڹ��т�~[���Iȳ��TY���(�<D�]L҂DM��~e�-���%�P���TЇc_"��D�PX#ͫ$���@A�`H���b[���{eD[�wc	D"<� ��i`8��J��l�-�|�1j�y  '�)PQ�Gs�ǳyH�倪 
k|��JVj�J`d ���_g2c�q��O��t���2T��]�7�h����cJ�hDɒ���]���/P&�.�'�t=��zIͣ9�#��v����&L��	�C>g�A�Ϻ'�jӧ�����jC�K_|���@ qL�%4�鏑d5P��5�d���g���7sN@��S�:~c��@��n|�6d	��i~;�0���E�i���'\DiٍH���fFm>2�q3ϼ��o*@�k(��u3:s����Wr���ޘ&�R��d}g��<o���MGM}�<NN��F����K�ik�ao��7_���m,�]b���8c�˃A�����RPG����o����\I�7�R ��2o3�����8�}\S�o�^%�2#y#�.���"u
[�]�NH!��a²�sР����c-iZ��8m��[�9H�=:�Im0�I}����g��
\�~�@
�l�P�P�jiȀJ�@�˳g���)�o���~�7>��ޡ0a��|z��>����~�����H�O���5�΁�D���������7������������������������Ͽ���wy�0f@���J���x�ցg8�I6�P���PV����g�1F��n����.8�s1/������t���h� F���`�Yh�6�ڝ.����>d�)d]zE/_<���S�3٨x&䷯��-V~����I���>��#��O���T�
R�B)]�*���&ʌVE�ϲc�8e���Tl��L{b<a\m~�4�3lVx���`��i7�|D*Ʉ��㺞�el%��bJ4�_�*l�
KV�*�Bx�{l  ���c<���˳31J BJ�8>U�EA���J�-1}A��c�Z��wrk��Ld�;v�׬��d��f�Fy����"~Zz_����� V�����V�3g�ֻ����D)�
'�gM<�v�Ĺ�J��Y�]���I�z�V�9�z��D�AG
�q)��aC�3o&��V�.^��3��]���0�8�C�Բ<#g����)|X�I� �<IW�^��.=~t�߻O����]����/b>��Q=��`,�[�!Aaz�r��D=w��Tc��^)
����e�+ �� )���)�Dۭ�?ء�n�ڽ&�M>WQ���x��cF%�59|=/T25� �V��kx�F<���1� �p����E��Y'+a�
ْ��e������kE#����)�W�"�g}�)V��:x���"d�F,�|!�q$���Wl��(�Q#�!�y� E�$i�x-�M�ӥt� ҂�"?����"�� �c���w�U��k�/�s! �0�Ŷ���F��vX�l�&��Go+�ل������e�]H*�����ȯ�z��</��%�.N������ؗ��e�z%1�>�d������3(����p���Y̟�TOxy����Y>��|�,����^;X�ՖZ���wh)�R���H��<��z �4�U�� @ÉB#��Hq���!���S|����J6�����w���6c���GY�#�c�Χ����{��B�L�qg#+���#=��^�����;��}��>Oӱr�������;ʝ/����Q�-*I�b��lR��2ݗ]�GZı����v�ҫ�;�M�(��K:���k���i�����ܽ�����}�i�$�����6n=�w�ťlf77�l�N�E#���_ͥS�����a���n&�j9��� /ʃKD��02QNJ#W��B[�,��Z+D5�#���,��@��,���v
�i�W���8<\��u��b]� J�:�^z-�]�g�RZ ,�L�Ѧ�m��D�5���Q���B���ߡ�]y6����o?�O��g������Dl��t���m�5�w����~�u�Z�JD ���|��bB�銤�{,���(%O<mhŝ��ld�F����=�ں�#��l-� ��\�IX'�bCHB�$�١����G�'�޽czp�=z�^��]����Ͼ�&@T�����A����Ǐ�w�w%}�ɓ���Ͼ�_~�%������[Ra��W9�i���4��}��KH���B�����Y��z���tk�vT���Vq����7��	��8Ja}
���I1��{̋Eà�E!S�Ւ��*��^AjB�y�Qk8��vQ�.�5A҃ɂ���CÊ��Tiݔ��l�n�;�ɝ඼RAc���&��6f�����y�{;�{��J�C�4�jS��WQn�*1����*x�}��h���ȋ�����j��1�K��FUhl}4U�,���aרW$ eaR�p^���*X+]���.�.��\H�
yo
��!��f��_��D�@��fc��J`�z�����c~ߣ{l�!�U����x$�!�G4����K�}&Q��FcBw�ZU��;"<,`ct�e��,BЀr����z?�л>��{{��5V��h1��gC���lV�ZЖ~EȕE]��ĪTg`6��l���iP:��P!-�3E��[�޾-2��H5�K
��"��/�! � ��|���J����I��:�2�hd���^A����� Eja�־#�|lA@����l<Xͭ"���h�]���~�e�kF+Ip
V|e���4��>3��̇/�D�)�~1�z	(YW���VT��%+a����g|��)y{|��'�O�2���wʞ`��`�M�����ym0�qDt+��W{{TCČ���7ϥvf�Qi<%�u{��M�{��?�����vJ�V�%e7��Am�'hp(5l�N!ז<&
��}���3�Ϳ�k:=�P����8�5��"M�VlL�`��H���(���L�f^���d�D]*���}�ؼ��_rƞ�,�*����/6t���m�*�k���LC��f�F�J��Y�l 7��E�y���7F6nDD�қ�]��n#/�B�L��ېQ�n������_2����]>�Ҵ+{��|�WΈN�wfi�9�����(g�Z�����2�ݿo���6��N���CR�]�Z�d3�O���E�Tg߉! @���UŮ��+(��v�{�a�\���kD���bI��f���(̄Ś D��RY�R�\��V��kDgg'|�+iDr0Z��>c0�F£�DlT�_D|�ׯ_0`@o������]�p�����r�KU��m��NGR�0rݿ��dB�фvv�2�K����R��2���%>�D�2���L5�'ݟ��㟰]����������|��_�a�l�|5H�Q�`I�7D<�r�"J��5`�zZ�	<��[a�� DW�M����d!G�^`��(e�=�d���8�$�vw�E��P�S�	��/���g_Q��B-�æ'h��2��χ��'O��O�	=�����;I�`�ɒ�O4[B�ya�~J��y���H'recf��l�Ąp#���'��r]+sg�y����'��e��	�B�� �w��	x7Ѹ�������L�Hk��l��1 A� {V�]Q6N�Me�+�uC����WR	@Ɗ�P����CAIbo
��g
B�bٍg)zʚG���<Bl �8��&|���6񌢵�Y��C�	}�x��:��ኅ҈�~�-�胇By�� `�'�(2�"��L�l>���S� Pm-�6�e��a�w�`���DK
�<�U������Gϐ*���1�{p$E�^��a��BL0sF������xM�P�䄍ε�Dw@�-�RǣRp�Hہw�bR��?��-����A��I���~��?آw�Q��@nO�٘K�<�����,���!RQ����y��k��B��jhE����К7��5��*�5��%hP��͝��*�R(��.t�N�'*�:+���M�K75 �v�DƭC]g�����D�=D�.!��.	9��\�[�Ƌ��� QvB?�.�X1_4��c�vp���z!y:]�a�CI�Q�Xe�=/$���Ƌ����Ѭ���Vk%¬T|��ܙ������ 1�#���{߯��N�� �=4X�-�K��Ijr�*w�Ti󜗠�����fp|LgTb�QAt �ݠZg��W�g�38?��{�Y�Tig{���}��I�N��H�*�9W}i��.�R����������t=\P0E~6��0�8`�䙞@F�H�'��ɖ�,	�m5�r�~�=�"�����R���Җ��������ԛ-N2��������U�w��xyN7K�E�I���y��}W�);�U �a�l�I{L
����^ҙ��M{v%�h"b���J$1�y�p��(����ye6Ӕ*��U-I�H��\$o���^:9��:^��)�ݗADv�}��I�����[���r7��I�eӥa� [Dk�4��4m��|�r<xK؋�����u���HS�=�ȭ@�l�Ղ��&l�W|*�|@�FR�2��<����Z��à�j=D_$��1`{t�z�~���\��A�h8���	����*6t�k�9K>�ɗ���O�f۪A�n�$�����%ɀ�-�r�j�{ ��m��k��a��8
��m1���C'���˧U�]B�>�ի͏?���|���?�O��G����_��_����������i����"��;b��(�/ЃJ�����f��ޡE�� 3��$��D�:����q"Q����bH<(h���B���JՕ��{��H��n�z��)}��4��};�v ��j�b)�j�z���~�3��J���S6�FR�e�"^q�qI���zRf�4�3'�ҍf�s�J?�ɋ��M��ѭ�A��|��#����l������c�� S�57���"��Pë�62E��Y�7��h0���/����B���9��N}�\ʽ�J:9ڸ�RNzs�V��y�k�;'��S.*!�^��3,�-��E>Ґje�`kCb-ĺu�n���҉�Q��@F=j
\5�*3X����4��ᨳYX��ZU��N��z(=[^<A��+�y��A���I�p4�y������L��W)�:/�~Y��D�ߣ�s�f0>��w�֤Ē�]�Q�R`Pb�P�{h���^i�h�`�z{۴�{s��d��۪<�!Mg#�_��9v��H�%l�5��x���
�X�V�<�Eߗ�%6r�sH����/Ui��*��-2ƱK��@���XrX}̹T{��G���=~/�|��iZ B��������|�.�	(S0gE��&`#ۣ�D x6$�ԷD�幤�a��X*deA%W�l�A
�5Ԥ��	�k�>��S��WPĺ�� E3�K����$y.�D>p�e�cE'���&�q�rQ�jgׂz�Qc�U���Jt��3p"�B� �'"�FmX��|���)Q��2X�f`���x�����@��g�QB�&�b�Ҵy>.��[����Yl�䷈�;E�#}���|�	U@������Rm��P-��ٷt6�5�(�0���)r�`w&)X�B�P�w�Ӗ�C�k����ۢ`��rA��3�_/Đ����8t.��JGk�?��T���J����{�D����wاǧ�{����@Ē�lx��6.�)����y7#�'���˴�u9}���nDG��=���(g�:�1E�2m��V���Ʋe���3������i<^�ZĤ|�S�ق�H:\�@��1e���"�jH�����c�6�]�G���`��0�m\�pTjd&���ct^�|�k��C��q��Gk�F��T�p�����n�I��!�e�P�˹E�F���iκB��u��A&����8XJ�?�p|���Tkvhk�K�rW�)Q+���v�+�$�P���4>E��[t�>6�ܛ����W�G��[��h���uw�Ț*�&�c�}_�"��$
�T.���$�n�`�=y}&�Q�	0M����D����Bz}yE?��ϥ6���g�%�*M�>��/��H���O�T���$�&k2I.�]�������Be�s��ի7�	���) OwI����f�]7@F�vRq�[1>i~dI~��h�M�7.��P|�.�((=�`�8�
��j���-z�p��h��wN/����}����B�C�
L�+P(/�/^<���|%���I�r�G��1%�	���.�M&�sc�9f2$6o�sSg~���;����;q�ρ���W}gg��g}N�f��+O6��g�6췝�D��ڃ�"g=a7�P��4��M�"��]wz5��v����Y�p��E ���실yꦐ+�ye�$UܷA�e�2�A�MSp
Mx tG�?׻1�y��Un$�{�6�(��p"k+&S|�9N͑\�Hl{bؔ��GO�'�n�Rh�� ����[��y��BW���m)ep�5��g��?���+���S.d~�����+6��4��c�Hy�M�e>ӈ�!V�� A���\@}�O�;=����v�?�5tGxJ�V.S�Y�R�*9�[[-麊�����Z Ü��p�Z��|Yk���s���k,,w���Y���9�� �:+z(I)`m�_F J��,R�ʆj���(c6dYP�#V
��G��bB��بY�����U�x�q�ǔT����h���*	�ߊ��j�F�
n��M��b��!�T)�iK?+G�X��R]�P�F��� ��Q�K`b��r/+ԣ���W�.�y�a]|AH�i��g@���ʴ��Yz�q݁woE��t��`� ,-��/$��2"K�G�|qeO)`.]*�,�~W=�`d��<! �^$�RJ��H	�5�fp(=��u�쓵���w�G����Ua��1xR�����^�΍�z��|�Mq�~�V��W�j��������6�M�^����]R�ڢn��zc��r-k�{���у{�tqr�Ɔ#��i�@)!遅
t���g������V#o`	+/��r��i����/ٹ�k�D�c��3鶑n�&�zU�ж�*H%�K޿�NC�=VH2����w�h{K��K�1^��#�:����.���ϓEߑv����Iux��$�b)���Vǌ�#������Y��%̵��,�d�J��8��*kh^�P6x7�G�s¹���Y�#������L��^	�)���=�<s��-��W��8�����\6�0Mj��I��*����Z�(��g2%��*�ʺ�0(@�on�X�`|\�����+� L��u��{�����N�ud��X�$���������Ͽ���`2�KD��4B#��b��dJU3�@�VSe����*�m�KD-�X��jT�d��H�P��]{��W����GTf��z7� D�//O���%}��Kj4�B4�� ��E�U �5���>�i�[*y�=E��;��v��s�������������w������/�����''',\o���(!��u���Hv9H��#a�ܸ��-%i�b��8ƃO��TX����wBu�I�w���(����X��4�����|A/�yJ�Ke�����0΅���&�?6��Sd"t� ң��r}1�@��poN8�Ƨc]DYO	�!0*��"�o&|l�V:v���,�|*�X�ۨ�ܡgYW�xf�e��� Js�y�ESɆ����'#+��$�}�8��.!�4�Me�[-m~sp��6����sj�X��i��p(�h<cC0��^�t�!@���'���,�\�����T��� �e<�k���{b���D�cD86���� �*<x� p����2֚>��,|C�k�oCܠ�h@Rhf�iY�*Yl<���-"��h�A��E�9�=��+��?��b"�!T�Ƙ@��	�~��5ņޥ�u�) �k�XI��zo��h��K?��v�v�Z= �i�HM�RؔP����j�u{R:ua�Z�2��t��)�X
uk��+�%j6����	ۇ�3�]N�X������R��@`��@!x(�?�T9�"H��EvygQ�%��l>�q��)K����H]���B��&�R���O;�{Hmc��T+�x$�Y�� �c��#�����=��Eoy�y�búZ�Pl��֚��������]t�_y}��Gk)��zR��a,d��Ԗ � W9A�_���#/�9�k�_�}t<�x`M1����!Q�hxY�j|&x������I��U>�/Ri ���(�/K$:�Q@���_K�&��`Ň~)5>���b��k�v� �c%^X �%"߬Ϩʿ�=��+:�;�`J>Z�R�.S�ӥ�E��9�??�f��`�"��f�%��9�(���.��邏-���z��T�H�u�-"k(�9NNXJu+�͞�����Lľ��ۈ�����I6���U7�FD�SW�T"����$F'��~ &�^��M;#+Бu`n1ә:TrM+{o=�C6B��6��9ۜ��}ǎ�i?oJO�+BbI^,8r�0����OGy��VH�蔾_Nb��6_Tb�D1����)6�b�C�̡N�)��-�Ki/�g'eN���_V_� U�)}�+;�C7�w������_��o��u�S�F�E�V��?ÿ:z[Me��=i���E�g��`?,�F`� 2��&zm�_z!%4�h�B?�1�+U�������`�)4��E���V����_����^�8��ˡD2P��r|��k<�U����D���H�E[�j��:�u.<P����ur"�
�{
Yk�HF�Iz0��:'<�?E���%R�.��/�Rc]��R)�3 �y��%u�w�����=���2��rY#IBlM]ʁ����G����?x��w=��?�iX��_�~��ʱa	m���8B�<�L���T��έ����=�V;����BƋ�8��� ����yt�Fb��0�c�Ê��p�����J��Sz�������%�]�2�����u��
/�zذ1�F�DG�@E�Γ�B��h� Ұ0���P� �i��<�����fP�Z"�J�6[�ȈSo�7x�G5m��☬Y���3�\#@�C"��~��,��~~v��PQQw�oȆp0���x����</h�#h��x9��/��rovy��=�BZ�q�(5R&
��D���ͱ /UPq:-i�\Na�7���~��3=�1�l.�KY^$ja����J?jٺ�K��9�Q#��N�JW�3z�m��@�k���x�`�<髯.�'���B�� �@�h=��F����+���{�'�4��D�B�R��@�=�mY��Ԩ����$�f
ч?<��{{��;���hQ��A�QxpP�=��0f�^)�5X@U�%�4بc�ޗzW�+"_�e����T����!����΁��p�khA˵6�f���
�&C !D�/�)�x ��H�	�h����-)U,��B[�kh-)m�44�W�z�ѵQRu>ĸ�� V`|��y���Wti-��%��t2���E��+\��D�@�?4���)xT��T�)�c�� #b��00�M�!rM)FzW!0t�E�[F�u"�jR�Ϸ��k]��k�
1�.�](�L}��ue@ ƈ��6��%S�)"���D~|��I�LD
�#֡������� "�{	%�5Ҩ��˚��N�KՖR�C���|ӌ瀟�ШS���
����<��f�
F"ӗ����e�եq��k��gZ�Ϩ�-����l]̧������4�Ş�����D8�`Wu�Ci�S��8B�t�|�@�nC�N���Gw9������9oH���D�-0�쉡s������C�Nd�g�TFn[6F�u�ݸ����,�Y���c�ܯk�k�)kh��� b�x�ٛ��-/k>	�0�V�:�?}i@B%mr��8�}"���5��NHF�1+��tn�$��N���A[���m:����'Fˤ�:Յ\��_qz��[R1������e B�_�1��<F�fHCj�)����h�"=�pd#���\�H^�D��g��һ=��pH,�4� }��a~k��g.Y&V���y��#zx��f	Mئ����ӓo藟���/�����zM��T����ݦ��sb��:�ls^7+� J�>X,������!��m+��Zӂ����J�B"C���$}Zc��n5h�ۖ���1��$�(�d��V�鈞<���?�{���}:8��{/�M�kV�&���9|�$G|���ѣ�������	��o�3�#���h��K�J���lʫ�k�"1+ec!���.�\/��Z7�ܟnT�N6(Qw��v<��f�������>�j��cz��g���_���g"*�R�"A�P��b]E����T��zkJKv�����$ �$f�!�}���|��5��TL޾��s[��#Q"�u<��v�	����)-Q��|ka.Bx�r�Ђ �kj�%1Fj'�A����о:���6b �Q-0e�\(j�҆�# �<�Q�F/��zǺݮԁ�q��bg��b�����5u�!�j�����y�0�I��|��F���,�O)е���Ҕ���*;�͵�FA��m/�����K�
� �c�fŦd�90KHi(�F�52�Ȣ뎬A���}�4���Ɍ���� ��GH���{G���d�`��ڒ�jA��Bj Lq�#6��/����Ń;�H�0�%2�y�#$�\P�2x8x�G{�[�� ����Fb4��{Ȇ�5Y@���Zh�*�y�%W:j�E�X��BiX.Ƭ ��Dw�N���Z���>��;���=�\Lx����Ų�Qi|���$�=a��qLx_6�9jABu���|��Q��Qz(ƾ+�(�xgy��K�{:������"Q/f�\ҡ��PC/T,~3�q�@�E�e4$r��<E1�"kL$ �piF81�Bџ2_n�*d���� ��#B�&� <��|-��k4�C��<x}� �"O�!��94eʑ��,*ݴ�T@y�ޭ�fN��ŉCI�$*�)Hkx�cD!j��gV��'�Aמ�h�\A��׵�( ��C	�4�y����̃�$�7���ˀ�|������P|�� �f�rS҄g�%}��)Sm�+� Q�g�P��AƴO��^���JT�x��T�j��
�Ǡ�+�)��	My?͖+
M��"m�XSN��:�Jr���kف���/~l���L7��8�O]`9�u5 2'��R��6B.rְ	JW���>�u
)չ=�ª8w�.������s>m*�ϒ��1�UX�,K�~@_&6~�c��p �JI"lf�$h��8��5�+rN$�pL�sz|b�+VГX�d.����[}����7.��{,���2K=���B9E��;D�n��̶k,�{?�t"!H�D�S��>.��GA?�cD�5�Q�eG�Ѣ��R��6����[���)����,�x��J]dn�Pґo�������/��WO~AϾ��.N�FB/kq�w{m��k��g��$TԈ�}B��P�U�OGĒ�KqA@
L��I�Nv8��v�dR�	g9l^D��_MG�e��!�lcDH�RK�Z����撌	����~��|�-z��)u;M��٦��L���A�::>��bi&,2jS�@� ֗�z����!�}��ǿ�{����|��_���?��?��?�������C�q͊ԭx�n��QZ���8�¹����oI��"�&)Ba<P�D~��M�;[��l�����W��_����z,����`�)D��Z�X��y����PXv$C"D�v5wyьh1�I����}ڱDV=�# 9��9i��������Q9��\�7b-���i�H?2D��aQ�p�f�&�í`�"9�b��m�\2�=�6��'{�)*�j���y�6���hK��F@{�`�i|(�G� ��p�1�QZʷ(A�H������FQgCC�XV�4��GBSE\��yIW�a��9�x96���i��FN�l_�l��|�J�)�Y��"9�k:��dh�Jb�j^7�Ky�?�>���2�~!6s����V�0�^WW&tyէvk�z�;t�ۥ���lHg痴d��� �R���z"��T(��_��	1 A$tz{;4������K֙,��к�8��pH�^�z�H���pu4�c�������P��^b���'�@��">�F>�D�Z�kW���"�6=x�MG����Ӡ�N�����є�nSd�V�?a��8^��ϞS��P��@�Kkå:��Sb�#4����5<����=IMKȜ#J�"x�+� 4ݯ֨q$�	�E:�����Q�)I�L�����6����Z�!��+:B��)���`q��uE`�{j�����(�g`������IX��g��g�@�v����:��/?bj��=�3Y��G����w�(��y�b�����r�@6�CS3�:P��ԓp>�4<�.�q�Ra�PI#T��*�Ӵ���x��x!�����"m� �{�p\����$y� ˡe,?�R묆���42a����dz�@aFh�g��jZ�@o�f�N�_�'�Sr��h�{��ޥN���S�x怕*j�jtx�̀H�����6B ��d[��i�M#ꦍ�zoS�
�3}���E�՗���XgW�DkdA�%m�N��"r�UY/��$Ǝ�~Q����/�F%\%[KӨ�C���}f<g� �u�>ˢ&���Wb�g��-Q�<D�N���a���S̅��L}���f��o>5*�'��e���!��1�z����pR�Z�+�i��a���a#�a�m�w��qz�Z�3���	o^˂��5�����b#�I�H��v`��[!�`sEj |g)i�p�R��;*]��Hd�ǲt~q�rg�i�,Sf�{T�wL�����u�'�aXD����V���pEu���'}z��)�~�%��|E��%M�v�W��a�T.���)��%*I

>��DJS�^c�i��0�8ǣ2�c'�!D�B��b��dmF�6�cz�(�-?���gQ/��أ�O����y�t��?Ͽ�zE�n�^� ��;�����y�c���${������"�Dy��N�m~��������ˋ�������]i��IP��*�51���Al��+�$�8��qZ�_b��u�Z�m�p�r����z�`Cu����aeP�b������+ZF��n�� ��'��n�wr�\J�Dr P�̓�:5�L�3i7Cs�XJ����&����,`��].�c����"ߕBε��T,��ZZ��A����a�&'�/R�AJ=�
E3��A���qd"�pJ�A
u�Ta �	�Ỉ\���k�k��7�d������B�i���8����֦9`�jHM3��ؗȦ��3ʛf2#oD@ZM��ث��Fl\_�I:R����E\Gn��W,Vk�T7�M=w�+搥8NW�@Y	o]G��pC�%
2�;E�E�q�P�@7��0���=1����Iw�၏U`��I��u�K<1�p�I�Tqb���hox���1}�˯����Z5�v���r��_�5�6Ы�%����s�É䚂��k&`qzzB�z���z�EϿ��4���=�n��s�?�	_��wyɀqܧ+�} �ᵤ��ښ���'O����@�2t�n�k>����*�+��:��ο��Ex����������?<�˅�ހu�YgÔ��`�E�����Z�8)	�w�T&�E$+� _A��.��l�H�*�m�c��U�NN� E�*���[��JȀ!�j�$���=����ܤ	Ʀ�=��+��"U���C����J�	GuM�
*|��X�>5x�<�	~\ m�b�5�?�s%���lu�>�V�\c`�n�5I�L#�8I��1�"�h9$2�R-Q�����UP\nk� ���P��Z�~��J��1ZK7��_�m�:�
� �����-'+Z���R� /�I}�ߨPy�J��m��%������b��/�:�Z<�2���y��h���8�=\,*��K��x���t0ќ������������)��5�i�e6���K2���L��
+���]gH�l�5��ʧT�5�F9�kQ�������5"���0�T>;����fU}� 7�In(��$�y
��H������w���^���;�2Ġx���T���5���/L)c�l�Eplz�ƥ���T�I��`*عfoD6��Ωb6��l>ǯ>J�.H��l��$��Y��2�J<B&�����}�R��jq�&"BuG��}��DSY��a�M������Z�'_}C�;;t�`�:l�K�h�OTǫ���>ˎ}��K�8I��)�笧�"��wK���:�) u�r��_Sְ��8`K���)����BI�"F͵'��@�m�%�
�ǾLl�IB���s��8���Q���.�,�c��'}�٦�ӍFKR��Ӊ��0\Jo�o����S����>��3���#�����}�����PHi:,ck���������x�v�_w�ww��?�����������#�/u�`B�F9
����.7'P��MQ��v8�wRБ���	���4iu����z��}*��Y��@�.�h�C�������7�)��z| ���� �!��`��&�s-E8ꉌ����d2��`B��X<�DPG/��l>�	��Q�Wd�C�.�+)��(}'ө�;L�J�����8����y�]L�6���fC�@��ٸ����ȏ�f>���J`���©�e�b��U�k2QQ��)-6�Q.c���c�G�Y,�.&��(�����Ǧ�t��W��#
T����V[A��~cci W��%��S�鬕i"0`�ї�2�+͂6K��	d�Mhse&Ƈ�~=SΞ&S�_��B��~��qLNc�� �S�M���Xr�،��u��)�B,�{�N���lRe|��1���k6Jcz��ϩ�B��c��
�k�xB�z,ܾ�f��-��o��4���%j$�Ъ������R���^Q�z�ۤ�N���{��jR��B��g'4�_P����@�zN�b�O�%W��%�#����)�.��%/�9Šcf���S���7�5��7�b���7Y�&W�`]��/!���U����𚯕�wE�F���&��g�JkO wd�!-)R&@�+Ɔ�J�����+�(1�t�S�Ҥ��Z	��u�)6>����K������5����Ld-�("�*	�H�z_#�4�� �V�i�
:�"��:C�JT1`��-�U�-f+��X���N��1�d:��5�c��8T]��`L�t��W#�ϱƋ�h��QpWe�h���n���� �^� F�O�?;��4LE�_�
b�D<Ǩsr<M�
����p���Q�
�,s&�|Zu�շ�T`�J��Jt�K��P0�w���G;�-�x_Qt|O��)[�fC���*ZU�7Mz����/.i�:t�U�RwzJ!DX�T�������л^9w��$y3HQQ|�x��HF7[�Ek���nD	�9o�U��6��e��
�Ոb�lRsq��Zi�ǖ�v\3��P�������5��Z��FQ�1wQ�;���0�������ACZۧ��2,�x�EV��ׄaK����g� ��O��C�,��L�J��|���@��s�h��w���~e����$�똢��Խ���jwho����*��>���E!��V��5�GB��ѣ�	.���D����a���d��>;�����s:a���ޑ��6��ЩPُ�����	=��	�~-����>X k��Cj"Je�7H9���u,=>`�R�Z߅��rUlV�+px�3u��I�
�ңK���!�D��RV_KȖ���F����]��z]!�)h��N;���\b?��]�e�h<��W'��?��/�����>������`b[l݊ԅx�s[�X[B���d�8I���X"�p2�<��]�cC�jw��[(�6�U�B6􋩠��L�^Z{/
+�R��E�������po��<ƌ<<8�J��l����h���bq��*1�6V�Ґ ��D���EKJX� F�a��@
����K�=�0k�D������,��u��T��(M��e`���X������E�Y�?��t��MKa+�M��\�3��a��Z�a�IłF��g��]���wM�W�д6�Q!���Z����S����/��Q�|�<��/Bل���Ij�zC����3����,�\�❣I@����y�o�RX�^C,S1��%������< @�Dâ(1ŷ
�D�h7�*1</)���"����ي��qҴ	52��cR�L\R=��\��!0�b�4=�^I�"�l�$ �5*D�'�9��Q�6-�<��8%3����Kr~1�����+QH�w������'B�ݬ�Y ��g`���y�x�G����lL�� /x��Xxo������ޥ��.u�l�!����|L�}����Ų+�����KF ]^ŋ��%�!PCz�1�����0��2�d��ϑ�vݪ���PɊ��D�fَD%�ӊ"t��%���b�1_i(Z"
Eߤd�|��`�@'�x�SQ�DI��(I��z#[�%��D����H���A�)8���6�b�ny�r����T�����v�5U��w�6���ł~��x� �=U[��[�{W*�D���c|�-y�PT������W�WG���p.�!��3�fŲ�}�\h+C�Q��v�����T���C&M7c�59@g2 @J��+҂�����" ]�/@��b!��臂�(v�4X�XV����|�,��ڲ��ƫ�2��j���=Z�~��)�b�:X� ?���2�!�g�E���g�i�kpȲrL���	�S�4�>�������|(�v0�!��w5%T���P'�R�ߦu�2g�N��+߇"sj�Α3�S@���5�c�+�����K=�c�8�w�Hl�"�nj�C�Ύe��󫱡]�c�Ҥ��/��í� +}�7�n>6�ol7@L�yf��i~g��y��q�-SR��n�9�'���r�~1ћ4��7I��oI�#�����ޘ��ow?���ӟ��O2�D��u��RH�׀鸐��R���x4x�~���G���.�lo��I��4AM"��͑�h*,	������KJPL�}�`7��A�C�3O����ڝ&�����:?�/?��N_����%���D�;�
봒8��]�L���JE��a�A��5\4���0�#6���t�u������C�M��R�bW���d!i4��ܴ=�%�5�v�c��,�&��PA������d����u�h\��1@�b���.�����B�������g���e����~J?���[��[���>0)`���8��4�� �Z�_| 6��c�:`D �-����
`�-�]D76�E�r��DM�l.�v�z�����_�����G����1�j�l�hւ���H�zxǵP�>�"��@ך
`;�ÐRF'WY��X\S�4Z�D�B���蝀���18����м�)N�ZU�.4�ʄ�
"�bq� �0��.i�XI�8�������XB_h�Il����x�]�H���z�R�T3���c'/n4�C�?DRp�O k��C���Ҥ���x�ib8r��t2pGO'r�*��H˔��3F#�c�ȅ�O���f~�����Qog��e���7a,��1/�����H��jWDN;�WlC�ځT��	���4�a).s>2�l�a��)�c ��/sr�7u�$f.�3oC�����\ �W ��)���Ň-ѥ�b�.&�M��mmM���"��x������(h\1��z�hȆn�.e����GR�\����<Z�Q�i�`4���e��&u��T���tlQ�I�Ug@_��ރ�g3Ȣ�:�:j<���Fxx�;lD�1ho�J�4�MH"�s�P]H��l�8�6B�����A`��5|1�����������5Y������n��k�/�HM��H��(4G1%<�
v�ڶ��.�y�I�c5�yܗ����iw$Wr%h��ؑ�D�܊d�,��G}T=3G����c}}�FR�6U��&�d�	dbG��>v��s�@"�Uj)x@$�_��gϮٵkSݸ�KՓ] #����,:�����Ү�y ���(�(!��3�Zд�� C�Y��\�Y75c/�8Φ���ٟ97��#��l�:%��E��Ӊ�d �A��a��n,�Ռ=Or��.0��V,�d}S�5v!�C��C}�Q�G��Oº���s�V�L }v.�uwf~� �[! ��c9�u�.zީ�	��R*��e��5y��*/���#2�4\kS+ n�=�5��bf�U�f2�-jȡ΁��Od��6�8�Ɗܾ��@ȩ>��S��c��
j��1fsܘ�t[ߕ3�7J���
<�?-;~u��zg�u�w�
hSA�~}!��~�Ttר��[[H�Hx��²���/P����t�\��NӅL(6���J��?(J�U�kǬ�9�>��|jha+�!�q�-Y  r[.������f�Xs�:V�UT!2	q�0C(O\^h�?{G���N��|��{u^�^�B	D�k�ǫ�+�y3(W�C �@�(|��]��^�_|���I��Z�S9?]�S4�==�����'s�ۃ|<�2��q������ִ�6�Ŭ��k;�MEo�1Ϟ?�=Oܗ��Ƀ��B�b��~[�32	���tY;�FS����V�y������@�J�T�t�͌?9��.�uOꁃ0�bfao�͜��E�����c��?4jx&C�����>���U�\�``/0W@�]__��������k�/	���������z������nɭ��regK���*� lU�99�N��:9k ��e�%��(�)]-�Ֆq�[�y�X$�4���d�M�
S��v����7nQ����^�:��5i^QGG�eW7���UF2ɕ�k����YA�]G�4�����1c�'�M�43
Ap�P\�b���6#��)�
��JO�lmmZm�=��N�뤴 <L��'�b��\�ʊ�mf�~�H!��������|��a\q�9���=�MPԭ�/
`q��d��vTN^t�F6Ê���
h�eH9#��x�K��6
�0� �8�
�iK���lf�qO�j"{`�� jT�P�1�d����+���������#9e��tV�t�:�ؼ`Gk��~-Oj>�𯃆W[E\�V#y�m0>o�8�>
�+:C%�������'GsF�ͪ7�؋�Y&��K?:RK�[:)?�~Bd B�Q��YkJ�"�k�($6�&P� T[�в6z�v�
�o^ߖ+[�j�7���+Ҍ�To�'���ۻ�{wWV�VI��9z0���g�~q|��ǆ��E�{���{��D��鳝G�V���*�c�t��)0=QЀ]�y��껐���:j�0W�إ3R�� #ؑ!{�y	����( l�L�T��cN|1*e�9�tfL�J��M4��T�8�� �U蘳c�U�c��}&�D�9�3Mi?%9���ڒ���c�:��}6p¨�����}��mn�A��0�y�c �~΄�GĐ�׵���y�"̛�^f�l�Y�Xک���Xw�/
E��5Cc,8�
L�S�����2@���2P��Ou!ED���&I�:8���������V��SJ21*>�����2ƅgx��u�I���h�/=�� ��s������з�w4H�<::��H���VR*ȁ��f��U���N�N���tr��,hMJC����2�/�dc�y�<~�B���)H���Y(��!Yjc��|��8_��r.�X�����ցE��M)
@�F�
�����P���K�i-���w!��9�b�=CY'�)B��������gZB����%2�al��-9ڥ�}��_�*j�����_�#��Ǽ_������o�XQT���R��.�).�*q���epp��]��׏���z�ٯ��w�J���O3��3�u#��$i�%��MY��8�
Yk���Z[&�-R��	�ι?�e�NO�2NuT�l4Z�H]�������)7����􏿗��}'��{
0�ݞ��~
`��`3�ܲ4S�q�����/�c3�[�=w��0e�瘀��78g�p쪮�/�w�'��ӛ,�����m��RdB��<�=`���9;96!H�7�:5lPp���N�ϕ���E�4>w��{��������䣏>�_��fC �P��s��֩�84h	_0힐V$�>���&16kv</�m0���䩦�܊����Tej��#��6-f�(���ȭ�;������WG���r�d"��t:��[]}��qTV�{R���p�!Sj]x��Z�hgF�p$I'�0�	n�e�b���U֌���yhm�/.!7��v��担��=��W(E|a#�*� 2&/�����)�,�y$pa�>����9�bx�Œ�a�ru�^r�Ѓ��O3J�Y&���"�_p� ���̔��
�T�M�� ���/���%PD�X����P������e��T���ڎ$�5kV5HyJ��jCf��'pmעb�	^{CT{oi�2��9
�$���5J%�����moo���)j���\p�Mb���Fr��E٫�6��d̹41�T[CN�����f��s"�3
9�4��N����g�s�+w�\�;
8v��˝;��FL�X���X���c%�2	������sy����!��:�}u�6�>����º7f� bSӴh���Q �[p�"6��y [X��F� y[��v��Q�5� !�i��MF�{(<@����Є!G����N@�	�{Ц��A}�����-(%�x<�Ia�/"��Pd�������!���6���B���VĢH���"=u��|��]���FK'r�P�Z��A��(�+��h%��h| V��JO�x5��j�(�I[��B{�'A�B(nA/���Tq�� 㘢YV���v�sU��W9]�pD�Bؐt��pp�F�SP�@�B](%�=�iba��:���nBY��Z��4[�`�r��n�ٜ):���"��=l�Y �IZR�@���6�`�Ɩ�L���}D���^j;M��NO���+j��?9Q;u6�����k:<�kW�����|������L�	�C��[v\��0F&�a�ehm52�5'2X�0;.�m��/ �����bpߒ�U�\i%k1��X֢`�#��F�������γ �(hP�P�y38�1� 
��e�Z5��J��6F	��/}�[I9@Ņ�z�9�,�e�+EE�:���j���=Qw��ߣ���ۏ\i.��ʏ�W����-m��_�.��H)g�`��HRʵfCA݁p
��C���u��=݋�^�2�ӹe�!�M5@��!���і�&�(�hg���{����ߗ�?� ��}-��������������;�;���X����t���/;Fs����,j�|��4B�n{Q�Hh�,�LZ�0ǞM�솔�`Bළ��AY��X�p3z��%�K��f� ���A-=	�Y ]�?�}�6��#� ���萌�����ͷ����/?<|(�|�|���r��Uj�uؽ�W:�2��A� �h<�Q��}�|����ҏ�P �E���D�h�-�9�z�
#�;�U����o���7n�[׮ʚ:�I1�BF(F1�$�%�OZ�t��ʥLU�}1d,!�s�`Ӈ��qA�f~��B�5D��Y�����C}G�2�i��J���^ڢ⡀(��٧da� ��YQ�ɷ5k]��l��'0��m"b���yHL�,�Z�O��T��^���u�+֜[V(q.҇(�����Ŵ���2"���.�#7����Y��jD�����Ky���<�Ggᡜfr|:��)DWu<�1U��)�ϡn�{�N^'�6����|aK˽$6��ء�f���mmn���֦	�w�g2����-�EFݘD���4Sa "H-�� �Q�f6̃JS���)��y:ެ�䴎������;��;�t\QGj]n^�dã��LƧϥ0�N7��!q{���p﹜���jl�������t<a&�9�8�l���l��7EmDҒ�:��J��d��h>�6��vIA`���HO����2��aӵ>��� ؘ�H;�� �����W�N�Bsg�Yp�:�fS��9�0
rd8��ք�nP�ff��D���ENǃ�H���f�"텂4�S@>THԔ��J�t��L����g{�T�5-���8+X+蟝Q  ����iҍ�NSF��)�ex�M+R���E�� =:���It�p+��f�,������~5�X#HS(��K���n�ܘA^W�æ7愯��=6p�� ���E Q��IʜׅM
Y>�J E���@���T7���<<���պ�" hb�U[hR����\�o>0����'�'#��:��<z!��YM�̨�80@����`]��~tmsM~���r���	�
礇M1J���Q>�5�"���N�2s�6��T���y��$�/Ǝ�rƫ0̅�����j���ŌU��R媒��.4�EE�H�v������ޥ�EJ�P���S��~F9L~?�LPx�G��屪��x�<��\��&
[�2|�U�cyw��>�ϛp�@Ǻ�N�e��" l8�+���{�q�����Z���5��N�m�<��n�ް��Fƙ}�؃'�.X2���Z�p��hp����V��,��y��ܿ�P~���Ё~���h�ߧO���%�ǯ���mkց��PŃj*��l��N}ؓb����%�۱e�E��Q-�U����	�@����z$���}:�'����xՂ�Ȯ@��R����� l��9m��?y�}���HZ��7r��j��������% �2�� ��m��� >�d|n5Rν�ܚ���R&�P>�bĲ�`d�'@4Q��3�i�[�T;6tH�uu[>�sW>�}[v:( R���c�?��:��V$q�q���)d�з��Vp�,
e�J�"l
0����F���o�3�T��@�K�"��^C�i�H\�k/?>@���E�ei"3օ�u�&�yt-Nl�嵔zFU/LL2Kɑ:�^ �݃m�pHP ���0r�
�ʄT?��� �2EA�1���˜�
W-#.t3�L(��z�� �o����3=�����t�@��#p�a(O����g'
H&�d3�
eC��(�,�!��^f�CieT�e9F7����N#.� ��w�0>1��D[�n��[W�O���NDTnBqبK����/2�k�)�(]I�H� �ӊ��c�������>�o��խ5���&�ӗ���\F'��ґ�(r	�sY( <=x)��HfjD0�ax�x�%P��dhN<X8PI���O���K�N�w�����#�pN c��JW�Mf�f4�A5d��u����ǧ(BcF�W1k) �����6��[�6.d�L�-�� -'ώ�j���S!Ɛ�:�(f<�ܮ�@30��Mn�2y���iǜpeț�p�ǪO۞g�ϼ�����e<Rf��錵59��N�	��b��{B0��`�N�E�B�0�b���1��ް��:& a-A�B�9T��dZ�b*ׅ7�H��9ȇ2� ;m��H��9���>bNӖt�fF o	yG(���
���vj��
�#�щ����:�5�b���Eb��3-����H��P��>�=	(���4����3�#iXztDL�Ȥ ��dV@����ֆ���:�_�Af~�ʚ��P��\�O!g��A�,��G�8V�0wܦ5�_��w$�^��".z��Jy�ĳ Ym��7��Q+.ǌ=2�k	Ȁ����$G���1�}��w����_��H	2�! X�'�4���u�#�Q��x�<�,[<���Z��������������� ���Ra�,u-Qf8��BS�(�>�]Q�jY��?w������ "х�<�T�<|�X^TPڳ��<EpA�h�R@;���e4��`�
v��A=ғ"�IK��c�i���E��>�~����	��{�ɽ{�嫯�����J��C ����ڮ����F�
��>�z�������fv_�ں��/���{���Ǫ�(
��k����H��B���[���>E����������3�(�$lnU� wq%Q���	�@�~Ja����:�[����)����y���������s��/�3y��7�m��p�ϭ�2
E�#�xB��ĩEW���(���2u�lԂ�S�(Ld���Ɛ�$N\Y8�=�^�-�-yﭛ���w�4w���&V:-��7ڝ7�46�K{�Q�r���Kj;g�$8(�x� ��a4��xV&�kV=%\u*/<rc��L1�k�Һ��K�AiV� )w�*��<lr����ȳ-������<-�%R�K�C����E��p2*/�E�����Hb`��Ms�|H�0�1k:UDF�%�i?D�1�ܝ�����[2�g���<x�R�Y{*��9��^N�ĝUi�6��+��F�u��+!�TN��e벐蕿��:wѣ����SD���F��HC2k���\hP��1޳i��->��S�Y���"V�Nw�ţ���q'8���6����E�ܼ*���y��:�WdwcU�W��"���ǲ�I�M	<��z�35�GϞ�����X�����~�۬]��AP^�:��:
o���gt�bD�0z*h��RG��paJ/�0Z�!C�N!��fL#u�Zj�Fjtft�S�(ثxa��Xp�#3� F���c�N�oY� ���zd5 *ZE�Is�٘*TP5����fH:����2���&���Y Y��eH�f�\)�jh^ۓ2�/�BAE�)�2:n	ڛ�3�@���h��"k���aόFaQ�fG�7�2�1�9܀��u̶�	�~�@�:�8&�şcf�l�d�HFQd�-@��M7��!�p����ye��%ّ́qA��u���1�	R�^	X�(�'�\���1��ԡ8�y��Xt�Թ�S`�][���-yq�)�q�g%�-����_Q���Hk]^�<P�2���;��<:�v4_��wLу�ν��SY_ߖk�W�.�wu3�Nu.t\�+\3��A�Bl#A��4!h�2�.�TE.�,վQ�܇}-�#�hP�z$q\s�ڐ�oBv8Ɩ��5dg�(���:�I�ŕ��Kzz�bN3+��Y� !>���h^��uq��k<�B��d18x�4����M_�iKTy�B2�a˥��+z�,�\qT��')"�!�y��O8�%��*���{]�P]�9[~o�/�OE���>q�lep���)|���إ\#P�B
�5[�*�� Pܘ�E��g�"���I�!�ʙ�T�ѹ<��|�����O���O�������!W����:c6��N�Ե�d�F(�>ef%[X�S�~h	�����2w�>����A�H��1@�B9TD/<�X,�8�պ܇�
aqyX�vD֦�)|L�>R_��?oY�2[��Dn}��Ŕ�n�5/{� ����2ȃ����L��������O��~������?�?���q�.�0����)/d����xD�!+��G�&��ɔN"�t׍'�t,8��bb_eR���n�P4���ˍ����;w���鯴Մ�d�!T�����p��y+j���Ɏ�T���'�B�W�Wm2��?��C5���-�3+��|�O��X���y[�Za&�X�����rgp6X�&UԦ(/�Z�n���Ax��J(/�/��˅�H�-�Y-\:�5p<j�������ل�A�����-�6Hp����Y��Ù��K�}Z	Q�p��/�(�8K,�r��.{X��i=��NN��|_&���Թ�E�++�-|Q��k��.���j���W>��c���6d��r*L�����ۦ�AN	��Ϟ������� !"�/&�p�H�(krL-��bKA�Z����s���� �_p�����ݝ����m��7���-���*W �^u���<�A�<T'u��c���	�l*@ɋ�|<��ѩE:tl��6�[�������QH�����cC=�C���` <�ɧ�ul0��G_D�gӂN)�HH�Y��1�!�'��Y/��m)��R4/�X��9١��c�Y����'���I���24���&CZ֯�!�=��JX��2�EP��@�;6$v�G�BL�*O����x�!G�
`7�x.�
���f��R3���乕�+�h��u���P������'C�iTp�LT�j*�j�-�e}k�e�I{�Z�~t;ou!oX�uԔ��AR;m �L%���A�_4������:�=h�j���7+H	�-d������/���|���ؗ&�j`H7��@@��s��S��1�0A��D�� ���n_�:F���5.ĵ���ٖ�:m���N��dC������ =RpcR� �I�)��/�����֓wn���ro��P?R�QM����Df�H=,��pUPdy�� } %q'��Tdq(��Xwh0	�����&d��	=:��T�;�<*rBy��� \BUCT�W~�S$��������"�����"�l�� ��zeWw
����q�-��~��|�kdʀ&������ÞQ��'��+Uyu!
�/��(�S.ǻ�6����'w�
b��57��t�%��_�o������sE���I�f�X��Z�=&��z�E�	��7.)��y�ѽ��jt���g�b��@>�����L�����M���왵��b"2QDZ0|Ed5���όbr�t�F"�n�DTc�S �y^[3�+�[|�EQ	ڋ�\��pV��ζ����Ђ�G`��JIȦ�% I����"B1�*�Co��:T��B]��o�w����@U��ӧ�q\F�ň�~�M�i|�@Ǣ�5A�C+�\���l
����B�y|��d�߼�@f��s��M�#�#Ӑ�;k�Ν]yS��+-��X0�	�-����5�"�������u�^=d�$�=���'O?�7o���#���r��p͂S�������^�s��[+��|�mrynM\�v��u�}�u�c������Nt�C
������n�`��\^����LB�7Ҙ\��v���Im�CtE�����5E���Au!�jQ2��0���J�o'�J1�� &+�q����(*�?
��s�ƾ1Q`-��:��Q顐�'��Uy��U9�q<���dA�'
��yOzj��RJ��2_�nar�ƐVFϮ��Mx�������I1��P�e��Ω���9`�2Τ��\��6Q��Q��`�n0B>l!�R]N?G�X�/���6�͕����U���m�����ͻ�rugUV{괢/�٩�����Z��}���7ьI����?�������%��j��;��A��t�9kFz�\���P9g� � D��AJ��9� taC��eF�q�x&�(Q�4�`�:� �'s2�����o�&�Lf�'<�����`zeDK6��r]�	T#��bO�ǁ;֘�9dfͱ�[&7H�2��(��fxh��T���)��B9�l|���ԛp�(��[=�}Q�6��A.V�&�Y>e�"�/�3ө><zR�4�	���3���QO�����/5�7���|5Z�	��Ȩ�~�&��W�bMQ)'��wf�<��L���y��o���^o���d<g��&d&�(~?	j�@�C�41*�-X�M*-��F#�`MGǼ�脂;�:?�����C�����1:>�=_��D7���!�m��7<:fa:�O��[2A A�d��e]�~�I�tt*�қ
x沲�"k[k�ymG�<�@1�T�c<\xХ�榢�bo<��M�j��@U[h4���"� $d�cW�����d7�b�e$~�*�vN�+d
ߥ��[ ,Z!�ǈ܎��D���kX�8*�;�'Ib�U����u�X�żvX�8�����X�u��R�����eIʠT��VU�e�(?�.�FE��(#�g�*�`O����ǟ`�Z�3�{�]��0����x[m�����^�x��	/?H��
6u�"�=譃�G�%S��D�mƺ�vī������N�i��O)b�W�'�?|&���s����g�^�!���Qߴ�VȒ����zp�� 4Z�7+0GQ��fC�t��Fo��^>�:�Dʹ^fkR�E^ـ:����}Q�{(b�\�ŅgA*��Ua��
�s	`��g�'���EA�V�P}j���T���6\�O���T�A7E������'5)E3I��Ɋ��_C*Ya���w�#���`3��Z/Ŋ�(j<��#׷��ݷn�O޺�q����I�&/��Ev����$
?�`�D��g�b��|��W:�� ���,�ٽv����`�X߰��	�Θ_|����ߗ��3O5����Ȧ�A��A/�!o߹-����I�n�*@xtT��	���3�R���/�Tp�)w�ܑ;�o�͛7ټ0qER��0�<��i6���#�ŋ��`| |��q-��&���<z����}�a̕�;<jp�2U*-�P��H�h.�9~�z��w��*��!ZK����W,��^�מ����N�����ա�\�ɭ�TR8<:���c�C4^0�K�871��,;f��|��l���bQ�$��q}Y���y�h~_�@U��T��ƀ�#���0����q� ��U5� YA�����l1��ժ�ݭuy��y�ݻ��O��իkl���똞ˡ����I&���1[�g�Sg���Svxv$����K���(���hBVu�h�NhIt0]�߯6cY��i����H {�ϧ�#DI�zdrun#�����E>�t��__�R����!eP�z�v3�S��Iv�ꆃ�����*�������ݩ�JG.��,J��i�P��q)�;�]?w><����S�����'���=����С�(�8d"3�_�
K-z�N@�S���bJ���t~�/Pl�(6$w!�ՖFX�(X;��4/��躜еt��y�с�c��_�cD�z�]��n�B{
N(��G����&�gG-˛"����,&�C8�C}�M�98�Rw��� 4��I��=} �,�B�z�@�l<���/����\�	���&A�<�@ZS�An�0Sp5G��~D�F:�g#��L&�V;Hs"�����Ȃ�7�2Q0y69W�ߒ��+�s�l��rx�s�N Q<���M���[���j-�cZ�����}��0�ˑ���y?V�����T��#�KԦ��KN�Ӳ��`-�Ѱ[�\�����߫�u�:���ˌ~,�/���*������Z}�e����R��k_�~kW����1��ܖ��l�c\�}���|	�&��-�D*U� +��I@,�ZB�mK�����? R�_��W���η���X-̕�	��Ü]D�S�$cm�/����щ��fe��6m�d�9��v�+��Q$���8�)�8���:��L���;=nK}�-�s}�����6|��7���a���%���C@7�e�����8ogYE�FJ8d�L�;!l����q�@9�ϵ�%d�6͞P`���(� A�`>4���X,	����:}��fd�`qL�M�_��}�KSlz�$~�����B�Q�NK�{/�M0���35�G�f���֏@��\X78���؊�so%���+�ru{]��l�Q5��	�yО� �7�*�Z��aT���{||̯���7zzzʁ����*ŭЦ�""���L����o�;:�(�h��� w�Y�/0��&(@���D�Dnݺ#[���p&TN��^�̿��W�h���[�ч����@&�������^�:�x�Ϟ>������$��� �w�Q��S���KJX�]�c��<6j���o����5 ��ƛo���/~��\۽J�jqA�U)ܠ����^S�z�� �/�&�yp�x��J��J-JI�5�hr��VBJiy��[���W��-�o]�
��tO�Ɂ�Q�7p��٨��R�ya���Ux}G�n�Y����HHʨ����׍� ϝuBq�ØQ�(D��J�]� �R�A�#g���|�����@���P�X��I�˝�M�ɭmy���dCN��� -sq��<��yr�Y�6ek�+뺦;
>8��0����}�28<��MS�Am�b���ӑ9!���I��fm�ZE���TBa�ΫVa�38��Et3&�\7�H'k�����Ôφ
DչE$K�5��^j���y��	v+�	G1[�Y,X,�:i�sm�.���Xq���l�ڠM�PC�L)��A�u_?S`y|~���vv�q�2 �?�����[�n`��n!
ϕ���eS��(2j�IR��z9�9��jR��)Ș[�����:*��|c=��@���s�Nϙm�Xbb&9D�y�隣bb�V���YdQ1r�a��:SP~*��ጊ��&�e"��R��l82]�|�G�|��=k�f��5S�se����A�kbt>`��|8�����&d�������zџ���
A��A�U�Ր�ʪT]���s=�B���l^ےg��@�i7{�>��l�x4%�����7�ڣg��w(��'�1�� s36o,̎�!VGq��/U�3��*�\e���Z9t!Rnv�x��	��݌*>w�T�+j�����?�LHlA��~��]��bAA�n�+�R~/IM,���^��)�kR������W�^^"Qu�9F�5�dm��,���12��?N{n�a�*f!��+? ��t�@D8H��G��|%�#E�}R�LyA快�V�w������U��ǫ������,߇ݾCMMT!��x��`p*G2��.]ӱ�$�K�7Ϭ�2l.��5��g{�{,*�ӟ��O?�L�>�й�`zuu]����VI�BM��/&&���u*�������Y5_�l��n��䫣�_
���:��>��! 9���g�,e��@d	���;L�ʆu;�v�R+�D�9��,�*�h�79D P�ㄟ15I4�>V�8�)������n�n@ɊRf-�zu[��� G����>�C��2�8l���y���+�R.-���?�����dG���5�X[a$N �P�w�aR�,�!�g<���80�s�� ��H��K��kkk�(���?�$���V��z$z��"��n `��9���; )H!���:�#s>3끁T�s���I�������?��<�T�ՁFf�o��o�^�$���#3��2~.��Ѱ���edR���A~����G|H=�O>�D���#�a��a�sA"����Ϟ˿��ȗ�<�Q'�����ם;w�y��6�+ie��lT��("��#����cv�|��	���wߕ��{O�z�)9�f\D.�g�~u��}S��Fq�F���lo�ʛoܖ㓡�y�\�hA�"eVC�_�(��ܺ����2�㖯���	UT��U� X;�ia[����b�,/�A�H��,Ṷ�O�VeB�~���+sͥ���2J�I�[mB��H[�C��w�o�;7����U��?Δ;��>{*���B��su��hoH�Ѣ��"��S�:��
<����*ߴ\}��@� 2�S�9�
�=j��@�Ɏb&��槣��w��Zg��6���nRP�,m��ʔ�(9����ņ�������%6& >��7�sZԌ�.�>M��c��%wA�,�4�^c+�材ML��U�>���ʒ��x�}u^�x$5<�Bm 0Q0�Z�4���b�lټDFf���v[���'���ܲgStS��,#�ss��'B��g���`�g�3��8fo
�q�/3��n�@v	=��� |����z�P�Pь(.�t��P5kZO�bQ~^L�h�3pĚ��kI� ��j��3ңX�1N��� @7]��u^ӹ�:� �{�k�\w��4�H�ºbA�tf��x$8d�u^G���b��t|��x��z
�|��''�
<v${�:�����]��+k�>�~�@�)�
���k��7q&�ۂ<�$Uk���R�~��df����PP��J��JVU�[�l(��=�Y������s�-s�T)�d���+.B����W"�ŲM�.F]+�6*�V���[��C!}8�A�R8��9��[ȫ�����T����{t���1 "��$�'F����c�I/<;�����njs�u�r����v��ku����nT*�z�u,��+=��:!���_�;�@ ���<�/�ޒ9���O��\����\v��ۤ���ل��G�|�����g`�ܓ�O��x4W����t�+|����� ��b/��Ͻ�ty_Q�R���*\�-4�+�{Q	,�+��!XՀ�9�-�]x6!s%��^"��&���� ٵ_|�5 ¹\X��5�`dA�:�2�~`7�~�`��lou�����ɱ�qG�ͽ�DR����FT1ئ�2�n�my��7壏ߓ�w��������?}`\�6����Τцl�,��g�!�n����ٽz���[ԃ/�Q7��^%�J�3ײ�L�j�O��/_P�y_�~�m��{]���7�(ņ��8��Ε+W�����O~"?�����?a�8>�/��/����ܻw�@Nx�8�� H�3�1�����3���d�'a 7(浞)X���|@�B��(�~ds��± D��(؂���
BV����i���έ�����> x��o~#�?�/���?��w�23�V�&��`L�(�<}"ϟ?��?�\��kf�Pp�c�|��JZ�4���Vi���r�)y�����ru{S�妼Tge�ő:"c�@
^����(�"��S�s*_@��/5�ir��Zs1 W8�I�M�7n,LP T4�꛸!)�D�ȿŅɫDq/'#���t���1
�9F�bfu��r}�'o\��{���ͭ��*�4Ps0�A����������|'�(�f�{�� c�A^{x~&gj�i�aD�M� <��Άz�����<��_�B���qQ �#p�>@P2�n�漲 <e�[3�M� ��%�Mx�86P���0�b	� h��+�N����n�F��"����Og��u���k>��0�4�欳@C̎�]��Z"6ʜ���))=a���xk�����e���qЀv�<�$8Y�n�̊��9�\l���7P�
�3	ծ\�{"�M�䨅�H-�_d�&��&%���St �&�rYF�Y�C�~���J{y]"�5`��C��!�Y�Jc��ٝ�2&�&̙�dZ0��}���c-����N�̡�WC�4�qޔ>],ct'���_��T
�J�ѳ:72j�w��+��Ku��f�A�m%�����y�w����!�gC:��Z���Ȇ�o���Z_A݂`y�NL6�[ݚXtI��8�
�5��PA�����ECs�!��K�Βɨ�MPש��R��#�C��i�<��ت��η|����U�T�{���C<(���g�r`^!��~��U!��^G���а�^!;���j���g.�^9�f�"��i�*���`	"���>�%�X��]��`���/H��K��PV��b������Vz�|��|)�8r���A�5�bP{$��QR�7V_r�g
BF��P=����bֱ��������_}uO>��K��?d0yU����i�o�	Mf��i�ЂX��ZJի��VД(˻��i�ђ����U�Yĩp'N͏�x�@ ��b�=��f��^��XB�(ENĲ�AY3�'1f��p�X���?f.*$�K{}
�Ȩr9���l���?ݠ#s��q8T̑y�
T��.#Ot�7߼+�(��������A����7RQ�`ҡG�-�9�xQ���ƭ;r��-������n|�nE�q�Ի�۫�;��d0(p�A�B��LCF��ԏ�9���J�D����ŀÏ.��k�v�uЯ_��>�w��?zL���)at��XO��W���k�k�c!s�`�ǶwH�6��'םOr���qn\�/��/Y@ �����	F <��oܸ���I��Q�me��՝���_���{���?��`  Y"�dL�ԅ������䉂�Ͽ�\<x@�ޱ�^kz]��&��(<�%J�� ŲNK֊*;l���6���t���ع��P����<V�Ǟ9=%>̅Id����܉�K��ՖU� /�S��%����ɺ-��E?�ynAq#�u�6�E��=`Li�2�&n��3.������Hf�Wn��4��^K~r犼{C޹�&�-�T����f�x|z,{���3�#�rs��#�?�:���i��ь��
@�GNl�4ٜџ�;�@�;'����7�M�	�I�D��=�o��A	+�	,H���lx�Pd�(B� �f~����@��b2�9��Q6�F�m8��t/�~��Pn�����e�u�PD5,����]��9�̓�_1;���]��e�
?�ʟ��j�R(xnS��`��̡��lB�>�N�4Գ`z��e|ʉ�D���xl�E�W)̙o�c��7
X��%l��x��z�:�: jh�^!k�mu�YČʳ&7��	�{K�AiI�ۖI<!�ͷ@�#���)] ��V/���>�6��FǶ�tc쮯��@�mCC�����0�#� ��|4��4�ט��ۭ�DP=�$}a5���4"P���(J@ �$%���|�]O<� �D��B��뒺�������}�����9��^�Omțo|"��})�i�NȝNL��5D[!1ق4����{l�Q��#�}�2%�'� �_�W���t���n��cR���������~W�G����5�ޤH���Ut7\�E)�2��$��YծԷ��J��WEE[$��ե4���k)h��o��Ep�]1����Ȭ���<X�R~?KW������m��3
;��@�l��\r'K���������Wλ��@�[�������8	N���a��@�Z��%��)�;���&�f2�[�"q��`s�9��=|�@}�o��|��}ʿ��՞v����ڜ�Y� |���c�����qkېUʠ%а bTwN��w���0A��,3�~h�֣�(lɼ�1���Y�Ga*w�U��E^��Z������mޣx\�,\82?���E�eu��,H�� 0mV0@TM��m�j�=~t
~�5��رV<b�����$�5�38&c� ��M_B�n�������&P,^H�o��ڒ�
<�}�]��u��1&"y��d��OVKE��&yq�B�UpC�� 5p��H�N)���!3�LY�rV���\���Ո��q�3 ��Н�w�^�ʌ�E 3f;X$�w�h��P6Bd^��`MW~����m������q`u�V+�0�Gz�О�
`�����"��o~mҿ �������gR���ܸ~C�}�'��G������O������S�.*Ԕ���j_����]���y�@��,�Kx�;?y���:�.�ʫ
�Q�����c(�bWm��h�c��
:�OD�(�<����2=9��Sօ�-�� "� z��E��25�`��ԭs1"�h�/��BE�#b��BVxïآ��2�I;�,�A������4���SW�=g4\,���1��\6�y�Ʀ�?�-�7R�h.����<oS�'�Z�0�d���T��@�c�a�+%� ��-��HՃ�n�ȁ]lXA\X�>tG�kl�(N�@����@�E��9c�l:f��l1F�Ō��%H�;.�+�w��X�X�����M��5���@�V
:��W�x����%��R֒`�H��	u�A��tXЎ�Ɔ%���6�97w�ԡ`��	��,'���M�Z 1���Tؘ=N��>0���d`3�smw�F~��NxH�(�	��*8�� ���2��@odҰA%-f�����ұ�d�^��J[��?��}0�P�"�+j���S{?�y���.Л��@�8g-�X�ጛ#���$S��؝��,F���G�<Iۍm.���7܂�6p��4ٍ�5�E��8�m@k:���; Eig�^ �;ѹ��9VV�x�-Rp<�����ae��x�ߣ�.hZ�؎�!�.��� (�=ޖ��B����d]���L�����P{��am�ǚH�H˔s��p��� �l^x �AF�� ��"#�G) �Y�-�gA�=zlG^گ*�#���S~�cG��<�(�ryE�^��de��4��>E�j��[��q1���~����
�E^$�3���@��p���e���J{^3~,D��wA���Ɯ�%��g�^|.�B����*e����˽��+��c�*�A�0L6�-A_��?W,￬{����|�vR8��{���tM�h�NG��<��P���ږ�0����1)�/����⋯��o�Wg�Z�mWVVu-�JGH#m���M�H�0	h0d����]-
r�p�w���ol�ZQ��_X2�����?��,�����Oa�� ^_4[X�<��'�(OX�hD��*�z���K�֘x��(L�X���� �&�gI?�3�&<��C/���نTߋLL�!χ{�b(|����is26���_d:�QE��L��&���Sy��Ċ�XY8�2w�>23��	=�����[7o�Vˢ���,������ �ԯҵ�eS�������馈MvU�Y�B-㠿9��W�τ��j��Ѭ�*�h��b�4�0�=�hl5��'��Q��"m��V������`N��
>PbM�E�r��}�֬��0��cBkH��N������Y�������p������A�8A�ʍ��孷���IO{�B~��߱8��*�T�P�zǰ� �@�;�`w�x�4*p��g\�$Qh�s�Q�sO�=*�E�Bⴑ��؊>�ݝ�
�N��|2!g�E���~"�v��B����%`��/��:H=�6ɸ6H
�M��#MJ��T��n�	"�E���yQ0�y��F/��+�(uhW(\��ʇ�ܒwo��Fr.��@�ơӞ]ÃC��������S���H'N}\SIt�G-u��iB3Q4omN"ƈR#��L�u�j�.[��x�Y����"5MJԜ����LS�tG�<S�8cT�j �LS�0*$�J!����h��g6��t0��X����X�7fۢ�<)���LًN]�����C�r�kP�XO�E�RG�3��\�ߴ���k�wڒOP��@�,(-�Ԛ���p1c�>{$V��H87YTuN�)L��f2��J-fP��~��Td�74��T�Ā ���3BM��A�����&������A�v���L�a�P'��v���գ��yhx%o#�05
�l4$��di�o�1�����c���������A��U�7L�76A���#���h�2�(����S�� ԛ\A`���JO��ybs)�[S,�!$qS}^z��Nq��2$��A{F�����Ln^OY�s}�>��I���XG3�5����Q:|�F�U�\6�;yx)C�������E��֝�P�a�ۂiu�ֳ!(��Z��4�1�ɮ�A���&�@Ы�}���˜*��x�BU}O�;���P���L�%����W=pE� ��DJ�V�x����nfH����rE�qi�� w���M�^�����W�:��E.!�y���� ���(8y5����*��A!ˁA|žw�ڲ<�?��������|,gl�ߊ �eo_����Ǐ���G���#��{�����;��V�K��f���(8P�c��
DE�e�2�NC�{��?��Eb��R�f�6nY^H�B�q�(КeFN�20��<��<��^b6%l=�r�f^�}>r�w�p�rUuV��.kN�oaQ�����ތ�hj����i>�D����^D�#g<X/"��ǘvZ=P��P��
�x�������^�{���DN�^�`xfQ\���4�7{ѹ�P^�^�uz�^ݑ+W�0#� ¡E/yk���f��E�`��0;��4'P�Pk'��ݻ
&rs���k��&O�o  #(��$e��:�6A���
���k
*���"�,�=���� [M�+꬯����ӧ�������ק�.h0x�L�ozV�pPf�pB@����>"0�u�6�{{{��wr�殢�&�ϡH���֭�r��my�7���駟ʯ����:� ��z�>y�: '�;	4����x��Y�~��f=0h��ξ�tg�R��^�\��y^�
)��ҕk;W�7�rt<��ӱ:�/-�F�j���w��#���EK���F�!`��J����1#�Q�x���)T��p��g�{ࠫ{�j��(f.��\��:g�"�VX�ęl��r]��On_��^$��P������}��Gr���OO%;W���j�N���\M�m5�3���^��ʔ�xhN֣�h�����/{v��`�Q�
�!��:�jWf�9�lb7�'�I+̙�;��t�&��:W��I��)L�A��١�� 8'��;�x_���{�4ÜQ��b%P�C����l����x{����-����-t��f����!�����=*��s#2�@���5�N!m�S'�nGQ��EeS*g������1��4#�1��	@eoAU*3��2t� ��F��|2��!�EYSՒ̞#�}��=��Ϯ��0�<�	$��67 ���߂?��gf
�&
^G��kY3D��ĝ�C���������D�����O��׋-�,��&��ڭ�J)�y�o���b�Ϙ�V�:������:Wөem@�Bma��U7���L�c��c��i$�:j똭�����>�� 5?�lWV������5*�)�3�x�;sȣx����!�Hv9��������V�����9S��V�Y+B�?�=.�=��p@n+c��.�
f�k9�S�����E���f��,ϲ�Tl� M��e��.9  �eϤ��g#��]���K�;��%�/�\鳇`U^�)��R�Ko��ͣ���r����e��>�p���� Z}�e	�R)����"��i��\����^����������nW��fm��Ad�?y��'g����������>�h��n��(h�ZH�:���=�=�4G:g�>I*
�sϛ�Li���X� ��g������yEQ�0J�nch��.X�1'��� �8�����k�j�g*@j�bbAB���� *�#���M3��jd���//�Ph0p7����Z�a J�����G1��Q�ІoI�D��F�-c�!F��Ԁ�,�����P>�#�N�D�cC�C�l��y����&�.��\�do�aH  G�g���TnM�zi�VN����0�����At�(ЕP� ����ufX�7jiBD'��0�B���S�{����@ FN{�F��M�)A=2@�S�|a�C��E���7�Я;��{��>�_~���xȸ|��bo��4��2Hg���F��΍�Q�QYk�ms*�����"�yГ��ƻ��b�o��F���|�<��a$������;fUvwwI�` z���czXME0Z��F�nY��\d4�B���hdj02f��VR���&7w����rx|.gC&��r�+<P;qQ�Sy�`$C�Ĝè\p��"Y��@��H~��5��I���L<"�ERX�92�[v���:��wK�M{M�坫=�{�#�䥌O�ex�\�T���q0�c}�GϟJA@mǠ��Ƴ�,����*�	v�6�c1_�� ���B��;h�*3u��)����:�5_בկ$n�).)۹;���-�ٍ;&���l�Y��|n�wB�o��*\Ԡ,����� [��(x�E��ዙ���Xuz-i��P���
#C Yj[�Ȭ�c�F�#�H�i����q��_Ѭ��O��td����K������g̠�F�<�BWM� t��8R�~��c�;:��/󎴲6�����ЁB6b:T����t��d�e�#��������v���g�6C7�E�p80�]��5�p�Ng
Z�%�E4���l�!%�G@*1�M'4+e��h�y�r���m��a �IH4��"iG-��S�Nt��
���\og�Rp�I�����*�W[  ��	��e�sdݚ�P��u����~���ζ<���L�Nes���|��y�G����v���*��kw�߭9�!�!�͏<�]���2�g���|���q]x��z�GgV�2�n�<�K��w�}����gu�֨^��Zr�G`!��2%u�0�k6ޜ&{_�j�)�U�l��;�*��g޿f~�jN��$<��ː�H(46(
]��@�5f�����}o��;J�u
_��.�� jJ�q	�ԃ����}]<���>DV��\ �(�[��#�����e��c9�,��������G��K�;ԧe̾�::�=A���#Ď���������t ���/�_�_74�o�sGFS�|P@�z<�� ����[Go���|FP��{���F��79\�0�f��H�B��Vs[����B�Hn�,�%)A�V��e�ʫ,�H�ν�������(�3�0��a����u� ��(�uX8�#�;|G�!� *����v,��7���'"cT�#���]�����E��v�m��I�x��1u�wl�I%�'�"sy��@��X���>`Bd��OK���b3U"�ׯɭ�7,"O'Zx�p^х_pn�T0,�����K]��>;���ݺu�_7oޒG:�}�5�^P�ڹ��z��-j�@����S��{��D��4,$d!�U�F{x<@Ь��|e��A#�3T%#��Bm�����n�$�BZ�=ԃ<z�P~��_�g�y��]˶�������g��� w�kF Dn1ϫ�Cn��Xp�@CB4bD�ׂ���zh0��80����x4���
��]�y��=e�z����i�[ۘ�2pb��5f��@��|[�߉dC���[�rs{]����N�`G⍜j�W�dg͐�J���|Pnϵ�z���pA9 O�h0w��ʙ���z�8'��	ߣ�]�������v
u
�B6W"����bq$��X��Cu|����r!��1Q���-C�[��)
�P&����T�Rk�7UGJA,�S���տ+ i� ��0�M��+
t�0�l[����}�SS��Mf�[s�)s�n��MA����/Л��� W��c�;pL�8���}֞�vxhB����##7_ ��CKYƬ'j$���4L����`mH�d|_�[5�@O5܈���m�wԀQ���dB@4NYD�����S��6
 D��DJ���yn�l�h�QPv ��~> ��&��y�^Då�'j��!���n�s�c�1�O�.�D�c�L���]�q��d�_�K{���'= ���Y��(�̐�P V82[pt�V��06�u6���l$+;��@�,w� ���<�u-�z�4P�N=���ӑ4z+_��1	�s��\Q uΎ���1���|��Jog
g`�#3X+
���̦x�=_A�d6��������HLm���i.׶�d�7`�{3)X��$�����: �v�:B��'
>��3+�ປ[��6"d�C���(iPх�٬�ȴ XY=?��u�^�b�]�}:.)yT�@�(�s!Cc�Ge��t�<�21��˽��xyxMvc9K]{E�Y�p�����eD.&����ߖ.���" ��&baoM��X��σ���x^��! ó�����x*�4a�AQ��RՋDׂm�"�W�X&~B �^�\ؤ� ���x �r�^�@_� 4qV�jVj��a(܎�ȧl\��J��eL�d����K��O�����i�I�:xy@
���p�t ��L�9�+P�Q�qv~�{j40��T�L*�{�M��*2�g��M�m�2�'X0+ 45<�}mem�}�0�Ơu��>��h<����0��p��Ō�o��SI��[��<0l��-��L�-@�����l�S��Ҍ�?X5Y+�m�#�mB�K���k�Q��f�F�$�QOz��9P��^.X���\��rrj�ؤ3���ϭ��"�x�ߩS���NG~p:a��Vd��ڲ�-�-b����6�c4�3�e�  �
|��7$|�eԹ���y䏎���B��[�ـ�5P��F{p����!��M���� ���P�P�����w�a!���ke������&��$d^�"IM3���{�II�x8h�ܺ}K��o��
���(��κ�OWn߽-��9��#���!��s ��z���G��2�74�EUj0���P�ұ�r>�L>����@&��7���SH�˷���9��,��[7�> �|bδ��2��73�E�J8r	 	�~�R�!��� r�ݎ~m�[rK�Ǟ:K���B!(j.�V�U���2dH�@��H���y���o�b�'�h>Sx0�q�3��Ct�=�(!}��CΆ1���N��J*��ޢY�@&h4�ڤ�.&�g&�p��H��Oέ�?�ɉ:v0����&y��Wd���/�Ѽ��oH�۱E��9�s}_�|�͡a�Љ�-�5P���x@l���^x��	žqSj��3C����z~��� ��sJ�9�ql��:-������zi r�Z���gd2E��v�V�q��#�`ᨣ*����MF�7�mC�G��AGAx��vO���=z)��-����o���X�%U�&�rn��Z���ܔ���)�Ez�Fj�2�$Xf&BE����)�;t�I�S�i4�D�t`�B�Y�$��I�OzZ���bľp��T����z�$6�Q�� Mkha����v�}��ծ^2��<vf7��YVN�P
p%	��bO#:��#��n�(�c���iC�����x��/Sd�(b��d0d�jp�ءs�1�<�F�Sa�óB���G�G�ܼ�@�P�u$^��z��W���^��k�Cy���D�
F!錽�Ă�ھ��-{ ���%�v�j8��"/�O����G�vS�5�jWN�)��xY�o�9�˩Pv-![�fR�q/m�%�+�<�.-�����Y��Y�2K}�j�����G?���1M<�; ����:N);��n]e���V��+��"������;���<���7�k$�ӌ��s���{O�&Eq�-V�,+$�}p�%��|8 �����P�����=��/Av�0M b���پ��F�9�� ��@$�����+��/_ȟ�8����r��v��k����=��? �w�H,�*hWP��/׃߳�B��P}#�+�����]iR6[k�����m�Q�4�n0,�n��|�u�ֺ��À.�=�
[l���������r|r� o��mu�j�Po��"���zC8�x@�T�+�LLX�?>/����w�.ap������޾s����z�3v����g�����u=^��!V��lY86�,
z֡�p�M�wQ��iY�1���xL]�A:��F�`@���yvv.+�U9Pg&���'L���b�7��l��������$ �k��)6,�X8�ɑ~V�Bk�fS��~^(.����֛o���/Y<{���p��?ߣ�^�t�<�x��?�S�4@Ő���ƍ��~�h&ηXXq&�ݖ�2��	 ����d�I����∜���7^ǚn���O��������/:._Q��ɋ����?O4a�<W���@"q�;.��1&&б.��@�*Ь���
> XP�~��-��U ����(���?�����c��G�/�����},u�N�5�)�VY�:Yڑ�U�_��f��,�X�%�~td�۔u���{�ے�L+S_�W Hq���~]�}�Ǌ�_Q9�Q֬���aN�
s�[txZl�CUR2]���ήb�F���ͫ�b![�=����/8�C���Lǲ������m]�>��9?�t8�܄�m�!"� ՠ�_����y\Cp��iM:�4{��'(�E�PO�O���Yͯ'T�""K�N[��j�dV͂*Z�45��X�in��&��=�g���9{�.;����FěsB& 8$HI$%j�e�r��^��֪��^�Zn�*�\.˲$K�8�bL ��}~��/��zT*�o��g����x�3��Z��F�-xQ�*��T
�Џ�a��t�.U�\��Kb���\���(7C�m]�(c���DBT������GbN�c0��b���!Qp|��cH{����)n�1[�m��@�֎2ۘSH+6ӑK4�T���x�@���9��=�[��n��,e����hiv�����m������_"�;�k��-C�
2|7���N�*ݥ��)����O��}���ȍ+��*��z�*�+�e�ȳ�`o����$���+����Nc�*=;��+c�%f�}߭PC�j����ҍ����ѫ_�G%�ii,"I!�����0���`@�����,X)D��rs��Aؿ�m�ag�{�
V�X����X�,V=�E'�k�V��Y
��uK!_Yu~���{rZ���Q��TB��W��j�ۭ���PӸހ��;t�7˚�������;5�g���i�~�U�]�S�}�t7�����X��Vm�G=��>���h�	�׮�Sw_I� �@��k���:)��Xŏ�r�Z�ɤ��+�3~��.yC�
M�"o�ޝjCU��Ǒ�������8�=��c���U݂AU�d��'� G ��ip��B%�Y�u���7X\RO&ZQ��m�
kL�U��Zy����D�/��J�mN�=�5�������V�d'I�����fx��Ga &.�S]8��헛�� 81�`ޛ����y&����=�	��7�����)R�/&ybe3Q�H죪�uX.�7��\�R���$��J�l��>���������+�nbS�1��TV�
���'���Տ_z\�T��"����ש��j�����B��5�
9Ik�A���(e?���aΏ��̋�P�W��/5W��L��J�yS��Mn����j5J5���@|S�s��l���-�*MW�Oڇ��8���nH�DA��^TzZ��]_��2k;�I�<�ņg����.H����)�[�5�U�{��=�s:�q���k�y�;�	���J���~���|8��������l�p(M�b�N��-2N��g|�/�Me�S�mq���P��˟�\T�_��_�O(���ҟ��O�z�)�c�#�c�⏍}�͛��L�e00����u��?x��p��>��ǁ.*����������x���Ò� G��_��������E�������[o�w�}'���~^~�e{����I�m�o]���⣀G�[5�>.���(��6F����y88/\�p.l��\f؝�P��B�p��0x�f�٘�.P��]����.��SƸȼq<�xGRGi)uڭu ��t7s���\�7@pqۀ;�^qVO!�?ш����!ƞ6N�k
�e�	^���A�����h�R��7�C�**�íkz����2�}���-���r7x齝���>;�yT�ȴ�d��+!2_,D�!�Y �`<�Œ�����gKo��\�F��T�[@�Pw�zȖǕ7_##+
f�(�cb���m�ŧ�/VdcC<��·���b�N�T6���M�k3v��'v��[�Ϣ�A�9-�~�C���E?�9�`T� �������7&v?\�*��iي v�4q�9`k�&T�
l�#�L��W���ܫ.Cی3�v�}�rג/$�3܅��r*��I�k���*���̡2��W{��sz�[D�\-Ǫ�S��R��,]�!�̊����Ď�>��yG�^C�'�v��Ai]���ܽwO X�E����c5���#�*0>m�o�q��y���Ŏ������2�sۀ{�-5���@g�jͫT� �[�3�
@8��k%q�4���@�zV��=Z��c����uK]ʲ����k}�5g��$����h�_ٙ������|0bYL��K�C�lm�͚�y<��u���>ҩ0t.�ß�w��cJ{M��k�\=1Q�b b��~GU\�n��X�N���s܃��V�����Ʒ~O�z�� `N �{G�ZOZ�W�T����>  ��IDATt�g���ϡz�F���l��!k���Y�Y�;I�Q{����AA�RU�j�KJ�u�(�T�HX��i�-��LD_0��F��ĭ��N1�?ݫK�LUKO�<dQ��$��C_O==Y���Sɋ#�(A���υ���Ν��.��  pq�R������U�/�r�w��ԯ*� �SK��V�r��
l��Ѳ�+���̽�S�½�}�s��&lV������Z�΁�=O~N��TE����a��t�\Fu�Z��$�����߰V��Cǽ��0�Sƨ+�'�w�%8#
Y�q��넀挧BA�7�����"`2��X3W�%�>�-�R����L��ԋ���Bx�
��.�wP�9W-�E�)}g��k��2jl�soX9��vm@����B���^{f��,.�Z��u������{����9����ax�����ｯ�Fi�c�PZä�e?��Z�]mnm7���#TQ�yO����k�e A���H�
@@�\�#�G	,�(L�����L������ux������B������E�����x����5>1@� �G�sp5�4�@���o�����7�r�>�H�� A.�*�^��K��2�&�R�^"@�2FQ����Ur�G�����u�����RS:�-�$��tU�x���۔O]��uh��h����f�`�c��a���0�@���=g�8>.nZL�R��c,e�-����G۠���|����yõ2�1Z��Em�U���M?_�����r|*g����ͩ��N(�;�������oX�\��^�*n�T�
뛥��@��b���Q����B���l4��x-ċ����4o��U@�_�a3w�@�O�~�=�Xy��U��[�{�B��Z��UG�l�$�1"���l��-�9u�f�J�ĸ,�̯gP��0 ������V�
kU�Ԗ�@Uޯ�<W�o��,���҃¾���y��0<�g���fX���};]�O,W3�D�p�ܦ�@����3)1���Zt����Ǜ-;�A�Kɋ~�դ�Q�����!�o�/4W�ր��>�Dio� L���zU�f[�������Ra�2�f9�c;V�PD��k7��&B�����r�6>h��}<�=�������=��E@�c6�%ƕ�Ԯ��]�ͨ��)8��nP҇7�&j�mv4;+W��2�����;w��g��� ��B3�e�5�F�b�sڜm�_-��"l�I��ds�n�~�m�ln�7`}.<��a�>���4O/So����d��"����Z5�����N3�Ǥ��T1���#ob��L�2�i�묢��iωK^V�b�.��x����$(�E�ӂ�T�aa�(I�d�-�v�����������M�u�X�]'��e�� Sj���h� ֪�E���q�l �,���)H�b-A�����K�8��5��8�j��o��	U\�`bX�[��>VV^�ș�sWʴ&��J��I����:
b�q�y�*�o�t:��:
�����B���DbV����QOr���B�s:�G#2�cK�s��S(�ǊH��(�f�jg��[|���~�6?�����{2���=/�Q���l����?ɓS�e8��FS��������ė�#�3��~�4�T $ߦ��@�i0ҵ�̋Bޓ	74~��	Q�fS�@�ޮω�c넸���#VD{Q-�=X���IJ@�����<��]�7'��՞�`��9�.L��O\j��IV�u1ag�U���U�PW�j�5��^^yT�*g*dq=*Ct/Tg��%ĨlL6��]nXZy�5��4"���fy~O�9�0-�RR�U@�Y9�?U�{�o.EؾIhG�_����/���K/�û��_A��*�{8�x��g�_��/��@���4eH��lD9����:���gy��U������{-㵤������LM�����x劔b=x����������g�~�c$��"����A�ʆ�	ܧ�|R�b/A	�,�q$�q�6e�@�q+�/?'Pù�|��c�Xh�{D�Y�� �^���!���樓����;�9����{�}k����u����7�)�md8��;����3������P��%(�`{c5Q��xmX=r����D���7��Xr��� �1�y�Iٕ�=��-���W�$g`���k*i�٣��j���j"e����Ȁ��V�NF�ͪ�	dP�d��x�*���P�X�U%��\d��THPWR�L��1|���.W6�7�,��S��b3�dm���r1�'ŀ�V���N4���v�����A����y���'}���� �af!�vnb�=�$~ �:q#�E��"�H�"CL:m�wsC�C��6��J�ۦX�7t�*�h�\v�@{Mo>�9�L��T���͈
��A��+��2��PC��9U 7c�Tw�jVvT��+�y+�у���x�c_y ]�����о�N�Z@Ibsf��zV%e��<B�!��,��-qk�ڲ�pϮ�@��<��d�4�Lk���Ta�8�i�4����Q�
�6BC��<��W���Z9U�Do��9��<����(��6_ֽc|�6}��s^���x�?���^������q���_zN�_@� !s�u��ƝP,�\N�a����<�"p1����duw{J6%��yl����tq?<q�B�y���@��@���yLOg����L�AJAx�W�+"'?VE�Y���]�PW��ԭ@�܆!P���}�Ҫ 2)��N'^g��DL֬�ݪF$C�Pv���<�uS�H`K{BU7�#1��L\�]�#k�Uw�m:�?�Ru��"��1Q�B��tn�פ���Z�S�0� ���%c3͟�y��|�Y���eHR���/��8)���*Lh��>"0��3tp�pB��k������b���d˒�]m��BUB߻�b��{M\�.�U����H!�p�]�s��'�2&UH0 Z����e���4��������.���\}X"}�7-t0L��1y?�h��0���ww�þŞ�/*��]��.��$^E��l  Q�s%S��S>�ۂT���ƺ��5��k�� Z��}�oUb؎\�� ��pPE��>�e>w)]�(B�B�:��b����s6��'#�� ��^�����p��ǹ�ݞ� ��V�|��OI��l�>�X�f�)y����E�
q�y϶bMUu�9��l�Wb�$ap��^T�e9`���xS5�prP��R�ly$d�;=#;3.#�\f�mHkn%�$�(�TQ��F�+�&:��D��:��_����@��P�ȱ}���ɹ�~Gi��o|<v��(��R3�Bk�WǍ��qsc"�'*�l�z@U�O�+G�T7�9w�s ����X��RVȵ�����SmP�����<8�1�AO��&���s�s m�r�����jr��*Y#����`���'?���,&*�[RA�c��e�(��ÂA$J�9_އ����A�q`'YŴ�5n)��l�m�a�?$�ٔ�s�V�Vb:ʐ4�>7�ۃ0��aT��j��$���l�9�zm�u�F��V��ѵ�p,'�Х �h%4t�G�w��4\�O%�)~���g˩�
�`��G!-z70�#s;��ll `kP�1%?t���p6�dG��M�I���@**J �A�3c�������* �d��M� \}���3��ਞ��dtj��XH � @m��;�ŉ�҉>�V�$W��/R�L��%!��0@@��S8/XH+�T�$��$TQ�[�=��"5�#��M�Ϲ�C��� �Z-E�A6Q!e�ۀ�`107(ɾ#�{j�aj���`Ms����)��d����B�Ů＜�9Z-��譭[��"�>	�7�-[z��k'��^V���֎<�A �y6�	P*�A�c$�Uh|��T�=T�C�u��[N���C\�륍���#���}�]�p��NVSn�jX��{�Ɠc�6'�S\>p?%e]Up`�2y?ivѧ'�x2����'nz�C5c��;�ap���V�,�e(h�ÚF ���fG'��H�W�~���I�S� �j�Ai�$?6�t:�]�A�ZG�����o��3���ll�ݝ�����ʚ�p��lq]�FR4�HHիX��dެ����z��K{�;Tc���9<�|=�j����щ�禵�Ceҿs��g5�� ���ݽ���)hl�y��!CWhd]��i<)���~����|3c����X���b(��:�f�<"�K�M!x����An��y�$ӣj��/B4���L4����q=kc��S�h�u4��b�1A�r���ǻ�ŗ^PO]���$O_�����'�]_~u#|m |nk=g�ޥc�H��$z+�'$��B�ϕ�K��S����NҶ�������a�Ț�%ʜ���W2s�2��2��n|n;�lo�s[U��VJN�2�w�4d,=J �x
�P�%�_��]��Ò)�N|Zd��jA���֡�e^qnTU+U�ɆRks�x�В(iiN������� %�3��jf+hQ�G"��
c���R�C��
�ܬ�ج񢑧H�	��Φv���!��J}wZ;2���H�N����׺\V�?���Y���t�=Gӣ��`���
�	��D'���m��{���і��V���0R�6N���-�6՜�Z7�KW=��tׇ3?7�J�޴�Z�<�H��.r�9���,2/�A}ʯb4ry���uy��H�)��8(偲���W���r�Ep�$�}t��<�lczڂ�����qPq�1�{J�$��� %�m�L�n�
������O>����h$�������?x-��ʫ2qT�TYGt>	���w�o��^�������q���q�'�����e/f��0����u���z��MU��&��^�=����2]�1����6�l���ꨕ])(�b�n��O]ذqz?�*��a���r�yX%Y�{f̥b{��=򑸮��hݷ�sc䔨�E�pI��.g
be(��o��� �b�}�nX�8�j��|�JO$ſX����楁��ᶤ?'����������y�e>�쾪*�(�j�#e����C�qo8�,�aFLI�xH�F-��^�M����C��
,�s9C��JOr����g��݈=����}%6V��J,� �`�.Z8�r�0�M�9�"�a�6�(��p����
�D�#��mF=��3(tA��bRy�
%d2:
���+�g��"�Pnʨ�wf�.��P�T��F%�Y�C3{4�AT+��H��c0�֧�}/ ��'e{��;�صY��6)u4����\��H������}.9&=�(�����`����{�+�����w��r�>k�66*6�*;����,��{-�3��c��U�@I
ժ*~������<��*�Z9�y�����smW��& �d~�*�*
3L�̙�̃���z��o�[ga�����]���6>7��%��P	6�ݓ��_;R�q����S%��k�F9?�s�-�̽�s1W�C����s7T}��yۀ�CX�uO&��K���'�wЍ�ڞ����6��NW�M�y���|l
|﬛�7;�]�fѐ78�=� �Y�^Pq��gz�#Cu�� _��M�&�n�Ҽ�{]���\��5X{����Ń�˃��*A�U�X�J�^S�p.4�Ž:J�ȒF_%0��,ى2�GZ���M�6�v�ҙt�U
��(�[��q?|��'����ó�\�]�Sr��g�����q�s0�ga�֋��w��ԗE�X��u�}$�ӄ��*4�<����.E�*�n�*����%���"g���TW���Z�zgM+���m؞���aq�f�i J���Ɩ&P�G��L�ܬ��I�I�@�d�<\�CV�����Vpf����c,6V,gY���)|*A&��\q�t�,���c��s UM#�2�}��� �����y�yԕ�I�)U�۹V�_�j��J~g��b@��ޥ��������<ʸF�G*�O���;o�(���Z��Ft��p�$2����*6 Z�Q�^u��J��ֹ�e(u���t+�i��]
N�Z+���_w��̢�г[��.�	��(%
%5�$�k���k�3e�����{�]60;ך�T��ؘ��L���{=��c���y��x��o��0e��.?&�㰷�+�j(bG�\��p��a�hд�k�O<.�_�*X�Ȥ~��]���ny��GM_OY����򡙀�{t��&�ͼ�Y�s�I1g��_}%@3���U]�	�f��W��|:3����	I%M���Egs�o o.��ύ��Q����ZƲ��M@��`�$�:�롭�y�Wcr�S�p_��O>q!�b��������`�JA�s$i�m|��Z@��`{���۹�������[a�����T@>>1���F%@�1h`���J���y�%�<�?��[Ɗ��H��aJ�;�2��z�cѣh�e���*"�f�B]>���֗%�3�<�o@c ��B���@��sa�*¢�*C��ӆؐɖ#_+m{j�D�x%�)�U�I�ֳ^e3FsyyP�x�[ �I��*��$��p��Y�q\��X��*:@�f.�����8?���y�F�h4B�?h�����y�5�t�]����|,��<�B��x_��gji�������e'��-=��X��a���ז����2�䫽�J�<�-D�C߱ �U���B�	�����*��Ն���3����i-z�Z�rG�������\[� qC]EC,2g��=��/e�+Q?r!�BUg�O�d����K�6(���-,����	��=r�]%a�B� ��q�Qx����}1K2��W��(S�i����
���C����|F��U\0/�1ܲ�1�����!J��R�ր�KV��V���������koH*8ET�JO��B��n���j��Ǡ���3��Yrf5K�#�͚�Y'�<(�3�c���l���� .�f�A�����[{4a@��z�-���?<���-���#emU�*S�n��>t�i�"� �
�Sko-ϣ��[����woEW�V����y�ܯy�a��MoH���15-V
�/�o���XLp~K��M�s���<�������;���_}��Q��;����8��]J�ԫ&i�*>�+�zS9�1����k��{V7̏'i�(W�z�!Q=%���Ƚ�H�mo�*<Y ���<�����S�'R[Rq�* �&�΃:R�2%�",l�*RE��Q���ZG�'� �/�� ��6p �N��D�^Fd����Oqk���x����d��,�x��V֙kU�.8�?�d�_$zcq݈9ƳbP>\%-�iu�z<h��p&k�����0K���G� ��/r-��H"��C��~�͉�V!49�,�O��Ȅomm�wȍ��9������ϐ%_��Er��o��+�^��̎'G�&�����S��Α6Z���	F�`�Fe�S�~hR�q\EC�,�=�FL��̣|f�_��<8ߗ/?'�Z ��ds�K�iO�B�v>�\蓙D���i]�x0-$�ap\�{SD�N�[�u%��\ ����K�1Թ��3�"r�ڠ���fӎ�^���c�*Φ@[NgS�ǋ/�`��q/��Lw��n�?��{�V�:7�Ay�_�>Ū(PJU� q8(@Ο��́-N}Q�<�#�:IE��8�G3�D�ㇿ�i�r��8/�p%|���a�����i�Z�*��X���[hR����Ь�n,�O�'���*H��l�=������}��1	���B�'GzO�>����LmLRqY�>�캟P��ʂ]u�����#G��Wt��L�
���Y�4K���0EO`g�,��(�C���~�x���̆�{���p�x:5����9~�@I�,�h��>�1 ���F| I�[�j�A��U'P]aⴐ9��'�e̋$P�+8�#��y�����7'��c{[��;�0��J��}^j���U,_k}�Y@��I�:�.V J�6�J���(\B!i���=w��Q�p�8���_I�:��6�\<`�^LI��>���˞'�5���MȢ�%�k]�Z����S_� �ٵ{r��F�T��s�o���崙g�{1)QИJ�O>����Q}��0A�w(������fn�J �$ǚNE�7
c�Ǐ�_�� ���a����!vJCcP!��ߒZ�ͷ�S��{����t/��͝K����~8�*����5���d�z�q���a2���ɉW~�n����d�D;LFd�5$�H� ����GQ�,5m%�G�K��:�FO�π����g/��`'pyD��f?���*"Q��W8w[Ͷ�99f���zM���T(��M�=��sk�����y~c�:�,�v��#�K<�^(�N" 2_��b�s��*�8���k��3���p?��A�9:���=��E���ǡ�YP<�Ϳ���{9XX*�S�������k����a�~�fx��w��o}>������w�K�z���D��wEu���Xe1���,6Gj�綎,���N�TyHl��ࠠm�1�U��;GR���#E�%kE�s�����M'xx��{�k& ����!R��Z�:��i�x��#[�hHg�oII4��x�z���č�03��ֱ��''�Ceq>�|�'��F@�s��2������d���V�,Oqqg���_vm���t|�TUb$�Mu/�H�9���/Ji��Ѝ����y��*n�)
d)
j�M�ķ7n�й�$O`kո��Gw���xX��DMI��q)͜I�Bupn�O �`���E�&�tҩy+ez�Ⱦ�hF�$�"ćJ9[4pJJ��r����3�8O���M��e(T�xghIB}�]�f�#�~��'A}�`)������9�D��V?G_}�(�"7������A��*J���-�b��|�:�RO���y����oZ�Я���;	��^7MD�#^߃��>�����e���E,��5��4���kCŇ���NC�Jz�����I9v-0��B�Ǭ&�썇� ����"@y�x��u7��%��������)����n<��s�G?x%|�ʳ�!ߓ37R����:\���xC�/��e�%Y0Cph������
W?x;|:�z�+D����|%&�0�'��>_���2�w��ٜ�87_+�U�;�Z�h$�r�J]���FZ��T*h�d���"	��#_�,�jܱiDf�`&�������N.j�b�
���r1J,��{<g\mQ��׹�_T:\ݪP���h�f�{xh���m���Y�~D�9�׌�bf�:l怞���Z����@��x��m��6���ZB oZ?��=�2^�693*8��uh7�-�W�ZE��ʯ;�>'�%-�j���RR�"g#�֗94���\Oj[;��@�z��W�"�V}�0��J<�g@�9	�j�
n�I��H�V:7e�K�=�q4�6|��2�ژ���P�(`�&�LBǾ�N%������ci�C�J���<}gk���1岱<bIG؛s�T=J)���R�.�m\Xn��9���):�� a+�F(�A���'�#�m����7^hT��yCf�$�L���g�K��Ζ�){Tk,����c�
Wx[F
�LŢL&�$����lI�r1b��W6�6 8�����6��1oʰ>�u�����Z���CB����\W�b�_{�+�UXzԱv����3��s:` ��giYy`��y��M�)"!9����JG�u�j�x�D�g�bhU�
�'(�����A��zY��ώ0m��M�6�]������5�(�T9�'�'qp� �2���g_��� �����_��7U�������*�=��L�<�ׄkU;��:]Ϭ�A�m�lNMTߺL5'!%�[�ʪ�*a�*�V�����(v�BT�����f�j*�Kxg��_f����+�n�d�_�v�=�b6��;�o�Ͽ�B<O��x�鰷��>E1b>߽{Ϯ���/�P��PR���H���\�-[;�X���:�ǚJ9��ׯ��>�$�/<vQ�A$|	�y�M�_Ĵ��"D��"s������K�JU�X����A���W�����O����.^�d�Y4b	)6o_�ί�]�/��\J�������=���<T�J6ET�U�n���ժ񉠩��wߓf0�ϑ{�T��U�و��ɽ�yN���T�)K7L�)[��1� x"�K��s�a�s��#e\2�GSnb�'h�q�F�z�+�1X��{�j� Be1���xn_d��q�khK������fs���j�M��޾�F��w��ޓ����Mv�(�+���RY;Ѡ梭xyR����p�UM�	P@�/�<Q�x��7�qr�����D��s��T�W������o~��!_6ιW>�uj���;�iy���W^y�Y�M��L��������6%������K~�Ѩo����ӆ|@�9YT��͙bG���/;?w�o<T�l/����Ӱ���Bx��sv]�|\�ى�~j�%*D,�{�]����9_�c乒�g?\�p1�ۛX�u�S/y.n����T6u��)�š��������P�������ݻ�U.��*R����j��w�����!��P�W���\]��/ "5�q��j FT�։�S����n���Bzߵ|H.Bq*Q�"�욓�9A�{��!߰�HLD*衒'�J�&+^�M{��S��d:�E�C2��bJ$'vl+�D�Rz:2W��S�� F`MS1Y{�s�"�}qzr�M��^��;ѯ��𸖅�r�6o��� i�*�i��ܻ�ϕW;�����tb��V���BڟM�?)(@m0��Z4,�B}z˂a�8bt (A��^�l��{��z��noN¨�+�K�����y�d=���d�7PK&6&
��/8�z� ��
��D��"�����J3�zW��b��Ю��u�;U�@�}f<V`�U�JU�ʀn)��6�Ő��j�L�)����w��<����a㭜X�^i��O�T.5�t�@��^4��{�����5ܲ�4�u�ysn{b�
\o�C���
.~/&���%�[�n�Jɞ��JJ,u��,ʾ*X���y�2��>��*� bW��!���׶D%���K=Y�&��dW	����e���;��*�>ܧ�U�I�P��6��g~����񨿟}Tulx���8��M��Ji�K�돸G��DTK�8��#���c�Վ�$�J�_+VA��>�րQl�n�#�D�1S��M�dd���O?�������W�H���b�m��O�*V:�ǣ�ID�D?^������z=�ߥe�ǭH��*�WZ+����Z`�������s[6���:QH�����-�Qؚ�m�9�G�޼�|�ƕL���gGU����߻wOj����o��(I ��ݶ��'_Ď�L��~�U@z��䪄l��m�vCM�?��X?��?�u�d8��� ^���{￧���?�A�я���Y:Τ��.616�ʻ�k@�p��5���qTY;X"<�E��cW�m��R�=����}����=���K�Wo�s�zyӠ�X?�w�	��_�5��~%�$Đ�\bi� ��%ۋ�]y�L5�k`"e����EaQIϕ+y�/��p�K���&m��I�E�9
'i�U9��k��)+=$�6��������r���E�s�N��o�=�cA��vC0٣�A9k��6P�����g�E����_I�@h�_�WU(5�������N�r���_��ɜM�'Y�h��/kZ�@I� ����%m&S�� �W_]����������c��%5�U�Br��7n�7�|Kz�%p(qg?0TM@��.n��0�a����3O��������G��W�L^����B6a�&���y8:��y9�ҕLJ#�i��GwQ;�)��Gn�S���gd���}���=�����Q�q�V8鏶���5�l<��vO�! KnT��4nAk9��;၍���{���R�� -4�ݹ}7<v��RM��]�%�V���Ɔը��nL�>Cƺg㰚���/G����f++XU�G�=Qe�j&�M�MU�ۻH�@J*�T)$�m@e"�,����oXQ��j�}�ڇ��ʂ��,�jr�3���ɔg�F%�7���L��9��>c����,z%�F��䮹��E�\xO�j��5�ɦ*6�/��ƘKL';��p_!T�B4��`+�_T@BY� ��h0&��]2��.U=
R��b/	As�K��Ȯ�]����B��|���R�HE5�I�e�=?�!@J2�6<��8R�("g�|��C���*�fNUn+���℻���'��s.sw�q�q����F1��}�6�f���gҨ�`��i�ߛlH�
T��,ڃ���B>&vzQ��FȜJ�́�8W��<<�0�,�O�y��!���@-DCYI羴}�D4VhP�&�^89:��|���@�����<:��\!�3��Q���z=�U>=��x��1�L{�Q�j@E�ҧ�rZc0�k��U���������I��x�R�Fjuz�Nj��Z$���q_Ď"��}սVM߄���g*?����o=��o���Sٙ�In�)�DM��Mp���Y��@�5�M��ߺ�ގ��4e�ᾡ��,J7����ޜxub�{&@��GT�R�B_ܗ��,޹�y�}���\�<����z.%B��$Z�_���׏c� ��}J
V��DjS��0���JUe^�W�*�K�,m�®�[�'*i�;���k��c9s��_c�)E3��v��=�T�́���}�ć0F0Wv��0*�:շ�ER��Y�q9>:	_^�*9�˗/�瞻,
��{���܆��_~~����VY���g}y�+��X0OI�˾L܉�����'��=9~)|��uUc�~�-�$����WO(���LIth�?��/����ͷ�y$��-���/H�-v��=`[a��Dbœ����pt|(����2������ ��~X4I|��	š��Iʲs�e�Gm�u(I�r��={��H��N��6"[��d% D�ʃ�JՇA1�M�b���g��r�RG֔�����$x��d-h��AU���������xܸv�.�B�P�t�f���tGG�1KD��M���ҍE��g��/</ r� �v+.��pr��~�m�	�uM���|�o����s�P��_.�s��Gz�S�����)��9ج(9�2���F+��/�G>��9���y��� G9��m��&/�A�@> O=�t�W��wޛ����z�M�������F�|����DyH����>h"Pݜ�Xp�����k�&�v���B�hko&.1ƨ�m2�b2�;�â[���7��������
�}�%> �x�i���LA=jU�	�6tNn�bq&���ٱ�+Ib�5�g���?�g�.�cv��i��}�v���X�,&�
�0,@�rVJ������7�/����,�Y�9cW<)+�(�ױY�>��`�fRi���o톓�7D©NM ��N����k:�J�|\]i~��H.�{���X��N�"o殶�UU�8�@���k��]��B1��E?��e�����A��婠P�ڟ�R�BT0Ud��mǾ�^P�\�d)ޫ�5�]�)W��=���.I�+u$�Vj\�Ǥ}c��Za��I���#��I���+{Ρ�����xM��P����%��嫡�H�cգR���]ǌ,g���h/(mL��y�X�{N/��c2�lI?��d���E#���<&�@ZX =Jdӡ����Үcŵ��2���M��,����N o�@�4���] �0��W6�O�Ӱ1�Qa�>���I�ɱq���b5?���u����~u������t�����Q���O�ew�1@ǻ��I��p6�q�KD����	��.��}k�$�}��i)��"++��e��|�ar/ ���nf����m?Mfl�o�hz>��Jjf_�3:t����C�ih]7������-�e3��lj��sq�7
��@�o{0�[�^������bB"%W�Uv~n�N� �g������hq@������[�õ�Q�����w>�}|5 �����Z� J��e
�z��I��͹�T�&�˓�z<��#���T�'*�oQ"ݭ|ss��	z ��r�Tm^)Q@;���{��Q��i��R���&��������:W ��cd�dMom��ހmӏ��x�{6�������.ї\����_�>z��CUd˦�Ё=�[$;H �i���0��x%�r�(�y�F6��B����G?���,|a��g����}���/6O�A_J�����/����������}�����;o�g�{.\y������d3����ի_�_��JZ߷�f�B���?�Q�������Ȃ��֮v�dp!�(�+����99�zD�=5,;�(-0�$@<≲�,=���Y�<K��	Px�r�YgB�ޢ�9��L��c,���7�?������o���t�_��\���3`@|/Y7��
���>� <�Y�����U��?�PN鯼�J���T��㨎ҋfQ,`7�F|��'��7�P��p���������=�5pϑ�otdO��1�E� ���no�|x���W�a#�ch���>��# �x �wꏩ���� Q"{Ү����g;��u^L�O>�T�<Ua ,����T��νzt��~��TkWMI��{�1��`�~��dS�ZR��̥>�M�MoQH�d��}Ө{���_+ݎ��<����&�I'*i�|��{�����G��p+|��=#��G��7g�-�s9FSIYU���ܖ�ɭ~�l_�K���C�n9��v�Q݃^��r?����}�^�>_I�>�T�*�&_L��&�+�R[A��H����b�\���d�F^T�z�Q�۫O����I89��Ѣo��}O�j+.=Z+�<9f���О�}�*�n��'A5�+G�8�Hl48� ��",�Wt���S���~OC	A5U�f�-��?H�Jڵ^�t>����VS�L2�`ٹ=��H��0u��Q�l!� 4ܕ����^Л�opkeXf!���i�#��7UD�q�6.NIJ���~R�Y�]��[A@l��Gzgy����r��IE�U��[��p>�1kAv�D��L��+w��p�`���A�F���`�!�u�gy$}#c,0ŹF��K���j&�&��r����͙:O�����CV_�%�'�ڹ���- ��n���ޞ�U�l�' �_U�GY,V60�t^�8���v7C=��tT(s$8ZIElD/�=o��j5[v~�T�1���
�<+�(`T�ᜳdP��1/+����Q�o%�b e���j���ek�{��j��YZ��q�V��m2x=�c�<��Պ��<M���J<�z�����W�����R��U��$�}y��`�HY��6N�.�@t��C���m���}$�S�e�{j�!�>�ْb ���K�G�l����(�UE�="���c�9��W�l��Lt��Gh�Y���E�|`{�;o��G�C��a���|�2���J��
Q��^���K��LJ��j�G����Bh@L��#6�4{~�ޛ�\'HUbXr>�����2y�Ћ�����H�ׁG+w݆-pj�MLx�{2�������lSa�"�0sBh��Th����/��_�~���������k�j�CIz뭷����������k׮�+W^����}�3�W$��NNU��zܸq3����:oh�T!H�F������z��C�����"���[2�~������0�&v���-��lF���k����ǟ|n޼~��߆��/�l�uE^oP�I~�՗j>����;�c^1���	_#|���I����$�S�T�hTW�yqи.����j]nWq1q�	�Γ��*�
�E���r�1H����hi��kA�Y���#��#�  ����5��O
�y��2\��/�����O=-:���v^Ъ�㞬���EӸ���X�~`�w���Çv�$P� `"�9[xh"N������ݼu3���7��ѱ�J@n4?K�
9���,���X�L=̾ ���q�@I� ��pa���\d�x��[�4� ZT{8g�4�,��q\���i�Ĳ�]�(�: 	�Q���Se�96�s�N�r:�$����8E��>"C�لB��dr@Va{s'lN�ĭ$�Г�U[��h/���o��Č���;�V��T��~����9�nl!�:N�Z�Q�(��YozF���:���q��C��6���B=��aÀ�7�[�:���8��F�{w�9�l�&�^��pK��Pه�fGo�ԋ���c1�f+���/S4i��.=�PoYF�R�k�p#���x����A�@��@|�j&�J�S^�T.����otwx�]n10��P��L5���Q����ϳ�J�^&_@:��%e����^QUY�����jd��۵#(��׵s;��L|:ܛ��n*pg(�J�H�F�RpЗ8C��ձ����7)tUq8VU�x�ZN�{I�H $��������R�߬�(�u-\Y��ʎU{�z_�A��������1U������ϳq0f>و�u�,/�Cs)�ǉ�V�gh��q��8�^���G����W8��=<��Z�Z�H9e͟E��d��)�o@n@y/W�5�����d@3�oJ�8+��@!8��}���������DЀD��������㠎��C�R��n���D�mC�}溍��]��]�1Yn��9�i�%�~8<9#06fbP���v�<B���J�õKQz��2*-�X�Б�'ݲ���U�G��^��FѨ,^��c���x�b���r�y�EO��������+��<:����AYI�膜Eu�
ӈ�4��-��#�"���G=�n��wq_jtp��x4Y��X�����W6]޽p��,��i~�R���b6������*|̦�B��t�4P%��RB��n^��~x��o���]S�'�YC��,;�����y#�[G�H��	u�����u.d{�;�h{W��S�L��HZ�e#0q�|���D#������D�c[���h,8p�|�!Q��Ǧ�j+2u�#��	�qӃ��;�L�$���wD�� Hv�x�`Q=UB�����z&8���ޠ�G��&b�������4.߻9O �)1����7*>�z+Z6H3�s�
��v
񶔦l.~�0/���ާ� P�߾h' d�|��ja�u�V�q���/�f��=:>R�4���+W�O�S��^|�I�W�'JQ�q_O�q!Hz�r���dgr�̴��t�R���};pԤs�`@���鐞���'ZUg����N����pX�8�3�,�|��g���_o��Vx�ɧ��M���=��Q/J��1�_�� M�2�<0t��|�wl3�2u�z���~����?�.�_[[-,��p� nʭ���<ް���7�g��JE��xW���� �y�K*�Ix��Wlp�������<�����+��q��&��dס1��@m؈.�&.�\��|��0�ɞP��1I�,VS�<t�q�o�#^��g��ȯ�K���n,�d�҇�� )`6y6e����۪g����;��n���,W�/�����6����s�@o��w�-��GaA���l>C�|

�P(��C)A�дk���1��{�,�_IV������T��}C��{�ic ���
P8=9����{W�
s�4�>�V���h8��j+H���J���ߎyf��o|��6Ry�׽s2Q���${��@�� �M���q��|�ۺ�w��c�Tx#m!�ޕ���n�&͸�Pٕ��tt�Fk���.��p�+��l+|W��Y����c��)���L?���7�Zy!�2��l�L���l��#��3��(4�캿�*=1�X�ڤj���8��񱞒�OM�`#�5KԦll���J�$U��̍�7s�E��.�6�ww�:� tz��y�h��Tc��\G?��νoB�a�A����j%���4W8-0�qUT1h��0�i 	�B�Yo��-E�C�w  c�~~:yp������q�l}���"��#�q[�n߹��u�q�k���^Z}��P���m`od�ٯT�ȝ�Qs��S%Җv��ܸs+�ھwd���:/z�&�8�}�ƞT�w}8�;<��^��A�v7+t�� Ѝ�}q�^/vԱ �&c��u�г@�e��w�p���I.>V.��Q�Z�P�5���}��F��*o-1+"�+�~'Y�B�N���2�x|S��Q�#Kh�U��H�<�Ar�x8���q-�֍�2��� ߓ^���ceý`�aD�t�J�T���{P\gA����{ͤ�G��\J��4`��ƵE�#_��Tk,�޾�5��=8��U�8�"K,�D�%��KY1\o�[7�^�5�'z��;�ܩ�v��xO���/�Ń�MLp�D����~:|=HX�4��#��ub�,k=*\�����nU$x%��,$���SȞ�g/�Ђ��=�$���"��@[�2q�;_��[��������)dU�*ç�+>Q���ºA�A/��S�9H��!���ϔ��I�>m�#�ׇz�����zC?Ǯŧ��O>�D�磏>���U)�8o���,�{�B�
�����o�H�0�Q咔��K/^	?����_��_���<����hͥ�z�d2�\A�]9����\R)L�Hd3d�\���mjVE�eP��B����'�}.��u��.�84��o����>a��ɂ�`� �W׾�f����$7r�w�7��Nϒ�@,1�o����P^� ���?�ݒ�z������/<�x��[0Xh|���^טֻﾧC��w�JAh���n�Hq?�BPV�[x`�+U�?��G�;\�D�D!*�`��� o�Gd��w�\�\j3w���K&������}�ys��+7p��N��K���$�ĵ��������&=zì��Ij2*��?A?�@�u���l�揟Fq8��eMShzx|{�#n�k��v&i��6#��pP�[(Y���_!nmO�J��y6��;}e�s�,$�:��|"�V�t^8����X(�~�'T�x���-��l�:'�u!_<%�A	aY��І�A���*G��8���x'��]�����|�z8(-�Bd�e�Z.	#���3Ik�)hP���3���'c��H.-|�Q�<IWH�Fyj��� ����^)���THɘ���n�!UVq���h~���?�rY�ް�~���2�2Y�F�'o�-~N�����k��)�S��G�j�6�~�Cʊg5t3{No�Nu�kE�+�=`�e@UʽD�����ͯH�d�;8 �@>�t1��t:�!0ٜ_`����'A��$_��T���'�NbB�b,��fm �c+�&5 {��M٩}�%hTM�/�d�m�T~&?��
����cd(��B�x��	;ny�����.M)�VQ8Տ���*��f��1�2\��)0���$Ӽ,����3v�2�}s�w�o0>Jc �������N�o�yPߢ��΋�s��i������zoO�?t�v��*s�Q�*�t�鶎��^!��I�GZ����,����Z�ֳ��I�:�M��,jNU)��{E[��b��V�}3��|�c�<6��<}�t��B�a.%��N�k������c�
�>
T<����jG�YkW�lňdJ����#i�Yb�׸NL�,���'X�{ۀ�`��隆��G����ĐL�ȵ�eej�$��'�NQ��zY9ET�����f�U|?o:oM}w�{��į_���ek��}�%n�L�':��GTqM�+�B{��A$ �^���k�d�W�s��ߝ���qm���Gs���uef����P1"ՎK�]����"ܻ{?lonkе+�e�*���l��k	�1�3�Va$���T��J���֦�A�.��8b�2�0c�O0w�/X �����������?����qS� ��������ޘ�&)�W�Alw�·�tbBhRI�K"S�p�H����N��}`�(��>��SJ�_y�U�س�'��v�v|���4��sq�ڔ��`5�Z�W�L2K����H�*��#U�'�#_�<X!��vsn��>[���j���#�#0?v�1�=��SB�\�:q3�u�QZ��e%pW�ڰI�i.�#2L@b_<@:�Q���޸/&����K��PՄ ��o��k]+�Q���'Б�Ӧ��"��~��JQ��x�0��2�j�{5@�Hz��W���{!3�`;g��}�2��SUMpl���'A�d⠂&I���rvj�rl:����;e�D�K���#�>m��f���2�ٕN#s��!�J���  �ᠧl/4����J�W�?e�Jǘ�BNS�h�.]�?0Α�%k���C��k��:}�7�@�Ɓ�D�e�2N%�h�!	k��?�|���n����4�6��YPn��|V,o�BŸ(J�ч�3�K{�1U͕˧����,�4�o��\���/adb�(�=�I)��S7��\
R/��p�@�l��Ӣ�]�E��敲^=�A{��Sm�s��Iȭ������+����
�\�[��/1x2�qS�O ��U%��L*K��^*LıB��6[&�[>�����]��" ]V��P���7�z���I�lg.�m�H�aF�E��3��՜ޜ)��S����~�����QrU&2rې�>�=@�B�X����b��\���,��|d�J�������*b����㞽מ=�� M�\Ug� ��Z��A�.E�"��0���;�V��P�O�7f-	(z�`�p�V��X�^ ���z}W���dtQ ��5f��aW���}��LV
&\w������2�C�]�665G����^\ۚ�^��{n��c�����P@u� d���Dk��h
m���BG�<�b��p�%Ǭ�SƘ�E���3{�j���E���!�	R�'d:��#v�YC+I�����|�y��(���Iԏ��A��iV��U��$�XY�+IR;PU3tݯ���zpN~�����H�K��tN��ϩ�,�kP�yM*QdkOl<��@R��*�}3�"��W�r�b�����&1��?R������C隥�'��U��_����h.D:��U��F�'1�(e���n�jv�x���=��w�m��K�Ϋ��/����y�"���8H%��,11��|�����?�ll��XE�j-��zUclٍ��4���]J��,
=�ފ��c�G�D�^D��t�Y��G{V����7�=������6��s$��5q2R��������Ӫ����K��^�!4����\�G�[w��)�t�g�> ��/�n���*8����JՎ�p�\�ݫ����w����/�R��.]�����E��z5����?j����{���Šω��D~�c�S��2�(��;wnG���J5��?h�d}�D���9�P��ԟ��(9���ʲƳB��W7_/�`I�^K�� 9��N)������(emk��ֲ�L��r�A���
�oO^��U��+�UM�FW1{�L�(?=��b���Ց�� |�g���.�5��݇~�����]+�NlL��:W"j(��I�;(��>��#x|Tyh��������� dp��@|Nr@O�~����o\���s�=@� �,��1qS#�{z�� 6�"�T�΢ĳ�>�,r��_ݿu�D\P�o.���֗��H�N���T^�"�?x�=l��T���=�da�_��eV�mm/�n6�Yz�*��g�}�D
W��Jep��L�^k���^4�2``��S�MÑ���2ǃQxlw?�"���@L��>BA;�)c�G]+{�t-�4I�.K��#���тZ<��)���Q)Y3KQ�z�L�f��̠��pA�:SD#���(]��6��Þ���+d_ <�W�����dm��*��.�*�!�Ӯ<.�zE�{���9�����,�f�VQ���h�We���Ju��		T�&c6)+5�)sgl�wӹW80I拓�ۗ�t9���������y^�6e*������(��G.l�����G"8���8WZ$V(0��Xs\�
��mȵ��M�T}gi����y��_\t��d#��FI��jH��fa6{�C��\�i���jY7`�ֽ[y��q��!�����nU4�RO�$����
Q�2n�������-�gM�͏!�`6;�Yi��6�����w�pjsrn�3�]TPN�ˤ?ҍ��(�Lp���	Jm�0�n�r沿s�S �� �®ÉOS��y(���T���S�.�p^8��iK�hɤ����
1j%i�^��]�|�K�hh�{�W�М�I^� ���6������J�(�ɫ ��9�,��E�Mr.|
���Ƚ�V��b��}fg��џ����r��s6���J�8y�n��R��^���lv�K�/���km�7E+U�]iJ�Ϻ�h��t��'O�*��+U&�׺{nT.�]G��h���`k�0�R���H�2��UV�5�����)^�x�ҙ�1�b�Fi-����������ln iz��W���Ɇ;}�PnmR�c�&��ҁ}�� sG롛*b��ARYǎ�kngg��1I��g��?qI\��������CJ���k׿�z�ēOD�#����)���DV�;&�E��o��7��/	4��/~!�L�W���˯�E���ŋ�(�^��KN�/���î��ۈM�&�K&���A��Y�J�o�����EL����T-��{|aׇ8������:���;��^��������z*�F�E9Ky�G��h �#�&F.��7EGK�U͔	�{�l���E���#�)��?�`�InJHip��F�Ԟ?ߍq!g������1姧ON�L-��ʫZ0c	X�xY*��zn亁��D��]+�+G8I޽+*�X�A�jT�t�����0��N3(�pp�@re����ǺA�Z% ��t= w rd� �����=#ܥ���W_|)�����w�a�s�(pL	ҷpz�T��f}$�A��/?gh����he�l9mk�p�i��K �k��b�������%����B�}%��ת\Q��RAV�~x촟�>�X��C��gU���b$ύ�6����㶪d��·[�g\*�2�ړ�E�1X*K_)�e�`A���0�L!5;�*Ȗ�����d+�f����a�O���SQDxn��(^M25S��'2��W\�w&[����޳�s�����X�$�,j�&���z�p���@rI���YSz7
�ĲYp�z+<;V���Q�:M����M3x�T�S�0_M����Q(s��f����]��[*+N 8������C�:Vt�se��OI"7�ha��#�ܣ7���YѬFj ^̴��1�Nv���}�&PO�@�,&L2�ąU��8�R�:�B�M�(5�&=�������z�Ͻ/EY��I#��\>8��}��U�?�U�=(`��Ɖ�8��4T��ҩnHL�녎U�?�6�U/��h2�9�>��x���>�)��C��I?�}VߠGU�3J{���V���<�K�T=��v�2�]�J�j����9�bI�fF�wԸε�_�Ve�����0������D� {�p�Trm���9�����)l ������_й���N��TBH�QXI}��8��%�{��*�q]Z	�g$��:
�Ta���֩��lH��oY��"�x�	������M�y֚�1���I�����S���>��k���$ћ�+1�[�~��P�jΙ�J�E:�wgN�9��oVXL�	���mv,��>h�eq>�G��oE��)	����u���w�ԯ�SS��X�{N���xTnPZ�C��rJlH���,:��H>�1��q]�m�\��6�ᅦѶ���50��uɃI����Z�Eю1������vč�\�����#c<�)�3�G��ȸI��9�uN����J%��H�7�Mx�	0�Cn��>��`�`ڏ�P5G�� ��I¢2��3τ-��p)'qE��$�{�bK�����ǡb,h����u�?�^����2��y���������>w��_��tl�x]�"�Wٵ"V�jDL���%��E�F:==ў�zJ����_�`�=�a૯������zRT*�`FN?3����al͵C$�׾/K
*?.6�KYl�.��1G��_�V�.��Q�����庀E�&s�iM�9��n|�Z����Cw!�~g!���ߡ8���:|��g:�����ta�\���!ɕ��*_.��:	m���,�ݪ5JbӴ!$�>�O�������u@��Z�Z��m��<�(`���\��j��{Q	�Z����Ӯ���wB��1���vMvw�4aQC���������;t
�Y4�"���\����˗]m���|���W��UT2Ȭ��>s�o@�8�Q��*[��0S�!V��nz'��Bg3io}���{��j��s����0fe�����zΜx�Ǵ����)x/�giB��7���:Ȳ�D��={��V�K8:C�Q��J�K�\9���\��~#L�.|��4���{ 0�䢄QO}Q'���qz%x�}0L��s�9���7��YO��\
�3{�ytw�WY0:/��~X����=q���_	����l���k7��J�a['u@�u�=�җ+oGyJ�u�4���noDáJ�D��kX��Y�x�x9��۹�?<��4}2H��d	����m}ʩ-��A�0��`]��賖�72�4�d�T5�+�X�ڔ��id��Z����G��C�u��뗏�,����]�)PPU��1�����W!�t�<}UD�Q#���3Q{����P!���8�1P+	�,2�4��6nX�J)f9�I� �q��c����w�}C�g�>���T�Έ5
O�s����S��̂k��oA/�/Km��vC����}n/%
]�ՋR�q
hR���(_�b# ���:[J2xj`fA�&�����^LZA����/[��}��ذ�K��b� �ɸF��z�P.H%7��ql�h�֢|�6�d�v/��<_ɝ;J�����u�ڛ��f5{�~��]�J�$6T�f��ʕ^'��K���q-o9���fM�#G?-�R*����Hի�{��n8�i����b��C��o6��z=μ�y]�?u�&O�r�}��^u#��D �2�C�,���D�HT�-���&鮟c#y���%_GU쟣
��X��"U�>�C�Y�oAp��u��8{�?9����Œ[m( ���(R\��Z-Y��ݿ�L�_�����n˖�K���)�HPk�1�{�{���$;�T�*3#cy��=��{N{!7��M�o�_}"Ht܄�$����1�{o�JA-	[nk�����(����}.�g�o��}�cg���'��8�/e�C��9S���u�����݆u�_�	��|P� �O Κ�|����i��fE��;�_���꫿�� )H�v5)o���>T��b8�{�3f�^���K%�%bds��B.]��~>(Sĸ�I��0H���:<�Ն��PO�a�Ӎ��%���Ո����»B9#�h|�_��5�4.��$эz֗�����K/�W^�ex�@�?��?I�����N�������s��ܫ|k�].�yP��N1w!������
���Ce�j)ܬ5��N����0�@�x�=���}4K'O����c[V0�S��r�������W��N�(�<=9_y�+�V��i���b��urb��c��������8��>�'?�������o~��c*�]�rY ")��bf�G���A��t�m�|>���v��g�:ة*(yF���==)'��*y��荗Ҹv)#��X���������o^U����,��b�.�?��3�L{��5���i!�R|(m@�UPL��������R���]�u��#��M7��BG#��E�����5��w�~V�?	m�K�o���[t�L�?�W](�����L+a�LO�p��ɂ�u������H�W�G��֐�$���69�����q��}���O|a���ի��?�i��*���Gl�j�g/��#�`t-�}X �0P�c �2�<~�(n4k�Q��s�պаݟ�=
{;�aa��]=��ۂ�4�(n����-T	�yP6#:��?<w���"�~��©2�Cb���-��@�k;����:�lsx]0�Cc�����X||��Ypi��R��;���׶`.�Ǫz1k�*E�!�+(J;� o���1��(&�8�����>r��;kt��US��wk,bE����^�=k�Qe�:���]2rP�e�{���r�Q�� P֢�b4�w�&��RU�����Ֆ�����'<דs<=;	C�/��,�GE=d>����v+2�\s�K�� �!�� ��:�c��+[��a:?Wh��b@gUA!8�Q���n�7?���P��r8��r�J6����K�������rb���9�F��ߩ�#�휮��S�l,+<�R@sS4h\;8-s=�\`���{s����Y��RP�l�	_/�Kԗ�i���f]О>��nn��f�[p�Q|R�I���tX�؀k1��|l�O	��H��N�I}i�=�ͽ4H*���'��C�ݼ���R�c�qQ�;�a3C��-]+�#�Ԑ;�*y�]�+�^�C������D�r����#ʚ�(&�{I���wx��}��XV�=�?��纊���JT,LO������6��������b�V����o�kAO\����\o�b���%Pj��%౿�^p	`�M%u>Cݪ�q��E$�ʁ�5��W��>�>Jg�佢U�^�b�T�L4t�?f�_����S�[�o,��"	�����/g�7�
_����׾�5�W:w��.�gJX�9,P�"�>??S��u�H�(��a���"�_7D��[I��y�n-��9b��T$~���g Ķ��9$�8���G?R���r�`���w�g����W�|\i$ix��u%����/�'Q&��y�=��&�k]�"-�[E�
��0�]��>o�n/�ʱ+�:��u�Ac�""�,�eqEɢtc�H|�6ݸ��Ҁ�{�~7B���|�tc>*��/�G�!LS@h4� 8�[�`���	�ؐ��<w�[�:��.��fA<�&���7xP
$�_G^,�����k ��S��z3&�x�F�O�Bq�0\hR���d3�1SƓ��`a� ��#�k\#����-_�;��$��m�|���ce�=!���㏇������x��P9·\�D��!bӨ1֯}s��}�c{����7���c`�c�F Jf�Ľx��6��F����"tKXO����ߩ����#�,""�",�4P:�s�Gv�{�)�61���z�E��]�v`F��$�4p�+�d5��&/_��]=ZPCp�}�6�EF|a?��S����*ۣ�Ku�{nN�-
H��N�Ei��C#�'<-����%`q�fE1�@/��w�d�A�KN�R���w������*r����z�h�N�ZHV+W�✉�'Yԗ�Ye@'S`�'_�U��8Ȣ�]e0�!;���
դZYB�]�e(��9����AeLj&
� �`�@����8�	�q�V��M�����,�P`­~9�Ɠ�MN��M�����T��#�XBO�Σx4��N���	p��ta��4�#7�c*Y8����Ve2�c�,A>C�$����Db��W�����*���L`"S�5�jV�TUp<[�?��YPa�t����E�YJT�g�X��m�?e�K)�VZ���p/�*�qec�cnԹ3i��8(���C/���*�MPs�RR���dܗ�]]���D�'y��4��md�;�����2��b������h�9]�	���Yٛ{��v�1\>Z�
�zt��3����=ٟ����4�
�����B�r�ƭ�5=h�u�9#�,���Պ%`�4Sd'����e�6���l���i���_|{Y��E�������>��r��X�V��}M����U��%E�ƒ�p�f&ߞ,����A�,�)b��^�����q7u^�R�E�z�y�zR�⿽�nס$럎�ײ��׷����~ꝣ84�R"8o�ĜT��M戤,��J@M\���A�VtT�����'�:5Tn�)W�7$>e�{o���f����~�$e�����-V#�𐠥���A89ujb���E�������?~O�r�!V�M������A���JQ���s�m8��aq �Co&k-�( ��~�S��p�{T-%��5&�����j��\`@�J���9�G�\�B��u�}���wb�����]�?cMl�*VDm�Tr(��#*�{�=���@)'��V��u�l�(��*u٤z|t׹�r�ldyI�ҁ��Xċ�V:uIT��B6�Ӂ�g�e�4a�I�?H���ˆ�@�?�a���mC�?�����Ă�K�GU����x�&��J)8U�(���%�ZC������'o<���/��}�{��SO���Pq���>s��������}�i�\��������?�^�
������V��ƶ(�朽L?!eL�C@�N�-�����H(��'?Ŋm_z�!w:m\�����`�>j�}i�&"����M��7�ɱ0�D�Ie��ELU���	����~*=�.CQ�mi��Wj�%�]�<3�k7��ᦡ�����>g�b��7�z�n ��Ã}�9�7Q���&E8س �|�*��Hs�2���dw��-�������g��\޷	��%eKh�=���K�7ۘ]��
<˰����bb�������8]7>��&Q���6��]( S�V���~L��L��\�!�B1�!>fQ���Ugw-i��ى�N�x�iܵIr6��E�,9��ŕ���l']
Y�V�O�\y#7Fr!�K�ǅO��leʮ�q�eޘ��T$�{X[�9?��;2�C���<(���n�3\Jbw���X��Ol�NV-�Q''ʼ�(V&��>5�*i dw�ܮ��E3��gp=~��[��0̅��+:�������7^� ��l��5)H\jq�;6J[,J�w4N������R<�u��@���PAU����`_�H� j��}�ռ���H�y@�Rdy'��*ժz�9�J�.��n�h�~��Ǆ��a����M7�9��ro.-���~�nP�;c�ҙ�6P��b�ϏC��K�gH�Ms 9Ȭ�%�*���`9tGc]��I�|��'J��򰿫JUեA5�#�����TQ���6y��w�L
ַ%o��8R~B�Z̳d��C)�h�6�(6]���mbD@�LYݗ�����x���]�6x���M �W+!�pyl*�r��p쵦�grX[��o"[l�t�`��ZX�5!�����`l�Y<����,�^�害Du�[�g���&�Y�綩��G:�Ɠ0��ǪG@z��q�bK�J�.O�V�4iz�m�N���|�j�Cc��q�C��RѤz+g㝱��bR����\����]���1q�q �ITx̣Ly�Q��@ڸ�[����M�wSȠ�헿�e���gK�������*��d���@��^��0���]�O<��j<�܀�|��r�q��g :.���8*-r�V�8G#�����Ϧ�1I�?�H1��ɩ����Rǂ��E�_�$�8fb~�b��x�?�}�����Du�;��m�q����l�E,��3 �}���1��+�I��7xJ��3-�gj��r���r���r!Uƶ`�Π"�a{3�OZyB�1s�\O��6b�t��~������n���=x��4�$3`@`o���>D�=��+=h�ߒ=��W�p\�l�LՒ�nܐ�GG4���wVF�j%1�A��W
P�>�d����T~c`��?~�f �h\$P%����pt3�QP�&6/%�_nn%�-��m@�=�ƓOJ�����ڗ�ա4���|jW>�w��7گo~㛾���!�`x�M�&���/z4񂦉0��M��&�Y�m} ��&�4�:�Lq~)3��S��X&�r�VQmk&��l�ݴ�{��g��MTl�14]��[�,��� ��v�v������s��W#a֪ad�Rj&���R)�������^�)6<�`��6��	��Ȃ�R�J�����p%��l��c�ǹ��<�]i��7���jbS���D��}!���@7�̭�`�&���ce�i��W�y�����X�j�ՉEy3��
�* G'g��Pu��+?����b�T��Ǒ���GH��c��rnm;{vl��?On��I�ė����W����(��־��Sz�з�~��7]�!��7gWvr�Є���KHdB�X��?8P3B�*�=㧢t5��B?�1��Ɗ�-�;dQ��*P*�Z'a�4����E(�|��|M��FN���ZcP~4Á�QM��x�w��c�c\���nQI*�",";a��1�����K������U�J�L+�Wa���\������������K�U*�\X3)�ȵ���Ɏ$���w�	$�tT:�B����<T�Ñ(q�Еۂ��^C>}�lmf��<B#}�����b����G"T�;��"z�S��7�e� +ziZ�1��J�4[������яRE��k��(�e�"RPC4�-�2�Z�/��
�'�艐���wuSmZ�S ܤ8�7o~W�!��ݩ� M��J��v�J��g�y�ˬāhǞnd%�
KQ��G�k]<zrS-���fr�T~�$*[�ҳU|��G������ݪ���-��CK�J��fc\v�k�)��h[J�V���9P{S���f���$QޕA��)O��8)�d��A��
V��˻�q�b6�x���4]�N���+�=��>��"��i����-�k_��*��#%�I</��?��㊧��b�b��Cl�8��_V���H�y`1 4h���uC��{�G Ds�=�+�*��R��������� �"I�<8��A,��~�e�'�x��y?ʮD�����
m�W�=�I�S^>M#����b?���0Ő�c���J��^��J�藁|�x��O�* @�X����T��R�B��a<�AJ܏U�IT ���\���L�=��&�H��e�Uf�J�iSf��~�T�@1��78�o���ɁN(A:���.4 }�ڀ���O�B>��Bs �v#�F}p�ZYxɋM`���'~1dx�-
^\!�K�)Ĺ����i�|�+_� Pf:sS:nZxt0�?���*�1��9<���	������yl(��5��ָ��߹�F� Б)��A�dQ�a�$�f�"�����{ٶOq�6߷9=��[��䤠E�4zȬ�N��A�M��[v�n���� Mߘ^�Y�,M�R�
̢�r�+{VR�8;?��f��yу@��^b�Q���F�|᨝.'�̍�h�n�I(���G�/^���n߽+S7|cF6i�Pw0���|8���1vb����C7̽����ƣ�3[X/=��~��&o�?
��8�����i���d ~+�F{Y$h���qT&/��M]��l�d���.v�hg"��*�\��1��l���tQ��py��!.�[�l��ҮIq��1` a0����)ٹ:�d�ίܠϫ��$6K�Hd��T�SQ{�2�����@3�R4� �U�٢��7���R���q�\<&�ЃTq*���kB5W���΁v]PF����2s�GՌG:�X ��Wy��ܓ	lKy�� n()¬��m�Q���	��n�H�P�%�_=o��5�4����e1�N}(�BeR[�I>�P�2���*$N#�#�g�3~TCPmT4v����%*c����͛a��lF9}��8ɩ�|wr~��G4���3�jLє����k @	�,��;���q��{{w�3�Wu��y����|��t3N���к����ԛ��Ǎ�ns)��Z��#I����,�g(��w��G���i�UT�J!�vR�ݕ��&�ݙ�F.bSǄK�p7?���g�,ǖ6т����l��ql����>5�IO?vW�rI� u@_-r��(��F�M>a��v������ՓJ2����$��)WMz�}l���;���ت�>+�d_��bL/�^N)�~��2ߨY�KH�\�+��09�x���P�{м#������3*]6��DQAKӉ8�Y/�Z��Tq�7�읙�ڳ�Zڍ!�5;��c�?U�֮�JϮ뀎�}�2J���{O>�����<���IQ���4��<��q{��5P�S� R֥L�9��t�wO��bA���$(c$���/���ZԨ�T��8lA�\�1CE�~:S���e&�LZX�(��TM3�g��vP�X!���Mũ��}��#�j'*5%>�2:�&���D��F�&9���ӠN|/2����o$��Cَ4Qe��9��Y��_x���(qaF�;��F���M}�O�n�B�x�NVU���PC��en��]XLf|'}ulK��.]��e�Q��l�z�2�1��bvhN";��'?�i��o^{����_<>g�
��YKj���:6�DS9JZEU�"6��LW��fbTM`%���a|"�ȃ�Oeb)��M����f mf��� H
�{�(�*Bo��Yp���Y�����g�Z�#w:%XC��F��j<s�qejh�֕~���!�����Ӱ�)�\?OO�D��q��;�I4���*P�/�'�!hG`H��R-b<0��)q���}7T�����|�q����㓐��9�Ҕg�|\�$��?��,���ϔ]G���#�W�][@S)L�3^�<<��Sm��1�a�5[�\}J���*,P��ܳ�2��}%eBB5+�0o�a^T��U:�1���Vn>78�J�Օ7FG.��"9)˝�)�I�_��p�p�k�V�BE��`n�g3[ Nga�c��z.ό���Y�l�VI�Pt�
�xF?�b`m�V�x-�q*8���i^���e���T| �)=�y�\�B	A�b1�y�2��~��"�jR)d�+�p뙨o�g�5:����W�g��� M{*;�OɺN@�>�N���`�B�`�H�Ů��睱�۟�@*sܓutW �y�����ީ�g6G�m1=({�od�+��i*��#���>>�%)��g��+J�%ܾsl����Ex 0��VӴ����1pjk�#�Uu ؅�r��>�3�w��a 	Cǳ��p��i�o��2u�� �*�R&��E+=�l�n]��@��"��A������.N�ch����?7�P����X�je�[�q����>�[�s��%���m�%
[�����7��zs�j��Ո��D��}l�.-���G'�����������X�K���e���)�WT'��*�Y��s������4���.�*��jG:�^2�?��7f�xb'H<�n�����\+�l����'m'^����h�D��<��h�����+����ꕜ&�����wէW;e�i�\ݮ�~e�hϕT���Տ{�v߷����Gz_:<`	Q!��]Wcx�+��u!��@�lY��:П��i�$q�U*ue��ؙd�`��ATKZ�Sh�Z=�kijT��=Ū�$���^zY��$ѹ�;�]Y=��l���ؕ�=5���}o��'ŘB"���Et�g7�y���~�D8R�Ħĺ�9!�D���b]�xh��淾���"e������i˰]����J�D	ӘͲ �eϥ�Ӵ���A��$���y/:�|���!�w�ڞtC��Nc�<`H��=����"BO�u2vĭ#��D�;�b���R7[m�U�dU.��``۸�÷�'��Ft9zI8����BH���]!M����n 䏯���� \T�w���z���^�!RR�7��v���3|������q���y�\n�z J��td�So��q�RͮM�*&�ۮ�ٚ��zwY����}����G�}�a�B���Kq�g�Ydez�.S�d����==J�f���9�݈͝��"H��v6?����ix��~��� ՝��������FW�l��RIV+pQi>C����ܕ�~�]	o�i�]�O>�T��S��/Y�^�k6��=�w����(^����1�:H�f��ږ��tml\��D�c�� uu�\}*n�ݽ��#Y�Yd�U-�����p�m�'ʰ�:����'j%v]F�y�^n��!;g��wgazvd�>�:}#��[�L���M;w{�[�1i�x:#)M��6�w3UyF����P2%^�8:?�s���o���-������v�q��T��S��֮���QA�f����\��"��C�@J=*s��Z� _P�*m�p ��|Y�<�v���[T>�px�Z�����i� יc���x(��� #�����5�s=s|>
��u]�	��,E���541���Vz�s�1)� <+VNIS�[�A4���D�dG�Z�U�̔�2�^>*Q�#�;���@��g�u8���+Ur��I���\���`'����<>=猡�G�L�ێ�$h_�?2761U�@���eT���%���zy��$=��$���PCXk�f+Vk��j�ǩ�C���w���'ΰ����S�:͸�`��M�K�_��vNɩ��9�n6��;�>��~)��~����Eс�:��H�7(ܞ��<|�i�n�@�>�DXӂ�`�5���:�$ʖG���+�n"���~�Y���z_�]�HsJ��h7�j�
�u�hޯ|$$�% ڎ���D���D`���2_�Fi'�0A��%��E���*�(��8�bn�{�!����{��(�G%\UD����#���H��iu<���<�������N�����qQ��}ʣ�q�E?���M���
�P|%�#�p�^�䃖�9��t$,���54v{2)T� �K�敪�g�m��t]G�Z �;T�o+P�L�bL��	�o�z��~+S��Jv�s7��rճ�<F�H�-�ڞ����?�$���?���o�ۄ;�K�O�)�z�����k��r Y|�u i��8yp���W�s���� 3�8�H)W����pdY���S�b��(�[$enB/0��/z\0a��m���M6��K�7��R�
Y��x� ���@R��Krl݀��*�A�S��x饯����+��RA��������#Jf�'A��W^yE
]���K �a���c(.�SO�� ~T�jo�J�"�����������;w%���8�-	ŃN/�^��R���jM8?7�d�a~U�v�o6B����}:�Y�׸�Ro.�M��l<��W�ݐ��X|sL�N�\�V�%ƪq�i��g�M ��������dҩ��j����M��'���ͷ�Ε�'@V�""��w$���C���M3�֑M���A�zd�e2W%�1l�������7��lL������@垍���>{:��"qS��D$�M�������e4ٿN?�0��hQ�ëb\g�'�N�Āͺ��-N��|p,@�☆����w@�kBpYN2q�TuJ}2)�4D�0��`����ln���K�	!$��e��
o"м<�Ƽ�*z���.}&��̾o�pip��,�x�el>ܵ�}~<S���ƕM�J=�%*;��I�Hqˮψ�}�fcUA�7������4������ٙ�DK:�������{�\'6n����+��\�]U�֍S �]l�[�xT���T-T���.b�� C�u��5T�H
YE-	i�p�>3T7���o8��A����1�
��	�S�ce�Rk>r���tjdM��HՉ�� *��'g�<�p'�������Kv����E�� w3Ƽ�j=�ך�{pMM�M�.W�M1PǶ�5������}�k_.�ޕC?#wc�+����;�G�w�U+��o�ͺ�×�-�H�����QN7穦e��js��~%� �� $�]�,G "�u���t�Ԫq_�(@�v<�,��=o�Lp[	�f�����u+����=ͽ�~�b�$s��T(P8+YY����)Uu����PH�w2�쉪��B�S���X���^ţ���;�T��̿�wl�u`�Be�����M
��wγ^��{5֢��$�?�eL��*y�\�=i�41U8RoQ<WI�(�:�����dk�=��������F�������M���x�Cxf����?8)E�bBY����#�S�˒�k�yY#�����x;O��<q^E������Y;��_7�c�+��bV�Өb�,��Q���G�[x;���?R�UHZ�D�i=��b��$9#���0/��=���J�s-Qq�2B�ɱ��V[B��+9I
@�*�L`�q�w%�K#y!�HKG��qY�34z�&�#�>1%Б,�Ӭ��Tv���?1�&b��+G��z���hڒNv3��G��Tj��L�'��<ƔAZGD�&����>D���� 5-n�'��!3o<���{��A/�(�rT���'�4�#�u��� ���l�C�U�&��R�g-������r<�������_���N����e�@���4�"z^�~�s�'�+�%���غ�/�Au��Jn����D�h�B��3�s(���^4LFP1�씦���u���{]�6fbz�l�Sd�(aW���Q��5��qΦ�0��}���&�Uu*��{�ʒ�;�(q�ZU���}����tV����:�ݺ������S��#gz���}��*{c*��X�6ڛ��;�ݝ�Pi	�#���B	�(IPxPt����	�0s�Ub�:���::̫�d�A5��8�O@%���j(��3�j�\��{��:���s6Q��/�ݥ2�y�;|P�#!���%O��
>��P>�`�,�k�>�Z�h4V�>�WA ��J[�n)?U����:p�������ݬ����ހ����GWԻ�Y �}Y$�;��Eb%�� �MT�rƘ�a��h`@hqtFp�����K>d_�Hfx6n��-���p�藪8C����62���J��2u�)�+�CP��T.��i�U��!�2^������/z2���fw�H��J�VA?R�;{�(]����I 4�PKѤ��yѼ�}��k��d��0�r���
���|?T���@I�>���9��\x ��\>���H�4��5���식�+=�6v�M��-w��qk�W��Fǵ^�ɥILJҡǟ��H�cк��Rc�{׼�߲��zkP��$�~s�RZo��66E7�H
f�X�����lU�\}�>GuǴ�,�����j��$o�xd����	���k�ds�W������ih}�O��.	��>�4�_
?jۈ�\Mt�.�Wʥ���\'o�>�QJW�s���	�l�� ^�I���U����6�we�6�o���zS���n���E��4+���TO��x�e���!RTc=�#�**x%F��6{B5�61e:Y��4!��P�����q����d�����z�So:��#���f�Xu彵�	�IR6ň����GV;���+"�=�.�  s���Ą�v���uޞ�:R������9?8M�Xb= ����U��c[�88>>ұ�wBA�x3Z'7�x�6��n�
��n��M�|��׾n��j0�u�����FՔ��GZ'X�D�d_ʈγd��b��Y�C�Ȃ\$��o8�38�0��t��EȚ����>�����S���2�&/������m5"�J�DTu�^����,�O�YȺW&�ঊmU��D��O�f�hx�Y�\P@P��*vv&�f����
8C�)o�)�_��~*�IB��T`��'�� m���9W5K��x�a��5��W^
�b�|hZ���!�&՗�n&�B��;��
����r#q������/�(�t1���亀=M�E������m'�l{�i�L��Abf^�D�X,cP⭀q;��u������3�x�e!z�(6yPN, e�arZ�W�@�@A��l1� T��?K�n��j���Rwl���� ބ��=eGh�k�΁�d���� T�\�Ȏ����!Kۯ!��I&���r��w*ԧq��(�����$�,H�,���E2U[-�j4E��B&��P�lL�Ex�w�d��.!(	�Z�|@o��p����_�����LN������e*�콫�e/�>�6�X��V���~RZf2��@yS�&{�_�o|>��!_��;NZg���M�L#(��=��d�LP�Jw����s�d�\Յ`�k.��hu^��}�u�K2R9s�����!̵N���IhV�N����׋}tg��zlTd���ĪG6i�6�̸'t+���ξ�P��)O����hnRٜ$M1y�*A�ud��P����8fTe�:��:��|���/1� Q���k��~F��pP����@��iO+��@���*�+Iz���O���źp��=[�N�zSK��;a��k��-�p���������ј��s�Z4Z�&�=;Gv��fx��8lt��l~#ե����|�?�Z�r�X�Re�S�})[�J/����AK/1�Ľ�)���T��AU�d=��?�J��,m!������������f�YV��uߞzQ�*����&ۮ�ak�Oێ	����?]�p�c땍f�=����{�������C*6��N��{�JO.�z�c�=5m嫳��ߛ�[�KN�Q�]�����ټ��?6�[[,; �2�I��I}7Y��q�޶�+������﹭)Fdm�}|�ĕ��}�(�M�E��4/��6���"�c����z>��s݂W�Uk��N�����.��6_�(�d��p`�������)�b2�C����g)TI�p�w����24&~b�@���Y�3i��P5 ܜ����Bb��ǟ�O]�t�طɂܝ���&~�e`�G�Y
$��NRS;��.��1�!1&�&I���;gm��N,�,��۟|�u��([���K�9�Lw��j�$�1A<����D�E�l̴�(w�5��Ń48m3�[h��� �S3Z�l>�x�x�PX��}�����g��3�ZF����&��L��ܹ}���S��m�'�����,.�@5q�d���bV���j�/����Bj6O�#��8���v*GR2۳�u�n^��B���Jua�������K��`�}�������w@0`������~X�T{��e4�l`2h��v��?��#9}�c5��mbRH�1	��۾���rޟźs�f�Ϳ�G�E�??��+F��R�A�K�eq-u�A�H̍3M��2$[4�6��m��y�M�_����(q�3�M��p6�q{�@����:�7�O�y�����դB&�2����������0=������pn�����`��s{�̂;' o�e��#X�ʷ���������@�}��]:8���x��}�*�jyXG�"NiE��;��
7J̳�4U)-��da�ͤ�)�&HQ"yJ�>��5��-x��?e�Ad3,�X�^�Ll�{�o�t�xS�����k��2���ܢ�4�U#�>$�(��^���eC5�#��T^a7,l�	��U|dl�j�V�].A�)Q4œɚh|h.H�("��+UI����P�rE
�;Ǩ8A���R��@�}�q �Q�
U����,DQ�Ճ���$���0��^4� jhq>����>谠7Ɠy�n2(0 c�^5KO�z�zmHle�����<d8�RՕLf)�9�u�*�T���`
/�l*����Q�j�XK꼗��D!,�h�ָA�p<T��1��)�$�r�TKfc��}&�Z�6#cx�M�$�G���.������Xc�* ��Pq���z��X��kb�ڥ�~�s�n(����u&����4��.]����p�>��O���x��4k�b ��B7���'�"���`�Z?h #��$y^���4GW��)�"%�sЫ�t-�[	���#�+=L�?��}s�_-i�\mU	"���hH����KX���]~׳�\j�'Z�Qp��ζ(��^�	p��̓`Kvo��½�6�i�<5Q�*Yvץ���Z(�AQ1Ft��4{&��(��ڌbƅ���$���u����c@�K�JRE�L��F̾�q��JG�<Tھ��~�[�@��N�p����k��!U<h�&n�q�b�T�y��Gt_p�$eʼ�Ih�~��_
D��⋲l����BL�gm�xzr�}����?�Q۠�JI�G,~�PH��'e�<xk?0z���A����E2 �d�� lߩX�Y�	�l�ϑ���$�T='�^��?�"���'�P��Xy�@�T�&c)Ď�+��%�đB,�Sdiɀq��y��b;�ߓ�������o���pݙhG$CH��v���5 ܈-&e�e��q״��y+I��ɳ���M�?z@$�x�G�*��E�N�]�ɷ|����&��� �t�-����c�t�2�!Z]�ݷ��U��E�^w��7jB���Rs�+o9�a�Z\U���RA�s�����ZB�t΀�y����C773���tV�:t�&%�lP��S�9??�Q������_�:���;���BNrxi*k{��t��Y�|7���?�H@6�đ��u�̖b�=<T$��.61�Vs�����Wtv�i�p�rƙ����k��5��Y�B��i���Z�����݅}�J�
��V�,L�K:��$w���, ::���15;=7зoA�N8��`x��2��G6Y<x�0T7?QB@�#�X�AfN�m�h [�}>�������$(���_�"���qл�8��q89�,\i���.e��$ �Zm�R�$H��TU%_�X��٬fq��
�*�EКU������Q/_N��l0y�[C�U��g�\�U�j��h���R�
���MXLW0~$ P�w-�o�M*7c�S�a�Ut�^�d������y�^e�J�>CH����e�X�zP���G&o��OHJky(N6��seUX9�'�'$�
���|6�}���Oӈ.�y��[�C�QDC)�� *%A{�թ�:�K�W�מ�UjC0L*�Ro��G�Z�u�L>�s]�/� �f�[X�����μ������˼^H��G��e���5)���8b=���:T�#4�B٠���Q�'G'j"��B� Yz��3���2ܺs3���h�w��降�ʀK�ʠm�p��o�m�޵�\�W糰{�1Ĝ;;>�T�b�[}4(xe��b�{��u���a�%���С7	'�ѽ��I,nvs���l4�G��r�q-M�e��T��C�*+./<��簳v��1�SǱ�"����;B�d\���B_x��g_�[�w���VA*oi��I}�����D��|$q���W}Iߒ�
t��뱎@�}��y��_n���{{Z:�?s}�h<Y���|�}L~��Z�>�Ne�qq r��;��Q�R@�s��#8K�#1��Y�����E� �,]�8#�A3H�����}�a�{76wh���kП����/~���W~��s>^�ϡ���M��$"��Y�۷^`�� J�0R�� ���^|��Z<w<H������W_�Y����/���
ε������\���<{��m��Sb;}�Qx�ׯ
p<y�-#�{�y��v큘H����}У��s����\���)��<A���p�	��f�_!�s�A�G� ����'�PMa<8ZP����M�*���������y��b�$3���8\:؏�t�zL7��������4$������ �}5� �VRG���{u
D������ur+]+�+wVU8<��!]��WР+bb�vgtu���{��o��Ȕ��!_�@џ޼)tL@��^8����4�<�P�l�߸���Q��O>"�����/���?��|��u�d�h����z�w�B���2���u��p!����8&����jN����o|C�G��)��1K��%��\]P��B���M+�뒴��N �E���%M�U^��?!��D��� )-�������&l�Ti��|z�2���S�g����x7��� #��RA���4F�W�8����]�Q�x��%w�&\{��K�-�t��S8�m�Mv,Z�E������r 5��Ř"��p���M.����0�خ���	:�T���օ�=�����LA�rEy�R`�J��&>@sz�
̗��m��W�?��Yx�朣��ao����|z�R��]�`������*��Q/�|��ej�]뵼������.x/�q�Q�}#zp�Os9��.-�W�I�p��8�R
Y+���qF��0�3����R=A(�QQr^�cM�6����*�Ge�����DC�t~f�j%0;�{5�snǄ�<�C�'�ҩQ+����c	 ��`D}
��9R��Z�o�*�R�П�l"���j�gb�yEkg<�a.,t-l�Y�u�U2v�j^�5�Q��Y���ZH��)�o� �eC!$��UM�;y��r1��?T�R��/TI�5^��V�&��1pq� ŹZ��L�~L ýg��d|饛/\xmA�(w�M�=� g�f.Eh`&6�9�TzV|�	d�+�D��~usN���X7u��������:Ũ��0��h.�zin�L�I�bW�6*������d�Yf7��N�i� �m�-4�sl7='�vw�R@�%�g�M���_D���Wg���N;�o|:�פy�	1�O��,u�TQ�+~.�֪*��t��,�*̢�(��z=�NŅ�OUK���؁�,toh�_�%:�u�#���+5j.W��RF���{��<�-��[������칻�o�H>	I�MZ6u�];ES^ �CI�t��h�'Y���'��ת{�c�����_���U>�����|�����%5Q��v��
ޗrwj`��7�{�����GH��0���ށT� q	X9�*u�x/q���]�}�����}9�s����O��cU�ӋMR�������}�������+W��} H%+��K$Q1&�\p �7��p�dЕ�+*T *Hr'�K����~p^f����DD�-���ᴨZ#�Q�pZ���ӥ�2QH�Ɯ�Ta���XBK�cBg�;zitH������^� դ�qAY���7��@9U1h$$�g�c�F�/�ްI Gݥ������g9��%!�T=�N�]�AC�w�i�F�b�������oZ�s������D(�^>T	岤�OEʛ�j��d�� ��<Ĥ ώ�WQB���E�ɢ��kP�.T��0��n"�����K_y9ܱ㠪��;o�Rڱ��e�ӿ�ݽ�-2�����_�F�#��w��u�z��{~H��r6.�n���N����k\�\:�F���!��+M�4l{ST'��(}&�M��g�v�=E6��g�ՠ�y���E_�PǶ_��4��h`�|��<Nƻ^� �Ev�F���{w/�
�����-`��9�{XS6q�� ���~4���X���~�u�j�ꅍ��½!���{iH�b�5�����R� ;u�Y������^x��%��%��
�T�#�GKWQrܖ�V�9V"���a���<T�S��g�/�D�1�b:�\�^0i]���՘JD�,,=(����R�DY��6X$��q52���:���Һ�h�}�*�<��-� d�Ik9'{/f�S���R��w0����9���9�K�S��,O�B6]��\�%JOK��&
(�8M���C�0 <�:  �l(��KY�#�_ʩ�ȵ|>�cO�S���S��{ytE.2Wri%Ey/~%��ͦrS�oLU~8�#������(p� 	jdm�أ���Kr��E�@�0�DU>�K�\�B�wH֌��� zh����PR��k�hVvG�YLUb8��&�\�2��
�����Q�4��@)V@�
@o��Ǆ��\�h&i^�����Mo����h��7�m�Eo6�T���z6��~�`�� �W��"�2�E����Nk��w�g�%;�KlmPl���H�{3�9��G��՞�xn�}�@P�8�]�J���J맨�|?>F�U����B�+����DY�����ٚ��dq�� B�X�ob�DuGڱw�������U^��Ӊ&�T Q����G)q�����E{��t�&?��+��Vi|<QmMl�����zT;�o�]|p�_[��뫕��o����b�|�K_
���o��xloW��R�aB��sE�-�������_�Rx�7EU��/~��ǿ}��$P��;.ꢗ�> Q�v���¶��џ��~�{{W�q����eg�H?a�	0�7���h�_����/\�gH=��u%���,��䘉Y�������i�
�t̟}v� ����Q>�Zk:��_�Vw-^LI������k�sA�{����ǵ5q�ہ#����w���(��ۚ��`�`0q���+�	�5�NL�����#�<E�7�A�͓�i���m=�ɹە|0�Vn�Xծ�E��TF�jIy	� �hyp��\����FB�I�-�ѕn޼e(���]�Ox0�1q�Ų�Z����'^cБQ��`49�q�����?�)��&6�A���}�z��/��˲�I:�UE#�!<+�R�M7�o�zTFN����}�o�W�f�Jm�a���)��ߵ]M�2��V}=d�WKѫ��9�E����c��5�jwbkw��l�����иr���.?ב��� |Q�!��r_�\�Դ��:�:��9��lM���{�Qա�x�R�D�J�#�1A:�ȃ�K���}`{8W��GVvq� �R@�}X{t���.S������QԗB�C�L������3?��ᕱ�,�� ��@d<E�Ʃ] _dL�c�l̫�{t7�<pY�K�Y{�A(eRfRv1�C�<�A@�*U�����.�m�@�����9 u.A�}�V���!�r��ʮ+�($\ !H�u�7����5Ҽ#�SP�
�iVq�<Ɠ�"��ݓX��B�$�����}�2X��c~�q{:](�U!�N���p�R�9D�v�/�/4��mEO@�h,�G/>5��ضe5����q���$�wT��q�����U��d(Z�o�\&�P� t��'B	���B�fqEJ7X��k2���=�9�� }.������l��仠��Uu�룤��C�� �����k�QN+�[�]����ǵ�pb 屝K�1\*�E�f����F��q�nf��Աs3޷���O$�����BO�Uբ�.^���%��~$���9*����n���nMM�����O|K�[H��v��ߗ�\~O��vZΒ�e���(X�����4�6�Pz0+r�ڶ�&���}������v;�v�zJ.m��(�%C��OuLK�W{51y�M1�(�*3А@��t,��^��񄨗�qA�Yr6ｧ[c@�Ğ��,l����W]*�Jo�Mհ�꾎^��&�����x�U�������b��-��-���{*[	DG�&���Mݗ���=DM�4m�ۗ2��Oq���m�쳛�k�B\�_�j��׿��J��uZZ|4?L��ˁ����^�L�̲y�����~'<��di���]�Ձ�W��+��NU�IU  � ���(�Ogs�x�E��}��\��~�@%�Oo�)����� �"�?d�{Z�T�@�=���VU�E��LNO��H~��ň7���J���y{1,�Y�'q9�Σ�C�������W�(�U�5]*<pa����T���H��NȨ��<>��i�l��'Y�6Or�cC*/fo~��[��
?��O��|]�_j����(���������@z,�TP#�;]E��t)�ut�E5�qXE+O�y5������mx�?�Q闿|���s�sw��gT�Z��gn�IUb�.�����~&�K�2<�|ꩧ�>��H���+��&�&@
�:���\�dտ�<�v���-\{'�-`Zj\���*�y����?�>l����߲{&�{&�^���u�0N6=0�/s�u�>��2�Cr�Y�l��6�G�w!-P�����#Ҙ��)\������h):���A��*��N�����GR���4�Ƀ.�s���r7��u������0����A�Ï>�z������M�_ +m�G	X^�=�:��tN��an�B� ��V�Pt���:W��FAA�2K^��$�{6W�2��Ξ�i@l���ӳ�}v�#��|B���Z}4v퐂e��Qҁ+#2��>���S�"�2���̲��R�K�eh��3=?�Q�.�E�Mڹ��ߔa'<7aB���%�t��QقW{"- 3��k�2��3<��H-�*P�RG㍩NW��p�3��7��qx����V�����Z�6��`V��<�5T$���?r���d�C���8B"8�*3���G�i5��@m��I���<�4���_,�H���bcC��WN�{���rR��Uw�g�[F���Ur�-c�S����q�iC��!��K�շBP`��(��`>���1�i��̺|tV��jX���׮J<�c��ї蝁R�{�=cT���*	�po��Rg� �Xv~P�v������2� ��떫���u��x�v�rQ��p���H;i׹%���]��щZA�'�~"�m����6b@����@m�.��J��]4� �+BZ;�/钒��\�=V��3&�$s�HL�9�����Ŀ�DY9�i6޼��7�H}(i_҇��F�Q�t�����8��ƽ*���Wk���ƕ<;�1䙏�����1�>hT=l�.�!�[�<��)�o�C�7۠��g�S��d�R�7l&Ss|j�F�m+wJ�G���}��Ұ'jF�|��ո�.�g�^��<�[���?I*/�$>�{����7/z����������ޥ����)zR��3�b�/����8��#~����5�X�X
#j��R$��q$�/�g
���3��m�`Q1I"?|/ d��2@k��7�qx�=�j��T�^�!���l�}�|�	US�~��򄣇�\���������ӛ��O?������`� pG�Bk=���t5��g6�޵��شt~|(BD��}G�W��u�W�E7��D�\��U<')9oG8О���R���d��ޠ3ހ!%)�1r���#�����P���|�P��C�o��,�&�XU1���'�AA �.��6�*NM�쌌e��l�Ȗ=��ᥗ�V9�'�,|fۧ���� ��.P2��������s��34~3h�y��Y�3UJ>��ƀ�0h6�� L�Ȯ���������t鲁�υ����Yh�_��_$�� ��R������̛�e�����>�ca�\n�n��C����q��÷�T}h��v;�m\b�K.�!C?�%�^QJX`�B��-�i��ie��ƭlK��g�d�vj�v4��q�#dj�0����{�T}�ui��j���4'ʛ�� 5�ٍb�"�b��g�K��B������4���ۤ��($7;R���y�p�˹�ߵ|�%^�� �Ȏ�w�!*(Yt�-��'�C��Nm��L��&8�dЀ�L� Q�g�v��B@"���3�w�^��������-�n/U���{37�x/�R���i�|4�h����Y�07R��$��@�h�N�J6�
�W�B�*����ιMy�����e��6���R����J}P8����k������=D�̽����������Zwc��5F�nΣ$�>��X�+�?���N��[}f	t�\&եLT=ͫ���봜-����+~���Ʈ�Z_H�:,���^�$ͬ ϵ�"��D�uc�o|��/�H�m<� ��c>�&u�s{μ�p\ŋ�r{�@�m��;6 �g S��K�A���ӹJ�P� W��S�0�D��Cx����SU����/Ot�10��᰹��-��}ݟ���4�ً���Zm�Q�L�� >؆���:��A�P+���B�˘�>���HAj��Q�7õ�f��r�݌�M"�-�*����	)۷=�&��G@��Mo�l��v)r�c��-�qΎ
2JpǍp��--��:�G���ᬻ;z�A�h��t/l�����~q�c<����J�N$vE�xۻ��[y�������@���J��dY���.RҊ�/`��,�6
���,&��t�C������i���3k����Ыxx��{)��3�b�����*f�Q3�q�J�e<H��v���NU��د:�h���,B�Y�a�B��N��A))M�?��c�	cr�8��{����R�X��*��>;QtIB?�(6ǚф�U��>6}�e�~^ )��sz�N�������G�8����G�b^��B�}ޫ-�%"�:� @�kD��
� ��_���x������U=�I����ѝ����?����x0�h�����S�6O�[L3�'�|�+M�H\�K>�vӠ��;v��al�,m��k�aqePM�;���6�$�g��^R�Z,�md{
�����l�ޤ����B��n�l\���$N��=����nK4� (��g��2�{��5��&�h���5���^���ɑ8xTn��TH�iQW[�@�2�MdPiTbp �F��z݂<7�{Z��jҲ�q�QU` Q#�����a0�� J���{ﾫ�v��^x�y9���������(�Q���O~�ޒӓ5��v&{R��Tݍ�T4����NRn���_�J��c�ђ}�Q�������{W�w���G7�w $)��K1*,d" �dgh�,=8e��镕���7	�e��=�i����DJ8M�:�����8�r�o��<�4�
XJ�g��c�[$�Z|׶͹��6iL�UIβ��޹�^ڱ`�ڽyV��0;>
?���xX��և���z����i�ۻ|IT��*xF���Lw:�p�M�d5QRT6��R�Ƚ�X*Dn���-?��S�p?�]R�"��ق�W��9���phbvo1��5=��w�NY+�
23e�q�\
T��֗�+�dU�ѣ(iuT�0����
���b*���LX[p�-�����"5Urma�����X�a�=3e ��=8gC�b�U�D�Hr6�Vy���閄\H����j�B�f���s�\�������Ds�lq�Y�9�< ���N�B��Ξ��9�L�Ñ�+���Y��
\�W��S}����]7N4Y,0��iM��QO}�Du����S���*��E(m��dzX��05p8��^(�{) 'LU�B��yn����@��=��'j�zp����z��}4 ��ȣ�_�\&�M8���ݎ�]���W��-�ǀw�8�P����B���6�/� P����2�\��~{���<�c"��g4���*�m�c�s7?vT�^�6N���<�n���Ҽ���qo��@�<A#k����V�#����s��8T-�I���MonocP�C����,l�u���5��Vl?Z����;��*ʬug�Ӓ��tAz���N�_���Q'��q����a{`�S3;sCQ{�<�`�QU��C<�����L�[uHN�>]�E=����r3�Y$h-�#�������C���ɷn�T��S��bm��?���i�f��b�H�NM�`4���Z��=Q�6��_xl���g��2��c��#�xx�U� ��]+��C�n�t��/)wWx�����W�i��K���qpI���pHLs��ZQMBƘ���	�b������9�uH���'\�����I������68�S?�k�]�s�}A��s���K��X/�,&=�sA�c�?����lW���Q�#F&�`kWTT����鴘7��b B� ���sH��I-d�Q!�4l)?>i�Qt1�:a��l>Upp�V4�L�LMj,��6.�O����MnBuv��J�-�S3ͳ϶&�r{<9ֱ�T�]���_������B��>�����qzV� �(���?x_����Me�28@���Bsb?���o�/�E}��GċS�P�)�����sb�2�Mb H:��Pa��5�R�i4�r������UeL����W��`};����B��3����Oj�'�$��"�4�m1��wl>u���~�����U��O��������9�s���xh�x�Iժ��j���%�h�`��{���-�$P[�xU��8?��J{Tn�����\�=����@ʞJҮ��!4]x����k5l�UV�W-,��	��{n�_&����x�`A��d����~d�b�� \��4�j7��;� I8=?UO�t Mk;��4Q�w��TJ��2YPqH>��u:�x����c�^�5+��?s����b��^�����B���$��=$���\c�J	��ӽ_�=TΣ��l���@�Â���i�"c?SPD���wV�\�i�1*`
��=$���l��m��̮��iz٠s�� ��/F��������ī�=y~��f �o7�,��4��V��1�YB8�sl��4,��B�N�s�9�Sn#O�	c���Pj���@HϜ�QGd�\�8; hGN�\�T*U/2�#ȥ�-����j�/��ܞ'R���0Gό��f��2H1�1؉">��%4�A����3]�X6u�2U솹3��`_�6$ 3ëWB5��8��chB/��+��$�jr�7�&7��la��c��s]Icg��ڶYKb?��-��*2.g���~=[�ɥ��������@f�n0�C��\��{U�����4ԡ���3P��{�m��q=��F[�����\TN�徝
�R\5��b�/�(:j���~0����ڰ2K�1�mB�6���<��L8-�w�Q%3
0�O%�P���+i�=�"Q���;
?��ʒ�7 ��	[���W&� �A�6��'�v'<�[��t�Cׯ���Y���=���sZ`b��㵧���u�$���W��bxT���������߷�����-�yTՏ���'�
TC��b D ��b��&�<Y{=� Ah��kU�ʼ�v��WY�sأ���[��Ar�����n�_���\?��d����g�)�5�ݗt�uo1�Лi���L1$N�j4��~��{��lʕ�[��I.��D*J�������Sq�5�ޣ�#�k�퀘75��cj��ňJ����RRxՆ��j֋/���z��ǔ@�ة��d?��	M��g������+jܳU�m�m��N��
�����jIJM�T��!db;	͈����g"��~�(�(�Ѓ+�:��Y�{;����R�ք���к[�����e���d�8�{wQ��,�\&5éG��9YGԕ�������/��.��5�b�����5�p!(u�P�IgI��O�@�z��s�=o���۠i��$��5���c�'9��>���z�`���w������7��y%����'�'���g>/�_���[
�������믿ᮙPh��D\ܗ�#C0��B���+������׿���o�/����Y�U��k���ޕ��6���S�&���>�݀s5�����y̢���ٍI�oDX��<4��"K�oa�=3�pZ^-�+>��:��ĥ���[^�,�@U��RB�lq*IP��< �B>in͈��+6Nw����G�����J;�v]�D�X2���4��+�b��E�7�UņI��N������X�I�$���T;�Q�

�Y�`l���&EϦW��Sc(���),d2�+j�vkeɧv�P���PJ/<��`߇bq��.�(\_�țg��"Ӽ��3�o�/;�%�)����	[Q����]Ϗ�6wM¹��v�G�g\�k;�Ӑݱ ��" �T�i�kIU���R��	��k��(�U�.�e�B�>���Qu�)���(��D��csɝO>
G_7P���7�RiSb�)� V\�_�vmW6gGg���Y��|?� �v헢��Z@ѫJ�~c,�zW9�kc�~�`�٘
�B.�IUEM�(��ga��\{���c�F��+/��f�i�T����n��RE��V�ef�E�"����U
@��� �X��:d�j`i�cb@� ���R�����⣃	�^%��#>��4GN��Sh݇��C��vh���ٙ=�u\;�B�"��sD� ��l�L&�	�E�j5��Y�����.o���&����"��lddyk�ִՃ�gi{)�I�i��~4)�"U��񋛭�=N��Jݨ��i
�N�&��_)	Y�|�זv�T,k�����n���H�S�Jޫ���RN����������sמ!����*.N��wm�Al.%:m�'3���V�,���x�m�#�o4yW�����iNᑜ��F)��N�&q�(/�^���O���(ԑ�R�����2�T=����%��L+I$��Rh�����E�I�IT��J.�;��a4־�q]�Q+�QU������_�x��+���~���O��\��Ï�x�JO\L��]엫�[�\�$\��?:�D�������7�xC.�H����/J�����Z��LTi��Q  p�O7n� �\i�u����
�#��y}���q@d_�
P���VL�q�m` ���Zqm��>`�]���ǟxB�'��%��/$��� ������,����dw�J��o�:V+o2?��S2�(��2X&⻹Q]�=�n��Mj	�NL��u�4�^0hB��p�G�b$`�*U#��tS���s9]��(��psd�$����s#(*.o�\��X�� ��k�e�F�,�8�J�=N;����>����QeķU�K�Eos&��h�$�PY����d��ܹ�J�TU�*}��Q֥�s��#^����c�L�Z�ӯ���nr�ud��x�ܽ����rn~�� 
`�ca��s���h8n�e���f����o��	��n��n\)3�T���6��hԎ�غ�[@�_z�m��Q�u�����@��\�7<_ ;YqI��~>����F��7�;�����g��������a.jS�d���}0��&��v�g��+�c9����HZv��w�P�8;=v�<�ם�K��;�K�*�M����J>���8��d�e풽#�	��B
O0��X�� �bMH��XP��YZ��3zP�F|������1ƶo����ԅ��)�����ɑ��L���&X���N��@��d�nsy>�3 Ҁ�um ��Eayn,�ǫ�eX�=�V�����%�u�y#��|��tU��#F�!RZ���?@�j>h�hi(i� 	�t�4�hWUY�w1�Ͻ��e5@(�Y��^�0ל}�>{c	!t��H\�7�v
6���N��  ��~�^�f�7,f�۰�����α���g����!�x���y���t��]��{F3���+Հm�˖ۺ�t��2-��zm�R�2����B
�hx�Z���H:-�ڸ᧔i���H��#%�7 ���.�[�|]��1M/���ЀAq�4��K�
Ԡ�P��zD��������pl�+���9�[5���_"\f�ti�ծѮk=��]i�:X�d^�/fM�G�N���C'�H6�7��_,���� ��꽲q�)g�'�{V���>4��:%W�ԨW>etҢ�B�D��E�Zc��� �.��^�*%�<H��p��x�ao�J�w�qy���$�s_ش��y�?W���AF�5F�i�O��dO���)�O?�Q=&���0u]���ګ�_"IgYg\ԑ>̧V1����s
�3y��~�yB D��X�'d��%m��$G���E��io�Ⳋ�xq��1�9�	>����6���&�o֙7t�ֻ��M�E��3],�Zt?ܳo����~����,{'*�5U���J���z�ǊUS��Bb�ľ�X�j���\p'�L�V���)�M�#�E�{���{�}`���o32�u�S9T#��8���E^(YA�R����* (\<`@¿���2@��$�H`�G����7��ě  	���Y�m���C��DҾP�aa�> ��7��M}�i�'���$ZC��7�!�p�pt%+�?��U�0��eTZ����8���\xV|sS:�<��i�/%%[G#��'cU ��.4�%�\������`��|ZdT]��K7ńXiٶ��ěk���ޠM_� �	�����z]j�̜g�l�D�y��ǟ���������6����\jwMʨ4�����x��_��A(�HI��|(QN�*T�p�{��H�טg����f�� S�'�->�DJ_@P�P t��l�g@I�kB��	��ޓ�y.����kr8jr>�)6���3��;��}U����s��Orƻ�ΝӬ�!�-i
�W��\᪔����[.l��*��H�jt�[��f�g��W|��Z^����������#zd�����9P�k���3PR6��P�?�[�,V^��{U��c[	����ˉ8�׷���y �?�1}����8X<G�
��vM�J�	�ٱ�"Ķ>�� Pd���>� ��RG�p���z����C���jX���p��* �^�B J	�kw�^��del�~9�Fe/���	=�l�Y�ݡ9����8ͦe�4���������U����k2��)*Q�h(��ٽ>�C�c �X�+���\� +xs*/Ь��u�K�X�I@;����l�c��Z�����$�Y@�m�S$� ��p+lN�a`�?��j�lq;G�a��8,ʾ�@ho<�h'����&���d2�/.���e8|pO���F��ez  �p!���τ<������K�&� ��~��xUa�|�S��T�T!��<+nֈ|%p���0oe@�t��CI�b ��T^i�|�q���2@�#y�Z��V�f��kz��b�p-�*����1C��ۑ$q.k6�5~=6�7c��j��}t�ј�m�CW�6,72z,xOm�~�ޘ9�/���3��8�IdE�}1���#�,Y�h.�v����TƱ�{K�R��*�Q�k�թ򦠹#(��5�⎂�:��J�n��5�W(��|��fu��:EH=Y�thQ*��GX�>3�;���ګ�v��)Ξۉ����Б�1]��;w�î���`\T��Q�5+�Ws��z����jr�L~4�̽��<�+�u<h/����Zw�v%^U��L�qm�%$�R�>=���*=���W���ߦ+�ޗ�[�F�̕�ҿ=Џ��8��U�J�1�	�{�����b2�����[��%q+UF  EU4c�z�n���(��(_�ASE��9���}%��?�����t-���g%�'�����[������U�\���U���I��{}u�ĸğ$���~�[�ߵ��D-��u 
Ig�*�:�G� �&��'�'���|�M1a����K�@����v��7��x��'��Pq�g�؏*���vc&>k��� �
��?~I����i\I�}�*y{t�a����D�빇J�G�@�O\mh��<�00$C`���S��
PoEey��@]2l�5�d�%��j��SƮQ��7���M��]._�����6o��h2�q��f"��Ƈ��u��/~m��$��HU�f��9�M	�r�,\p��p���l�����2���B��<y��h����"��5������k��9P�Bct�)4�p���+�K�	�a"i���w�}o���|��Ņ��b1� b�s,��x�j����l�=蛆J�T����d�~>q��$�x�w��e)��h�J�1�U��P�m-�[E܀"�w簏����7?w�粩d��}aQ,3ɛ�iAʆ��R�Hl��\Y�J�5a0G02R�C�\[`�T#s�ۄ�|.��ã)w�~�ۛ���K>�'=pL)iH�mQ�����z���=2�H����l#K��@��`���L�F��8�d���2��؊~f�/�'a��y����}�0���0��$���&*�`SX(�ugi��V��];R߷W��_ҽ�)n�d�`�} ӍYD�$��ǩ�d�f��E�& �mx�����x��b��Js.~�=$R�2PC��X Q�p4������${��ϩ6��Q�GEn`E�s�/�J��]J3Tn�פ�C̩a��ei��ƀ&�=Tk�@4��Z�_o���F-��QVN�b��]^�#����9��g-$il#��`�
��F#OT�P/�\3!m n�4�g�^/�A+�
��,����f���i���v�������R��_��C�R�v�ޅ�$=u���ݥ��:b��>��亟$���k�8�}�T��1	XF66qa�����Z ����F�Z��H!�;��>W�w|1��X��08�E#�JE�Աl��s�e�ٳ*�����
��zjoP�ޠ�YeB�l�z����=���gAG[�0������d�x#��L���(/R�N��) �����5�k���e�Z{����q���>�E_����7hS��e���X�(�J�nh9U��y�w��{����{�G�h�v"�'���0���x�1��#��1�����^I�V$7��ɰf��%Ë�Hg��g�W��8��TS�R�LV�^i���EӜ��;��E��-�;USAj+�cա���_�(`��B<��:�m�`�'SO�*k:�U
X��A{��MM�.��<� ;:U
~yfe����_n��ph�Tͻ���a���U|A��f��q�0`� >���n%�;�����ϊ-y-15�# ��H�"�ֽ���/�B���&�@r0=�(�+��3���xX��I ������e���%�{a?�ӟ	؈Jm��>�㨾�x���k��Ȼ���E�s�`\���O�Q�;2&z�N��J�<�iROՐ��AM�;��ϰQC��w��]�#2�R�I���/XJ-ut�ln_p��8��7!�]]@���S*@�I��?��1[r7p����Ws�]}l@������p��B��|���f�T�a�p�b����#�ڸ~JM��D)尛kAF�n���O�iR-Ay���s{OG4�DKΐIVn?2�I�%�T�

��$R� eUe6�IS#Q�{�a��TV�w	�e��q�(����A��t��	�M���Q�&s�5Y��W��b~�n����K|�-�����+ю܌���/�T�:^��M�>c������ŉ)ۨ`"D�I��h�Sq7ޞ�ht�f]Q�ҦXG�E\��?}�P {����6ś�X��W��0b��� �an������ɩzL^>���i��xΖaxl�7P/�,N�D�˨�Y��7��C��(W��'JB�	K6����S�U�.4VS%A�t�[�޳�D(Wm�5��fb�p����\��"8
���l^�^\��㥚� E�Q�=�KK��}�!< ��5���'���d.>�,�4^3oc�ZO���@�(����Z,�!,fvb#�g�0[{ŨpjZF�Iet[�_wZضn�4�=8�w���ݘ,�n4H@d��'M����=筭;+����8R!����T?��C���=,iD'��f�A��8���8�Y~k'2^��qu���*�2�R#�`�W�I��9/E�� :P���Y�jU?*{���A �t{kgkkEic�@�ޑ� �wckd�vt��$���Q�M��y\a��!�f�iWd֗���bl�uc�'�z�x�HT0��^/��v^#�e��_���2�X[��AO������D�	�ԛGo�*.��y#�|�6�w�� �JX<c e�@�j��軬���[�5�r�m�|�� C�TC����ʾh~�u�Uj�N��&_���E
�]�4���,t��ѿGAu恻��c湔�rݷ):e�(b5_T�D�s��,% y4't�L���W������T��B���~��W��n1i\@�/�zL�t/c�Ɨ�{���C+S��C+���ELp��
�F}U��e�]r]=O��Z�A�Z�ҫ.R���W>��,�u�L#I[�d+)VG*RݖAkv��g�4R�yz���{#w��7�k��` �8T�����'��RM�ۋ���ʓx�M�ý�U����*��Y;{{u�3S��U�J�/�R�q,I]�TA��9���'���s������>n��կ)F�/j�1�$�O��Nw�Km-v�R��E�#�J�PIX(�9�꙼�w�������O>�9"��zq�Ď9=E����vx���u^w��$�{�5"t���b���T��å�MC9�i*)��JX�^^q1��i��c��{"|q�Ѭ���^{��B��+�h2�R��� n��Nz4�n#���y-7&4a�������A�T�·��w��(|�ɧ�$�,�ø�A�WP�_z�k���@�4�)�4E)-�0'��l����QPA���&eRab!W憃u�����	�jd=��d���q�R֦n����OJZ�d�݊��_�J�ɓ�R�2�N�PP����]��[����b/�sz��@·c0��YD����gj&�;ca[V{��������ql�"�a\����^�����R�F�� ��$ט8�Y�p�.���zǽ���{E �-�=c�h��s£�[�΋o�n(�R�k�$��*;ae���(˕�4�<n�茎�Ue.�݄�l�����ah ���Y�<��
����y8���G'�@ �	��֏>\�ej��A�ο��� ������W�2dq�L!�M�]���u�-��Z�r��jJ�܀nH�]��l^I���l���+ow��@��vfW7)h�d�T!���G�U����K�c�nl�|zm���p��ǶP�����ĳ��H�P�JWn�a��Φ�[�R4�R���z��d"��m���M�x8�v^�~W���B�z��;�)PD�wy�OavM��,��N��I�sq�}�+�aXyU�����6�>�ӳ�hs����
�*�	9W�m���|-�ߺ2�Z�@ B}uW�;�5I �p���\���%(�gh]�q���(��8�o�)B����!W���ԓS���SE_�m� ��|T��"_��J�֦O$DP"z-��P�d�ٗ�^�׺�}���A�B�"�BF�T��e�=X&��ޘR6��FR��$��Y����0�֠0VJ��e�J9￀�7W�o�") �B,�$M�2
Y�څ�U��.�L�����k����P,�ޣ�U�Eյ\A{J��1���
U3j�"V=���gP$*�:6��Ž]g�J;�)"��5ލ��/7<��6��;�[ɉ̓kUj]q��f[�S���K{��iXn�9R�����s�s�U�d֭��u��U-WB3��U*�-Ժ:
��JG�|��枒�I�;��:j.F��^�:�ْ�ʒ���DZ�i/�@ ����(�h{�����A��\ (��?s��t�i���Վ�Du�ݴ�c��^ؒk�%���³�$�Zɠ���^�*�ۜw�G���}���3�����=+��ÇX����}�=�'O���w��<6�a{)R����̘�ƪ��zw������V���o|]tz����`I�J}�|�PF��^e΋&����/>�@���E�#�zH�#�����W_���1��ٓ�����/�"G�J��������vL��?�J
�#����oG��ң�+���I�:�E pʸ�� ��N��QSމ�%�7�i8�QV��l���+�ͳvʑ;xo4.�X|+(��מ(�����P�n���Yz`)}�oL
k~����ρk;���(|��ߐT���{�b�@�_�R��7���$���"�0�Ѱ��O*T�ޗ���5��],��}�ߐ���/�W����pyy!$��
�	A�������&�W 6���J���T����H@�����1���;�Ǐi@'�?J�4�Hp=C��87�� �P�7C�gy7���%�s�T'�C���	����!��tw��(rD5��4�{�P.�v��ci6[�{:Y����Ů#��w�&-�K�v�{���T�mU?�&J�n����m$(Z!��]'뉛���Z���~�jL�����Oi�z\���n%
��{Ð��ٸ���t���VB	��a^i�����@t�sa�
���p�a����ff���n����ri�tH}.��lQ>Uy�t�Y����\7	W�.�\��fh��)�8�x$�{A
[h��@72�2hD�ۓ�Q��*�qF��v&�y8;y��G��Iy�ŸƉ:rpʇ�����Tٱ�Q�D��.',��=�Ix��G�/���l�� l�=(� @ pd���`��r1�{6�{f��8��
��@���|xo�M�DLL���w�I�����"f��G�ӵ��6�=���������j�YV
�=��j4�e�l:a:e=^���z+&����\�{�N�"�cl���e�\��zk�7	|L��v�;�Bf�=���e[�����W�@�ʀ�1(� ����A�s��U�y���;ԃ�"��2l�y/onE��j|R���/m�[��3%;���k5�� �He��Grp0�&��_~4��A蟜��L�zN&�H��&t��SӢψ�Xg0�`��dϿ[z�����ĚM�: T�r5	+Q{�"mly\{�����������)R/F�x�xI4�:UZ�ڸ�*��M�!*�%�}�$���I_��c �zL�d�i?7��ˬ)��5rWN�U�p��5��%���Z��Qfz��Ɏ����c��� �B��Z�"`֩����̔�Cq��*"
��^���y��+��j��zSRU@��$�x�:���_Vt)X���P[#����R�2����E������m��D�c%L?#}3F�;X�nl��Q;�o|���w�w�+hguY7�X eT��\+A7�C��c���e�XK �i�-0v��K9��~��f�{����UA��C d6+7O�?b�������^���W���@G�jIh���&���r4�s.�wH��b�^��gF��E�,���ĀH�ȼ���^'� �2~��)�w��:�D�rۇ"�˾*+�0"��ŀ����( ��|qs�cn-��9b������������<�A��8:v+Z3R��:T�����c	!�E��o?�����m�,�q�X�˧�i���MZ$�a����*��=N�o���鮝��pT��[8�4��<��"[͆B�픋���:�����AH&�7���4=����I)��!�V	(��}��=`ʣ|$�����?����o{��7`h0As���>
��wR;x��7�[6�P<�)<ձ���e����g����G?���L�w2��5�&��C���
���q���S���/~>��3e��|��&�c���7Q�������_�u�������<�6�L�)���
�ᓟ���� ��O����;Η��nx�o�jr��z#\�bv!��~����9Q��},>K)��"�X���@)+^�<�ޠi��6Ѽ��e)+U'�u��v�+�oS����tr��U�<~(p>��܂�"?(�X];gUM�Y̦�}c�7�Jx@e �!�{u}��w\��!��S�K�';�8ç����Q��CA��q�az�
k-%�����Y�37T^�%��9��lݝ���8���v�� I�w��ʮ��!��88?	��Q�@wY{#-��6��RYj���Ɗgg�t<S˽�cJ����H�@|4�ۑ��a��O���q0PT�������cߓ˫pb -W(l���M�׺��-�hE�B���۫0�ܳ��D�"8�F�:멹�=L�x�l��uX*(�Y�R�7\^�p{Qx������L��q��Z�������<�^M���� ^T�QIX#����%[Z�0�I����c��~f&��P-msu8�hW!�����kAp�
���]�:���SYЍ:���y[#+[�[���F�jc�~[���Iu����,L.����e8{p/��_�8ZG�H��R�*A`�9���l3�O�Ѩ�^�lM��*��;���mh�w�����J��ڞ������e�{�:�Eh;��"���G�!��ɚ�W�g��>�_�I����8��d,�w���I��ѵ�QE_G�I��G�І�i7ݭ��A��P�R�z��O+D�d�k�E�b�Q��FK���:.����Q𮀤t�Kڟ�V�y�TT���V�N�ٓU��76_#���2�l�e1�@=I��g)�.�^�m��)"�f��TΠ��71��{K ����|o����U��B�Ǎ��D�<�ڕ�C�.�v}�K�S(�C'w1��{{�[U����}m@��V03&i�:���1L�:�;	4Ɏ��F�Ǉ@졨�`�� ��@|��c��z�@���91X��X��xiu���t|n�\R����ڀ�,�7r��8�$��Z�]b���@�%��{��W�^u�k���y6�B��D%/�wI���)b9����Ol�t�8��#��<Q2�����X�6E��F
_4ύ�+g�8�3Q�`�����Rx݀����t-U_�߽O���?#�m}��� 2˶��x��7�|� Ϋ������ ��u�&��������>�L6P՞>�<�������;IE ��8e�D;k��rٸ�\�s]R�p�B����le*_$8��ѷ�#�,^.LC5K$�.k&K��fX�8+���#����c��<e�7^]h��Q�3ӗ��e	X��>y&�6�/������@nn�5����&��R��`�gpO/�����?��RƦ���E#c��&�͖������`��38�ց@H��ַ�yWL���D95�&ӱ,�2�y^����l������]�g�{/I�e@��c�O�o�����@�8�My݁O�lha��]�*�y�C�&_XjbT�J,H� l>]۽��׃x�/��۬n����c���^���wQ��y�O1���F��$P9խ�m�t��v��e�����s���t1�#=,��Q��q��<��"s5�czf�}a�����d:�c5��x�J*�:�`/ts��� �݇硶@��J%� S�����ņR(y�/(Bwh�m���o�l
������/����L�*P�Ni��a8��G����؉=ǵSv$��_�Md�Q�J��mqz��!����sD�%h��N,��׏b&�+#ĩ��M�3(r(��R��l,��pi�m2�������I���v�]�8���(䞤=�+U?�Z�������fʶ:��C0��ݮW�}T� �^Š�G\QSpQ��4�/Q�+g��܋UY����͡�[(���,��"l����rkkܡ�<��o9�{����z�����K��<HQ�E����P�"�����(Im�Y��k��@ Թ��Q�DU�>������0��x���5�,T�� ���a��z</�62}@��?8��$�P��Hv:eC�����9��j�<<�w$���xg��K�HI-�8�n�E�%�=:+��<���C��&�K��j���=P�HU�.ʸ���h?,�]�*_�b{Ĕ�țo�7������U�[7�5-��t_�3y?l�g�����<<�R��z?"��%GHfW]Hfp�[��r���J���m��w����]�
���"ѷR.<���zIw�����U�o�.��ip	�=/#5�q �G䐫���T�S�)8u��a��DK��Q��6�|�l�U��_��ԛ����b�t_^ܛvw7b�z@��p�A/m�l~�]�,evZY3n���8Q��(�J�7�L���4q_Q�k D�ݶ�0�^����x�^ی�8�ӘOt@�ZJ��b�!!!3X�����د��w��,5<}�e۴)���Ha*��b�]��+%�Q8ϒ�Xzv�@�:*-�+cu��	�*�}�R�?Ϛj=&T���U�������^�*���J�� "��{���ԫ+?���~f ��Թ���*��֛W��ĪIJ���Z;b� ^�ya�`���hY�e���Tb�|��O�/�T0�
Jt�T�\���E��NeRe\b?��V;�{�k�$���7�2���\q.e���f��L@��	wY��!4�;o������ ��㲺N(����K���XܬO~�Ix~q������{e���2��}�:��Ʋ��{��Z��{��:���c���pa�`�9�O���֔GS.�՗�\�&��?1��A�A�P�Ӂ2��9�O�Q5A
��(�ҥJ@P���Z��wz��?�>.o��F��ޏ���C5�pؖ1U�MháWK�T*�
Kw��	�^�K�4�K�K�F�'  ��IDAT� �z����9��0�i�k�M��n�����mjU��{�@T�����l^�|���W�࣠AѰ=RX�<H�#�����7'�y*خ��[�:���	�������܉Fj6�����꣗EI9��O~��}m�����C�:�f���r�+(r(;���i�N�ftrl�6V����;���xZo$;U���"����B���ųp�֗Bqе��z>���� I ��=��Sm����m(��J2_�`��*�BUj��F�UPI�0Egʼ�N�y�0�ml��kQ�N'�,��i�v�P�h�Ga�����W�,�O�ؽ2tg����'7�_x�S�^be�R�q)�:+��b��&}���n"�c�>
��-��7+�hԅ�����Z�P򷥂y��9U[k9�OH�Z���J��2���<�\��O��Ê����'{��ۡ��A{@<��w��;;綱���*����Y����d}�Lq#_�E\-��񞥀�bn�UԒ=^
|��Æ�2�T����puq�������r{�Q*�L2��-���EI��8����IT�� �14�
!��
ic������ 8� �a��`h�ڞI����������=!��#UغR{��ݷg*�L{�k%c�rv�y��2>�;�{�N�R�#����FTQE�L�=c��{LR�D��{q-K�[���-�X�<�5w�.���j���f{�=6��z�G��x��%U-��t/���w$p�G��:&���ގ_����Ip�����;�)�(�X��E' ��Y����j���~��J"/){����}"�s�c����Q�:�Wlxl��ƿ����$�7|���u����7!5��) �债I����ھOI��7�"�I+�[	�H��"�_���]��iԉv?L�+���Q]	IW����	���V���k�b|Ў� ?]�N"8%�%Z�
�	dထ��]4�kw�;U3"� �K��})#HU8������Е�V�7�QU	�8 T쎽���>�'-+U>R:Ju�����$ZW��`�i# ��2%P�ͱ��9�D�o4�W���F	n�Rġ �?��������*�oq�vզ4��B�k��i���rTQ ����(�O�� ��
����t�{	��O6S%��!Մ�(���E���ꤖ�p�\�4䨟�s�|�E�B@Q�P��Ž�Wؕ�v2pq��}�����E�?���f�#�x�th��ԝ>x#}�d����!�K�����1y����^��EK��!�w�5x&,�	@����=P�3 C� Cܷ�r.���RY��µ>|������ >x��	���)��c>0 g�2���$���ɿYL�(eǱ�fQ)��Ȟ�����o���?������,f��|(����oy�w*��k�{?o���ݼo2!I�����҂��>?ӱ;�m�<�fmo���_D���W�U��-���&bU:�j6��:C�{�p�M����"�+s.��-B�B1�	�, � �L1�Y�Q�Z��B ӇF��������G�w4
�d�i�XZPԳ ������ϔ8E�t1�ʃ�,�%|����H2��d��z�v~���E�f����ͩ�&L�<��|y+��n��������g�qa��>�
���,ج�2_%8 玑[��f����04�0�clʅ�M��kH���3e�fp�*[!j�Z�xu�\����s�$�Z������վ��%�����Z\=�	�y�߷��t�C]��8�7��mW���<�hU��'�����KAl$@׆�R����4��\Fx���hlm�NE��E�Ă��|nn&R�b3�J�\DQ �������t���E��>|b`l6;�	*}3;��ݫ��[�RC!It{i���@�e������)�����t.Un3����]Wekѭ�50��p1�-���e�,�:�O��&�����7�@s		�DK��`&�7u�"��fܷ������i����S����(�6>Uu�SU"zv�:��h���t�83��:1�;����Y�h��:%R�|ݤ�����R��h@�R٭Tq[�3��%�-}1N
��i/�dQ��jI;�@�����@)�k�Xeѯ�J&����8x��ک"I�/Ĭ~�I�i��i��Q?���%���j]�<4&wM�*�%�����W����Pš�)_%�$��*�q�w��g�Ck����n�
Zjb����^�l|�����}�� ���-�C�y��,Z	�2R�v�*����z���?_M��b��M�{��h�X�3�?j�Ox�}Ӄ��`!��W�4�|�#�$4ae�ļ;^#�!�1"PΛ�A���6�v'��<���1P%Jb؍��TZm��m5�PNϳn����W�1��>L���ϩ<��2�*Id��QD琀]|n	HJ�9�;U<��&ީ"iW)�] �S�V�Ѷ���?x뀀�0_'���%�K�Р� y�90	��RBl*�s{?	�/��e���e��s&)�l*��:�Ӈ����_�q9�Y �NG��?���Q������6��8V0�b$:����m�C�]��ѢBU��(4<�� ���M���'�}cTv<eB����N����ˏ{���e� n8��j�����ְ8@�n�=��\��6!V��Z|
93j���j�E�_��������?M�������z�����+y��|'62q��)"�KC2����`�B櫬v�"<+����Ȁ�gO>SS�������X<x�t6р؈Nyd�3��*U#~����� ���`���ޘ{v�Y�R`�J�w��.�фd���f���jey\��+@k�]-�� e>�2�ܧ�{�r������"��[����;�����.a<�E����>���p~�@M�~ #K�Þ�v�c$��e1�[2�j2t6V󵫎�kƳ��u�ε��C����gO��ߙ��#'��P�lj&%ՙ���GF��C��DLp�$Ic�ɅH��bA�p?�۹6o�Z�ظH9;�M�L��摍��-2��pac��m�O?�4��n����T,�z�v��P@C��-@�$��R}H�ne���h�#cL���LT6�1������<x�S@Ѳ��Ϣ�"�-ȩ�0�����%������ٱG��T����)/���*�<� ��kak��ak�C6R[�,^���y�Ԫ��a׫�Y��a�?xb����ޖ�ЎG?�bj���­�I4������#H�?{���ӹ�配�ՅmTŚ�@ti��p�N���J4��(�z5���J�f��mxI"oK{�H�ֹS�f�p�t.>���?�Y�?���9jV*4r;g��Zuܷ�U�Rl��ޏ���1�vΓJ@���wm�]�t�X��7���L�GOKmZ�lN&���vssc�t(ș]�� ��ƞk����j2�ءB�dL�k;׮��Qh���M^9k2��pt�s=v��m.��s�s�(�Ɍ�Y1P6�� t[mD��eA�!�z��%CԴ�M�Yy�n�"(yreQ�#�ꂫHz!k|<�W���������bMy7�q����J&�ʁ0�t�R�
=M�E'J�6�t��4Y����b����{H%�Ih�*���ޞzR@�]�ג��F�����M�;o����W�]�tCҷ�ɢ�H��K`�ƻ�����퓋�=:g^��(d(�u�5xٚTʵ�>{��{j�����{�4��h!��=�&���*U?v�����?W؉n��>�R�C����ќ�3��ӟ�\�� g}Dۃֵ�=�Á](S�؇�jT�{�صnN7�s$Z�&��r��:�K|Q�g/ᘅ�]ڏ����?Se��^�����ٿ Bb�@��=�(�>��SU1��4�����;�@���Ik���D_"���I`���;�7 a��gϒ��RN����<���#	e���X�����r<��q�S���Pɵy�w\��,�wz�&0�Q3�c�(��؎I;@'��ބ��A��@R�A�7�X@ ��@��dO��������zu4�f�7S���\�}��%��{�]�4�q@���,ѿ�h����EPI=eP�h�x@�}������|Q��7���L�7�i�6�UT�;�A�8CG�r����i lwMI�1�
�*-h�W��d�W�s��;��2�+)#�/�fHz�{�o��͕;��b>o���&9%7�Z�#P�'L�4l�ɐ'Ѿ ,��f��T/L���}�j�ٽ?y��=�#��Y�6��ě,��JL>_�{�6���u��1#��JM��Wwr�ĸ��̵)�m���'�ա��z�1����r��*����A)�J����$�@?��8ʱ,bY}�1D͇�����-#���G6�i�D���^W��GS<"�"���@�����խ21@V�;��v�þ6�}�Z`|CO�����-@�~���Ȏ�S�r��U'l����A�:�RȷN�^��tt�������uwq�[�*Hk����%jQ��lլ������D����5�΢Yߡ�#Ã#;D�ӡha�k[�b�m��ʈn��@zJ�Q%��(B�l�-Ը�3�<�<.Ʋ¶5�t B�p	5Ї��A%U���ؙ}����"�^MՋ#ű؜(pV��03 v�l;�M�, �&Щ�,WU3����x���'�еM� *��W�������>Ӏ�|)V��gi�:���d�;G�W�&L��l�K��e!���1Q��]�+*;o>�U���]W��
�p�����d!$1WE�V0E��g��l\^��G���=��Cɡz9�v��:��yE��[�-���o�
{�=����'>M�k�/�v=�m�.�z�a!e=*A���mCG�O��j��¡���zmk�tSȤk8�bI��|1�}GQ���<ѫ��Ҵ&��J4*�JR�b"*�)����z�f�����d���t��+����G|8�4�|QC%����1]�� ��y����.���]�G
�j����U[�ڔ�z��z�y�?����U�T~����U�r/ v�h��v�������M�!sF�7/�>ںa���Igخl{�de
��)#�_��=���3���5$*]����X>���_��_uV�m�,y*��9$�o���7�JO��E��b&�{\�kf����&��e��hji�ݭ_��#J�
p����瀡$|��J:LK����αvr{_�ӿ��1H���Z�X�!L�[ҿv��"�yI �1ys5U3�cRI����C�Q՜�Ie*�?�\��萞
�Պo*TɦA�W0z=~$�!�߇�k�~I�D�HX& ��L(ST*x�$V��]���^�����:���Ԝig̽[�+ŌQ銆�Р9����9�ZY�����y	��v�|��2!%v(��}%eT�`�!D=��E'�de�؁�f	H�-����$X ���[��b�8�~��b�^�V�#�":O�V�a�+� k���5�C2qS�(S��8}cƂd�,�JUH����\n��������W��(�88S�?��PMT,��ݷ�Q���f�C�٬���²`,6������IA�џ������Ҙh�9~�;$���szqB��hio��v�	�:�s�L�fM����:\�L-�Y���#K�����Hm �:v�} �k��Z$6�@x��@Y dj����\n�������^HT�����Fv�G��#8����8���Wx�7��lh�e�[`~b0&zE�F����,	/Y�tn�����p{3��)�$^��¹�����a8������JU8Z,�%�Y�ae����0߆�����cz�l���tz����s���B��}�wvF��Q�Q?�{kq��re�ye ˂z[�1@��X��YO�a��=:�Nܙ?.܉�
fq�.�­��R�$J�J�����|�fbvma��|��QyW�)�A�lp���K�ь���앁�)�mߞ�0W� ��JҴ��P����u�g��4J�������ۭ7Z��ö��Y\�=is}�� �>�/�:繎ͭ�:����^
���qE�c#�t��$�f������i��@�t\�(W���jf�u�^" ����q���
ff����s�����/gD���Am[-*]����{>'�\�3�3Xi[i���-7�;��[�����uX=�e10 n�Aԯ�1k��Q���k��m�������3_Ǯo�˯�m׳y�Ӝl�Ċa]'�J:{/sY㉍·����ނN��CTRË>=�z`�bd��n��<О�i卍s�Qv�d����Y�{�_��d#G���z�V�4|鷩�qs}�dkvJ%J�V^�Np���"�\��#9*��a�9ı>�r,��	���j|<l��Ot�Tϕpp3����(E��X�Y��!�'���3_�#��v��_�7����Rg)�+�fu�:_�?�
�oH>l�񸻤X�ȧ�XAs�~,i�i@H�9�Y��܆�γpx|�P`m[���"o���=@ �pAUcM �B%ɥ7���n|����a�|����� �
�.���$�o�(Y�c�s�9�D)�	"!�$'؝H1lj͞�O�|�� ór�y�4�����_/Y�@6��|�P���@�q��΍������g썍��L}wJ5Ci�v���8�ҐL�����I8��$R+�R�s�f��u�$�U%���7�:��u�3�w���Ǻ��2�������@��x�p�+%�J%�a�$%��q�s���
��g�B��_�Z2�4�㚎	"�͹3B�������g������o���o�<���k�+���0�q�z�؅�f�[�T����_�=���/���ծR#��ʛy�W͕xt����"�Ώ1��ghMB9k�nS�pi�:62u��f�+�I}h����)�l���4Ԭ��m0���ޚ5��zo {�^h�ʡ<f�g*���voo�	7l���,����Z,�f{p R�� �u��8O���V/K�t�V�?��o���I���X*���u*�ƍ�Q/�ω	/�_�l��@G�	��LRk,���	���i�#{���3�sQu�'U�T#�j^��Y*��D뭁�{��Q�>��=ش��BK�:���%�/��־��&R޴ב����=e����F�x�H�5�"b/��� ���4Ff
$��}���A\Wn�+�L��]]�|�����>����{Dv{d�ڞ)�;�8$~71�v}y��ү���N��9=<	o��x�QW�re���:v-@���pP`\7��'��߅����px`�n��>{V�7Rb����Q�	AboБr�+A�j9�/�Z�9���׃�Q��ԏ�)cCh��*P��[��O0c�TS��znnnU����D���d��hP6G���2Ѯ��oԢ,P��kc���8A���jf7t�clː����ø�c��B�L$Un]� j����Z��k���Q�Oc#�Fĕ��M�>@B)�)�`������� �0:B�J�w����hvT��GLO�
�a�b��V� n�A� {�nN��6�c�0P���Mx��Տ���b��`��%� ��f�c7ٺ����˅�}5�� ���%o�9����'�m���D��ABF�����@
������k��@��	�=�l�l0�9�����Y8;8�k�b�v'gg��A�<���%@�������w��o�+y�5�sCi�+����=O�=��%��4�,��1s
M2t��=�/�Z����t!�:V�E����⃟ː��)U��V�w��Ɉuh��%6���Z��׿�@���;������k�C)ǠR����1vq��,��6ޗ��PbU4{~�T�U����q��s���r�M�z7p����ߒ*R�y�W#]*����}���=��lZ{�n��%3��;��h��<�����"���@��C�?�K7�P�#���/4����'�5b!1��h�X�4^��R֪8�Pǝ}�.�����K��X!�h�
g?��mq������OSJ'���Dq�Pm�ɺ�����>օ�兄��Ŏ(��8�����>iŋ�_��cR��;����3�[e�qH5 ����[��G�O�b��<�WP��o���:��T��/�2|����/Pg� ������_�����d0F���g���۱{4���e�v�>���O?���{�յ|��[�����½������9������
�$�?����S[_��U˥+������6����>
?�яt�h!x���W��W��	�Q�V嚻^G���M�6����N�/BҢeSBJ}�a���k�<�V���e,x��#����ŝ��,�0���ǪK�CY4�i�~��Ōҝ!搀ǝ|
ZU��Mu����T��h��U���k�#Ps���ש`wj�[�S)˳�B�/�v�x����_��������	%���r�V�:~'�ļ�XF����q��(����Oy~�?s��A������{��v��xp��ҺWW��3QO�#������e�-���{�R�O���ܝP���8ίf�n�N|���ng(�N��8�,�i#RF�L�j���>��B��G_ ��hQ�or5!����{zD�@Ԫ������=�{��"��	.m�?z�>���%]{N�Lvw�"�!�|unl���q8<�����ٍ��.y��m=����ðo�ۆc W��PNn||�W���i8-2��[�ue`�p`���Wq���_E?�B�z���b.�_�W^{l��0������_�,���B�y���B�_��������mA�����+;�Ix��y8�œ>�N1x��۩mlæ�P���76���[��˳�Wa:# J�9�,�ok%+��y��<�Y4l�JL3a���ڊ-T��Zj8[�9א��^.=J�R���z#��o*_���=�� 6q'[��y��/=��kb�N�{�����ϲ�U
ȑե�1��,X��9���|ԫз�p��U��F}ж����/?��6ϙӺ6~/$.����^梭�eG`f<v�⳧7v�	xg�fɭ��t�T��㍑�����X��g�.�s�T�ِ{��g��C����s��P��lm�n�%6p�t�����#4[�W_~���6Ǫ� ���h{U`8R���2��6�����?/�&���{J��ф	p8P&���x|~���|���ÐMە֠c�"';T^�?��	�H���g�IjFj��z>�u�ӏ?O�ٹ���G���+)�g=~�8�����_��_7�|���\ I�����G�Z���H�r����,%ڢ�B��f�Tbٓ�BU�@Rɳ���s��Q�tAg����Z�Ez�36�/$��o�e���!c��a`���{�=
��X�LW��'��&��;���
f)I��LO1�z�� 1�.]��9�EE��.t����1��=�MZ|>T�S׮n��$��!�g9 �b��xMBk��ŊGb#�B�o���*x4����&0Q44�L4p%.�'��܅ �����>���)x����:i�����B he� ���y%u˅b�wb��d��Vs�N�b23&R�qb_P!i3a�D/�
�9��&�,+	� H�+�&��(�.�Eb��K3�8(�C�;b_�>_��Wԛ�~N2�t,��vE��������Te�������P���,���aTZ?�𷶟�R� �$V�o���|�My�=}r!�A�!�����k�����Y7zQ�	�w}}��`f��Y��PϨ0~�k_��?��n�� ���;�Q�X�Tv�Iѳ�Q�U�UDD4��v�֋��]��8etن��z���B׋�Mm�N)|QE$�C�/�[��n�s��6��H���)�Aje�3��#6��.����z��jIk���ݯ����i���
�B�o����'���3�E�T�B�aM��(��ބ)8j���Q���&� �MO{��㵥qUk�u����z���+��L& ����-����d�Ƚ�ˉ��ZPz��ǜ^����?ۥ�tҾp{F<6W����c�̭K��v/L��5�
b�H�Y���NY+V�j'Cȴ(�<�K�l�W����c{.���7������\�*��m �ŇeȂrz֟�7
6�@d��
�|2���Ce�m\n, R#�F�y���Qf�}��ւ�M����~�4\�����sB�#)�0����)+k�YG��g�`����2l�ǂ���g����M[�����'9A헙S��7��UW� �4��4��-@܆�}�J|��]۸�j�[7���7��lc�.l�x(��T�w<A�wc���؆���&��P4qa���Z�_*��{ 3rWrӷB�H'K�j]�����6�/>�S�0S%5��U=��^A-k]*��E��X���IJLj}��YT("`_.k��m6s)<��Lr��yG�c6������ ����i�ѧ�e�W���؄�+�Ȱ�l����V�5"�4p�g��0h6����
���Gt|Op�nnc��hO������T�.�1?1Prx|��,cnzy�  �ml��E�M��v^Ǿ��<���ae����l����I���j�g _���h^��%�Xg�l��Nl���~!�<���O�������x�P�$ךL�ǳ̬��ⲻ ���mn��\X��F�=ӎ�{*cK��L?��c��T'z��u�sdV)Z$��\�Y��?��k�	����%&�\	���A��c���ї��%*� ���0�� �����rA	�*��nI�I6�꺔7mpd��~�rJNL���Qm��䥇�X˾�>7�NU��.߃a_IPh/ 4��*s�q�^���188ǧl-X�P�ޚ3����6��3�E�d�宅���/�����Sˬ���$�}X$�K���ZR�.5��Վ]f��/�z߿�6PuT��D>�jW���7����X}j���^�4�'	�:Ɍ�����t�sרܝ�_{��ש�����@1����h��(H���=ޟ
ZA�����c�����]�l����o�MBp���J^L�/D̿��[NO/] �3^1ߣ�5�>��7ߕ��yk����|��SU���������v��?�s2[U^e�P{�zjVל�8S�9�@�[o��F���'z�|�5��Ai������_~Ob/̣�����������<�=z(�)�bL��}=#�|�z���YC���������	_��W#�;���M ���fՎ���~>I��1C��������ӬZh���;��n5*�df'Jfkx0m|C\r7�x;�MY��_��x��Lz�_�xOp��}]��7�{6g�L%�� ��\�gRK�҂�k>;�����*kO�`�x`�O�Z�ɼl+�b�q"�%�̢� ���\	#�F�,l��ຠf�B�ejl�ӵ�}���+��P}q�`��4-���k�����n���j���˫[m(�X�c�5f�c�9M�f��ݎjU�E1iP����dYIR�F�#,h��(��{Vn����q�5ך�R�ޜO.�[��p��N���m���ht3w@��&�e8}t_�*-7�/-�����^
��0�ǁ�lƗ���b�T�+�TAC���%G8���ѧPzR���{�Ε2�&ɦ$����O�'��ux��KRy;?9G�c�1xo���턓�N��EՁ�KhU:@�������Q�)�R%X�*�~`]@�Y [�se����a �_����=�~3�E}e��,� ��ҠI�����XZ`��Pj�3���)O�T� M'@,X���'V�I���B*L]�4�w��N [�U��:R�*P��eK��Yl6��>C1g�qݗ�=UQ��&������@W'�QG�U|�[7/D^wG/��*���b֑*U��ҿ�^P|���.&|��C`��oo���UV��=���q��mv�S�\1lL��u=^ڷWf{�X�����nHY�a��"�q�U����ĮgNթ��ǨZIM)W��h6rhbY�i	|Aã�|q�G�txb��H=@�m���z�y�,��at��{��M6�K{�W���1�KO�H��9�jw(gSgY��^��)�G���7�Do 3hz���J�&�ۼ�ĉ+��}�dG�w�[�D�!3�?��"`�U/	S{����Վz:A��ٙ���_5�@G�7H\J]ǀ� }R >RA泅ֹJ�3�[���F��7B�pq���{���X�IB�	�`zKRj�"��^��� �7BcBP��{�6��瓣S��iT7ꗒN�N�wT�:=)�{鵐_�C6����qt�(��ƛ� ]�� _�8�;#[�
�s�g,Q�TU�,5�W�Ǡ<O=����	�u���=P�����my�6�k��6�(z%����+�uOF���d��|܎^װZIѻT��9'#�T����I�5������-������R��n�A����v�J��f���Y�a U4�"�m�X4IЬ�������~��C����o��}�k�WJJ�__]���P����H{7�H� PBE�
����������F2��YcB�el�N�~�M��I�I��C~�y����C��?�Kx��+�_���W*7�%�}�]�������_�O>����B��/?��������bk��v<���}�P�&
�2*c�QM�e��>���D��"�E2��♘ۨ���z��vA]��[�U��<A���vm7������țJ���5q�As�f�b���"i ��?.��C_)�N�jh��!�@Ӄ��rtߝw���TA��/����J�,�i�hRO��5�sq�������i�������q����bݍ<_J���,[�l!e\é}u{��Iڴ�/���^�B����ެ<�s3 ����u��Hmf�&wՐZ����/k�cv*.�\�K)���e.����Μa"n,Z��(d�x�t���:$����yJP/BEh~3SS�P`��a���,��{���3of�0Y���g'�vl�iX_N�.É��d����<T�wl*Y�!H�S�w碌�:Vox�������.�h\O�|ƷW��p�6^N�O-�(�=��؆��0@�$;-�z!O���Z�o�ɭ-p������җ������z��9���.�y�Э7N)�� ˷�u�xt�;����}�(����`pn�2U��=��u`���
��M�T�B��������b2���=�*���R��j(�-h�H�3����< ��/)�р�uMwb��m�ñ���< ��H�N��+)��D��#��x0jsAEl�G����!���A�`�߭��Ln��y�l`�'f{V�} E��%+�@��_4	�<���~��M �JU�Niݱ�=����۸$C�2 4�Wd
p^���J��f[)�m1��$��Ζ������j ��c;V�~M�FP}e��Ս2�4�c����Ka51pbǸxr�|����ༀZUž�FJypx���!'�]zA���ϯ���� ;{��V�6NI��~�)7J��0����5�[po�|Jz��_�9���KF�4���QR����Z�w��{���Oܩ���GS��dV��k
t����rZ�&�Q#D��:����l=��(Q1!KLe�`�5� ����B�1���5�׉l6��X��Tȭ	�o�B�2ΕC�+)1�E �jO�S�����ʫ���eldEvA��AXˇ���ٵ�z�r���9h�pY���a�l=9�1<qe��5���~�{�e�6�]lӰF�o�x�~l4�睽ko�no������z�&�>C�Z�e�^����݇Nĵ@	J2�Mr��Ob�K��푨�/�fꔴQ�(o�=U�b4R�R��}���~�5�������g���I_�d�]�U�{Y���D`�{��R��2���S*����W�g>�Ur0�~C���(k�@�����1Y��L�E#ܖ�&]���I�!��S� ����I"��/}I��G�.|��'�aG�J&����Ӧj�Oޗ��Z��W����'�
�N�c;ƍ�P��s��W�k��EмX��ُj���ZA�X�=��,$J���yrXT�4�U��q�q=qrw�j��¤�y�2m�|i(��q?�|M)x��e �C�B���z��i�V�פ�jO��#r��9�����g��C:֙/!���OK���e�i,O�n�ԋ1?��#��"��GE�$o�ddq�͖t�O���r�
	���&R���SX�i@��3�`�_�:�)�a�g�7�=K�������ٻ�lw�f�B�:��u���{=��J�P�[T��,[�~w���f8��NM}U�Y`r$���Q܇M��R2����0���&�]5�ms��qU:'�G�Z���iXٳX�3��X�6
��kUPA# `�މ�dJ5X>��P&�l��; d!.��c���:�/o���u�P=
{
�����m��Ҵ�c6-+U8=!�Yzc�����\h`������3��Q9<<�qEY��[?ݕ��Ñ}v��fd����ex~���CU.�}�c�Ϧ���F2:����x��u՜=����zzrߕ����VEFfiAj�*�m9�۹���2ewl.�1T>./��ԛ��N�0��\�3���f�L	$�AC!^�O��<:��`����v`�j 5:�D�ږ\�˷�?8���A86����q��^[��E�fh�}���^�eN�T@����2p�BD�T(]9�şW�GUjPJbC#�>��\߳{rm�B}6���ܶ�@ɱu��G/I�h0���exv�,\\]X��vR��%�_[�KI�~!�W�6�5Y�2|��"<G�b���݂�ƭ*�As�u2��/h?��g�۫�����͵��^�E=%22;?�4�F���q�!{�T���
{�l�7k|=e��a2ݞ�s��HC	/V$p&�[U��N��]D��
�ǿ�X�P��O>�X�ߕ�g�n�Ϧ����������oR� � z�m�q/�ʅ�ǣ�d����+�	�����`2;�c_`G�ƣ��t� �����' ��)H�+z'�
�s���1�N'���u2s���s�j>ye�ރ�l�$1C�%�b�,D�*~��g��97���|%�&9�5cL�)*կB'�}��/e�W�ǵ��������Sq6[U�����_�:������H�#$ZH��H]vU�����I���v��8�����=�n�{<��=H�&�q����is<	/�A��6�&Fl�Y�����vI��`M?w����֊T��I���y\\"8�/���5'9�n7����A	$}b�C_w�S2u�����<��.��90_>�����\��$o�ؙuEʮ�8�MlE_����g�7�RE���6v
�F�Z��G<���,1��ր,*5׊=\��j�sxc����淿i��\)w��d>xp_����1��X	�'��u��pÚǜ�2Z�&q�9��m4�a!L�0��v;��I�/f
�!���>�P��-�$�Di �Q�|����Q�'~S�H��p�qb�AP�M�v����ARa�٨=��q^l��[e�_|]��*���������N���k�`OJ�$ճ�Z4R��A��z Y7���𔆾>����������L�W^~Y�w����Η�Մr�غq��s���� �V��������h[7�Y�>�9�Ι�+p�f�q{������[��V����sjJ�_p_��J�u�,E��YD΋L$���:�~l�r�_$����}:�:�=�2�U����r˓���@���G��z
,��'�����}>���d�'�k�I�A�!����'���m�����y9��}n�X������?�a'�?<��Bt,2�eS�i#V�*�y8?�c����``�Fb������c �����-����+{~�����AO�n0����lL�S��{�'��Wz�|td�}n�2���p|��,k���6zz6���:��=�w>Ǎ����S�5wV�H�X����V�CJ�mς׹zG�9.lq����.x�l�^"��g����6�ϐEr;/ד1/K�(p�о�rN�&�o�FL����$Ɏ���:��ʒ]�
p��{�%gy�; ��4� ��Kd�֡�}�w�=w��j�ódgVdd��'�]����Ɖ��%��Y1�7��R��0 �p��+-P� !�YK@~���0�*�j<n�A�t9�Q�ŝD)L�*6��Ei+#:��.�G+�I�Az5�ZN�R��O��|���oé�32jC�GL���8K@�#L�=��k�~{�,����gx,��Л-��:��Esf��Gv��T��C�;���<}4H�W��؝ښ6������fl�뚍g�w^��Rط�_���l�mE)z���9�X�x ���C����%}ckn��|��+U
޼9�:��-dhN�iO4#�E����W�[��;���"�,6��cG�E�77��+YJ:_�RY�q��g��\��\.Ң�c�Z�6�	N�_��k�4{I���2ފ>���b��'p&ը�+}��n˾���Æ�"��Z��r����u��(5��i[_�@�cӊ��|R�d����<�;A�f��������{�������cs�_h��:}��(��q�*�_������uFlSz��,��x��U�Ԁ��A����ʞ�x���i���]}��Uw�L2��SM�ު�3xň`~csKɝy���dj�(Be��t4_e�c���5�j�i�`(a=wj�{�3����Τ�䛎%TY�x�Y����EMϥ��DkJ� �����O�~���˃���$� �&�&�e�Ns�X
1�2s���s���hMvn�F=�\��@�R)�<9�j�  ��	��JN-^���M�螬p%EXMOjZ��(��$S���c�V�;�z:QDC�k�XU��R����2i<{P-���;��|����"�/�59a��+<�F1	����	q 晗+y
��"��`bFEж�>��;�]s�Ձm^Q}�߼�<�R�$���%���>��~j ��>�ydK����\��O����fN�!Q�R��A&��없�q�Y���g���;e[�: �_��W������o�rb����_z]W5��˗�j{m����H�=�ʠ۔qzw1	U#5���G��{�"G�!�u��E�����N��l0��*�R]�zԼ:�������e�&%�!��"�����[�d�l=�׊͢���GR_�x��'��I!��vT��`ɢ�XF��(H��h>;����vؼ����[���G>:�����N\���A�����i������n��*;/�m� 7m��t���Ӥ�ݎ�s��%�j��<ͷ�oTt�\m�m����AO�Y8z�*�}}?�mo�!���c��pt|��g��i8�`4��aS߃�H�}[�760ܲ�� �,���؞��k��0ٵMGR�B�lZ���jJ,�]8��R ���أh��UP�L�L������Ge���ld+�7j�t�g���x�;�� �3��]�D��e�L]d��J� ʾ�
Lf���
Ƣ�m�d�8>[ԩ* ��Y��Xp�^�E}��	QXZ��2X�bB�3N�UԬ���Z�t����L�C\�e�XʣC�w�C�j��/um\Q#��I�����J����B�x�.3
�E��n�+lDT�ַV5�.�����\�qgW�m�,J��̳�_�`�64��898<Q���"�#"u̼�J�[	W��\�y_�WfUO�t���M�8���7�	���@������)j�ݿՍ��iL4=�As}~)A����0�wO�2��Bف&Ւ�YZ4�=�$��;�� (?��L`%�6�51��{��T�	Im�G�\������ ���V���V��"9\�"3�Q/\�(�HzrrlA�z����{�y6st����!@@�@��p������{>�T�y�&��6�Z
*���T<�s��J������=�b��u[Y�\�E��)^\�rQ�ޟ�����x�5���d�{������8�������ŗoN��ȋ%2�^y��J!B"�ǒ5Ϣktj�ބ������"��BeI�<>�7rM�)uY�	"R����H��2ѭ}Y��v��w�8(r�6`r� G	��dvSe �˴�&�ʁ@����(�7��R�S�,?���gP��m��Z��߈2$7v�{�4����,1c��]fɝX0���t�A;A5l����;��7�Us8=X���0�M���Gk���Biy������M���Dq�7�c�
��x��UIU�[ۛ���i��dq���K��b�pzz.�]�7�-�C]�~�g�I	���$h�<R��t����H�L���w4��@��s~�����Px3�K\���~;9�~�������΁�D�b*��8��|n�Ѩ�B��ZI�6J�X��~� ��@�\z�z�&~�{>�9��{(w_��?�/����7�[/��Д�m��D�.�{'�r�V<���"Kj��]�F��_�2��&��,,�V$��`�ئI�w6�����Ԕ���D����������`��/������
����C�TV�Q$I��^���x�(֩M��;�2&�/��<Z�mNί��խ-�jv��<+e�^��<���R��uuTe�R�����z�{H:���d�'
I�P=Q8��0�h�/)�L�s)�����2w�d1��*��EJ��:Z0�][բ�d���U���
�T-��#Gl�htrzp�{�����A!��zJ5��P]y�*��������r:��2ub����T�<4JU������T�T�g6v���1���������p�ӟYPs�؆��������t�)�'X9:���yj_��m!���r6S�T��n6o��C�����%���AG}'�aa���+�"+���=bB)�Z@:�+k<?��Lo��E_�QC�>ykj�ҕ���[�+���쮐T�ܣ&w��8�&@�J��[�ܽ�6���-�$�d=t�W��er���`���V�^[��.��ծ�-@�1M��#�[Djl&�ݙd���ޓ�JVl&d��+���?=L<_�,��_� zU4�C	���>Sf�6.�����TIHl F�>���Tce$JX��_z\6[�JJ�h{�����@8"Ն��g6��S}�\�� !ǌ?��K[�N..é���(d�iE�� ��l�;�4��C`k��Ź�3�� ��(�Y�S��Gʸҋ5�sf�����a��y����"�������s�)��`���5V�xLֹ L?��ӥ�U��Mݥ�1X$kّ�r���g�D�%rrʃ�9���#$T�HP���;�2ISP�N�.�?5̛�s���4D���Х׽Y9���"p�ަ �Jr)-�) :�,~.	ۛHz��W��k��9��ݸS��=C����A�pW2�ɰn\��,�x��;�˅�Ͼ����w�k�z��Irͅ�P��Ѧ):�i�W9*Dl�P�_�DO�*����LF� A�5�,���iUυ��jT�}+y�T�X��*�U��^��sU���T���Չ�? d�d��WY��:���h�c���#��럓O��X�#w(����sK��g�} l�	��>��tZ�XA���J��ϰJ������}�v	:���Դ��p�?�����D
a�W����g�w�ݷ�VX�y=׺������_��z����Q�Ͼ��$w	�Ii�(��y*��������ᑪ��&��#�����]�D�g���G�G ����Zx����3�N��=���2��f��5�W�����!�Ae>bcW������P���QR+buB�Y��(SC�2������D�̋v�=Z��3/�|ލ�3o�b�Me�f(��H��t/ߥ������fN*ix�,S�����6M�f�G#���� nWu���7?��� bA�5�� 7���D|��-c��m�3ȭ��?����_��_h��ksf#�q��A��7���ʊIjl�������]��P�������h.���@	}}�l��H�^	IuS�G^gz��NC �9��~�qWBH3GE��F<ڮ�gI&� '�bUl{�W��#D�����,��P�&ۑfc\xi"]�Ts����(�g�۶-�ۏH�v`[���I��]�����GOՠ����z�����iPÝ���Ƀ{�;�Ǐ��^��A�g��r�-Gڈ�3@qpW֖�fY����J%fo�Q��ʯ^%���IX߾	[�re��wDO��"/��N�G��#8�P;���o�/l�6@�ӷ�{*�6��@����̮O�jI�rq7 �i�fsk$��t~c׸��UWr�n�	�3�4|Ӕ,�$��ʮ7�OF��� A���	��H��Z
�XCgH���8�y�E��~K���y,��B��@�uc#�l�U�����|�5W��Xtj��`Z���_AE���I 
hp��TԪ�۱�F!����á0�g{����1,d�p��z���o�m������'@����~^1�@�� ����u7�����z�N���	�f�5�*���E�ߑ�#_H��F��F�2�����@��rDudE�! �Ó�pvym�U�����\�Ƕ���&ʤ�?&N޾��kL	���{���Ӱm�C} eێ�F�d��mm�!iW�����قm��y��;%aY�KS���r����	�R��ө�闵GҨq�#�b=���'�n�vuJ2��EPF"<�v Ʉ��FI��^%�8A?`��H�&$b��b{D�ԓo�S%��˶+v-��{���H_�Eb��z7P��i��7���Z�{�y��C�4��ښ�����_*=TVX����X�!����q��?������Q	�B�?�ִ]�����>C�	"%5y�4���tuB�$����BT߸��q?JU��/c�?��XUЯ�TB*����έZU�I2��rod.���*\�*I��3܊���.Y�����i�C������Y�tRh�
���.�`�Pђ����Nl�YU�I{b�Dt�[ND6�Le�BDO�q��'g���z����j�>���P���?���\�z�� �X�~��@j7�[�_�� ��3�<y�fu �@nno�7��9�Z=Ic��Z�VE?L�(	W��F`�d�o���ÓǏ%��7�7Jpo��������rhV��lmV��Vw鞗����k ^H�s��bϣV9�'7�E�^�|���f�pX��zA��\��%�J5��RP]��Yj@�D�W_�9��71�:�ؠ�N �2��j�ƲD=��\�^�25q���y�Q=�<��3�ʬ|������o�ZjҾ3��R�K�Hc�*@���Q�0����d䫯^}��B��2hW]"ne�A�$�����c���'�~*��������_�>|��߲q�[e��&o�2�{+P?WV�p���&\⬋V�-,�G6�-�8��u��ڀ�q���^_�_܁t��]�n��,	|,j��@H��I�8,��ɓa'�&��ؠ�%����	|��1��3e�y{W��f���S[�IB-��1����v?����@c*x|�-������X\��cx1��9�k�pC�;���6�zf�W�;�Pj)=I@LF�K�cI.��$C��mL���(��a�-Û���о�?�	�m�}`���'���[܊�v.�!����TX�:�5����.N�pt0��B_��]C̥��OE�i�XK5����P�25���o����"lﮄ�=E#[��7}Q�VW[R�$RO	�[r
/�{{ގ!�[<5px�4B����^㻭YS*Y$w<C=W��]	�?$�G��ཐ) K���/Ԡ0C�\o �A�ׂ�T����%T��s��UO���E�}8�������ᨒOo*ϳz����M��)n)	�	����������������J(�op?V0��nK��@��U�F�¥�J����J�/5�&���`@���>o]r�d�_Ri���0���[�Wo ���̙*��'�v���W��󬡈t�+�`DE�����I�:?; z����jC�����SUz s=�9;�����\u'�z�����W��=.%��������1�:/�{ +�������v�cA�+����A�����(�N�{��WZ�Q*0���H.K��^�'����sm���+@� ����B5,���qE��]�<&�f�m/��r
UOU��g�I���^UZ{n�޶g�.���1�O=�m?Yd�-J�+��V��\7>�������O��3����J������ti��E���R�s6� :"���ƽ�2}�
q&Zj٢l7��y*k�T���|��q�z���=��٢�{PY7��˱@���M��JG@���b��J*�s]����s�P@U<h�?D|c�T�p���[���Uz-kY����s �$m�xAY�WI���0ɛ|�+�j��{��J"WI��"�ߕK��>��?�J����U���R�����}��O~"0�����?x@Y�O��e�铧�� �K�E!�^3�G�v�������[z[R59>:/,�K��E�(����n��cQ(��3��=�� �o}���w?����g�U�˽e� T �H�~�{�h𵧧�F��<��%i��=8�綾�����YT/~�˿�� x�T��$��ENߢ�ţL����\)Z ��hS��[�Hn����Hh�
����i.% Pwԑחŝ*�R����	�d��ܱ�n������R��e.%�@���/�5Z�|,}V}]���
IN-�m��FC��& \&�K�I�J�W/���D��o�;*;`d1�O����#�X��ߟ��()�|��M�=�>�.�E�y��sm�;�\h��e�\���ZeyTd�,x�� {8�������˟���z����Ƣ�z�OY���<yt,D�o�7�Mmw�ͣL�ԫ#����ŝC�'����>"�2�x
\�܃�C��z+�:g���&Vt�z�v���K)��x�ɷ`dǕﮇ�o�L�^W{^d��W�ڛ�^KΕ�	]�n���z�Bs][�˂묽��AX�;"h�@�iQ7�+��������vw�¶n��u��pr8���b�͂dq��C;[���}vn��U���
���vD�_����'�"K��:N�p��
 PPzOMz[;�������	�XpG�k���LT��NK�T��4�-�'3x�S�$F#n��=7楚�1w�^Ҽ�( >�P%�?�	�0/�x�����뫙��Q|h�[QOE��p��P��	|���Y@E���T.�Sϊ�y���]J���������1�
ȒhD��f��^/�6<l)cM)%ڥ~g�}ۀ,A���/��������O�ݻ���+�7g{�jN�HwB�x0�X���j��Mq�7��z��o`�0���(�f������;=U&0/l\���q]��s|k�|;���8ǘ�;8��`���Q��ydk��.н�;��^��Q<��>�㸵�pd���r9֤|���$'K�-n	����>�"]�{�X_镽l�k?�듡�D�$���I����WF�r�d�D��7�����(2L2�2�ii�e�w՝�H��*��df�������Q�aO�$��+]�=X�!�Ĥ`� 3��O+*W��0�O�ϫ�'�� \ު�Cgj�9ߔDCޓ���Ρ%yp�<
|�]q��.fkGvO؇Gp���3��2�j�ȈU*c�m��.J���f���M���P�j��	��V�j��/)�UD�� K���k�JHJ��d��-Q�B��pJ���yM&����E.�1Q��I+��߭(?�D��<ދ�v�F��Lo�:.���Q釤�Luc֝�rK�{����1���V��iq�N?���Y!�;� 4+z:�i(g|�����}��hV�~�����c����c O��S9���(���:���}Q��71�Ϸ\k޷��**T)~��߆��{Wղ��o��\����z�ϞN������/�#�O����� �ZOx$ʧ��u�����׿�b�/~�3]]�S)��rt��`.qΩٞ�"��ŋ�Nqn�v��P�Ǭ���Լ{@��ݨ�˅�`&�PV�`:Zh\S9�Rg	�$sAwnΪLs�{��Ԧ?�fE]��:U3M9��x�,�7��K�.0/��ԏ����~�1p�'� ��,�*�ޤs�O=��[u�|�J8�(�H��}j��6@���/5Y�nln�-۸�|��\K��F(J{�V���UM��;3��=�L���"�n�8�:�\�&�*����Nq�`A�k魛�Q� �����6�&p���o��,�jE��w(�:�{�3�>���R�T�u ��G5�T�(
L�J��7�\���X�<��Y�O�2����|`�LآL�8�%�;\ȏ�N�,{|~6v��BtxqJ�����ƞԭv?
cNs�PV���*l�aek%��?�����|~}������ ���Ù��6�R���1.l�yf�y��W �A�2+����a�׍��	z�H�^���/��7_�{������ٷ���I���_��K
[3U'�w/�5���{;�v���6�yf����������-�\�1 ����BM���+e�����C䭮���дB6�7�\�;�X�E�fA����Qر`d�![��!�`-T��|��h2]m4�+S+`oZ�Kn���J��RYH݊Ͼ���h����ms��w��W%C���Wn�>G�G�BPY�z����hT� +E^
�&�p|�1�P��,eb��d�� ��J��mcf3<~z_/��I7�<�� ���4�g6�aS���Um��/�6F��[ T�)��?��b�ҵ�nԭ��'�clZ|�S���d�����%ٚE��QC���(R!�|}}^~�Z�����1�*#������46�1��Cgܵk6T/�|2�4���[;�8�o����T=N QAEk�>���^�vn������}���.=L`��	v�_��U�^����?�E��g`�v}3��T�<r�� ��쓁d���۸#y��K��"�iPm�j���Ѝ���Þ��YE�� �>��Ђ�?��6�O�8eHodH�m����W�E������3��b� ���ᶳ���[qKXTq��M�� ��w��]�v˫G���k�2�l>��������������ځT�n1���*������2؄5e�o(&A��bݚ,\���2w��<:����W�u�e��ǝ'�E�X���t�V�zTY��^֨4��%�	Ѽ�n��1Y<����0�+�*J]���mLX���?9}v^G�X�\�}���L�:�E.�O�ZwB��=k�0�Q�yϥ^��ڪ��'U}�Yә�T�- -:⪒�P������G���Y�=�ka���T,��h>�添������P���/���m��q��G�_�vRm6�С�BuPtt|�D3k/ ȕ�\��7�8t.��� o���x��)�Ɏ4�LR��0��m���?�y?�q��'����{%�퉼����\�Q"4Y�Ԯ�K�ͣ�*1�(�P�A��h��w�(�$P�&�����J&:Y}�����x΃%mg^F�D��\�s,����ww�"�;�ҹn�A[�3����Բf@���C��1��Թ���7g@���*�("U��E��O>��¯�������	���e�����(2W _�_u��j�c�*�|Ĉbi>' B9ao�~T�H���/I]���iH�� j�����z���776�ϔ1���t+4�i�M��.�/������"YYsl��G�ٯ���L���F���F㘅�q;�T@����OO�J����QM���]���G�	Zl�lA��	�����E����^��M�=���-���pq5���4�]O���m��9ۻ�-�߱��met�Q��@:[����B�l�z.�]z��V��AmGw�e�;_\�;+v��L�W��?)cK���=;��ׯ����.�Ԏec�>����;w�鱺�x��@�������,��]{o��>f����0
K�eБ���ma��������B-�on�����
7���F�39JS+�w�B��4�f tcx�g!�۾R����E+��.⦜��Np
��{a�?��\�+-��
����MD���O�o�W�PE������ʚ�e����x���٘��	99�ȥC�ff�r�g�<ܶ��ax����st:�I=���
������[O�?҆��o[��6&	b�^2�������Ǫ^������zӢ@��$fhM&���p��r�5�E��,���`�+�{�4���oHsP2�$�9��(���݄����Ѐ�l���?���A��{���ː@��ЅÕM�(a�&��R�J���-�Oy$�U���J�?�K$���?����uL(߇K��fT�zϳ���፥��v$y�'�֤��?������`ԩuߣ}ow�`W�i+��5�����K�F�F7Δ%�����h�-\�EZ'C�R�7l�>&���ud��e�2�Kl�8R�NLL����P;2`���*Di�OU@KO�'�i[�e�����[Ƹ�����F���ѹދ������?Ϟ}�>�(��_����K;�S�@�-�z�N;�<�{�rI�fuU�F�?eiO�H��ʔ +����vW�dilYJn�hk��׭��!��ԉ�\�h���J^�/Q�l��kԮ�5��^7�J4�k�g~�(7�
u��8���Pǡyp�j���<���C��RÊ��N#��̛��zG�����$�f���:������%�������t�����;���-�T�Ji~�{s�^0N� ���D��I`އJ2�S������N��&�ΟJe6�<�ے��!�G�Cq��R{���K$��V�7����ɑ��׶��O��&;gxP�f�������Qsy����1ָnm�-I���Ĭ�zHͣXDI]G}��y3�^����V��Ci��G��A�Ɉc�vJ->�k�U[������ev閷뛔e���g �{U�v(�REYO�o�vT*�HP"͔�Π��#�2K�S�W��#X��%PS��_��)�|�
�}�X%AP1\C�~���m��%3略�BɔX%Ө8'�9�N�I �˘`��7�䔛G���Tqu��YJڔ���y̝��{��ti���εW
^����v���,W��$[�.��WS�oVĴ�Wܧ��BsM��`Ge�:%?�>�ÂN���o�^��F�ne s[ ��(OZ�����2|�@JW%��{�u�x�V�c4Y@����2dv'׷�L�փ�ae�&�G�ŗoÅ��o-x?�`�	�^��>���#Xs&�Z���/f#U5�\��y��	Te2t��|���vE�M��ѯ��؂�[��\��dr��_���b���������h��wb<���>JS}��v�� Y yujn&��9�������_��7 �o��7Z�D3X��q����<����, ��\\#w����5�B� J���ח��h�F�>�jw-��ۺI��o����[��p���\d������d�����硠%�Y+	�_`^�e\V���퓕�0���7����'�9���B���S�"&����hV<{d��#Q�z�(V�X=95۸�<�8V��?��=�|�� 4W3�çrӅ�|rz�.n��P�aws�6�m��Q�V�,�8U�]T8HJ�=�������^���
|𙪎\�Ȑ^�j�%���'�`q�_��3IZO Ж�g4��Y>40s߂�]��=�r0D���T���}'+N�?�t�H�ɚ��~W�qum��d��X߈&}k�P�@H�g�Cd^�2�b@�l���y���8қ<H�+w�yd2����NIaJjV�l�����)�j`��������٩T�.�~%�->�J �
�F+1C��͝4�pP�O�h�ʤ^?�E��B�"IB0AvU�A?x�i�~���˟���x�tOҿӰnǶP/]�J�=�\�]qN$� �=�~P��ȭ�;���}�Gau@��u8;9S�Е��*�^VՍ�����J>� �����fT񩥪Gz�**�����V����=C���|}�����(w�.I���GAr�N��M6�77p�1��W��I��81dBLX��!4/^��t�3ʳ��L�Q	�׌�`��ZR�������I��_�$3k m)�-��n;K~7<�)b� ��ܠ1�;�T�Br'Wr��>�{h��Gl���p��.\�3�q�����TE��JZ�:��X�KT�J����_��)	�1�T����g�e+x����y�H����2Uoڭ�|��pn��|��S��L���2�^�H��h
�̻��T})����2�� �2�^�S5@Z�m�[�q�Fw��JwNh��oT<��H�t�o%M�����\%�[���dh!�Ld}��|ݡ�8����GѠ��y���bqh9]��N#���_������w��Dy��ZTδZ��z�'�߄�soH��	
2xt%��)�@��JZ�=M�R�<�?e1�/
w2���͍���p��ע��ͼ$dj)k_U�\J����u����su%�ކ��Y����\�H��ͬR�tlDia ؐ:�]W�
hY��҈���*5���-�6ί���@׍ͽ���rj2�k�Yv���]��dնo�A�m��TcJ��k������+���}�P>+d(X��`}c'�/�5զ!~+yX���]z����9S	ɺ���V��п��)���5�qx��+[�v��OG�.�^����z��I�dǿP��؝�V����[�T���m��Ӌ�p}e��f!����+�U�\�<\��c��gE%�8(�>���� w�����Fc���j�e��K��p{Ŏ�g0�����1��� �e��1���M&8���P�`q�s��}�q]�|t��^�@(�)��� ^Z`ME�l.*LQ{��E��P˥�E���==����&�j-)$���0q-9P����nس��woW�+껳�2g�Z^1>nP'l�f�X�������*�`���@����~-����µ���3PP�&NV,��;� Lf.�9��Q��ޏ���������7�*�e	/��쾎�VV��+��7t��\ew;�D�}ٲbc��mT=Z��;m߸���?��G��|�*���6�N��B9�����{X�A���DJ�A��N��r�o�����۰+��R ���T�N~"��g�A#:�B�@�{������@�������.�-���Pp\y��JU��A�� V���z��^�5��AU��sѩW���0��8��q�=ƘW> �E����ùyC�B"�uyvH�5+�1��N���P���`Jb7Ut���V�� :��gO�v������a:cJ��"�SRQ���=���b����)ꉒ��«�e����	8�ϵ�x��,���k�:��w�X
�1cEO�"�r���{���欪L4w{i�H����z�D�ϣ�.��t�+;��z�+w'~��/�x��.;�����f�ٌ��V?�&�	�~-�
�H���b�"�!@_�"���QRc��[1���BY]�f%�`?	�@}*C��?vl��$��{/\�P��jĥ8�J�9"%��W��������'����:�h>�
��6�XQ-���E���@�߯IN�Վ7>x?G� �_\��K?�������>.�')����Nw����Y��-�XSwoz��4��n޵m�pC�4��$��mjxN��9H����͌s
�S�!ơ.!Xk��30�1g�n�(ե׿D���ߢ�H�nw2i.�G�%E���c@�=T́�����J�l,�_�x!�B6���+���\O�E�q6Io=�b �^�Vy�`�2A�T\*�@}�g���T��Wx�t�~\��N`sm��)J@��<�Dٴ�"4���w�ʥϪnp�S��W4*"	$U�5-�	x$�nXBf�7�3m�䒡mn�����2J6ǆ�Q�|]�<_��\Z�$Z����G�"�>x��IM���������@����,�����Flm����!Ԗ��pc�h}m'����=���!�d-�A��o�
�����{�����ƣ�4����t���Kt�-w�U�����M� d_J�G\]�eX��Z�u����x�?���&�9
WW�Ahv����X@�o d-@ú�<�@��i��3A�HUU0',�8����j�s�>5Ʃ~�1�Z[�|5�<e����2����Y87�v{�*�e�ڱ붽zk}w/��Z!���;k6��+B�3T��|7��՟������^����N��D��J\�*�Jo�2�*JY�ȷ�ou���pw_�Ǚ �� y������t�a�n�HZ`}rJ��:�'�!�����H;g�������Mg� ��k�"ǟ�� �*��T(�>{���($x�!%�����kJ��rrr����޶�����4�տ�ZB�M�O���#�:�6v1-�0���􂭭����a���J�x$п�r�] ��ȟ�^��M�������7ñ擨J\�!���[�^m���&{O� Dh��G��Ҁ��c���6��8�~�m���g�h����U%�hZgS�ٸX1`�����ioe��c!9d�K4�_(��:w���BpNһ��I���}��b"�t�^�j� )���(�>[�	:o�j.�4�B��W�(� ��k%8=��0��<�? �v"`�8G�}������ؼ���L��*�WWnr�Kzj�/($'�]hܜs���K�5͓�i�����$��a�t�F�m/&�B���E�wcc%��u�L�7�
UX_g��6#����S4���@)9��&�FV�>$�R�<~��ߧ=0��W��D��E��,����Z�"�-QT=���yS�I젌@5�7e�T�Z�u���Y����B(�<��̸mz��soEѷ/�,���Rr�2k-4�g���9W�q��ݾ�w+�U�R�m�'�&����0��E]�P��q�ܼԤ]y�MS����TF����F�8W�t���R��󨌷|�͇�g�V5ga[���S�?��?h�̣? �M=�\sO�t1����/n�}Ď��J'�<V�'xU��wj@r瘲h*Ӹ�JF1.�xc�
ȝ�~�Y���D3#��,Z��v����X,�&^[�9�s)U
���P��:A�lY�M(��Hx��	UW�2,O�*3��H������le�W�+���u�O��ٳ���
2��_�`�s�K�҇o����c��(�M*�q�o}��" MK�l�Qe��F���?/WsIc��o���t`6��E6R<ƅ�q�����~�X3@rv��{�S�����A'�c0�6�:��˲6�-�R%�Uej��Vy�s5��E��#��t p�h̦���.������
���h<������a��}������伽����8,��܂22���g���߿^��-��8���v�����ѳ��w?��&�S���!+�j|���as{-�۟�Ó�0�]��pGaz9�(�3e��|���Σ-0�S4�s�xD`�6-���7Q8��W�Լv~~m�ԍ*��m<��q5����B�\&E�g\��'��[���3W��Y�����lhe����vX)z
zT��0̎q�0�W����.,P:��V����W8�{	����(��Od9��dpo	dm�_ڱنe�(����%��?��_�F�l��󕰘YP6�dև���p,�qn�����TM���]���]roẻ����n�Ӑ�r�bA@ ��!�������?��4p��}U�D�j�Q��|Q�b�**^^�����������A�������4a�J�{o_42ۋ����������/���9�
�`�6��ˡb��﯊�s=R��܂��X5��򠞽B��%��a:�P����1��kCU%a<���`=� r��p6:Q����0��*N�J?,^�*x�.J��'v�
�ٟgEroGZk��,��)������f��)Qo<�Jo��q�I�E`�^�6�?�A�(�j}�)^Y~�U�)�B#%�I��)-�AΉϠ���'�}_{.tS{�+���݌7?��!�wQ� ��ʽKڞ���EW#�b�B�J�OU@�(6RT�n���VYϡ��e[��'��+]�C�b�+InHXʤ��
p��CO�����Q֥��Y�o^�%LB��M���N.'�s���x���_Q��Ɂ�+�ꈜ���GL^�y��5@I���\Y�+<F�$>�d�y,bKs��&Rv_U�,��1w�+���7��O��9ݬ���0(���yܔ%�����������Z��jE`+��(\��rL�1�O�q:�F�x��S�e���{N�@�V�����'�ɯOL�7�9����h��������*#�V���E�|Nʶ"�dCY4�B�Z��哀"��~ۯyi�ծ��9�.I{߈[w$�(�s�+���R�r��8Z'�gz|�WĂI�i��Z���\�En��w��s���\�,B5�� )h)����t.��p�6���
|���g i���ZP���[[#�:�M�����Σ����h����A�>8������R�ƃ��?���v6�dЄ�9�k�OT޼y-	���ӆ<�B�;��w���|=0|c�Ǐ§�~>��#P����&Mz$4���f�TI����T�8��R����s5��9���O�~j��t�� >΃���u�"RrB��;�H��X����M��F+j�G�!O�������*�Q��μ):�t:5é�J��J̔�UN��y��?�n�Ʌ\�l~o���Ʈ�HY�/��=[�|��z�z�:|�?
���W�yA�h�E��������Gao b����p�ǯd�Ƈ,fޘ|u=	�XP�6U���������0X˥(���u��=��"<%ņ=���t���~�6�L���p�����Y�y?|��'2���_�s��R��X����:<|l�>k#�BrƬOзz=ܕ�C��2-�2��,�'���t��ެmLlA��r�,���ق��}��A�bq*��3�l��}p�;�Q��#�������>��Cr��c�PZ 9D�+�����v���[���D
�'��mq�/�]^"�p�j�xB/K)pE*��DQĺ��Q����D~dy��c(�3�d�zD�o����{P� ��>�a(�Wʈ��wsCJG$9dL;v�*��`^yqq�O|��������U�L��p^|���px�ʮ��6H(����U����E�T�9���O�<��(P�:�HQ$ mm[�4 a�C�
\��8�۹��\'�dd���9o^��x>9;����u[S����ө�Oc�+ŴB�'A=1[�:H!���?�M�l�[�|2�[0���T�n�\[�$�u���Y���8^��\1�Ƚ>�TИ�g�3���Օ~핱�V�D�U�� &p��D/���&�Tӻ�<9TTJ��eYɵ�D��)�M�I�
�{ՙR�E�9(���As���:9Ȓ�(�P8�+��g��P�k��������7(y`|������'C�Y�*E���qO���F?$�Rj�N��k�|N���5v�fɾ!���h�����4AAx$J��E���`(��(�hU���ɐ�âhll!Ƃ�����}z99ˌ�D5J��,�(4�2*	7@��"I*�ME7���0���V �y]I��}����Pj�6d�� �y��h̹,��2��;�J/Ȫ���QfJ�'e�����}�K6�N�6��<ϫ8��4����-Q?�R���o���֒`����2�@�<%�.$)��)�ϣ�jri����3G�8��x�㐮�Td�f���;!�~�;�?$�z'�OՆ�����笜����:bjn����4C�8�́S�]�����/���z��»���� ��>��NU#��g���ݥd�%�ńܕsi��t��b�$�^��kz+��_���d�?�&�(Z����+ɹ�m��я~����K+�ͬ��:o ͲZ6j:���"�)�p�����rD- 9>9� �L��>{fǳc�p��(,��@�ro��j<��!Q��=UL���� � �~�Z�c�3z3!�I�Nr�3��)��Y5�jޟ8u0d�Qw�:��tӳ�Nfg1u�l,�̀&|y�U2�=[F�)�|�2�z�ߞ�z%������L�v���>�}���a��~���*[��m�+��_����	TB7Y[�c:.�d�������WJU:�|�<dW���F@!*o]��k;^�6�X^���7�E�"�������~��@/�}.���n���5w��C:�R�Bl���UP1�͐C[��� �)��қΡaLl#�\Z zi��}�Z�^�b�FĖ5/�85� ������=Uv�v6�Xza����T@��\"��U([h �j�ֶ"Jh�u�M�#ȣ:!� ����j����f8�9"󨹃m�+Ƶ�-�n�e��>	+HT3�P![�u�%-w��{�W�ʄ]���7��D������;��� �2X�������:�G�^e# ��4'����T� �C#P �;�/�\�gg�
�:�9��X[۱���"q;��ӫph_GOlܞ�:2�M+�!��(�.�w��U�< �LvK�YQ�@��x}�f���%�}��k
΍l Ɲ�������p};Tf�-�jƥ�꾄	yeXĎ�2fh[�j�.���=f6w�}�l�v�R+R��xn�����ny2�k)�KE����7� � ��P�ѳ��+=y+f�K� 
8��-�O(X�`��x x��Zs4�&UM��s�38�{��_���*����C��!���E���k��s����Q��Q�NG�F�G�u鸲[�P�"�d6�k(g�2����jo$�BY���-�u�m�Wg'��,�2J��^��u�Z�7)>�DY YܳlZ��WG� s�<�"EǍ�� I $�1QVV4��;�G_c�V�8��Fn5���C�3��mU6̣:����El�H�7�j�
w���je��S�E|A�L��"�9��i�]�m�U6�u\�&!��W$���hf�L8W����5
;U��Bf�J<��Y5~�����j�����Q�b�#���w��JOH{@|���x:%0`��;�s4ۻ`EY�C�s�/�S^�/�)�<XkX��-����-%�tb�����Ibfa��#��zDQ���g����i�c�J� c$W��悦E�Se9P/����+Q���˿[nO�_6��{�mYF6iMe�L��.��?X}H���w�x�Ξ!i~b�e/b��MN�n�u���/�k�u�;��4?��ӈ^��1xh�| ��.������7!�����u��w�IIg9�4b�duY�!��8��\�=ۘRs���YI21��1X/"@�r����NK�L�s��P�ʗ�,���9ݧ����+^F�H]�(��My{1R��Iֶ'y�B
<�9���_��;��2�}M��R�?��xa�ȷ�J{��-UDڶ�­�� ����?�$��W����aV�8|��p���ᓏ>������~�����W���l�S[n
�y��g�I�u�ޏc,~Oٷ[a0+�`N�4�9:�5 ƙ�n/���#9�蔹���ފ.3��y��ܯ�|�Xͥ�G�.>pC��&ll^˭{k˂ȍ��ǖ�Mi�ne��?�����M�b�� u-����"��n�N�}�[��f��Z�s{�R�����6 o�͡�9�de	�rWˑ ܷ�	���z��R܌���vW�ܷ�VD�x��j
�+�߸��fN#��³�B  B+�2�=��R_�N�ᘩx@Ϣ_��؇X�& O�^̏V�=}��͐Ү�͋���pi���f^'�����H1�����pu~�j8�l���	�P���*� ;DE���G�tYkn#�%F�۽5in����Cގ�ف�ۋ�ppr^����Ht�E
����e�IƜ`��A�'��6��n!:�̀:Խ�X��m���3o�J�1{�����wBw};��򏺢������m }U�����^=����牉���m�l�d�+=͙EA����֙9L��Ui`�z�G
u!�C�h�5����S�mWK�獄d���>�~���v�xH��Y]�C�]���댹-����ЎmE�+�9`Hԫ����~?�B�DM�u"]m:u�2�P�����ֆ0``=&�����ID�o�,�r8���ٹ����)c�k���(X;�������p��}`Ƕh�\m�\:L��J��丳2�Λ�\�#�(�����$�T����JIr�WD)��J��Lױ���&��R���7�����t���IR�� ]��4��YJ��8���b������P�u¸�w[�n�FTSVc���oz�ʠx�ݹ $��B�4	���j:���]R�h�>�	Dޓ~�|}4)MMvN�0�ҵ�W��D��ڣ��[���~�TI�R��!��F�1��I�=P�Ӯ��п�Z�P���"k�hV6� 1xa�����������R#��Q5PI�K�j|����΢���8�7.j�RY��q��\*�q3�L}(>�&��=*���je�$Ry3� ��n��E�^y��5�H:���xweＢ���n�����Y(�'�����wաB��He��7�_�����c��ٵ����u[ԟ~�����U��?�%pAF��_j�!�a�B� ����~WM��m��j����@qs�C��Ƶ/Cu!e'�.7��v��F��'2-�	q�޾2����I|t�Ν�'�Xth'��@�0ii)� �.#�i�Z��T[	(-b�R�ҥ�Т�B���%�<�S���J�P%پ��15~��Ɇ�ͮ�7I,��j���=/��u>�)��Þ�����}-J����e�Y#U	�����!3�Ƥ_���͙q�,��7��|�qX�M��ӧ&�8I֍�;�7oU�@ju݂����>��[�t�������vS?��S%ͦU�T=J#y_&| ���ȂǷ�U������Hɞ��D�oU��[qnw,���9�>�tH l��\d�1	�i<[1�����$�����q�E��mme���P]:e��xq�>1R��2�Xlmݣ�f2��?�Q�e��7}���n1�u��6��K�н^��
Zy�SpT̑�D�;=��@� �V���6���+�T z܌�菓��f�zO�S�J^$��2�3 ��o[2�+fSW��t�¥�{mm3@Gyk�6sv�����U���>m(�35\S%'����LW2�t�"�&xB�Lr�e�g �y=�R��o�i��غ ����^qZ���0�e \�n�h"
�H>������d� ���@�ٞ��r��Q�:	;[���?��<���pf���f$����=8��q� t�	\��+G֕�3�i�sd�}��T�����\�uz��]����4�6�5�g��}��f�s�/�i��رP���"�)!{�xj�z|�J{>>�&U(@�,�*$��Ѧ�L^�:�H�<\�> UNb@sb`��'��z6�0 ��Ln=��
������,U|��\����3�5�zFp�\�Wv�6�7��j���t}����B�mȘ���O?��ה���
�%�4C@Օ5ֲ�4S%}>KԖ؈-���x�Z�z�Aoݬ]х����O�T$E�XO��u<���d^���
���wZ��'f��ؤ��*R�<ޛIR2�B��Y�����*%Q�,&��E#���Z�Q���dC-7���ȝD��&%�tᙱ���z֝tl�۞`��-d؇�{������F�6%���_��(�&�<��zU^Q]����a��{�b�cK�^w�6+N�B����W��"$�������Z�)�:�����?�����_���@	�Br��5ke[*CܜN�u�;�8�Za�Ŋc�K7��3�Y���y`:U�}^Q����oH��{�!���r�Ht2�v��ٺ��d6�}R�h_�c�Y.O�w���C�w�B-��<!�b���^]�ox�f��{��=�����UV�YV����:V��I�dސ'c��k6���Y*� <m��,��ڮhX��>���M��Oj$J���B:�>�El,'#�**#�FP^O���i�FGo���nn�辭)kYz���Ѱ��	ȪB��mG�J;V������T���{���y����d�F��K	�	���q0g���Z.�˦;Q�_(�Z�o�Di>r����P-����ј�ג(�]��p,3�3�G�2��hX���(-P�hZ� ib�6��
Iς~ ޾~^�|b���>�DA�7���40��r||Z���O�ự�*��婚OW�U�O�orq�U��Mg�����c1�cM�qcsU%��ˑ�h�D� S�i�㞲Wl`�'n�/_(�
��ѽ���f�܆���ԛ��d�Y�(�쒔�pzj� ��vX�5���
��'��a����p�]�`U� ��+5d^'6N��Ivf�S�X���r(:3����%�$9^'�Zw&��t��B|��,�ژG­nK���z�1t||.�ˋ���ڑ��&J��Z�?&*Ӏ}�m^E
y=���^&Z�O�q�����Ymm��8�j�w�C�*@�	��P�˯�J����{6ַl��h��߻g��� p?n��&R�C��TF���y�>̩���JU�,���n`�ɘ���$����Q���c������?�4�cd����D��s՛%:Q�� �V��JF�s�#�@������َ��<��_��g@�c���J��cR��YlE�� i� ��{��@��%a�9��d�^�}f�5�sf ��=�^��G����1���@ۛ]�Ű�3��b�
��H��'r�P�:jY� }�á�y ����E�i����r��O���4����S�����q@�H��T�d�����H=͓��-�m%r�����͍��_XB�s�8� �=<���_���l�ɠ$k��"d�&.�n�z-|�;����m�ڕ(����?;ۻ~��`�mA��X7���6�tu�*��Ⱦ*���So�wCK�3;����;d!&/��އX,xޛ�s$Z��`�.i^Y�Z���V��.��,�yL��� U`$�V�2�c��p̵��\"����*��:!��:H�]J���&
g�9mM��H�
Y���tR�.Tq�b��c��$�#	�nׁGWb��=+���4=�2���*���W@�:��?��[��g�l�~<M�/�6��s-��Q���g�$�QT��;�}�����'?ѽ�[IBŢ����g?���7�Ze�:�<�\�e������I�6A �U��,$!��x�UR=?�� �N�&6��'�+E�ZRY�lO2�+��	l�˛y�e�f�Y$���L���|�KoЄ h�����X�2`k��jH�X�B����F�P�ǝ`?M��Y�,#�4�� ��,�����:`�Ҡ�5��Q�ׂW�$�V��Ȅ?������i�K��F8_,�fuPЁK�kU�V��t��V	�d��ZDN(���qS�����@���vAF����������ㇺ�k+�������(i�
S���X٢�퍰a���uyu�ŜfH6��l��VGx�9�{:�`ߒ�ky�Nfw<��/}&�N�2?�L,@���k\f3��y�-� �]T"�� giL�j�뼗R�"G��MU%�U
�n�<����u���?�	�����Vf��pk�����y1��슂�jA¹���X�}|}�6����߱dS��T@.��P�.�
����ە����= "��){�;U�y�6�6w-X���s|��>����9,Z&�i|PX[]�q�g�-�������h��t�� �\N��O/�gG���|��D�h۵i�:�LL3b�
�EtYiG���k�
c�Fҝ6&����li�$���@�h2��;��S�� 
�0Y��J���H�:JQo�]��E�% �����f��Ojg$�-࿰q��J;z/5�ƶ@K�M�8G;�������)=�a}u�rCK����:��z`T��mm�ڑ�ɱb�G�ɛ#�K\_y�
���Jj�eQ0�/�5��ntVd�;��~qu%���3.g���Hm�?����+y~����/���T�*,��b!@�&�RY�=����-0p��}<��1P{�������჏>	��N��~��KUE�NN�A�>�<�^�PI}����i� vKk;��/�ro^�/��B�Օ�:O�����o���Z=��"UW�#�^�I�Lr[��������]��000���B+���1#�P�}@���u�պ�����N�{6�6p&����O�˸���$�nc��"��E�-�b�}.6����־C�,K��xxp��nnm�"��
3J�#��Qea�.$?�3�i�^�v$�1	�.ޞH��*���`<J��,����;��Q8xy޼<��L�G-T�C������˫��o,�RPS�ī&�G穷�p���l�}G2$Yl�.�>�
���)������R��&D�����r�;���E��������'���X�XJ���X��_H}Q2�n��l|F��F���*�|jl���ؚ���X��8G�J�����t;��H-.�?����M  ����:��O���﫚�k����"M�vd/Sa�J����j@���9������' �!H�>{������BbB����"��8p#ʨ��R`��JY*(#�������~Y���e�~�Ł���#�[��eN�)n�e�9����يj�s�}�U-lh�ۡ����0��~�a��WW3�S��V?�#��厝5��z�$�^�;ot�n���e�t���[�&�.��%5WS�U�r'�f"���iOM�� ���P�(����|��/^�+ |�u9L�.hP�����V�8z2��d��Dv��H���6��=4��XM�k;{aw�����m np_��I�<�ڀ�XT��9�-��}2�q�<��o��H�Wⴓ��i~o u�Fy�(O#�0U�ρ{YY�<K�k�+��e����{Fp���J�����j���ɓ�����ʂ�o^���B��V�������Fp��e�6�y�Z��y�:eh\��X3�6��-�:���+�1��n�B�T����ptxdA���V\�\��(Z�Ni��q�x��������C&�����3tq�'���A7l��B��8� C�c77C*Վww��ӎ��d�	t���~�^��E��K�cԬ���K���Q�y:Y���uU�z�z�~t���VF �F)��C#sҵw�sw��)����G6��F�#��X*.���k;QՋ`���ׯ���g���tu�l�h�cD)s�YG�-jOH���8�x�Y��N���W�a|���e��R�#s!eC7�jGj!���-7 T������#�����,%=Ƴ2���k}&S�����@��uH���"ߗ����$3�{Ъ@�����ٺ|I*��*~�d�ّ̑����J��. ���p�
	U�M;��G�'�}+|���ރ'�����^�
����7����$��&X�D/,��0u���������JkT6�ã�prv�uF��yOTE5U�W�M��!�
�WUI)j��(��q~~�u����_ۚ}Wo�o<�q43�Z���E���j����'헾�����Ӳgl�U6��הk"?|h��M���t6՜mu�v���v��~���%� xz���~��Ʃ�2�el��H5�I�ިF�T�Bb�E�ۖh�=������@ܮL;QGb�A��Db�:���w~�]�#'R���3_�6��GL���P�{תd <1/�I-�J�<�'f�ˁ$�)zU\�<�_����P]��/%��ঁY��
��r��e#N�c�	��qX�����z'39��lY��B��-��t�N �>k�2��p\4�2H�'��UoZ6�:Q��J�E���~���| �N��b����c1�ZE8��	����`�S��}��w�t�fߴ��I�����\��4���u�SB����S\�o׿���x����I^�؆���*�����ϡ� ��,n#�v^���ȕ�y�&q���F+M�(G�3�)����l�A�U#�Zӂ��(N�wY_{�N4�F#_Ȇn"4��(��]�y�T�[ɽ=�]H�\�Y��|��YC�������������j3$�xx�u5/�wy�<���O��\�:��P�Z��k*��<k�"��x�#�)�E���^�%YY�ͣwY,6`9aƪ?�}��%y(�0��[�\V�ajA��Ќ����I�u�
���O��=}�a��[�(0���mF��Y��M��~w�
����q���J`$�%�U2<T抆����*���4uZ�ae�l��x�{�BU���9�� �Z^~_j�k���c��Ċ\�;\�m����yo{;�@o1��X�h�Û÷j����vض �ٓ����76goE�/<�����a<ȧ����X�V��0�����Dww�%oz�q8=���+���^.B���6�Y说�˂�Վ�Ut��x�g��1����v�����	Q�%v�j�j��l䥚�+�_��Eo%l�@�B����=cx"�TY]�\p�ƻ#�턃3���������,�
�a������Yі�z4W�M&��,Jmj��,V�P+��^ȃ2�>���*�^)��S�1;G �
���5�:�`��K�|��@�ɠ��.Z�!���WQ�<���}~{m�j�mv� ���0������ d�Օ�4!;��Gþ��3�7R���LU�U�Va}e#���Dʆ{Q��]���KU��/n<�O�ջC��z*��*�1[d2 K�@��}owWU ���?�޳G�,�3�P�+3+Ei�]��G/f��K<���$�ܷ�ٙ����]2�������ճ�8�6љ���~�^�&���l:6F��G�L*��5!HHA�&�	+�&'���"OV��֭9���#���O�ɣG2;?'gݑ��ڕ�x|�����5;g�K��1N�����!�T���M��4��\�y���7߼�=aO�>A��5Y�$�����Yy<րbvv�B���m�`�����S�ԃn�3�T��;��eEJ1�� %{ti�,�=]Y����G@ ���gh��TЃ������+�L<�QԿ!h��5��� �Wa����̗���6�Z5��3�N�F=�M�C`�+��<�Dkʠ*&�t������׿eU���i{F@4��d��=V`Q���=���zKVVWd��2���j#{���3�;���&y=����c-B�
׌��Y�Zeׇ�ǜ��:FX�MP�6�Uh��¬8�*#?�^M3�%hP��ņ����\�m����(��}5�Sb�Հ�HD_y�d�AE�p���uש�]��G������gbD�'cE��q��&��65	���F�?�ê����WC�����h|�kc��
��_��'T=¿�0��g���g��lnn>u��¦�'p_��~���S	���ϊ�kT�0�Q�w����z�3%d�)�YDP��I��2d)�XЖ�f!`L=����Ⱦ���߆Eq����WH�`F�2r�W6�=�z���JQ��>�ܡQ9sc�&���t6����������J���ߋ�k^��?�(�Xᒯ{~�G�G$���6����ð��/��+��Be>6�m��j�$��M��������l.©�w �C��ne�*drA��
�4�����M�-�vչ^]�R��qG -�Ѡ����ʚ|�O��}!bc��؜-8C&bՒd�����<39A�����X��c�1H�n�7g��G�鄽|��MUԍow{�26HDM���
�0 RѶ��0�Й�2�P�|X<�?�(#c�����#�����cY�w����oecC�#u�}�T�5������ٲ�k�|8�Ͽ�����3�Ϟ�0U؅�Y���~�-�����u����t|z�mI�"Ӡ��ۓ�LM��'��'թm7Hg��a���ª:����&�mpb����m8"̬ݶ9�/G�g����\�`'���H���GE������#ڱ���C��L|�sl@mW}a5����n�;�)���S̬�	f̮��0�Iy�1�킽1Q�:!�����X�"G�˥Q���rBJN�&7��4jL�����\�<֘1� ��s7<~��\���!�+��,�![�����0�B�G7	@���$e]����%����y^��8t�Z�-��Yo �gp�&�24�/�����3�~��랳zsv���Z}jpt:}���I������hu��a��ch삑X��l��z���2�,zӜ6�O|׀��y�s��E�4��������oI�qcnN�y����/�_�+�z�'��JT=0ͻz� �:�� �T7p�A�&�5��w�H��l92�`O2�kN�a�a�kN�R��p�A�=�Ye�f�)�?:W��>3�W���Tp:'́Lթ탽z&S����D����ᷙ%�Fz��<_0x�����d�J�+(!��=��ȴ� �	[_���Y0�58�Q�Z'�Đ�:�3ENSCR�n��a̪�+T~,�����(p�>^�:�R[�����m��s5"�g3��AB��Y����s��I�aJ�Sjg;jgA<����L��UY>���Yu�0h)�!��h^��=@P��> I�е>R���8�mH2��hp2�[�J���JG����2R�ug^!0{��jH�3��aV�\����)u-���o���>�%�۰9�GC*�����U�<3�k�I�� D��ݮ�}�i@y���u1�%R���C5�V\.=���j����z�}����(|HG�N�����{���aS�\ ��1�sxH?���ݻ$�XZZб�\-�z�%�g��W����BD��̹��'n�j}�pl���4'���T\��ze�o-@��cs�.�g�
�j�@�eI�*�W�fE��&�:���'*o��W�Z>s���n�Gڕh����M��;��E����p���'
AChFC�SJ|�WV���5��#���fx[�V�`pDJˁ;O�����i^���p���L-2�p ��r���z�2�{{}#:(>�����W��O?�H�G�T4ݞ�����@������uo�C&�,08�d�QH���=P~Ǽ��7�c���Pp���/�j6�g���@C�+�ـ�����O(s�j$�&�h|�j�F�3:A}�f�!D�1�pC��_��ޮ�φ�o�',�&�v|p��5�1�g��߭���߂:�f��>=M���I��+y˱[�}�"vSS�jN�#fĻ��t/�4�������aj�I���1�MB�����uHG�����l����ϣ>I�$�	�d;b��r�ȱ�{$/_>��]��sK�Mh�L�8�r�	���ДK7djf�`=:.[;�r|�&Z�<@�#U�i�N.腳q.�S3t`� R���8-V#(0e4�6��:�Y�6�ش_l��1�^���w�<8S�����QL�d	�6�Ӿj]Y�A� sO�}O�)0a��Ö'>���2W77��= k����V��>���>�ýu��ǬԢ9j��{ X�����i�y��
���y���ĀcjbZ�O����UO���Ќ M�4�z�I�mk̆�a�yB��'��j&��aCp�8����*��hhFO� 8l����01U�2yq<m�� V���O~�S�������2�d��D�y���|�Z�{�F�}�V:\���}άR�v�6[��rG�f�)v�Tj�ƹ%h�a�� T$��F 8�k��b����L4�*1+����m�1X�R���[ҥV+�uJ(��6�,���H�pp�p��j�`��K8�Y�3�6+�;�|o�	?���5@D�P-:��6�V��u^2��3 �k�sudw� �ĸ�Ι=G�X�k�kĕy�t'ڐ�N�Q��-��;�ߖt1X0S|'��5�+�]��32���I΁aG�����H�] ƺ�q���e_��#�#�T���f�:����%�)`�>(C՟���H��c�2��$p�)�}1�������I�P*�LxV����;$،/퉚C@S��2����A�a�	"��-���0��O,>�`u8.����*�Ur�g��m�z���?j�z���G0;͞����s��4+���Z�U��p����Ь�M�����*�_�q�?9*[�X��y�'O����ϙ�X�X'�s�	��7o.�m�DG�0ё� ��Ç���C���;в�A�EW�nR8ܱe�ǣ�ڮY�C�l�e�ݑ��8���-�∥���%�\�z�S���Wk#��6fN/1��@�3�l#o����q�h�X���mM5>�%p-�R�P�fU�j!�5?�(�
(>�����7����c| �(�H������ʪ�yQF�6����X����H�
���0�4���<d����x�w�������7���7��>���z�i���^�`cd��s3#?��<~rWVV���O�@��������q�13��(	����%fN��砆p�`����BD����cy��|��r<>z�T���7ќK���ydV�$�z�+\KN�X�`��b����ʜ*���8�Ǝ~���-9:;����r_r[�0@O�N/d��;Y����_Y���b��O��X��`���O7}l&̪g9!]�b�	x���`n�_��r�J<��]Vg�&:���9��ػ�۩o)�;�P�u������'�Y�vK���)�/C���zn�s" ��!vxt��jS ����gj�M�R,[lF� h���yfA��ֵ��w�s�B�����՗������Tרk�ؓ9Om+�G��a<��q@�3�bdi�p@�$�F=|�&d����p�9�ج �ݯl�Ż���O�^N/�d3o2p�3K�q���)Rn�Ee�� ظ1�%Y�}�Y���9Ն��=�p5BO�C�s"L��5�	@h��	�cQ�Cc���a1x6)dk1��m8��W�0��*�a��$�Q�DQ�%��xS�BK��&`:�!2�� �9�8�4�><���!a�;����u8���?`�{��Gr��=}�.'��jp���F�W�nK�X�w��	�go.f��?�Ү6��놂�:��TL
�!9N�U��9h-�x���;<�Jz����Q��
_iU$�	l�D8��θ52;�S����;1�?�=���U>S/��^c�r8+8��Dz�Ě��&�g��Y�w����HH *;5$�t}F�ZU�>C`k�ߠ����$��AQf��P}���P�
�`&��� �*�c_s��g�S��N��j�3�8-`]S�)6V��g��}�����^�'O�/~�9��󲺺&K7x����y�X�Q�{Cv���<dl�x���M��;s��ϳ��rxp_�tx���נ����Ev(� $4r��
	D�$A)6����nx�d�^��	�3����z��$��9q_O�.�� $*�ި����!�R��I���["�k�c#:n<+")� a��s���;3�K���|҆4��z>��Snԗ�'�߭��2��_����JƲ�Tȹ�@h��?�-�; ���s�\��϶��ʄ���5s`D��,"�c3�4I��� ����7n��9*����c:r���R��zu�o�(�n�*�:���Rq�J["�?5��F>�B-��� ��*2C�υ:�p�a���r��ZF�x�$1���"�lx#�xQ9
�P�����sw���/�<����{]�����9\�]�i�K���Ւ`^��xo�j��`V�ąBc9�1��j����M x^d=p��7��NF}�:�'�S:(=}��ӳ#B�����f��I�ީΫ�,�ސ�[hzmț�/�����$/����N�g� ��!����k�<9>ܳ��t3<ڷ^�l<4�K�������_~� ����Ā�B�l+�nk����A��(�grF��� ��f�~��6�47�/+ t��j �}p(o67e��]6��az=�R�����%�)�Ց��" $˫rzrF� ��A��E%��!T������q*��3��N�<�[��A�c61Qg�ŉ~/���}]�sN7T�P��j4S��>��j�3�qB�4���v�ْ��9�g ��$2����|[И��W;;[�4�9F���D ���X�ƴ-k�3�y�P�1>��ΐd ���2�Jt�m���`�`B�6yVLBr���{�p#B��IJ�R��swmm�����ֶt�Ͻ' +��A�ib��T�BB_yf&1�`�t�g[�	2���W�X�.Xap��ہdN��F!�
͎��iV�@鼝mH_�&���0GП2=I/��6�1�	>P�A1���'�^k�(���u^+����f����W5���	V�i��D���Bp:D���ѵ���u���	���H�'a�s�3`��t�zF>x@E8��9�l�z����m�;���<��9�*�U��3H�sMź.���s��S�'E�D�2���9V@b⛀SjF�zBT�-�u��l�=��=y�?�����9B�;�����k�5��N�&O�+�*�=]�A�
2�AG�������{[�0��Y��|��?��̈f@���^콆�;�p"�|�������@��@sdp>��r�ׅ�#p��Ӻ�$<�����k@=�Ǟ��d������-��0c�^�В@�ͪ����2z�������˟ȗ?}&��6�I��w/^��%��6\�׀�`��@z��j�s�C�1��w��,j`��x�c2}<A1�&��H	:-��Y!,f�FV@���!遭�+$�p�M/+D��fK���,,���<���[�c�˓��t�(��!�	���!���0����C�����L������`#������Lx|�ӻ��]��\y��H51������z�.�6@� ���o����V] Jfu�Ec9��y^A	�&L��G4H�!�?��7����������7�`�B�WhZ+x�AL�L\2v�rT��B�f������}�Pf0��F��y���7ÉZC���܍�}c�E�96YQ���� 1`=<�N�G��A߄��v��
?�`���I�t�%�^>����?W!����J�X�������
Q��z��%�'����`p�T�Sۡa�Ɗ�0�Pe�~ ��pp{��� �[J�l�l���`8��;�nK�j�D�ed��N�������w�eogS�SR���ݠ�Ƥm���8�2�����1�V&�'��2%D=�x��w���w��O�`���T�&Í-�@3��fy��ĳr@C��fS�a_n9Z� ��)�}��{��#�_��g�*���}�����;Q�Gr0P�z%w�ٝS�~Q�(��ٔ��#��t��EF-Y�;�T'�qM4m�'���^���f�	7�;wרv�>*TQE��Pw���C[@�Z^P_���X��FJ�Z�(4VV�ل�����l��gj��{�pcD���srtr��De ����0���s����<6d������:�'���͂1�cu���M���!��4��&��g�;v52�脵�d@��8�J[�O���uk�,B�ø���8�F�
��O�:�G�J �dF_�T7p����I�("thiy���x�,�U�������'�|߽Y��2#kz����7ږ�g�=��������
�hx�,`��H\�i���A<�%aDf�y�9�3O�f�
�'�<�0�Kkkt
c� ���9Sg�@�#�)h~$d:轪E�q�'��Ve�U�:������wV�ȝ{XY!%�ށl��ɹڳcu`�4�9R���ߕ"�Z��@i�<0�������U��vP ��,��ˉ��È@L T�X}RC�nk�}�҇�Μ�H�� i~��9�S��%dD�� �/Iab&� �d�#Ω��lCܸ�`bP�� �i&�9�6#�F�P�FV��`_dT�pTPYp�tx�,oP(wl�5��K��m36zݑ�|�;�YSE7�0����[B���>�H%�U�,�Y�6Ф����ȪC��QE���)���Fr{�m��^cPC��F"1P����S4�~��|���Զa^u������;6�onn9]r��|e2#v�� c>��Wb:+H�,,��sqaIn�Ab�ڙ�tu=��1��&E�OJ������zd�-����7I\T	�������|�����Z|��Q/񽏇΂{9�_���z̭B|����^�[�9�Ưa̓׮�S��w�X�*,	�g�׳0���
��4����J_�b]�����ƿ����^ID��Y��}/�S$���KV> ���O_B�����<�s²q\·(.�6�Y��`����o����o,�����{,�x��zbXx�?I
���?c-a]dY��%A(U$&en�Hnr[y��q]�1^2�P�^w�����Բ�4���XX�*�0#�9��#��ᤌ&�	���~/�'�Y�P��]_.�2yU�ˇ�X�+�"��d)]��T��|\&]s�W�t�<�)l,t�AMx+�6�C�a�q�\����8`Px��}���aNxY�bg�Ҡ��=�A��	XMM#9X]Y"����-RV.�ݔ_�w��L����Y]ɜ��'iP�yC��Dj��b::��ٞ�����;�����:�������c�-�R\��W���Z���#7�h���=]��x�Ԩ]��5"���`_�&���׽}��-0���]9���^� +�LȒM�����ձSђ������pl�R�Q�{��;�����O�*ow����5㹹i�;�'�25���$+$`+�tG�����
0���:���Sj���Q@og�}6++7	�����8�I�����ClnW��C���ޑ99�9Y7��ݲn�5Fs�Yp�o��VV����ʮ?p�G`LCi�k�x�m�κW�:5q��/y/N���Vlv�4�������ER�f�$�v�SS���&
8C�fE%��ޑ5�]�zI��h���v��=2��W����px)���Bb�訨��gG�4̥��3]}hzt�/Ƞ8x����ӳ@�5��]��1y�@=��9��_֔��G��zL���Ë�E%�:��n��X\���C���y�����w5�@�9�Z\P��8Ä,Ey�lX�*gZ�ZS�s�o�-�*4�Q��k8\����(*�`�i�.�?� �����Wa����g�G*u&�P]�Ӡ��U̅��T]��^�Uqfv�4k�[��=���K�dZD�`��^����]T"`�0F�
y�'
0a�����Bm����̝��7�(� �ef���F͙��5��'(Aolk	�H�����_��!͝I3�{4�P�b���X�3�~�9T�_�0����sm�y'� �@_
�p�$�ۂA��!���?йFf5T/�^mږș 
�a�j�9m��'Oʽ�w���7�<�����믿f��$*AK��� L���"(a�n�	�ql8���ثP]�������ǲ��.[������ho3�C�\�
ܗ�]!�iB��xB08���rn��S[�R��e�WlC�j��Lp{�5����Uy��S-�u�Q�g`�d"
�Ar%y�4'�b��H���
{c��l�w�����(!(���}%�����#TZ"IF$���ї����T~��5@\�:w��6Ɉ�����H�a�e	��W/_�?��?I��?����E�/~6?;���Q�tY�a�6)��Q��yBG�xg�"�F1����Ci�򑕮�(��������*U6�)V�"V7��ْ(�lf�^bk�66�xd
��Z�|���Ng9����WA���7[�%u�/�(�T
�ʫWnay!�a���}��ʾ�F"ůyu�z�c˲��U��KAK�(`1f���f+�P買�ϱE�����z<�ȁ@�g�������������C6~��Ѯӽ�k�A�n�d�y�	��p�Ѱ���w���]���@��3�P��w�`�P��4y�a�O����=��"+��A�/�	G)�YP(�zW��O�c���<���C��@)|F6�&�1K�*9ä�/W=L*.o`�ጫ�pxt,/��^>zp�T���ߒw���g'����ݤNG����nTsr��1׬^'f7�#�	7�322hb%Bf�3T��:r�FJ(���M2 ������z��&�5�M� $g���8a���P߾A��\z8$Ⱥ����	�Y�*�M��6gj�h`��]P�툔����7v8H����̄�"F1Ԡś�o���������`N�yͦ�K-��p��@ZQ:�tD� A��s�
2��۷9�(?�Uα����[.���* I�,)�n$�����xݻw�Y��ڻ�&g��3� K�kywk���O<� i��葩� F�f8�tN?�_=zH�m��XA���ܛUΚ9�W����#�FN�^�5������${*�4���ݗ=uO���
d AP����d-�6�Qm���a�n�>A��FɈ׎@��ԙ��@��3*�ɵ����e�j�}9���v��GU�4�<��g&Ը���$��	p���^	HIS�;���T�������i`�,ck�i�!��2]S粮N�50��e"�*�_d�a�N�j�G\Ç'�� l3��z�m`�)�UD��E5�	�ce�8+`�؏�zs6O�=�p�|�Z�ڠ�pԡ�����}+Qܸ�oV��b/���g���/K7�ۻ0��Ί7��,�� Q	Qv������5���&DIǹQw(a66�C�7�n8�w�ޢv����_ɟ�����h\�����`��L�4�_@�}��l�w�c#ӫȇ)�I@Nܺu����ܾ}K��my��5�a�{d����W�T�X��{��~�R!��}f�B���:�����)�]���j�pU|��G!4x9��noe��D~\��FXU{
hx�D�ٓ�u����]KN
�y^n�_�r
��*᫯\I�;<���µ�+c�WD�:��Q2m~�|~���@=������\��C l��y��Q��	������W��W_�1��N����������O���0ϣOC�W49f!R.�[8+�|�Y%�v�Y�$
"%���;XBl9�**�U����յ��<R�Ƴ��S��\�"(���22x?i<OM��ba !F��$�vljY�R˧ a<ܻ����~���&B��@�>x|���lB.�WU���x3��� 4���JЁ����V�JX��29A��!~�K0��0՟����L�؋��<�fZy�2��JDЁ�`2��͟�{xNHاb��<{�T~�����{������!ˊ{�'Wd�p-hJDoĪ>1wwt��F�Z�5'})�~�OO�3��h�:^�|)?���Y��G��5���ß���{��nE�6�JҀ����Tl�G�T�#�\��郻r��m�������d��Ѭ��U=�ʜ�s
�Q�A7�K���oAx��F�;↉�J���X������97Rd ���]���
�&�}�.L3�A&����Ĩ�3>�(M���;7���l����޻����8��㈪�@��6=��"��AxU�*���}���)�XХ2��Fj��t�  �|�!kk�������;�k��N@;CaN���.[SY���^ǰY�N�"g����'� ����u�c�v-�ʶ����"�\������Yq,4���38~��{�}��k�~'���g64��b��<�mߍM��P���EY}��p��:_�q>� &�l�?�u�D��1�(���蘡��׵�����7dmq��β�Y"ڐ���&NwHR�}����⃘��çf��@���^8�	��� r�엹��@0�`���c��$�Q�M�;��� �Z,���Gp��J� Ɍ��V��q�w����	=�;8���V-�f��Gƒ�>"��uO2�]`<��l�D�'TFp|T����:��6���󷲹���h�t�*�^���u��dE�E�Ãcy�nS�W慀��Ym����#[�۬��{w�eХ<��H��J	5��o�oi3ɠ�l^NTC��?�ҁ������'쿈+ɹP�	;W�����D�{���Fki�s��M�� 鲽�G��8%c0h�g�h@�51�4=+s�[�U���	�,�����IK�^���9��9�rg��\�1ɁJ����9�b�	�H贘�O��)��������d6ynv��o��Mc�ce�FpK|��#O�#7	I�2q��H�a]�>1��P�{z�a4�'�T�$a���uT��d�*��Ή
��&,�(���Nq�ȡ�Q�wZC}��G��OBlG�v���>�'ᬞ���P�³��Y��r�]��
��ү�?���ȇ`��>b�6� v��|�Z��O^����~�;~��w��a	���CV���>�A,�V�z�������h��MNͷ��=]L5GLx�f=�l0	�]�>ʗp�&!�z�z��#�]jMgV���b&)B^N*)�x���7�D&�F1ieN���D�z��
Eo!a��*)�8lx-�d���EM��NN�km��@f�q��q�J�����_���J�?8�ʨ��\������B���Rm��S�Tʼ4������ُ�L��4v+��P�4#`�P��8p�ؐ�^
��9:C�#̑��U\sGxL��C��f#+���x�F%{d�{�
����_ӑ[�F~��q���79	LjO���Zw�Q�	�c��*�7[l����m���!!%�o���P�h���U�xA7�S·�Wz�x"\(�)��[o���Y�P��䴥d�*'��� n��w�N���ll����Yi�L���5Y�x-��3֧�0N6�2?�N�:{B )A H�8d�n�c?�@�,�%�ր ���$��ye�6+(ggG|�Q��W�@&�&�NkU�9��:$�z]������r*��у�y� rd�/p�;�Ʋ�NƔ��7 P7/K��:If�)��5'���
�e.OMq�rjn.-�54�[/Xά+�ؘz�LLZ��U8hj�_`�	�W@jd�1]�zEL����J�5c�ʦ�'���G4��|B�M����؎�rg���yє�n�	��_�s�[��#��s}Z��f�W�
�z�g�����C]��b,jp�zs�ٮD�6�^�P2�q.�޽�#���#}ϊnJ��}�dD�fp���C)��?��c:��/x�z�jzo��-8B� �[{�r������A/#��@��q�~�$u�D�R�a�t���Y�AR�Zb���=�����g.?z�)�f� ���g��n��2� '�"MO�F����+
�z�f]>~�1�qW���h�ͱ�Y�8<9��4v��%[�V�M�	�~w�j��a�7Y��#�9�8����Sq��t�QӒ"N�
8uZ}!`�:�^����pA1;Սv��LD��M����tn=aX�ޘ��3��
b�UB��W��ȭ[w%����S�\/�z@򱳳�5V�4*����|��3�a�wc�Ӎ��s�b�(�zFf/��0�zd����q�M���Ů����da���,쑀� 9S�MPh�]Y�5����p��*j�� [��K3�އ�^s���R&˶��䍎���x<u��冬,a���ʊ�q3쏱*�0�A�f�R��܂H�_�	����UnGf���M��?�sƪsV0����k�E8\��*W���eP��"��	 B��o�c��:���x�q <B�\#��|8�7z�J���p�i"�S7�/S��I���,�Wο��˟������z\��������ݽGqr��%�s��x�@��lX���oh�@���2Q����_b�H�(��g��޽�_�V�4o��~��9��r�����6��؈���FR7jD�0ӛ�X�L�Lh��?�͂�Bf��`,�d�-
Ydm�m���TF�L	� N0�.gZ1:�0� �(Jo�m���K1ʧ2k5= q�3ˮ��,���՛i�\[����|"��G��ձ�+yx�yA{yV �O��Q Qrk|�.�7
$m��1@B?�T�Ǌ������$��.��_Y)ٱ�V�[�y��C��W�?T��:����Dꭆ�f玏���@�׾:��!3����M5�m�z�Paa�*B�&��@��0#t����uA�Ѝk���Q(	5�w� ^z��9Nz���5d<�-�ˏ�e���6�ne��I�Fی{Čg�N@-эx[ޭ/������+���*��ܑ��]5�wuc-+�K�k�Q)^�� �8�uo�\�uN#��A�C8��?���P��Q�ci��A{C7�C�4,���]����E���6]�V��к���ʌ��6Bӻn��{_���&6u����x�9����k�n@pLh�3�:�7���f3���6̧ɩLz�a��:=.>�傎�Y�
���l����7IV�%&��o�̆��C�JAp�x0r! ��+!�T����(7���uw�H��s�a>�������w�<��y����ybA2�Gi{�[
��Jظ.�ۛ[�V���н 9�5�_1�-=&*�r��577�'�]��5$��9c�����c-���릮��=#�;�z�	���	.8����}�YA3d��4jQ�nB1���;!�a\�t��?���[���Dܹ'�t,�����������(��h���k͖gNSn}��,��e!����ʱ�]����(��w��� ���e��%8ఙ�EC]��=�q\zp��#���'0�#*�cVMuʹ�t Պ
�9�	�+�8^�����T-
z^$x��)�a�i��N; ��o���51�M�d ޅ5m��H���.2S�o��F�G�#T@q���ޣ�OG�������:C��ו��=�Dn"��S;Q��>���z�M`]7kP(Ge2�9xF���S~�Kk��O.en�3�.§R<����Onq,�(!�J��W��Ͽ�\}�I��W���+G''�^Alm���ޠ�Ȟ�x��{���, ZX�[�^��C��Ǐ������M�|GQ�+�d�J|?�����p�8��ϗ{l��8T1M3qa̤�.V�
#7�SՈaR͟�E�6Da�_B��0*�q��I�\z�?Y&\����ڍ�2�t�z}xX%5�u%�3ȗl��	=�k����j�q�9�>��}��Ǉ���1�X��a��|�٧�ɧ��7_?g#:�T��@���t@	[ (P�裏�����ſ֍iО�Q�}�F2-#��h�$��Y��2��D� ��ט)�v�	�2È�����^kH�261�N������\�1ɼI�����f��(��P4�O h@c�S����ϒ��n�O
�0c�Ƌ>  ̴����u!���5�T-P�����eG⺲������J��	�ϥ�9�1��.ʒ�R��H��l0V*C�RY�����-ֱFB`=�d�c0��E͡E��^��E��w..$��r�ⷌJ9��a����1�>�N-�����wn�0b����%u*��^Z�!���\���ᜡ8�n�Xa��6UpI������ձmΏl�����~P\����!�`��4	2�`�8�;�Ef��0_Z7�˰\��2*l���l��;;��e�Ƭ^�M�s��t������|zt¾�VA�h͌��pX�=Ap(�W w�^��36a���!go�@=~(ܓ��o��W'�U�N���T�&�L+���^�����)A�C��g/�H:+A�V�x�7�蜜�Æ�B��[46��ekL_��4��6�w:r���� �*��dj B%g]KIM�5���^���&
h:��6$F���<p��Ep{+z�(��?;9"��y�*]�b-��A Ϡ�%������S�N������z�����,)�~�2� ��i�逮�&�`�6��~߿s���A#�����q-B�֣D��-�@�x�-�Ǆ'	Oe&�aO��P}D�9P��:��L�#V'Z�	�CH/�*�85V��٬�Ȋ��w2�f�
Bc)�nTN�Fܹ{�W��>��O���5#T�kP�������[9<��~v"
�e�KC�1�E�����-`���6�s V���sN���Kj�rp������H�j�W��'�c]k�=ɕ3{]��Ās���T�΁�st*� �#�h��賚��RoYV/��Ơ�[5�����!��
.�}���@z�ߏޖ	=^�iBc a[�L�"��NZ��De���? �%\s�y_P���!��Fm�	�z����bT��v�D<�c�(������~�P�X#�"���Bufl�~�o�@�|1���|����=�Շ8���:�g�f��������B�b�D�9Vo��1�$pL���]k@tD����hy�Å}*0���u��֎�#���{��?&I���㎷�/ye��,��i%��Cd¨ޠ��0��/��l]��*��Ā���>nY���a�a��K���h� $���-��.�<*�Y=��z��Yq���/���,�k�~�8�.�~�������<�,��������a���W~|��8���%����
(��VHx����;�w��nll�ɱ���@e��&���ݻ��W��������=�Óȿk�&��uO�q�e9��t�uS+�����FQT�J@2���a)�'𘥰���R^<���`Vac�=�C���C㒴���u��hx&O��J�E>�#�\�I�|�����c
\�9D�Ԁ �13M�y�'�* e�	���]�۪H?���h���B�{,�]�#1��1:X�-F��fQ�,�/vV��N5�1hX��`&�ŋJ��\�Iټ?��'l�x�8�x�@�����;�8��~�(������. {M�L��:��������9~�m,+:ٗШ���Ƭ�o8�B���	� 0ݰ���Y莞�����7��>7���sCT��5�0a߇�Ț�ڐT���ӓ���bj���jG	Ǻ�8�����ٻ�N�bW�������:Xл�_ܓݭ]k�������ր�+� u/dˁC���,7eJ�w_��ƞ��=0��� hCed k��t̲,<1�c����QQ
�	��i�x�{��ݞ�Bv�m�|D� �J�u�,��� ��$�66v�!{]c��{z���k��i��p���b��\�@:����K�i|��P٪A�8)��(�j*P����$F�y�`�xƭ��¬�%_j��CO�9ԩ��z�I���M�Ғy���&8m�H}����7�� ۄ��g5RĦ>F�'�#������̌�c�����38���a�w�ұAcz����lb.��Eux�>7�����r�W ��Ϟ�`-�7�l�(Od�@�*��g�3�������E�y�ޗ��P�ǅ��@�
c��[���*�L>��3���/dj~�6|N��$[z={�,n�n�yp��!�܃N�'�>$���]v4{���)�<9;�Hf�qg�cT�$?�-��pG0��⎑y�Ԃ�[�zD@c�
&��˿�@�R�A0 x��Gz�f���a47��8lL�W�M��!hvAMlb�	ѧrsaY���F2�������ԫ!7FG47!2 ��*Y���ܵ��%Ȭ��+՚��ǁ�é�©G�y:D�f�әO	%����lLK��|�e��D�]�_V�0��Ե����԰zwTm�yv��k׽��-��`��a�k5�>M�sv~�����gC���Ao-��������d 'G�$~0��(��.#����#ڇ;w�꾰!�N�J�Zv��	����>;��[=v���[�:U��.�	�[��I;��P�:s�@2��A��)��}g���$�wU߳�w��?~\x5ΠJ&�@����L�֤�Ax�I#��0zu����1�üX���

�F���.;���\�U+"W^�������=��ޓ�H�-5�/���ٳ���u:���m�����b�ԯ��q'��G�{7'�Z��,-���&m>�c8���mѯ�����p�ͦgsk��@���*�GP"7��
OP.E�!q!���@�Ӡ	Y��2��"f�G���F��EF���������� ��h~�P]�ګ���*���V�Q��J�q����&����B���)��K�����T���/��7.:T<�t0m3��i�w<�RkjBHQ��~���,���z|,�?�X�ƥNv+d��9�2�-f�M��MҀ�Y�� ,��q��1��Q��F���/euy���۝��9"Hdp�p�v�Fց�6�GegkG�7�^�"�"{0��:�A���4�lQ@'�ẖ�W�OBD���u��Y�=���K�����?��lLP!��GO�y�w 74h�p4�Cͼ�NЄ�-��c���)�
P���#f,qϞ<}B��:k�3�ԸɌ���	���3�[�c�ileeA�Ed(�e�V1^��=�K��&�� �KP��#��J��C6̙@&*��5���`��< �f�:��zq�a����-ǧG�뭭��kY`�~o߲�����֙@\N�&8?����%F�A2���3�o%��m��K��ō��ylQ	>g��Ճ�{� ���5�Dd��]��
wet����~��`�s�sÊ���!��ɓ'�~�8��_�:vO@tx���Poɉ�kc������`�����r��]�#�(�V#gp�i���5_^Y�9?%�v��0��E5�飇t�m}��;���WR+\;f�y�[@�Ƅ��N�Զ�R$])�����^j4�UG�L����:�S��E�ʽ{��?��ܺ{On����uvf�	�_����^��z�k�vP�01�g��A7�`��Ni{c
(�,�c����+p��b`Lh' 2"f��S�{��L�b-����HE*ڌ����.�`{F?�#�sg��cS*�G,�;/*:�`��7 �p6SW���nK�gA:�?��^��S�x��U��D�㹳)�!+���|�H�Օq)�9�ϧi��l8�FŋyG�P,E`S:m�7k�G���P%_� �*����Y�X�<�k:8<%d.�ۼ(Ҩ�Y��.[�W���$�N�,�IHN�:�'�� =�o~�����4`_�1h��Lnv�x�p�aO�PXQ׹����1r�%H�`Nb^����	f�s��S8A�0w"c��\ף�d�M8�3�.�A�ō*S;<Рg�,}�.TT����>@�C��8&�b��bb��9�mc޸_e���j�(��ܸT��ʻ6�ܒ���9�ލRK��O$�Xsn�Y\F��Ps�u,��k��K��ܹp^�5��p8����!1���}�V�zq�5���ҟlI+T�[$U��+2��5�R�m��Z-o��ޚDͿ��m[�Q�<Z�"#1���:�l.����<�O��TA�&;�^�z���1���#\|�P���(���4Bm�� '�<S5F���2� `^�5��by�\ �;���v1�2R����&̪��K����Y-P(V�A")q�bT��c�����VZ�]��6L����*�C�X���~&�b��Ɇ���=
F����	*�����@.�ޣ�chY�w;���5�^�ТYM�pv�Q�ղ��m׎5�<5B�j~�sp� ��g����o��sh�4H�s`g�id��x!x�}����	�x��32��5�	��3�#6Z��!���So'h]���ɲ^Θp�$�[���<	�5�<��T�+��nEd�ͺi�Ë�4&����6%Ŭ:o7j<�y�MMKk�&'z�{;;:�Cۈ�b�!� M�ج��&�y������щ�����7/d{gK�ET�,,��ّbxj�aCַ^ؠP}B��	����>����g�w�1�6s��qH�6?^�fҋ�M9�3���Ǐ�z��C�5P��yxDT��4Pb�$�0��]@�>��E��l���.�����0���-�}�!���QA�^"`E���Z�p| OD�gh�̚Z�P�Y]��@�T¼")����>b�S�U�P�������=�����k���8���>�p݃(�ƞ4b�G�2�p��������D��_�{���uN�	`�u:rC����M���G�^�ZD�T;z�?y�P~�_����|�շ���;�G���ˊE�����&	z�fdi���e�38���3;Xcy�ʜ��)�B���i`����D:���y�3-.,��%7WorN@�U����Ͼ|����o��	e���r��\������X��@Ȃ,plz�o��XR+�����T�O���G{�?J�s ����!+����DB�Ǿ�!�}m�o���ʇc�I�q�� �q�I
]�+�1n�`=\{Wǫ5��9k�p�iT��3x3��ƬΛ�=�. ?E����6�N�a0^&'S#l`���raW�����]� 91��Jű�Y�:A���&�X7h�°S���D�L�`_B��g��f��7�+��<@�c��I<�F�ln�>	��0S C�(�ʡ�3�!�cÚE�o~~N�{7��[��s��^8�;g#��&����2�-V3  ����~˱- J�e?�v$q	����ǱUsXQ{ݩ_��%�5����4S���gȈ�8�;ĺ�Jҵ������>]X�OX���?#���ҧ_HLc�
��������^7�?u`>*NH�a��L[�H�Z-���K�
�/��"y�3�֏��zTB?���QH�A��ԂG� ��$�"�9|�8��>�#��F�֐��z�U')/Nޜ{8p�^�θUZBȕ��"����ȅ��Z�Χg�3�q���-$cj`
��S9�� t�+0�e�*N���-�0���iA�e_GcWt��2lr�!��"0��iQ���p, ѩ �@���Y�R%/6�����\4dsq�$�,��oq/���	m�y9ř�
�+��lP�*�(K����9?�3���q�.q�}����S�:���Yr���h�F�Ih��Eu,�@�*��s�)�}.�Ji�hT��!;ZQ�sd�t#�VG�nm� �d�{�:�S�Ι
�'粻�Gy"0��!�g�8G:�ͦ5'7�hbNGL��1�x�ケ�Ӂ�C�QwZ%�T8xϊ�\���_�y@�F��N+0����we'ٖ�FK�j0�k��&�˷���;2�Z����aQ�2CV"��-u21�q-w�ޓ[��︡���ҩn΋d� �׽�~
������͛�d�B�-�L����$������pWi�"Q/ʽ(�x�T5x��ވ��.�K�
�� �M0q���ɝ��ess����To���2�������񨰉Ev���B�4̓�*m!59�Z9�!Xt~XFt����o�I��A��T��MR w���P(��L�!1�G�B�V��e��È���}ڪ� b����Z�J��dxr>�{#� �������ѝ��|���
X�=x@x���,i��fu�A�poW��g��~��]�_Z�p!��թ�� q��g��G��'O��@��[T8��� H�żh��|��y�:���F!n
���AnMD|�́x��'��(j��
��s  ��IDAT�PԵ�x"�}�F^�y+�^�� ��0/}�Y�--�C��=ſÒI���I���_���k���F�j�;^;*�ye��=��!�_��ˊ>�o�f� !���JR�0���p�~����*C���2D.J
�)88z� ��9��D����X�91�"�y�"c`Z4X2����obu�a�d`���^���˾αÃ������>��3!v_0g&�wf}�i�b��VZ����a�[�an�\C2@L%��M�S��RI��uVRFtN1V�[!�'	�������^�E�k+���C��7Y�E ������O�!��Qٳ�,s#&8�����.�!�vH����Q�L]�� /���7���޵��� )���������Q؟𞫚"!P�Ԩ�OW̓0�y	�)�yqL��L��>i��I=�l*I�1��D�Kǯ�8��� 4yl�_�R��w8:<��uj23f�z��H^�f���%$����y���Fnu}+@^�`�����_5�c��@�I��fH�
>�H�o�Q����|2����+����LA^�%� ���
g�6]*�V2B!�3�$���CI�!�%\��!)�.ʳq��gT�KXL���GT�'���Y�A@0b���D�lX�O��X��߫�X �Yw��V��~�, i�w�7�,U+��*X�B)7�OEȌՌ�ƈR�f���m�a���[F��@9�y��힕���r>�(�~��bS�`�Ƞ*.l���g��p�z������D�'�o��zd�Bl0:W�}
M��v[~'���8�'&��"��O���'���[��ۖ+٢<(�Mf�B�;��\)���G�.�F0&�
��c�b�\F9�	�`C��Ǳ8,bjMSW�x�A/ʋ{��cT�v�2&���wZ�Y�A��c
����l�]�ذ��]� sݾ��缞��6I#HT-qzS7M�ZB0�*4Ȣ��
�X7չ;�`�"i�����V\#8�A�:;;Mb�����٨wL�G��Lqt���-بy��(T�rhdoХ� ��N�QD�-6�{�������d���͛u(wL��c0���⢫v�L&�&(�u��B�f��� a�A=�4g �_ 5@5��NSl�����[&\����͢�KRG�"]���Ŗe�śt�N��s%�1��Us'����D�O�y��  	�[�j0���{��ˎ�*�t�qao�4�8��OE�#,��������tu^�vv��hб��(�`�c�7V�#�gaW�NW�㱮������� Ջ���jc�*嫫��"���޷/�c�*C�StL���sJ.0@fձ���2h��a籡���gs��:pf͡�ҧ_��n�]c����Ρ<�J648C�$�,� '�
yG�J�Mʠ$�":$���u�!�B��^!�zsGǬz�&���@��l3(΄� u�w��QY�Z&����6N��D�lcg'�+g]�W���;�uܵY��;K�bL�b���:�����[G�eT�@��=ع�L�ڳ��O�ޕ�{�q��Ŧ��>%�l<ؓ���m߮$'>BV���4!�l�j���熆r�� ��M$̈́�)'�@�-���䝊W%�ⶈ��l�%��@��x���w���c�B��pw����?F@>��S2=}���ߨ ��pb��(�I���Yva8xu���������n|j���o�D������=����/·Ik�Nd��]�x��1��d��y���#��^�zWgw�� �$�������s_"3�J�|��č�|W�s���I�	�7Us=��B�j����2�������{H�i`d<��3�[�sΐ)e��<l\���z���B��w\�Ir�oz5�	�.@�*�"IV�(��@[���9o=��z�����ۏʿ����m=��yP	�̌E�Í5��c��q�\�l��j�cQ�1i^6�[`�}
��:�+x=�&������:ߠB�,.�4�0O�AȨ���_�Y"s�)h�]ݕt)"V�Q7�,}�||�ْ��(e�"k�[�R7F�<�%+XyД:�}&AO!� F*���^B���WS�͏��*�����6 ���w�U�I�y�~$��T��"��?�dHr��d���A�D&�[�ZubT������F|���7� �����=g�]u���!#D�8�B���Z�Th�i
��? l1�p�����i$ȼ�<�m�s)�Q��	��0V�p�X4l�1~}&!��C��8�
��"Yz_�D�t����6U��z��֫��vt|&��ܿ�&7���������*�!X�Р�8q8d2��ׂcܹ�J�.�G����\g%Ÿ���Njp���h`��^i@֌�"P�k6#�󢒆go8"K?�,�}�0����rcqM>��!?�}<_����6vd�1��<P<E�D����!M�,di��n��X�M�ؤ^y��du�A����y�IdNp�r��M�pB0��#"�A��9�`��Q�����ܽwO��9y�浜��@�4Y�@���F��������YT�u�Z���D�?`y�+�>
�*�#�A?��>w��GO��ֱx9���?8��Mn���{Z�yS���o3�/^��ZA�wmو!���P�LK�����p �m`q~^n��2�l�k~Q�:�Y.H$����g��{�gL�����5*B�YT�vv��|��/'�B���q�rK��Ş,(�܈���>Hkx�*5�l@.P3Y3���n���_vg|���K!������U����F\�B��[��V/:g2蝗��q�-Y��3a_$*G3z>mVX�n������?`�B��P�l	�'t[��	&�
���F-�]�.�u$�#R�?�m�͚�3fH�x�C�Ɵ�s?:�"X�	�6:@�"�>�.Ae���"$">��uJ�&���w�E<F���a���3|)q�30b#;�ͅ	�LKv7FC}��)��a�/�����7�k�޽�r��������=�[ռȃ�b���l,�Yj��8$HrB�L{�H$��B�͕������L��w�潶�}6�=�l6���ز�"&h]פ���w�}����W+eu�Xh�/J���e���9ʢ���gx9;Fc��X�Y�(�A�Q��Xr��$�>��[�n���/F��tE�r�����@���k+�N��ß+?_�y��xR ��v�{�s���������>ң�R��?�/�y^,srC� T<C a��Wo�|U�a1�r˂7"��*�"�_�����}%��ġ�bȐ[1�����o�

��<;N���^��PxolGd� �#��m��(�eq-+Jj��f�Ь�����O������JT,���a��+60<�W�q�*Fb�`��e�b�����j���{5��8>��{8j�wԧ7�9�g
CE7
V��=6�ed��2{!^���E���ӗ����)�1<%��FdF1x��=ՙ(:Pǣ��{��؀e@������)&Uj� �B���4�P�3Xd�@��p̒7y�k\��M���������c�7�5�;̵4	%��F����#*�N��P߳3un�b�iǫ2�4'�˳t��csѕ���3y:�Ǐ~� �v08�p�q_R�7Jt�Ù8g��=�2r�`���NЇ��9�$�.�t��b���8�[H�� 6�c��zi�Ð����aΡ��E�#`@`3$�'��ܽ%+k������3����eokǠV��N�T4Z�.nW,ǹtS��F��S�5�8Jx��D\��"{yv~����ޟ��M�
���tB́qᏜ('��9Q�X֚�P��fN[\��3 �9p�s��x=�d�˾�G4L�onPO��RbduƸw:�ш<�рv��A��k��Q.bu4㤚�� <�h�!z���k+,��cF����.+��`Bz}!�z.�G0�G29� u��������O���ǲ~~N�iuhf�gY!C�Zs����e�:=h�J�HV�<P:�1��̬!�}x|�
��*f ��?�n'����â"1GS<�kϰw��D�����,����'�\4E�'^ݡ�����XQ+�ݲ��R���
��R�f�*�:I���K�EO	�/1�A�U�o�0��@�!څуQ�;B���jT'���>[���)i��|H{�����u�2 vD���&t'������<K��߉�����^��%-�q̑DA��k89=Թ8�����P5=���	�Tk�G#4t�`_��n�"q�1B��lХ���T�k�z�<+��%���v�/��l
٢�I�� ��*-�0�-$� 	٦
=�c]7͉�N�w8����yǂ�`g;�9!a8s��b ��V�O�N���<���6�WPNq/,�s��R9<��pVK�M���4���a�S#�{&&��� i���|/�G`������c!iz�#�1�곺o�o���8l��*���GA��.~G���֏ӈ�4�!8̠�ž���ʗ�ʎ�/{�{�#cILX�cŪ�~]�p��C�Ձ\��_���&��<~H�ᇪ z����k�i�c'b
~*�K���?|Tɺ�{��#���Ɨ�^L=|T���i��翄RI����`�1ٚ�"�M�l���Ư|�{���{�F��?��`�[p�jHџ�gݡZ1�c�$d�O���8p�{��8�,^�)6�V�STE�|y��z�	|��D�`�AT��ZTi*�e�w��XT�������C�r���	Z8�C:}�z��dA�$�7���`���^��b�|*\�7�Fy��ܛ��t���MM�"��A4���\g@0k���d<%wn��ӏ�0ӊl*'�g��c���O8��#���%[���}��Jh���6`PK�z����'���{ݫ1uuز.�+���Y��Pc׃"9��
v���)Y�_�)jgg�;s.](R��N����h^Lͫ���)4�6u�fB�C��̌���3��Z'�
Yu6�/Xcz�1y�[�5��6W�qg�W�.�� �M��Ej\�r}8<T�'��z� /@33�	qo �P��ҍ�.�K��������|�v]����2�����<����#kX/��0��������|���p���wt�w0_�)79M�𘉄�Yê.p��;��Ed�h�i`{�1��U�}�Gi���n�|?f6���o�{�l+�q�~y�����k��������p�n,Ȩa�yX���d���k
�v/���462B���q�v�!�N>Q�����`vFo�$$�՛�t^����?:�@���6�N�(G��G��\C��w'�o��|n ���KdQE�J�I­t��j���@/a�1IM8��2U�߇{:N�v��c�9�G������d�
6(w8��M�1V����K5/
Q�D�v��%�*�'�tl���ҁ��U���5`�BMH츂�ȸL����n���YhT�r�G>���3�&�� 7�ƅOW�M�p��$�6R&6
��1��л2vf$��0���DoA^$�ҒH!7� D	A
��ᰫV騛�8���2�
6*���H� �7-���"�L}r��GT�� ��Y��)��F��Cz����Q����\w��ґ��"^2��K:f��t����CF
�s������]�Q��	��[����-�fqdd2 �ނD�6��I�grcX˝�|L�s$1���5�G^e�߽�_�^B���8*�Rm#��)z��&0=ٶ�>|�w�*ש���6Z����F�;���2�.�_@��Z9	�m;�{U���C�X��Z�Z�M��0g��f�Qa�I+����̝����KR��yR#6��7��@����Y�+��/��W���Se.�N�d�s����޼y������ ���j�-Y��c�lɎ,1��#Rkq���[( �k�79ӿ����F��1�>�m4kt7� ��Z������Z�#N�md�Y7�9;���|�������߫7�ʝ�`b�8��f^�l�`4��d$2;.���y� �<󛹶z��H�жf*#�&X��AĦi�x��`��+Sɬ���=�,�:�s^j��٪Ҍk�l	zB�@)3_��̚qq���B���Ѩ�n�ۨlq�1�^>5%�ک"v�P�?oƯ���l���P,�v�p⠊5��p��c�ah�J�1����������[9�����m0y�$�u�ƽ[㶁���en�53=�W����& *Ӡ��� ��O~�����5�;q�KfIӯ�_���s�\�+;��q������	� ����s���c,)^z�}i��	hYY��r��St!i~���M(c�z7�ra_���P���P1��۲��*�v��zztD*��hR_���'��49>���f6�]Tp��gpqc�H�^�����֚��-�P\\豯�:8����9���t���*�N/k_��W�� <_��@���^Ϛ�q0��o�q�����ۗt�]q}��s���V��.�e��P�$^��n�Y���c˚�����U��5�s����|2.ŋ`��u�Vr�L.%�^��BIM� �c s�b�:������<��'�t��=�N�>�L�y^眎�ue��P6;�w_��ޡ���>{T��{cVM�&�$`4	j�bf�����<@���<�9r�A���?ܗ�>"�=��u@%Ҭ��y ��zY��e8��+�G�g�?TF`1�}��ᣋuH2�a���PY0T�s�9aw�ì7��M�v()9LZ�.��@���� 6O�h`�+����;�j���x��y�yO	� �zh��z��PͰ ��
�L]p��mw&j0�'΀'E��[�ns�ľ6vF]{��ߔ��A��~^�^sC?�<H��k��̍�Rs��#��}tIuj^L�w�t�RB��I�S��T=�R�_�˵��A���5���+�(��f���9���m��S�Տ��ƀ��k�+r��C&@��A-@8��'݋����Yre~��=���ꄄ�&���߃���z�{������z��6q�Ǫ�Y�����S1���2���م<�{ہ�\��s�3x�\P�l{{C��~�X;Q�qĺ����
��(42��޿�c��?`�Q�^^Y�E���<��(^�i�7~[X_ k��I�
��4p�C�qQ���u�<S��S����T�4U��+"k�����N<V�A�8.����|���q���NK�+&�8���')�c��Z.��D��	�	|k�{4Z*晉�@	��tr~:��N�It��V$����|��oֈ\܌볬��ac�^c�5�5uuUɲ߽|��������������>�c�B�������k�ҒK�Q���˘|{kƶ��JP��+ۺpD��`tJG�g��RZ�pI���Vyc��u��RS�D\<$~d#L&$�Y)Mk�6�w���xm�]t8��N�@��!�A��S.�L6��r���7��<n���˔���X,8������ė%�m��ʗ1JjFBa.s8<;�l�65	��{-4LߏI��e2��9�����նF��^�2�e2�D��OU�&f�m}v@�*^���2�6��j�+�X��-�
4�;���s�L���m0�K�7,�3{�a�_�Tu�w[*f���؜P sY�5&�����l��>7o��D�#���C--�F�ڟ�d�8�"� ���as���,@I���խ�Ջr���ݳ��<_��� @ܿ�B�g PkN�.��ڀeG<0Gc\���g<l�#+zС�|mu�Ѽ������\�LR?��u/�f�Rw'%�Y-h C��{@F����7�U�N�mqp(/߿�����^ʹ��[krW��?fc����*aYhi=�yq��:�?V=zݔыM���u@����
�}���`���ύҠ�[�����ꢬn,3�1�\IG�`޵<����~)|�{��\��p4ӗ͹�g�T�W/^��ꆬ-Z��ǟ���}؟�#sE���RA�˸��3���͛W�L�ʔ`�>(���[�������ڪ,,-˽tO6}~�.�V�*��!�ycT4�B���]�h�{过%#E����I�A���A���5?��M����+Le�e�Fn,�rYaM¯g�c
?�B<�����z�ɂ��c�|iA-��� � l ���8Gc+��2R
!���vυZXe�
��I���V;����hm�Pҫ��Č7σ�)�CV�`�HTV����*O�Y��dC{ �n�vż�����Yp��[��w��@��EE����I��@�x{˪<�{*�"X���v��� {�X�'������s����=���+�@���sK����5T�0PqBc<�)ì��LLLl��"�wkt
bu�Cn���7��Lhቴ���@����T��u@��-��.�{8ꐺY����-�X_��7E��}8Ԅ�i�^[5�JP�؇�3^Y/_�b�#0 �4��Ɓ'^�=�R%�K����ح��ӝ��]�yj]5���f����E�z�h�܄W?�.^�Қ	�~x0��fO�V7dZwA��Z �s-�9�YO��-��W'т1cA�/����Ll4�>R)q]q�Kgs�G܈�ъ������Ӎ��@2�lF~t�k���W ��]�؏[Ռ���k�o��2+BT7㘵^��M��`���������?���������y����&����{�wd��@�P�"�.���w(g�QKR3Z���h�d�#"�.�Ǣ�ҕ=�%���Е��F�m�[��~;לי]��q��M�D�ULnk&�{>*�4<����������B9�WC��=J��x6/w��� "˧(
���L3Nc�b��vqP�g���m(����� p2u�&�ˤ2��,�揺��=qm&�;�� )R�Q�e~�����P||�7�էofn�8�����:px�nάއ�r��#��Z�	�3KH��Jd�R��zr< ��,$$xM}�$z��VRJ�j���-|�Tz�|D0`��V��uooޒ��<��k�'�M	_f�H[Ib;��g꺽��&��#0_�d@JwYA���ٹu�����=Ԁ�\O�|�=2Sy�YOA�2���-^��DU|=�X��'�,��5iLPʆh߽}G������H����@4(�CR;�Y�A�� `0w�HPK�3�L��P�1s��r���=���_��,�ݻ���>e���ǃf��0���aUgu�6q�]��\J��'��a>���t��US�Z]Y��#��V���h��`O��� ##�8jL��0,���PQ�
�
���go�Q�C\8� ��|�*99<������m�h��ͫ������Yу���o�PӍCM!i�vf"�NE �D.:LǞ0�B��ө�n
�*>�	��N/���{���Y�ܤ�7���}��ý�*�Y 3O�����T�u�0�=}�!��s6���{�&]T:@�P�� ��6�$2�����9��{�g��ʅN$��{��~<Ifƭ�$���*ɹ��\ㄽ9�u�l���)��I�R�l���������'�	"�)��TNP������r?�+*|]�ʦ���2=�(���杝MS��T�:�@�����M4��lfG�	�ԧ�Pq� ��!���Y��0�� ��}��/�:�@�Y b��c���Ԙ&�A��>}��}i�	�+����A" �3Ǥ��8�c��U
�k
n�z���Z�Og^KgQ縮��+��\��>^)b�&ne�q�u��7�26�Èk���HB���dj"+��U�Ћ���.?z�>E \��`L ߏ}s��K���g^��E�P�|~ЃF��ֲ륟#M�#��"�.����M��2U��ET��T��|�
g��0Q�̟�zUr��ٗā�&�k���̞�i3����	$k�2��_\�-v6��r/y��M��8�1�f��*c�^I����l���D�ITV�(���t(� ������ �y�6hY<��~���M�4��*T����KM�׊D��S�������_�~�����)�+}�s�%��ຩ~��Li�lx�([�xf3���ڑ��zL<O��*8�b��1�sd����*K
W�H|p�d� 7_�g�r=3�uK5*����a��{A<��^K�(������ ;�k8�ޤ�wZ���Uތ��E4��)6M.��H�����T�9��*��&C�מU4GY������k��F_c�T��lb��� �G�b,]�7����42-�OT���l���} `0&�M��/�)�C�ڌ��)���8d�p�;;l����l�+n>G���9�t��Cw^S��C��[�����×/l>#�^�5�{[�P������o���rꔝ����+��n6�mdc�)��`���;zms�Kr��=�R��|� ٸ7oeo�X^�x�`���;�y������n�����C�V��ƥ�ή�]������݆����GǬ��Nbj7u�Ɓ�xߠ2!�*"�&�^�C���`0*�\��5)hp������J��Sg��k ?�}����g
Fr�������*m�ⲓ�:(+����WRH{�]���!���p}^Y]�-��3C��o�S�smcm�c�J�p�ȍ{04��@,�,i����&oT�>{�B�m{��ө��A� �}i��ར����f�U�Bq�[��x��l��_����1�X�^AG���@��	ܑ��7�7���ٷ��E%��ĜN �����7��ϧϞ����	bX��7@
�!��p�����޾��sB:b���l?{�>3Ȅ�ɜ�L���^��jVШ�k���a��BW)�U�=Q�jd�~��^�2�V_�4q
����O��5@>�_RՐL�LS��duj�_dTc�c��^���4U��3�K51%Ş�
���h�O����:^_͡}*a��)eO����y���!٘�{7������A�	�^%T��:�+��:S�p���5�<�T�@Bo���L���e��Ѩ�ߠw||�c��������+��o��+TpG���	� X�l�o�s�?8� �
b$O Fp�Q@A	��@3�����i�c��Z�T����({Ĺ+�-�n������P�Ǳ�g��*(����tћ�I�e��˺W_���q�Β]��' <��aｼ8�}#	���)���� 8����뾣�g�iC�濿�ϸ=�^�����K�>X!�=�_��듉%������y�E�9)��3�� 6O	�©��-6K:7�|���@%�{��[���d�$��e�#��&U�Ր� �Z�w���U�Y��=�d���W���o�E��� �a@2����ǁ���X�#��VP��y`���6�������/W��F˲ף�\e����Z����?��W���/�(�@D�\\�*J�]k�jC��ŞNB�e���\BR�zeRx�R����Yxr;vx��<�h��.��t?K�%��L��I�B�G����I�k��2�����M���#OME���:���F��u��mM��ҳ]t���g�u*Ss^��D����!]�����H��vT�d�L���WE���8�'�Pe�80�M&� iR5�&fpwC%�2"��`��F�U��y�k3^�X��=��@�����k��c��-�S���l��	GY�M�pES�)�
?��,��^3�>���=ݾ���*+�t�����qI��qpC�	�v�l�
Cx��XEýdyz��/֮8�'�"V��b���@�6��)'L:3� ������:V�67dc{G�{N�0	�<�zP�9<<�?|����[rO�tA�ZS��w�G0����_0�a�Ol�8����hg�3�����Z����ף���k+9�IE�\�I�_�������P-u��sƁ��[r��=��O~.��ܗ��M��_�J���[Z�غ�93�a�����&z�z�o@ү�Ȓ���dCr�!� `�^�
m���wP��v��"�= ��/![�s[��N/L,u~+&;��t��>��NN��>(% !�޾���A��A�I�rb��� ���7?���dcg[>�ɏD0�9^PD�T�:��{G&�@����dU��PTz��U2��s_�����␤y�����,%ĺ�J��`"KD�HtOc�.��t��J�ju������:��4���{��,,/Z����lw^��p@n����R��Kբ	�\,�&��hG�{�e��1�\�Oa?�
W�c�f��YɟZt�
r�$��i6ȳɮ�&������9`n�W�<R�o:�^ХB�y4q�x@��:z=0�XY���N���ɤ.���Č_-�6�k0�޶|vKJ��C6�#��5 � ��k��������ť9ʠ�ZsxEe�pq��+�����  \�F��~��������J@��+�I@}�k�Y��� =�H��9 ⩨�V :�fr���LA%�s&�L��.� 7��(}� �jn�W�S���ށܿ������|�-�h�N���ٳ��W�9	`���������{E�u�����:o&�b�����wG�����P��~T�$�v�`l�u� 7�����iT9S���3�L��F�Գb�,����E�V�I|f~�����|+��d��מ�N��A#�K�k���Aѷ�Fq��2�H@U�4����rV�iX������0����w !  &w�(��-�3	ˠ�\o����F�����|�hiHD����n>�����߆F�#���^�}�&C<N ��?��/�����_���P�����:�Q���R6��BƘ��Dq������*��Q|k���<Q뾡&���t*d�"��`?������k��(�ŀ��Ѷ�5ՙ��G3f�dj}����DTC��#A+��=jI��W|PB/�\��(���?����,�<�v�WS�2y���I]q���e������T�kG�S��L��a�êR��� �J�Ȓ�{XoL��[�^�hU=d��Y��D^�����(�5�k� >��5ө��u�������?|)_}�C�q��x�>�26�F_z�T,̅��C�hh����8�����  ��3���&}��40��!^'7Z;�$����h*��@H)%�(�Mv'���]Ћ�����D~��2�K̬ݺ{O�ַ4P?��}q~�M�T�^�|'�G'
ʺ�,�+0Á��9iP�0[�Ԩ*V���ٜ)�+������������1��$z��(�T����t�LU 4�V�G9����8|���L���_|.?�������_��| ��h|�~�����Alx�6���l�(�qւ���A�e�.����@A�0�{�!�9�b"6�7��qkw7� ��OeemQAS.s0Ļ,Y%���y��W���{h_�I���\\�
a�c��L$�A�h�oz �.��j��ׯt����?�Kٹ{�.���@3?�qiR�5�>�Ho_���2AӼ���tX��K��E���׼
�suM�sq5d��pԨ4U>]�����iiF5!��ӡ��ȌI3��eWA���eJ���C���ބ�<���)���z�[]5 �t0�Pr�X���Ľ�s�*O����1ߗ�ύN����vy�^u0��q�e1���/� �U�J�lH�?�`���v�BD$H(�`J��|y���Ό�W��k�;ĳh)����3#� �x$PIZ��S��u�硠��²�PV�,��{"{/hX�XO��EV�Y�(�{Y�$�|�*gI�+�y ���� ��g퍬�ɀ{	��^oN�r��$�}H�o8ߧ�3DE��?����ȡ׉��1,
��:��v@�ʲ[��ЕX���a*:��@f�.Θe{k׼�0�S3/��'�7_M���������TP�{F9��Y�K]w�2��0�o�\A���<�`;<8bV@�������vL�"J����^� ��J�i�T�ܢ
nf���x5��'U�*;I1G�% d�pK��I�F����u�!�4na� �7:J���@J2z.�d6Ǥ�<q`��h�W��s&P�^��F�T�"^,s����n�=!೰��b�^[�$�w�����ty�D�DTC��ұ��F,���u��[D�'��"�u���A��n �\C�6�,�{��k���m�z�㇂|\���F��OM�f�.�~����DAi�q���*���O��l��ϓ:�o#�e��l�����(��|5�,���7�Tgh7-e�7���v���y�u݀���g�S�Y<+&~}��U��-|��A1�]=,*"l���4�����Y��!o֚\�5��ݹ�=�'&+%�MOL5����rY]x�S��7=������c�f���Z�X����2Ʌ2[^Z�Q����������������mU�@�~�#h�4���r��..@����"8�t�5��e�p���t
"@��՞o�8�t�S�YX�h��D[�_3��x�������dƠ�i�5�gw��)UK4����Ԁ}]?�d}�L�I;CS6�3�/��k��
��7�X��a���[d�I1��Y� Ғ�+�^;�rȬ�����j�I���8f���&�^���ƿ9n8;#XB6�8}4P�3� i������|�/dssK�{�GR�^�z-�'�j����>��pd2��"��f39�m�Hp�@6s>�ܴ��{��9fYQ!1��	�l<[�| x�|��	$���ja�����T�`&W~(�2�ƹ�2m̲uF�������c
�˂}/�:�HXg���]'��k��=��S�w�>)'ຟ����簺��y)C��W��Z�ڽ;�Y+ b����
�XEf�i���8-�.��w=$�ʒ ��8��~I�)یs�b S��=�+��"z�_A���<�#|Մ���.*�E��a����tt�l�vFŬ�&�u�F���1_�*�M�N��@�j�	�I �K�+L���*=�][�x�HЬ�:���.{�����[9:�W���J�����s��@��Ή�2+,ق�s`F�V����^֞��Ŀ�D��"A�s��l��#*�=&X
��&Q�}��E� !TUz b�('�z>�WWH[��8S줖d���|�g/�/"اM�b֭Zڀ���%�,��X�c�����������k�&S�֭��w�5�8y��p�G�m���̫� �N��7�
�:zOy��l���+wt=H���f*:�Ux�����^D$����d�14��A�I݁�K�8u��3���ƞ��<;==�1�=��<�?����	ԧ����`!��7�5��Pi��zqc6���Ψt�랇��x���T�kb��݇�X+��uR�mBc�4�6�4��D\yޞ�䪿�HI��<w�S����ƈuXAZ��^2�Φ�]c�Uɠ�_�}�jLDQ165P�G#�.�׳�+�8b̘ ��<��`��x'�p����h��T	����=`!�Cu���l3K�R*kΐ��փ�+Mb%>�gmk���Q˳�O���?���3���K�]�x�wt���#�gq�qC(����m�W����;M���4�V��[7��x��HB��^��&��	��.�NvR��!Np�Yk*{�&��8�� E��+�m���B�D��hJ��q/�f���2>*G�i��Ez�T�{m/�(YZ/˾>QX͠�9�FS�)���-*�x/��b_���YM�}qx`R��2�r�g�nmz؇� ����(Mȼ���r����� ]�yW҈ʚ�衿�`׮�������m�,�n�l�U��+s0'��^�!-2�����Jd�l��lOMA�Ԡߔ�:�Y�fwaI���=��0�jo����&�Yw���ko�>���^A2����0��*Vwnߖ�;��� ����U�uƌ�53�� !�r� �]�8��L�)34�� �`�΃e�eJ.��e�B��@�+K}|Ȏ!��:���@��:2�Ru#CP�Z���\(mm�0�txr$�:>��3�я~D���Wo䏿�R~������Ɨh:����YR}iZ��4���P@��t=���]�!!��w	|S^3��9*�z�%���x/4�#ۈ|�W�7N�-S�GgR]�م5��(�̈p��,��ysy�g33֠E�u�Y����z�q��֓�y�s࿡
�埾b����ײ��-�w��=(	�>�t��+�׺��A�H����J��k �q�v��Ɨ�y`�B���vw�_�ܯ������R���E=��� $�
��E�����9^S�G�h�� <&�_�j2���1�]��x=�A������ԃ��eC=1U'	�]ָe{v*U$�{�c�t�c�!Vm�i��s��S��<�D����Y����N{w1G� �}�{��\E�P��j� BTe���zYC�ƆGh`#`�*x*����>Wy���$A�����u�غ|
l��y�-s��"�L�8�jO���pS������h8LUF�H�c�Ӓ��<!I pOu3�v{]Ӫ�ؠ��>���)!���ra"O��b�92��]����y�⽐�6`J�Z�<Up��4w����Ϙ�������!�	#�Hc�9qrt̊9��ls��!{�P�g�ʁ�hR~I�d��� ^8{X�F
k/�2e��`fn̆��s��t��i�K�$�No�=}@jإW~z���AO���*H�*����ds��F��y�7k5��i;��hBY�4l�i*7)�s��ȓgY�܌C��g�'G�a�0�S���^���g��l��	�c	�T1HX�1��_篸�a�b�[%����1!��u�Y�7��W��9��x��i9M�Hj{���νa�%���8�(�.�c���?�����������Y����+�y>��n����"u�_ �d��l���
���LQ��.�M0��ֵ�'��2_�xE�N	=�5����|����U�JZ�$�J��w�?X���|γl�����HCjO1i��$m���b�}a����unZ���R����%�h^9j������Kw(/�q�/zO��Q�z`|~(����P��N�W��TΕf��0H�#��3����Uh�C�@��t�@�u�� ���9ծ�C
}�I��/6�N�8���V�^%�2ۏEiK{��1VpP�
ԯp�Ȓ_3�$�B��b��~P��z|^�.e�̙6p�Le�@�4 ߿U�2����"���%/4��Ve��$�����Ϟ�۽�rG�>q>~��	�c�.�Hj�9p�Y4��RU�f�yxxċ�&	�O���</� �KT�Afv0����uYZ��*FP��  hWf��@�d�)Tn�����@�v��1T�6�M�S����wt����O�!��x��ʯ���O��O�8��.��17c�)�4.����϶����$Wc����Yjx@
��s���
R��}kX�"���p#�@� � ��*�:�����_D�aM���e�x(�I�B�ӗ� H�w�$��� ���tI���5�egz�t��Rϸ_���Z�y����Ho~����]Y�ߗC���X��f���>�S����8�*���=�����蓂��ֆ��=?ڹ�y�
玾/hhP_^��u� �Ӏ�?�AcA�Ry�� A
�4B��q->x��U7 :���s8<gu�$�\�5s9�@vD�pô�~���=1�&P�I/6��6� �+�w��b�I%��9�	��xl	$��=`v�Y� ��� ��o:�/}����c� .���N,�#4ʻyV�r՘ �����	vp1S�x�@"�e���թJñ�6�H�ao����d�ԪB^g���4�r!*�WtȾ$�j�A��{��V�J�Ӱζw�Y-)�Q��{<a{��D ���Dda4���c�c�,Q'օ�3�-�1�kJ���j��@"����=�%�P�0���O�:��C�,^��bc]�si�}�����,�>r{�O$I �s���8C������u
���o�>cZ�Is�pl�a<3A��4�燊�A$�._��2�Q�`�OL�Z<)�T 
O�YR��y� P�$]��bj
�nf1o~�)9��m�=�5�O7yT,-ie	^��O#ۏ�.��`����w�Z&=�d��-���_�r��5$M���zF;�1�����+r��[.#��3�J�a���dTuRA/�T9��@��iG�tZ����g=>������~�7�ʟ>�u2 ��Aoe}�'Y:R&�2d\� �v�n4T.�Y5�Q��ɳ5��9�y�tܜ�F攢�Ɏ���WVN�R�tخfD`�p�j���D�ԭש��[p&��T>ɫt0Ԟe
���vf�Q��ҋ;u*ΔV;�@4{M�v�L])�.K_de�~���$t���
����t�h2�F��9�oA�	����G�:�:��\BV���Q���J*aB"tsk��.�PWz���ׇ��=p�K�%���w�J����ŌT ����`C����|��7��O�꠭If
PzpCj0�d�e��5�x��	�Eڥ� ����7���@�=!��5�H�M���T�:����ook��`Ҙ'�p8�8�M=�7�6HY_[�G���Ns�?C�c��n�����-�_0��ھ%V���V ����.�{�t���[��,rdǖiɆsݤN�� �
�3��! _� 	�'�lN[��\׻h}��?��ѱ|��?ȋ�����B���������Š���-9��CF�T�2�+����"	%��q�
�+G@L���6%4s�:P�06�L|h��!7���\&%zHXq�!��ք�>Wt�Г���Q��R�:V�?����Y�
8�nE`�3�le�7��>е���f�z���:?6���!�����>0���������~X/X6V0�q��+}�� :fh
�\�6<C��>.����P&0,X���I����~�?��?~,���/t����9�O'G���>N��6��+Q͈��k���*���u׬K1�"�^�y�A�m�χ�'ҟg�t<Q�Xt7r셠�+��=F�����.ϭʈu��B�gA=��f`����ν{�M=�l��И	hk3I�\% �ܢi�phi����,�5�T�@��3��rQG�`$ʜ��,���-躆��Q[Lr�e�s�����<��`�Zrˌ#d�7��*|�Zn�z
�+(�7��P�z71�~��0}��5#��Ͼ����)�U�'����S�I�^k�F���O��xf���L`s�*���ݝ]R���)����'��֖��\��qL��F��8ļ����O&5����
��#	گd�k����=�$��f���+Z6̛qC-&u>��ޤof�<K]���k1�2D��fF����C�������^)$0��fsʣ�Wl��5����P�v�)2��[��˕��Ʀ� D�T�8�[�E���zD�f��&���=��U�,؟4�ν� 0�'b� �������w�9eRޝ��~
q#�)��q�Qn e$w=F�� @��xZ�1'��LU�ګ&_=q�@����:�.����˯���3�+|�9��ŕ^ֹ�ɺ?�f������*���Uq!:��9s~,������X��χ^6��JA�P����MT#�2�N�ve� -����[n��]�--��>Ԯ�����H��*"Y���t��$Oc�ʾ���4�Y���Q�9U;v��H%��O�;��c�QN��Ǎje#++����靡�um.����Nc�v���3�c�q�a�a� \S'T��yӓ��T^iK�r���4=w�VI�(h��M��S&|��F�$Ee��?���뻽��)�M,SoBҌ�|Q��z�����@�� 3����۟	����~���tXK_x��o޽GE(��z��/{z��7�T�![�k��-ӧcQV���:�&dq�!(�Aľ��i򏣏�k�z!u�ecY^�2��du�T<�I�L�����N�����䈛��ܢ���%�^��o8�8�767�OZ�o�gO�}JWkRi8Y����+����ݻ+;�p88>��D9���T�F�5_�I[��<����a�9�m�c�N�]0H�gc~Eo4��A����QFW�cj>'� E�M,yc����2��{zU4$.��X��XV��d��=*���p�{x(=�q�d���<CU�w����Z����d��Y=�	uq`�kp���FC�A�x�������Z��.5H>#�P��#����v�w������;�pNO��VV�t�0�����G�H|�浬=}fj}Q嘩_���ˣ�툟{���,�T��w�,3qe7��<G���<�}
 ��d9�G_��2|�@�	N!�(C^�Y��o��}����M�`Y��ԯ�YtDU��J4wǨ��e����
��n��53��� ���q�p ������^f�\:�P,�rz��s	(D��|�`sS����A�x� �TNZ��c��1���i4�����ή5qϹ�,�؇I����db.��;��7E�Nf��YaJF!�ZP�8r����hvݔ)4:2��,����ˮ��-���^�(!�� ǐ�.LA(/z��@��	�s��Y�J�	2I�U�VYYB0�ދ.=D����d�f=�Fݡ�Uf�byH��8�۸#�7�o��t����x�c�5���e��K�����)`�����.j� ���v1��Es<��l����D�?e�C`�X�u	��涢g�t|���Cv7O�JҜ�"[�gF�h��H��S�jbqm�1f�� ���I�����g�Y#�Y�7�f7U@ؐ�X��t�+�V����z(z�1f�, ��s�fa��IO*�i�x�r�d�Z�L#z|���?}���ϟ�Nn|�9��|�t��A��n>�G���!Ec���5��(5)��� ��m�>h�q�A��4e�`�2�xF8&F��Dp鹁�Jb��LI�6�,Q���<Ǥn������%a�<�S;���Mx�M2�?�ֿ��RY<��'�S��Dȶ�ɡs͔̃���/��ic"H/�,5؃�dA�@`�{\S�UsqMY�ze��@�l:��C��r:�� G^X������ֻ6��wh�D	Xl��o)N�*�p��F���Hi�Z�M�d��޳�+fr��D��D�9l
"뛫�M��6�4i^���?Is+k�³&s�>����d��Tut,�`��z[�u�Dp���� ���	�E�vxR�oc&s�/.�0�xnњAB6e	���l*8Y���`�룉e/o-�ӱ�?��j����/�G<�2&�
|f��,+8�1���2���޽���w<��^XC�KC�i�P�i:�g�{6mƵ/���{�������k o�%Wޣ%��(�Ҩ��D[{�\�~N�%�A􊀳�漏�@�����]R�\�\w�T#d%?���L�>�.��S(�e��wB��f�!�U�]�\^Z�y��c[��ѹ��}��/+[2���u���UPҹ8�lb�L@���N�2�P�Bs���{w�A��T�P"�`�?�9̪'ͥ���#�?|��j��S��0`�9+�rW�W٫�J&<NN/ًt�>��+�W����{���:��޽e�Th��s��gu:���*vv�]�z`�A�L]�� �����4� m�]�Qݢ���;I�3Rp!~7oT,B��z
�U�-ޮ���9 h��5��ؓYef�ل�j��F�7�ˌ��ݟ1*�[X���y��A-(K=�uX��,k^����
�@G����nG�'��fԘ�%�I�h,���[0i�1tk��uԩr �o T�l[��: :B�ef��L��������_���D*@�����W}�BPy����*���?�P%��:k}�4t���A5a�����-����1�D�����:6	Zf<5V��&��0m�D?���lb=��=?�}���6 �P��4��z6�P�gF��j�\�>����F|�=ʕL�v�}.$w�:K} �=f��8(�;ZL}�4�fE���_�q&Nqj����	��\Sd��N��=���j�o���ޕ9��iu�!Y��%��FQ��M�3 ���8M��+�n�Yu��1T��'�0�U�����I�����H��]�7ϼ�&w�g��Ǟ|�<�͝r��w/̗ҁh�L�d�Y;c&�A��V�V�n@��o�~����G~��{�s˷g'i���	<����,+�1K ���uqf-s�0�˜c� �#V*���t���p�L�V��Ҋ	֪�`aSz�z!����.�6M�(�֓���J.� ��MV������>��Gv���G�US�.�~�l��4�^���k��Rt+3�2�_�)B�o���e@s$���f�f�ޭJ�r�95�u�P���������6�k��@�	*,Ȳ\]k�U��]��d��2(r ��v���Z8,h������W��e��� �2c�u4��u���꥕E��"{@W஍;�(E����
#~p�X���	��@TN<�YZ����(&� �Z���!sgkSV76H�:�{/{��3�y�c������W<���U��౲Ȇ��ԼMG��*4�s�b런�)��Nt~|8=����$l[�5)5��"˺󽥐���r���;����c�?n�@�!ha	�@B�mjM��o��]��ӟZ%M����Y�A�r�=��3��X�/<��7dcc�=lJ��ʭ9��Wq�54�[vi��� �
���|A�!�w�����A�<p<������ }�
$ȘB�G�}�����7
:�di}S64�]�g�u{W��O��՜fkjcY�؜�>�)����ھ���mHX��+2�&�;ee����CRh�-� �:D5J?鿰���gQ�~�i�te�Z�Xi�ͬ����+�YQS�C@� 
Q ��(༰�Pp�u��%(Y*ȼ#x@Љ���Jvv!d��s�k'IX���g��
g�h�<t5��ekK� p��y��5��&����H��n����yT�Hcb �1���36�^l��.������ܸ�i��� 
�(���?��������C�'��%��]��f���0�Ʋn�88��t�b�������3���]��C��s�ZE��FzWW�:�q��w=�P��0�<#؟_H�%ǧ�j��SS�آ�HI���6ۺ�NL;�2�K��G3���8��71�?��}x2/���o�W�,W�?�,�SYP1���*�*>gf��w� �����l#����]+0�Rѐ�T��x͐pOǬ �^��}���2e6� ��E3|n���Smc9�$;}���8�>������g>�괚�����Ly&)9W[�)�io?�Hr�HKz��*��R���U��e��~�'�z����t3*xz�^���S��&j+��m� d������G��� K�{x���E{uR�ˊ= n�P�9�H���L#�,�^gbB��S��S���O�o޼��ٷ�~���8�W}x�7���w[�37�\;t��4X(;�R��b��N�e���.�a��vY�<mp��Q%��E��B�j[�_�ks��[z�{�W�X��tw~�Y��72��,���Ŕz3�e	i6����ۮ��i���D5��,>�d�r��h:7����A�\�5��3��U��@Sb0�X�(\�|H�T
��Y0ᱤ�͇q����S/{h>!�dG��X���C�$!�i�;���V<�g��'Ɠ�̌^��n�D��c�}��Fv<�݋B�qj�t��nǖ��#J�b> �al����od��֚�o�JF������,�+���0������ U�}�X~���ɓ'O��o߼��o�*9�}O�Cf���z #	}�"�x� d�j*F��i��KVX�P��r*��C�n�:>hzG`�9t����*��?��c_�Ӊ^���>#��Ѭ����N�g�\��Ll١� �c���?�U�PQy���|�ݷ��ӧ̠��|:��F�):&�ʼ��,���B9���� �6�U˭Ԏ ��~8='ŉY|�����)4���Q�~��{q�L+���L�à�0i�'W�w|,�޼�9�6 ��2]���j�������I���=&+{�t;�j�}Q��`ps^S����Dg5j������dl�N�>�%������󳠝{���gwY5b5vj�w�B�gP<3��� ��⺵���{�MY�ɾզie�A,ewg]~��'�꟟�Ȼ�o�P�7�� !�8W�Y�u�ѳ���M���`8j�ɞ`s�5c�SS+䥶�Ak;�\��0�\evߚ�A�c"E�)���[����A��,���j|?3o��׀tw�lS
���l�P�.��޽���n(oޜ�G�M��o��0㗜� �} ��-3w����s�6fr�׬b�����ez��B��٬�5�o��Qvss��T-P1QMB��g��h|k�Ϭ�+�-�
΅j�+l� ������Ҟ�a�s]��J������D~����o~�/����-%��W<Oc������WX��&Q�4-����<����]3/��TгH�
$l �۟_�Ĺ=���!�_W�v�������w�$Af~<N���eOd�F�A�|�c�u�>%}&�LͳL���8����T�j�HD�/�bB�����%��	|Hj�L�c�V�k���w$�@��Q�j�?�h	﷨�d��ٴ�d�7�gF��QΓ��i��-K�,0��yRMRB?ָQ�욌Fl�c�'�����Ufl~��ә����
	(KU��������{����j+�����%T�~-��3�G�Rw~�1�y�����ȸ!S�"�Ȃ��cxX��� ��QU�a7?g6��VwFM˸��+��!�k�A�I%+7�j
Z�`��%k�;�-brZ���� Өd�+ *�4���zQ���n��L�<��{c��WN�J*�n�El*C��Z���I	m�!�҈z� `� �`�&q�q~<�Re�\�ܰ�u9��z2����-.-���@$��N���`i�6En�T	�,�$��n����n'#��-���)�}w�šVtr��ܚ�Ųg�kb#��$f�x�oDs��AdY:����}��ŵ��߫g~PKk�F�1M�6H
}�G�t^FvA��ζl�ڕ]��>� G�r|p$�G����@�ԍ�p0��H�4+�{H5��A./U|�*�똜-�K�}sg��`�@do ,��  ����}VF����kTC��AU�����Ҁ�p�{ə��B�W����`?�}�|��g��O~L�9��/��۷|/�ۨ�>� ���A�I���gS��Ν[z�tJ�D���1�(�:L/�y`���_.rV�}D�����iЊ3`p8-d\"����)��C�5�@K+{#�� m�0T|��t;�ȕ>���%9��G��i#uS��'74}��������2���#����#	eh�+��<�݉˂�������Z@
!��\��ǘ�ݹ�£��Ԃ4J�o%T{�P,��6�� T�Ͽ�
S�7�G�B��h��}l�Ƿ����З/~��7�sA;������1�Q�uv�@U�!S�ji�	
��~o��;@������eS�^3���[ö�7�����#[pQ�M|l�Z�����{�Δ�d}��{kޗ{3�,���Da��*�����O?�E�� �,z�@Q|�������z�2S7�c�׮9h�q��jQ�G�q]@�������38?�Եq"�GGVQױ��A�t6�VU��\�&<`V\��ް��-��Jt}��Z
���=6�s�/*��9+�;�%*�I�sd�P��ۙ�m����_��{�}M��W�es���dHkҩ�^<�e6a�ܳfu�Ƴ�%�� �k Y�ss8R�[,�s���snen�g ����"�i3���^7S�A�o��wH�6D��ڔ���}�@2j��0����UP��<��}�jvh?�>2���[�ۼB��߽��M�W���P��F��Τ���"�N�Qa��PUU��/W�k�K�agW���`_��x��,����4K�eq�<3��VѻA�`
0�s-�9e�WGĪ��/!�w��,A��z�����<�"�}��>��Q>�ۮ�:�s��0��䕚��f���09I�Bi�i-F���T@�`�čkL�\g�(���c��(�Z҅e~����v�F3�!'צN5t�f�̳��Qy+*M�z[�*�����aeZM�Y5'f��ݓ�=Dn�f-Im!�G ��k�bħx��HČ ?� �G��M]�����9iW��m��Lų�f+d�J�Ԝ�8 �q�"���5�����(��%Q;[,<8c��c�
�G�Y,�G�bf�t(�M�Fb/ݟX&��Z.8�H-�<���6
\W��$!0��x�rje\��`�[��u� �L[+�j�/b4--�3�]�������T����2V��5Y�'�&=���e�3
�t���&�c:q*<]z�����mаr��x�!����vIK� ~_�~�y�*̻wة>5O���Mb6�z��b#�p�t���c�K�\���/�҉l�}!���{���Sy���|��7T�¡��R�9�Kr��=��������n�8��������Y僢QY�S͹�sh��i�+�v���2��A����3ܖ�ysM����t���1��V�8f�p0�>%=��N>*��=}�/�:Vx���=E�9'�ʎ����w;�}f�NjP�e'�=*P����t-��_��
M�:��{'L `��.�١0Q�Up����_5u��2�*�˞q�C6�8T��?X����ڱ����e�ru��;L�Yԏ,���>������-�	@"����(�J�~����N 9�S��!�Eb�x�{�a�k�-iC5(�o�+�O�W���^V6�����B��Çc�e�RҴ6O�Pu��D%
ja=�����EX� h6G3?�8�߼y�{�y�5
�9��ϐ�L�y�$�x�� Hgc \�\�5����'�R���{b/���	�_8��{l�'=덄��%%;d5�|��:���,�������:����k�2���w��Z�gG�g��e̝�(~�NM*eA�k����xNM2��BZ̯b��/�r�dd�;4D��^,��>7{�����F0mF��d[72��+����s2��os�z>�'.���
�
UVYT���:�9�vr��ړ�#�É��`�A]�=qZ�*J�4�����귯��4���<7��V�䀠�@W$W��6�$K�!��}�����f�1֎i�"��6���e�X2+�= �,���6��E�T�H�WY�:
z�wJ�D��KrM�$���so��/���%�-�aI�.�|_V�-�G@�T��k#�`����(m]�f8�l������_~����{po��Q���B��>������h�
�(�5fSXd2��mF�I�Z*C瓍K���SÎ��`pg�Y�)�J���� �(}�AF��3_���kw6��E�4��$ �Ir�vM��Qθ@<�O��U��D0(d�[5��uHT�-m�OFs�ԍ�`��ld46���AI�6��;�x�0�v��l:����n����H��t5�d_'��;��ѧ��έ�ܴ��|�C��Y��/��Q��K��[��9gß����:W5��!����i���hH� �~���*�!xBp�x�F�ٞ���Awzz��4�{3��CVG-���}���"�B���LH���� r�+| ��r���%ЀN�������+;�\[�:^Kkk�Y�9���C8���opݑ�Y掼n(��A%6 �te�sfN���n�h$~��_��� v�2++
�<mln3�����g�~o_�����=�,c�?��ֶ6��}Hpޖ;��1��կ���`�Kl.v�s�ol��ʃw5�KE���ɇ�o˧�=�ϿxDZ
h<�}�CV^�ck6��!T'� �z0"�8� ���{���\]O�r0D�}lG����G�Xi�r�:�+.Ո�d�>� �R�ZK�K���swոԼY{`^�Ϣ�f��djdVr�;��uثQgNM4�d���8�}@�{4`�5ř��Ֆ6[�iG�k���^B�ū�{r0�p_X<c�*3�l�Ɍ��1)]��$��!��g���k����CcC��
U����S&9�t�ι7�Z�d�5���~E9���3�Rd �����Z��)}26s2�L���
bz����s�#T�D��<��h���9	Zҩ��OT��c��khL,Y�3u�f+��}��~v��׀��[�vy� H��µ����t�����D4����֌�\ӵ��W�&��}o.��4�a��wEU�L�ӧOYq�k�-�������B=o�b�U����8g3S�#�(���?��l*J)�M1M&Yk�eM�^�r+n�= MF��\��(.�B����W�HH��ɂ����d��4��~	q���3E���V�2iM�8�[�$I{����*{�yO�����-���I�?�<4���RF�+yĈ� �y�E/���X���f_��3���|�l�����%�G��n��7=��8��l��cڿ��5�� U\q`$��ΜmS�M��zV̀��d��D(�;�ry�w$�S��-w��qm��oH�>�W��8�%�Y0:n��5q���H噁sߋ��������������7�$���:���@ݸ����r��L��vʨ��0�#ִT���4���ZV��oQ	�L)Pr጖e��F}m�p4{H|��`i�	���x;��\4=�lyw4#R�{��"m��N[\�<���B��S��+m��������o��9�0�l�5P�MX����ӓc6O� P��U�����L���r��1��:�=�D�ܺs�t���ЍR6h�����_[]ԟ_�5��1���:�zL*�Ȧ�ˈ�8x����]s�-�����
E��3��t�s4�<>:�ˋ��^��#_Xl��AYdqaYN��M�0�
�=�&�T���$��%���uH��Qib�g�z8�MR�̱
J��:�W���i ��Նܾ�c��//ظ �m�}�E ��q�L �^d��`����DQ�@�	*�5x���s��@���`.1��=���*l��t��@��y��#�oW Ngr||,{�!A���߹Ovn��(�T��{*_kP�ǯ�r=��̟t��w�ޑ����l�Eer���<����_�X( y���>�����Ր��s?O����z����A��_���9�(T�A��X�d$cJ��K ��%��	?T�ε+��X&�+Q3�g(rA����i�KZ��a��렻f�E�|����TpR`���	�3��tX��74�f�Ӑ��G�bKY�����������yQ�� =+�X����) A��>�+������k�7���hO�{K�v��Z�ʿ�~�S�|��soQ��:�X�2n~arĕ�/s7��AT|�7^�M� ��o�5�B&<Q.:��[�'.�<K���]��\���_��7�V4q�|Lݻ�c���w��[���xtxD�7P�Pq@C�p��*~u(�^����Q��-S����ƅOPq�X��H��Zy��`��i�U60 F����dT4���β��7��o�NQ���EbT1T�V7�H�¼]ZZ�*\�cH�=��}_��Rf=L�210�l�K�F�Y�/U� �'��tYZE�2�s=�t���R�X�='}^�񩉵��c�)RE��j��VH��YZ�;�b'�.��1˚���}�,��JF`�#}��l��9}��2��MDE��_�d[Yō&g�Ss|cTd�\�S*�24Ȥ�S���Z�)!Y;�0��K��j�4�L��@���c� ��_f�]�j⴬��Dr���4s�ݶ=C�P��m��7�G�'w�#��i�Wx^����{
�hM}��">�Y��\�~���x6 ��g���O�"�v빸(��>c����Ԃ�H�/P���c���>xt������������v`ȏ
>4��>��_Ow{&�|�=Qo�V�6V{��W���xS��F4��'0F�~iڎek��X�����qt
�M!��I"[����y��*_�Qi DL�T}�R` �$��T<����)���#X��M�e]���a�5����U:�:��o�f�e�5X�,!PmH��P�4%)P`>�/4�AG0�Udh���F�D$�C�\�P�B`����<��ܹ}G�r�A	x����	J��!{��ܻ{K��ް������kj�7�z�#���>Ј/w5�>i �w�6� ���4����lWV�dg��ܾ}_���=2��t����!d�z�g��|�b����:=eI\�4��͖�pI�k-�I��o>����kW*B�p�!�1�rq5���L�����"��ہtbT#�Zq�s %Wfi�/��=W��)}W ���x�`k��'On��w�L2h`x&ȼ�:�*���� �p�A��	_�s:�`4v��P�eW���7���ٳ�����ʯ���
��D"l(���Օ[�o�����G�ۇ:���c�v��}��'?����ޑνc�������{�y�!ؤB�����s�|-�^� u�?����µ ܃&��t�ذ隕���b����Y�H�F���ݬ�(���=i�]��Fx�hpP�l:�4��UMY�Ȱɤ&%��;F����Ӥ�H'4$�[�k�����;ˌ�-٘����r4张z����rR�e2[��l���,�Hf��BL����@�uZѠ��ΉS*
�LV�������Tx�%�:�VMf�z6�{�� �����z�x�7س��7��U�I��������Q���Pe�1�.-Q����J���>�qO}��<z���T*.��qe��h!�[�L����4;;撋50��I�;����=+i�h��x����
���x�2٤f�y�};��O�^��W�n���DO �*��[;\��^xEu���X��H!�9C�+Az�3�p)UT>������Ϊ��/���w=K��LM��Wt�y��O���qe��������@� ���0wx�6A`
27���w�\�&t�kz���R�
t�.ؿRV��=e��n��^R�����h/$�ܩpH�ܑ)#�7F��G0�N��VT ��_��0�;�}h42Ɓ�p��ϝ�8�b�V���n�i�qR�>^�7~R�̈́i�;�͙�N�� ���HW�o���N���M��/)��iQ[������5C�6���ɼ�1(s@.ZPy��c��X�{��{$�����w|/w�+�ݹ>�����VE�uL��[���r�S���;�d�������w���w�^����|�P���y���S�,�,RkB6���a��-3''�.$P;� �Mkh�,����Q@=�f5U�����N�n�Vu�ff�zZ��߂�	$ 	�d�m��;�Ҧ�]ӥ���<	v�� - kln�O��xi�Ebfdg����=�o��ac*=e
��}~��MT����4p��B2��C���p��'C�B���G����I�4f%�-x`x|���ɓ��������o�o�1������� �k[�l�����;/�
�>�SR���(ܦ�5�v��Q����p5���=6(�\�p�6���������ͯ���}@���n��0����{4II�@Z���s۩:�Id�������7���ͮ��H�gIp�k���}�x��
DJ�A&��/!{��h=5�[�LtG�	�����0�FߊSo߽���,�r���m���a�BU>!���1���<܌5���AeI����`�{����۷�{s}Z�����=�
@���eay�Ք/�{y����~���[E�.�1����1u,]ʇV�L�W�^* Q��78��߳!��3A��3����qo���< ��"���
��z?�
�hV=8{_�� ��:���#la���k,�t�����D沥��&lzfVEG� 6z��̦}V?��5%���2<�K���t��M�*�&�qYr{ov�T6�~���K R�ַ�4*��l����VY�&cl�����ͱ'�j�����΍lr�9#�.U\*�4�=��/���녊�%+��N�DZ@���**}�t>/��l�F��U�| ��ۚ�o|d~��+�׬�h�9�	��|=,a�b<�y���L9M8ON\�>W����5=u�las��<����.D�ZV��u�/��TY��m������CJ� ွ ���x�u�׌�֋����76(4Q�es���9����5�+��x/��x��~+���ӺK���sJ��;M��Q�m�D�Mۙ�Sf�<�"�V7k2�R�ͳ���|i�/;;w�?`e|:�б� ���M�b2��/XYs����Y�P� 0*@&�25��$k�g��R_�7w�|��c�����ξ0�D�!�1Ǹ���cf}ܨx��dT�22�>B>�SL,&���?Ӝ��_��(r#�bd<t��*�%0�Kj��Ym#I�:�\jS-e�5�$�Sm&�g�bk?mLh���yV}	�]UJ&g�}����� ������v���y��laM3y)�WV�̜v��̚��2ō������9����P��]�Q��a��+0�E_כׯ�k=_�~�����` �`���=y�?���/�ts��=���x��T7���M|,����M��ڴ�GΥoO"s5^k�2a��|�[ e�a;o�hl�-��R�D&�J>��ļ�nL+�5�ɐd� �Mٻ��F�$h0��]����0x�=��n�R�bA�Ad|DOG(%5��񪫦zd��^���z��p���ڄc�Olp��_QXPYM4\���V�L" �Ƙ�2f�z�	`d����Nl�0eZZ�;w��_�X�ޓ�˱�x�J��ǯ�y�DN<UϺ���I�7�c6��hHg>�_XE��sVR6�7�	ւ�X��-�N?|:V�������KJM>��;f�s�����y./�2����@�d��@�/��W'T�� ]�%T;��9��D�s*�(�x�ᖥ�V���"�%c����v���	��1]���z��_\����:?����I�j[��<�Q1��y��/�,k ���� c ��X��
@�
pU��Y����LD�J��&�� {g��9�t���/#�X�(����`����O_�I_ｼ~���,��pl��xA���OdI�{~iE��s]��o�1%>]١�+y���p|��{��`��������,h��͍��sj�c�{Pӯc��F��j ���������i�l-�TO�N�-k~+Z�z�r�R�w��?|հp���M�,�&�1D�~�*P�W�S�bPrf��&��߬�ْ$ّ%�f�{��RYY������S��m�|��3G�|�pDzf�n�`�-�*#32�=�w3�9�z�zd&-B�2�����ڽz��=Je$�G���o�j��Gv�5�r݄��(z%k��I#��_�q(�0�g6��0�(��.�bry,�)��A�4Jd�����\�N���xl!��:�ei4#8���Q�z|tL�ۊl�m�m���]e�o�'vty�v:�6�P��!Ë�V�R����{
�՗�^�sm�	`�V��<&�
o�G ��1ը[�nmy��6�nu���!(�]|��5���v�n����D�UM@���m ���G-o�h����y���A�U߷p ̹�*R�@$�GW�����j��{����(]�!u���>8�1��>/+6g��cB)��|}!]�h���
�frt�#?�|E9m�BJ�� |��ms}S����U��m#{s�vȀ ����b�c<Q����/��/�o��K���������C&}e��y���>DX�܇k|�����o�6 >XI5�ʣvo�;����%l��;�[F���lz! 2�B���&Kb>��{��{�;+�;A�/5��-1��Aɶ��ri^��  Q둨i��F}������XfѸoG_zb�������yO����^ȨMa3b��Bb�[�O,j�x��D^Ǵ�լ�lI7�A�Y5�,<�
��Z%�}��������O��~򓟐։�33;�z����g/�� ����|�X�fK�<$��}ӿ���׍d*�>�L�N).�E��B�|��RBu�h����f*X@%����N�P����?�H�I��2�]�LA7��ѱjO�e�+/&�75�� ]�He-﫦�_7�P������>>˅�_��F�rs��t�rG��n�����C�o������4P)�e���Xxu�%eQ<�6��Y�d��"�?!�ӟ�c�b�0�����?��ky�v���N���m����(<P��ɩ�C��"����՚���"t(�@%dK�PS.)�J�(=5�8����\轀,)����q���s1w�pI��^(�]G�iQ��F�	c�՟�ٕS1b��������/s�����"�T����k��Bl���:?�W7�Y?:�q���u0�˛��W(}�F2>=�\���Fy��G�V͍�{xrD�K�g�N=��-6��f���
f؍],��c5nȨ�
7��띠�_�~-;;oi���[��O�v�yz��UW����Ϟ?�2$:Ot~�nW~������ip\d�.o�rxzA�lpl8���{��BL.�k��$�Vu��ϝ��ٙ�}'痺V��Y�o�󖹤�7NM��: cn[s��[��p�^g�D���8�kO�!��"��Ə�s�ۅ04T+Q+jO����n�Sq���� �"�l:�v�w��~E+9�5��I[�	d�K��f>:�/�͌�E
��V���t-i��[�?��#:������]M@�0�2�{��Z4Ҿ9����s:�mݤ���mٔ�(�f��E8f�����1jN�HN8��
�g��7'�Ŭ_��{��6�S�;9c��5�.�'ՙ��� {c#�N�c65�{��E�A�7�� �j�x�@��X�Cyn����>�p�Ȳ�uf�P����(SxkN��~Lu�(�x�9k;z�����@�l��^���K\�h��g�vPʸ<��WE0��C�(�A1A!�{�r*㵐ԕ��Ǚ��\�s0�t�u��I*>�p�E����c���7���H��>!��v����s9W�:Yo+\�)����ɺ�哳ki�Mh }gh�ќR�����s:}�pP�xl�y�0Vr����ء�m6mɸ5N?�&�/Y@^�Mj��҈
r��O�Zf[�Xx�����c0K�:�)FG�<h[:����8�eO���Z�Y�ˤ�%wULN7jL�AA#>$	�X`�T0���5j����u3�<�����yAy�N�� b�'�1������g�qI����2�P�km����n�Io��<5ʔ;;?0(��$�նܻ����������?�/���?�ӛ������w�x�+�G�K)׿d:@���YF�i0o�fC�E�ؙ��t���d`���X֢�6�(�,Sc��X)�?6.[�� [SÂ��L��R{Y���ܛ:'0�_���B���g!�Z�{�͒�%�I��CkL�P�
���{�E�{�!Y�c�"I7b�S���$VQ9_/?4�AњL������?�h�F6$��{��x������{�ށ�{2C
�U��#��_)���nh'��� �j�`c�b��	�!�j�v����rQ���?���Q�&���:D�!��x�7P����
ۑɀ~:��P�Ƶ�}O���bؠ�|
vt��|�ݻ�h�ӧ���Մ�����%iU���0�Z+�[ĪMf�0�;y�gD�H��\���F ��Ht��ݘ����?8 �[!�5�!���a㡒=�>d.��^cGۊ���}�3�亝BnԜ�\�᳋����{m�@4�*����@a�}�=�0�M���`�r��� �E��ܑ����aÐb�b����W�����@��"�Ɩ3�����h�����MY��Qˡ:�mh���^�ݓ}��gt>P���s��	�h�J
f�-����iqft��zX-̖�G!%,�H{�jD�`''����ә����U�}�ƪ��57�Fm ��^������3�A>�u'U�e@s Ԟ�� ��Bv�k:=�����@�|��'\?����"4U,���9��؛�o��<�j��
	z$h%�m�2��Q0���5��A,���u��� ��3%M��^��`�
~�"DV�!jlf�Q���_
�&A��'���Y�@�iym�C����QŞw Mu�iK�}��쑁 ~�sˌ8d�����5�=��*�hT�1$=��{(2�Sf�1�ڤ8�l{�x�9%�S����tvD���6���_�3tB��ƻi�B�M�Z.
�pW�$�.�9ԭ�g�̶�i6ۛ���z,�:[���aR����N)t��k�L E��S� �܀^��d$_|�@�쮰��}v��#�otu}SjC>��s���w��HEE_��@]ٸ�ᾤ�"�Ys�������qgM�ާ)i�:���?,Z?�p��5JR�x��o����^u�Y�BLN�jBJ���C0G�f���P؂�L��V-�.Q$]���3�pKm�9\ӆjo����E�s-x�B�e��`31$ePb�� |D�
�j�AS���mk $�:�t�J�^F����t��ҳ!�)<�`��3���G���r��/ot���o~#o��p_?><V��v��ڇ�GN'h��o��������
>� �s�e��KiV��H���i��&j@�:��=�z�q`��hY��с�2�c]�i�gt�h���/��i��Ŏ�áN���#!c:�6��H-�-��N�RU�5)s�W�&��ÌbMF��TR���Q�d�s�M����>R�1�̄�s�Q��Fz��MgT"
�r�=B�4�kσ�M�u����`J+�� ��N�9�S1>Z��[ 3ґKAL_�,l��4������������o�7���|��K���7��*(h�Y��@eQ$ꔫ㰵�MЁ����'��*$:��O��G��E|��N�;0�DQ\�N����)5Q]F��֩��)K��	��xnl����@��:9靎�+v���8�n���a�ųT-^'y�1���"5��ѭ7G.#�ْ��c�����Z��({�E�P2�]QeŎ��8*>a찡��b6��z �7.t�F��@7[��H��n�-ٸ��c�"S�Sk+hOdS��q�q��ڲ�6�2���w���w�u4���Sf\ D��Cq-�"Ș���ʣ'O��X6�l˩��佯.����۽yZ��ˑ���Ѝ���W�{�tt�Lc��g�SJ�
:���b�v�+�W@� �F��(��LѧjQ�?�I�pbھ/��rc[l��K�0nc�²+��ď[D�G��Z�ۂb8L����j�|إ^Lm��@�Y[�RmIٜMR`+$����lN����L�x�ya� �|�T�D��ř��X�G�;�����Y�M�,�_K[Ul�-�9��'�H�n�����N�em���Ӿb	�0ccQ�> gd��G�tv�\�!Bz�n�IQ�Z�:$:!k���w�(���oM矂s�'�L�5���}y���%���]�ds>s�}�GFv��Q�)��.�-#wQ�]�u}cO����#H���QǠ���7A��L�����G�����(ư���J�����1�2�%U�b�G��~�2T�����R]�S��)�*��e�Ĳm ���u���U�u�BZZ�k``��������O~,?��J��n��7/��ǐ��@F�� dW�etv E�oF����d�ƒ������U$?������#E�lu�R�!��}������s��H�,/�5��4�����#{���U:�_�/m�/�"EQ��2wI��T+��[�-�O�Q�2��i+��|�Fv��-�H�`�Q]�Ce�I,XTz���|
*(�V���(����-���a �qw/x����t�ɚ�ϕ��"�#���.��i��u�bL��-������?�z������.�dŠ������g���{]�k��^�����������_}��wy��_>Zeg�K)����։ K�#)"�Gt��G�S�f�*H�D ��i,8���[��0�:+b�%}�<�F���k&�
^�ԥg��NWU*��vdFRKw�ry��"dm��������ϖO�4b�S����kX�^��f���7���k��b��I�Tv���2@�����D���c�v6��#����bq��)2�Hf��� ���7=.8�T��'��P��g�����O��_�����|�5�B�,���;_�q���gA���5��E0kn>�П}C�1� ���H���*46A�� �ju}� ���:���{^����5P�07�T�*(عMwz��."tX��Ψ3��b�%s�tQw�H�<�H��������YM`�>DMH+��1�������uk�������l������;ᾅ���*��A��.񇧗���]J�";�(�޴�0���@2�c���+��JǪ�h���/_��?S�
�?�	a7��T�p,8AѣfC�	�����[������|��{'G�wt&coY����\D��\�M[V���ڂ�1���N1�
z+�а�����u[ʵ�D:n�)�����I�c1fd��;	�%Wӽ�[��m��#~�Gp�?����\$P� ^T���]��l){]
~}/wQ��Yg��$���z4ϐ�f�	�'�r^Y�3u0[]���GN�����@ڨm��:���"���>�p���F=�	ˤ/�s��N�;p�as���ģ�S/*5f�E�5����K���1%���E�?hC�AMD���U�]1�G�۵}@��0;M���="�wq~"��3���
Ñ�00bE�82'���w��<�@%����<{��tEZ 8E]����(lG0'��{[^��
�Cb82F���>#+�����)-��� M!��>O�5r
��`��77�Ԯ�+��6^�I� �Cb.�*-�9�P�b0�n��뮌�PX�s�E��v�����H���mf��U*���X�qئw������AD��L���:��ao�Q٫��������R�t �g�<Od�1V` "���ٙ�Vs����`�d�z���M�B��c�i�N�����mlC���r�/göD�e����;5�F0���w��7��a�j����W�F����Vd�˃T)�������9�Ǉ<�\Xv��I��莀A�S�,���$ K�� ��0ː����Q���I}K5Y�"ݩe�緸�:�:��Q�'S��������y�#�o�0�q}5�\|��s@Fz��]���O��m�z��v�v���������vgggOm���|��no�<������=-�fp��2&sdE'�O?b����:+��kH�<j��j�H
����\�*�C�g
ᄆ�5�5o2��}���8��_�d��Yl��q2�q��Y�	�O/�ٙ/��p�qb�&bg�4�|���đ�i�S������ǆ�&x�$d�ƌ�@~p<9��AGj���nzn�b~e+e	h�~O<tawL�mK'������g/��]���{��#��ݑ��3��k�gG��~�N�2\��Ef��?0 _����V���oS
x���Fa�H [D�`�q)ذ���֞�7��M_��@���.V��a!~�g�z����d��֋����jWՒeX�:�������u�[���Ql�)ܦae '���F���T}�����Gc�ش�bjD�/n.HQ�c�ɓǌ�B��c�s����#څkAl������}98=c��`��|�ܛ�"ñ��%_��G,�E�$�z���� b�Ms:I7�L�=ؗ�;��s�t��K�L�{jt���T*��0�0SYԶN��/�� ��^�P��5�VG6��tOn�_�h��d�!�@���
Myc�e Z�4�xO�y��@*6�S:�i�*
H��LB�6�ߨ�4?-��9˗ݶ��{�=��uۜ��S�NBǘ4�����k]*�EF�(9� Y~49��
g%*�짅/��yQ���2P5c3���a���Nd�)����V��8�=��l$/�����w&�t?a�1u����-�Ut�)��k =<X�/��Ԟ�G��7_}��<1�q��+A�\m������Z��% �36���Oa��,��^�	b�������hY4�d]D��#ԍ�q���=Mj��`,>|(��O]-vλ����1eY�'��M� �����{M��g�}DM]����'��H ������a���ĺG�.�u���';}���{C����B`�L��W?�`v�b�F��
�{� %������^�}g�N���T���#�8�c�:#�ê�\/��g�1�wƆ�Q�����C�@n��fM���{m�+`7A�n������St$z[ԙi(������~L[&�M�jXXC�V���{��Z1�Z@n=�w�^�Qe���K� �[�D�ă9��ʕ��"[��`�.� �g�H滱�uQ��r~r���,>�C^�׸��F/���x�dO�Kmɍ�4��ˡ�ށ��/X��$�Q'�Xڽ{�T�{����HM�(�������O���?��j����/��|��w/�l��������~Z˵G_b4n;AM��[nhvӚ��'1���v�an��9_8h0mp�]_:d�\�����I������l�=���H��H�?�ZI��~�6A	To��]�X�'��\z�+}�|�{.�M_F�؅�i��C���aC�4�{�+�ep�O�](:�H���|��1o���<�H���;9��Fc�e��7���p�2�O�>���Y��ɕ�����R�"�խ�=�9�x���N��}p���/ u���qbtM7Vp����v�����
z��f�W� =����㺿wH�ԗXF�͟'�9i�y�~:�i~}+��=a�'���(���2p+��Q���w�0��P�K��Ȉ���uC�z?��@����N^,������zYD�Q�ȕ����{5���H�F�?F���l���M���cF�N�QD��j�F�Wr�������+=Bр������mPۺ{�k~o�#4@�n�(��Fk�x|v"Ǻ��]�y�:��J��At<F��n�-RK"�� �=�j�Ƽ�s���]��AGat�)��X��Ԛ}�v9wg��m�#�>�C��w����:WZI������Jw�C��L��o�������i�6i�m}����.�ͧ4�t�$��Ǿ/�[�G�dW�j�f�C��L�[�z�Ҳ��ɫꃁ��;LNev��� �ߪ�בS�
W6�{����څ	mH�B�
vc��S�1衔���Y��X�q�1��G����>3�&eCA���=�I�v��um�ǨA���g�tM]B	�c�p@�����+ۤ'�-�0�Ƭ ��8��g�F�p���R�<}J�:d}���z3�9��t� ,���4Jq��E�g���:e�p|DV_�a�=D�lR|��a���l�G�2�V!��6P��e�c���B��N��3l����t:��9{^�b9��.W�Zl�r�����[p
!�Ʈ�%�יMnu�>M�������r|z�c�Ά���8`�]5uF��Sp�����=�K���<��D��oh/!���:��w'�I�W�mw���[��:�B�#f@�c�����h�b��}υ*����D#Ǫl��|5(� 4��X�q�r��	��K,;�`l�>�R&'���Ҝ'T��Y���M;ǠO���d�'^�`����ɮ7ѫ
� Je*���]M��������n0���n�a&)��;�{��؀���W�ѽ���P��:~�����cn�,&��^N�ͨP�ŋ��/��o�	�<�V7����������q?Wà�ث?|�W���[D3{."%�6��Q��0��=M������'�"i���'�lcb�3�I�O�����ݵ�&�N�",x�M�F�T���*2&A�8C�s��M����7ܤ|UZAO��فL
Ѳ)�D�O�۷�);Dd�P2nd�irS��n�j������n�b�h6�T��� �l�Tօ\^]Pi�R7)�#s ��Ţu�Q����R�-�[w���O�٧_p�����c�}�+��#��އU��Iډ�Ϛ���:��3F�1��]|='�Z�%C�_�������J�`���@�*I#����C��e/!��sGd���3�T��^1J
t�4�97ȓ��f�7.��ӂ�&{߁\R	���u��bx=4�6�"{_�k�{3G����<��8�"F��O�k�:�d�Ic�9�|4Ac�+��]\�����򸽽��-��Ţ�67���u�|�[5�G�e-�?{&��Uyw|L)f4D7�?|�U�&�v~~v���k*�[O���L.���CʎI9֤ə���Ɛr����}aP�{q}s�k�������[�{]��E�-wٚ��:�s��:
z	��P�/.S�����R��]`ߌ���ާ�ܞ.�#�,����f$�Jk>��,���RJ=H D��3��Ɣ��	�-��4g�����x/�_aT-|�y�����J�?6ǆ�����i]�����q�Fe&��fՍ�v\����C(B�utӞ�]E�Ê�K:���r�{��7j���<�smu�?Yة7����U��Tԍ}�Y�<Nd�A��Zb�{G�2�p2�����x'l�����bm v+��Z�����D;V����2��t��Բ'�������3�?�J ��Xд�ۜ�����d�ւ��y@Yg���K�M��c�=�����4�~8�3�T�[��0�*F���L� ���V)�������F�~̮Rn=_����`>�C����{���1)�h~�j�9N'Ǘ���S0N��F���:�5�-4l���F�����F޽;0��E�Z3�jp�kk+�Ϛ��?�d}��� ֶO,����﷡��y�ՠ�����aۖY��y�/�=��¨�Yaa���51
�t2M�b�����>�t֒.i�"�X(6kEW3J�_5T�Ĳ\Ef$�9,5��D�O�~�~ �SJ�SRMq�n<�P�jzs�1�˺ܪ�u�ʂ|�懺�[徴��'��	u��7;�8_�M�ό֊Z�n�=:��~@zK���|���];�OާJ"�W�n�ٳgϟ������po�ݟ>:�_V}	�g����X�l�@砣v�z��+���Q�Ǣ$6�@�Ѩh��&C ����L7�;�[z�m�8����\�oF4�ms�ۈ`��J��:��Ƌ-d ��N�-�d��ӋEJ��;	d��G�(WW	��)@`��@��N�h�(<�cӢ��d)"X|�2s>7����)�Ԉ!bt=�V�{�>��Ɯ�|��۳Լf	l|������y��	�;���{w��@��K���tQ��B!����-�k�u\�h���T8�=ipҢS�Up���E�D!��!�\i{zF���������	igt��P�ӏ=�Ɲ�|K�޽/G���0A�);� #�Ny�97j*��T���[ѥ[�~y,���#�0&�X7��c YHr8E㽚�:?f���ךm���C���w��Q?�QsD�`�n�ry=�c�q�׺A��p@��q(�{����\�S��+��grr��b�+��M�_dR��6'a��,��₼TR1��Í�E���v�ᘉԵu��ʆΏ{:o�u^ �f@�޽�:_J9??�^'��a���%H��t]�&���� �Ry$\XX��m���kk*g����LA�~R��(��JE��%,��+%���~O�\�<pO	��#HC�j�W/Q���o4%Y�cq��Y�Q�T��^���!�0�O��ù�G&s 9GP8�0+X8�:��8�NK_�x�!�������uq�+[oE,O;o |
;���l�Ik�`#sN�z�
�7���L(�a�t
y���g�r��鞛@d�<B��Qa���YG�z8��:�N�>)=�ش{9jP�,�.��`j1�2F�Sw����omm[1�>Q �( (�}���B�������Q��k�zme�mEő����=��O�G@�����>�|���b��&�c3vq�l͚�Ω9���&����Y�7%��}:�g����:��Υ�Z�E� D6s�(^�E�|�Z�ӹz���aL!s��j[��.�g!>��X�tnDI@�&�x���=��5H�"��W#�:����\Cf���v�����f�ڙ�|���Ů�Tas��k�������pz����j&ѣ���p��Z\s����0c/�E�����x�:E	���ϊ4'Ȓ���VU���O8��N�ʳ�l���x�F���ҧK���H#��#s�mf�J	6����x�+�錛� 	_��'���,��|ʦu����B�b��������`��T�p���|�D&z�c-�G�W��eՆ�Am�^\�y���#�dנ q�7������W���Y�׻�e���)(�v@���H�G��&��򖳔�D�)��n��>i��(��0c5��r����`��j��n�+�����r
��� �ݐnӠ0P�M,.ᇗa�+�"�+O,R󦺊>�Se�I21����}�^W�
���_���/�u�H�͋Zָ'F ��vm;g[���%�<�t@AY��+?�^ʵ:�S8W�A�y�#ƥ�s�b�58�m���t<~�(yuS�獼ys {���� F
�z�C�(4!*{Y`f �#����#W�|=~��
h �(=|$O�ܻk��0G"���bE�K�	zQ ��F����`N�zv.p,��D�	�ip,� h���A��Y:�����#w�n����|<��Ј{P�	��' ��(�������{��f�LE6�i��[Z���s��庀�Tќ�D����TQ���E������Ի�S�6���]�=:>;g���?��D�9�tÙ�Ϩρ��\��;t��u���x������'z��c��s���ٔ@��}�,8���=sT@[�+_�]����fԡ�J�� �G�	(+(V_�1nL��J��߳0��"��	[+��.��}1A狹�Y���}�{��� Ҽ�M�rah�����9 ɏw{��1?֔5�D5��zaY*�Ck��3��H'@켴κ���e��z��.���ys�p*�󢛜_%E�ٮ�V�U5�N���M1�蹨5�^����&� � ^��k)L]B.�3��Cs�LEO��P%�Rz� ���ۘq:Nk&�<�⾈�}��s9Q�4����kS�B�!{V���c>O�T���<���J�*�D`o�:�:0�������7��$ZW�
�A�¸ZHa��<������c-�IUUI��kN"�b13�$��C���Eޭn_m�@�ύ��(b�nU�]QH��ZZ���u\k[�[ ��?<<����>9hJ�n�vi���t�GI�2�� Iq%j�}������ڪZ�ȣ�3�ՠ��I*	'�r��}�V@���xH�7�W����y#�X�W�2��aX ��2�	{r�F�������"'��v�)��D�9W��.��ލ=�BT#�1���rP�qJ���y������Kq��JBb7Q�JI?�3�?l��g-��U�A"|���8Lb4SL������j��E�pC�&�8F�Œ����F�Ȇ�9�_G��@�	����,�k�'l*�*[/$���|��._� z+M�b��P��{��?�����f�c�˒�ˎ\�7b�m�/0O��Xe�N��9(����J�q�Q������ԩÌ r�O҈���Vh��Q7*���c����ic�a���d�A�d��[mг�;u�4p
D��q[�����gu�мvn�QĚ�S{'�V�u%�Uֳ@
�jX�z�Rjx,��e��$���D�]P��~��c2��1���ĥ��-2(�/�%���,E:�ba�Q\���>A�:;������ǕN��n
+z�}�/J�݄�/=2h}[8�5�
nP�p��u�J)�#<~��|D�1��P�
�����n�
��=�<]%+ �,"��p�O4���s+2��B�,�e�`��
=	R��|���GBL���l�41���$�������g�>��ڋE�>�3)©��b��ױE�F�o�SkFI�mTcw9��=<���mR��M�֐Jf%�ȧ���A����1V�l4):-������ȋϞ���Ohl�s�T�6u��9��V�L-�=b�&_�R�/P��g�s 3	��u�:�icA����!T�.�6j�,�+$��rtf4s(2'���(n���G�|����I�yP�CҜo.�x;Z��|�&��)q�}D]�MAl�yE�h(�F��xZ:�"��5��(�@�nݕx�R�\<�����w>'�B>ܢ�uǑu��ɭ�=�qE&S�������b�Eq����6 ˊ����Ye����{��@q'"���>���[��6�
����@X�z�q�:��-F-ဢ(�W�����;�',����;��;#�ޱ~
�t����J�d�~(D����o�cv����n�rU� �b]�k{Ժ �pL�8B>�Qd9a�ш�$�C�{�ǌ������k�F�hvu^��ݨ�U������j0�X�W��du���/�{�ak�j��wN�4ݱ�ͽ�S�z1�q��>�+A�!�vh���F��'I�̀Ǣ��g�
�}V�2Rpv%�������8���d`��2i�i362X�І��bӅH���^Z�k�=h.��en0������(�=&��=v�0sP�)c��?×�!�����~j�p�h=�R���&���dA�P��D�]fM�$
��ZϬ��+�&�d�2�i���6��Pms�p*c2���٘ Q�i�8R�J�ڭ�t<��0��)��X7 ��O�	��ƤYYe�3d~�Ge�y�L\�5%�v!ݰ�^;)^�k ���������G���?��_2۠�u�{mE�s^4R=<�7.�qdb���nk�E��Ŝ>Y7?7�]���&��+;5�E�=Sx�����Y*��$唰5���h4�}$%s�i4�����Uɱj����"��'e�Ͽj����Ft*=�X���/���~��N����d�lj���+6<���H�4ԭ���nR�`	�"�S�q������J��U
5(|��Oհޗ7;��D��@x�6�Ak�5�����C�~� p-��A��X�&Ӭ�<y��<T'�e�dGrzr"o޼a�/������Z�m}m��,����ӻ'k��v���.��7��ܕL��fy,���r	����_%�&vvz��V�Pr3bd-�?x|h���b��E����|U�`-bb�/F�PĽ��?�0�!�<m��4�:?n��tl��)F�>���*:�:���K��	��	�ٟ��
븧��tckYY��(kNp�{���j8������#�!Vx����3y������1�veyyJG2�P�&�^�=�s���{RN�tF,[ұϼVd��B}��g	Z~`�|T�,~7g:hq��������^/�����p���0I�ҳx$'��e���B&�#�M��������|��]�C�t�����h����w�!
2&�}����@�<���u�N �k�8wS� ?,Fi0G�w'&��	�+r���(���<(��^S{�i[�� ����G_������q�q �?���&�E�M3R�o w�l�k�#ߓ��)�t�*Ѓ��F:-Ԉ kkr�8?���÷h$ݙeg���,1�9��6@5����a��{t5Q�)��OA����$�ťGY��隣���e�hY����?����_�۷oY�eclc��^^�u�#�� ��u��R1�Iu���s$��#����BE�� j�d>lZg���sc�\�!����X�|�!�n���(��W[U��~l��ǟʡ�}`�j+�OQH���W���X��B����X=)h�<f���:�N�D���~�נ�]�]�}�oٳ�eϊ��q�����+>-�e@�<�[/�
I&��K%Q�$ ���>C戬�"�p�_�ҍ�\��A3I_��0ؚ$�R��Jj��=��5��8���a#;�lP��[Z3�.j/��l�l�1�M�!kyP�ь�Qm
ifg�Է(��!m�O��fr	`ّ�w��]��,zt��>a�>�|�2� *`q�:���6�,�n���§]��T���������>�k��_hz_;����/������Vg�5��B*��[�u�k�I��P3��̠Xr:��Q���i,Al^��ěo�ĦF�E��1��U5�(~�t�M@K%����g6P'��b\�@̖��Si��eg�g�2�[�9�f@H(Үs��r�%���}!IAK�čh�; �8U�7�E�%��M)�b�B��<�\<��d��7��%9�K��#?��p2����V�z��.����])ؗ��r~|&����M2�\߼E�5X�TH�Y7xD��l?�kؔ���o�p�DΎ�t�إ���w{���)�0x�#��}W��y�SC���9�
=�8O=��U��4�a�㳻��H7��6Gi�.�:��>&�ȟӏ��䌺;�ҳF�&83�)V/���������#�Q�-͔���gm�]K�o`�1��l�2��R�-
�o�P�)r1�Hyv�h^����*w͂�m�����%���bq�B��-L����K��?���Sy��s�w�;����?ؗݷ�
B�䄝��A��HS��3�=��+ʪ2+:_���哧�Rj�����\���:��&,E�����#�_/��ur:�G�t���<I��6���+Y��f4Ԋ��pd����Ά!Lg�t#A۰�eP�������ݱ��tVu�nI�����L�����}��,�
� K��,��̞�����U[����,�L�G
k� 	��y֕I�b���ء&�Ǣ�U�j?XJ�6�i4�����B���פ����gR�7ż�&+����"�-8nsut>��x��P�w �>{B9����ٙ�|@��(� F�$�ʲLw{2�0̎@���z8��� K�^��Y!��0����R��jV�[��q\8I��cM�ށ��F�K�C>�~�����KсD�ٝY�vV��)����O���tV�C)W�K1��[{$�k�lԉ�+�>��  C��'JK�),�_QOj\���b�IE[�}��jAz/h� d�N�С��� `� �~m}�u�m="���,J
�LF�e��v d�P��1^��-+�H��t�Efꬦ����F$� Q�����q۾� �Y����� �}�A�ܘ�3����N�ծ@:;�1��Xc���a��:��1��,(m���Μ�7䝹�q� d*S<��Y4���Y��
��<���Z�M,����M�~ɹ�p�r�ӽ�EX9�#��y/�zY���v& 3�\=@�h�r�+hpV��ECN�XZ���"k�q�q���wq�B׽�� �l8:>��s=����F�k��$̈́�o߹s�_��/�Mm�p�ѻ�N�.�@�1
ɺ͗�,����I�v�:9���ȃ�Zz%�@|W�ڣ��u^��$��Z�8����Rt�nϻ�w�H��RaT'~Eq|C����*��E�"���Q�P=�ާ#gԞ��)UHJ��l��_��ƭa5�~ni5�䳹��A�R'S�x���ƚưA�5/���G�\Mjy�c�3)�z��{�aUn�V�6d��cy���:�em������1%u'�̽M��}f-&X@s�:wL(�7��f�\���o��X�gW�o.����P�}�eu�<�E48������o�L޽ݗ��y���|��s�3�7:^:�4�b�,�U�"��Q�ddsGܳ��"0�C�,�5��z��A�����bJ��;��C�;��@?�
�=�,�������O;�4ܡ����z^�Ӽ��q�T��':�C�zUIV;d�W�jM�/޷�x��	�#6�+}���щ:Lw�}\Q'�fJ!��M�b�R	0�t�c�e��I_�.8W�r���UxtBI螮(���QXFdhه!nQԳ|�ew8 B�����!�����m'!�|!YT�nΥv��Cn��\8��ߟ��g�t�V������������������H=Pб�)ݵ;�g}�T�/
�u�m�s� ��H��@�'�RO�����.�E�-�3�g5{� ������ڴ����QeT�k�P���=ր�R�o���n�j�J�=��\�-������C9֍|eu�vr&�� c���:�x�Q�J�ͬQ@#�f��D�lo��z���� uDN�y;z ͠ێ�7�9����|�y��o�#����J�n��cٱ�ԕQ�N]���AM[,,8��rQ���P&��!���\�⩴Q���,@`�k=��]i}��y�~9��e�{2H��W��^^��D�����z�;#�뜨������gH��k���>��vk+-E�4�ͭw�Z9�;���C(	=~|�׍����<=U����P��}ckj��m8��;� ���&x��	�5Л�Ş!]Z��
���x	��U���9a��.�-z����8E��I�[Y�|��G������`�|�jn�`�u:6���%>������y7��B�s�ʖ�^]�s.�H5%u��Z-��}`:V#����Ee����_x{;� xDV)�q�[�I��@Ҹ��ZA��z�E��1�#�i
���GS��D� ܊үs�4+ǧrrt�*a3��Ecw��j^�~�ּ��)u��23�(YK��R�Z���ɱ�}7r� ���{j�M� W��(�_j2�������%h>(�Ba�x4g�Z��	��f���7?7�S�j=,��l?���#u�l��.&�y���9%�f3�hf�8Gj��������m�@ ��nw\=���3�eQ{E��+BK&�x S�⓻�ϐ',Y0gq3'�m^�h\dHʬ��6#撽�����!!7��5`dQ�� 	���y�����j� �!�*�
��Xl&5X����'�~$<a���h,;������\bS�!��Sg����*%�V`��-�`�T�@I+��u;mK۶KFA:j��|�"�ǔ�df�$8��z���R�}�ș�36�0����|R��D7/4�A]	�06V8�x/)g�:�㊢��%{q]U�;c�r���<�Ҭ��H0��X�(�T��u��"���&�bL~/��pXc���q�{�Ւ��6����z�=�~9���l2��sE�Y�}s�H��1��kA$y���y�]A�`����ږ'O?Q�!�'g�^�sr"GGj`Gc��D��i��-�W�2
<�׶>G�����A�s��Տ5w҆#�j#ck睁�:��Xu63���m	ƥ�w�#q��Ȳ҅d�����ĭ�c����";����'M��ڈ�<��_ɷ�_��7;���=�oߓr}[�we<��	L��ʚ���z�'z�ʙ��Ŕ���$ ����?"��_��] hV�X�褏kW����j<l/�s��N�N,�
G�)�p����n�kr���N��Ѷ�9x��!;o?y�P���w�z��e�<���ul�TqJ��!�)k�Hdaa�Y�����WP'�B�޾����	��3Y�k��h�9����4��T���1�17�ǣ���hl���w߽$� 7�m��cOZ[_UG�J��QEK�LR��)x���M!=Y�z%���b�c{ue|�#u�޾�帢��Ǻ���~_�C���}y{v� O��c5�}]ӫݡT73ٻ�}�v���T�T(������Ɩ�zK]�E\���5��VT&�@U:~���� ���M
��L��\L�����2��5�\w�Q��p��9�[eE�QS6�q%#u�u���D#�Y'8�]���u$��P����A�)�j�۫%���|U��k���3\eFe4���2P��V��P�z���A-.�kM���.t�݂�����#��B�8c~��fB���$n(��2)tҲ�҈����J� %�MB((�;���I�I�U�޷$���O��+]5�E�lG�cfjX�a(�����noO�Ǒ1�t����Ե��\DX�B(�
�Sm�te�۶`P>B�[�C��W,l�:��ӄ��D2��'�d|��ʗ���d�7��ܸ툨����-"l��Q|^�:w^��˓�η��Bd��wǜ6Dj58cD ��w��@����i;���Ѓ��G����ESZ�݀�x� Ѵ0!f��J�q�����b�!��U8�q�V7�j� ��V�?a�jDz
���B��,�D����x�����z{З��� ����ݓO�!�wy����������H@�F�$tA����q.3�%wa�4o*F'������/Θ�x?x�@����w��C�acu��9�j����1�kw��=�޺�zH�b����x�n�m+6��S�A ��aC�1$8�٘������(֢tf3��h73�K�Z��{�߿]˛L��ǀ�k4 @��Y^���7�S���H+��ۀ��l�&���NR�C���p����B��m�x�4eq	�G�� 0̧�g2y:�����?����:96�BQ8�@�;�~�c�uS��H�7�n3�}��'Rנ��Iý��Π`!�E�眵��h�GX$��Qoy��Iv��<'�>�;{�������1����]��\���N��́[z2|��(R40P4�z����}���=ܗS]룙:��F;
>���ޣ��Zv���K	�?�1���U�&��n|�,L6lɎn�D���Z6Q`�[� �ޝM�]����gi6�t�@
6!;	��4��P���9�W�k����ƪ:�;�ǿ;����9U�p�Ř*{��dmc=�m�������ӱZ|�p�r��v����ɯ��פ'�y�C
YY�qs%��:�1�hɄQNP��c�Rp��8�ɀ��dpMy�kM
��^�u���7��wҲ5��P'�x¦�&��Qm�=Y==_H'CF�Y����U%��N��W�� ���A}�~�Z�~-�����X��ĸ����L��u�����C鮕tĹ�ٚ�$D��L�cbM��������$������zz?�$��uK�[�ll
�0���^2�T����-��b`j��=
�V��_��7�W�5��i-(tU"�����ܹ�H��������B�0?Ƴ|��Z-ۖ �Ѿ�,ؘkb}����Ѩ��TÑ�w17k��M.8�m�xϠ؇���������g=� ��G.���5<w���>�	mo�l͙�.���T�ܨ3;��n����R���g�I	Y�1_x����m���7r^-�B���Ǥ�'��ڐ��KR�ڲ�D0b2��q��A<��=���P�0MQ�Ԙg�"g�#
+�H�\aо���*Y�|�/Kω� 
�.��5�H8��.:�$���Q��IVD��ky���V�H�Q�|oM�Y�~0�7�Ff�Zx�j1�͙D��u���=�����v��Rafp��i����bB��h鋺6�:���4���C"����g`�a��֦�E��n���s!y�c�z��MRvi_d�Qg�CZ/ۆ�F�E�����K#w��T>�+O�>�M����grpx"�vu�8�������{����W�)�	�R-R�)�"��~0�Z[��KuD�X���C;(/?��_��{���_s\��ru���k����񸺹dt���?�O?��i��)�y,ߨ�sxp���ֱ�����86Z8���D�,�1��ZƵ���E����R�J8j6�"�ܿ��g���~.�y��_�]s'6�>��.��yQ�2�H���E�w��RmXќO��Y6� @�,{��nO�.��Z�4�ڸ؈�|��y��ky��{y��nڣѹ�~+�^}/��{��j2�-R$����H�b-
+ n%�n��ϋ0R�8_�\4E��mӋÙ�K�]$,c��j~z�H|	)�~�s#�|��۸U�m��(���uۘ�P~2 �QnI`#���ٰ��}36S6^���H�;6��ٺ+�֊L�m�X�Q�R�T�@*D_��1�[�c�5���ҹ:��t���Z@��s� ��ÓO>�Օ�o&3
t�|ΘiF�i�3�}�|>���
��k�ډјԼu}��7�2�X��_~��y���G�'7�k9�<����k*���*�7Z,Ƶdv[�V�[��=�3�T�曗r�w�>G-'Gg~{��~�M�\��{����	��*��E����zxGV�mܻ+W��ad% <�Q$;1��X��.��+�A������Na
�`*��A�4,�e�� `��.���������G�t,����=$nt����S[�+7���qG����(�Q�{�^Q�����U�5�
΀��c��S��.��mN2�9���b,�X��gi-�!�EeJT��j��fݿ{G�n����Q�|,8�!}�h�^ưf��?���c�v�#�|�#[[r~vi�N��\�1�6UАӀ��C�E R�{S1wG:�s��@g���)�,�lB��_6=y�B2@0��U�9J�f$�S45��A@YE�TU�A$���B`��пC�p>_�߃bTu{BM��PI�������(kEU��H�Y1_|^TU�Yʄd4�V\����(�JWɋ�P\8�9�\Х0�)���T�4�ձ������3�0u�`����ZcB��,���)&Tt0�-��\P���[ZM-�{�OD��?>��?+ګ��l�NЎ�9
��
����R�EV��ͳ,�*<�k pv2	c��m�yQz6��>���f����@���5�	{������=k�F�2H]e;k���Ѧ��Eʜ�es���݊iP��MtF/*��]
߸fkdo�΋�;{?>��-b�"�e���q��`	�}�(d�Yʆ����^�VE�Ɇ1�چ��c��O�J��
����;��CH�Vn�3���-��jD��x+	$5��n>_Ƞe~*�1���5�_Pd2�!8�N}oHP�H�D�[����|��gO�'�������D�v�힄+d�'��+���b� >����ݮ�j��`=��Pש�~��2�3����e��L������1�r�O�V!���51��5,�j�ȇ��P(�k�}�0Nչ�����Z�%�`��U6�_x��� L�` �I�mҗW7
<~����+�~�]@䒴+��z9TNr`NќY�)��#�yLD4�/Q����=v\	�`�u�p������\�F"���rP��Q��'e�>�'�~���H6_��
�u�9[��}�����F��:�{��
��kdpu�!� F��.մ%3Ԃ,
R%��E�^X�kQ�Z}�)�\!�!^h�M5�5���e�Z3ubt��7��������󋑌g&s�sn���jDu��/
o��13���hmsC�!�u�u~����ڍ�|��+��Y}���&`R��$(�G���u W7�I���n�tF'E��ڗѵ:V�-�w6�]���r ���Ln.u�!��IS���A����m����t��A��h:&����M�m������-�ș�����j\��ȀT��<��N�.�,�!ܡ���*=���&;��Vd��9�;��k�D���:Q���v���r���u<��
��U)Wa��Jkm��k��
>�ތ"��r��v���2��!:��{��dk��T6��g�o�;%]]����t?}H�p��&��2��D ��cD�b���9�8*�]_k˝�{r��fh�8��Wrzr�l�x4�����\���'�I�X����U��?�aS6I8�ٯ2�^�5.���I6#-�<��=��/�ť���������2n]�/ 0��&jU4���c�� |0�}2^���(��$���	)YѶad@D�Z�`���]���T-S#%���z_αI̗����6G*��1l���u�+8�?8T���A�~�j���QE���,�_; ��_�����:���4y�����?��1�Q�n�ͯ$=܀����G��˺X�)��0��R��5B�6+l���-b�F��ܩ���1��w�o7'ɝ������8�8'�ζ�V <�T��b��t;� ��� ��p6�O���才��k>*Fc�6�;�L��̱�V��Sk�ğэ�;��f�t�յ�Y�����r��"uK��p���ȲQ��$1q��D�Ǐ��ӧ�����ry=fq��:f���1蚡NQ�0�f�,�Μ�ۧ[��t!��Mg�Ζ��A�ǂ@
/'�� ��j.0��1x��~7X�ђ��󿶶���5����j6�L+�o(EDP)X|Z�BJQE31���N���hGټL]��QA������-�;��u�������.hf�3�k���dE�Ը+��>w��8u�������Ҝ���0jc�45#��-Ay(�&��խ��NYæ��w_)���~��mN
���w������`�]F|1�W76�҃"Z�B��	j�b��;��!��:Q�j���ہCul� )��Ϸ��M� )�ɟx�N�{��±�mPi�����.��|}g386̢��6��z7c~�v	�Ҩ�p�j�9d4|ޕťڽ)28�5n�=�:N�F&���:��;���2/n�`��9�z��5�CY�L��*u��N
���"˘�Y���)\t���rz1���uS'j�T(������h��~��y�Þ��T��	J��3y{�Oj�Ω4�Ȃ!l>�q�������?�mS��膭���Ʊln=V�lK���tF����V�@}ot̐��c���c�S�hS5�r�
B0���cZL�ζ�ײu�b���]�R�����+�䆤-v����bh�c�/GO�zѕ>�Ll��~-�V�I��,����ޑ���䩯m�0 �������E&ʅj�?���f.W�3�I���e��-��{2��"���Yc���<�?�>P���\X�7�Qh'Z�IL���L�@I�'���=dA���1(����R��]�d�g�M	8��q�������O��a%���ɩlo�aSK\��#�57D08����*-c�Ǉ�s�I��D5˯g���q�>ja���!����B8tֱ(  }��k@�{�5����y��AԽ��u��+Y�?j���<���LI�泔�a#��,���.��+ೱTes��:���_ɳ5�gC�̏eY:�A�u@w��,�٦��pΌ�f��˗��>:<��g��]�AL���̨1VCSaY�1`m�V ��.��XCC����*-���Q('�}�(�({k_b ��/�@: !p�Jd�(��G��}k��IX���)埃I7/�l��̭G�-�AX�7�Pv���z�=��S�h6.�>�]^�l� ��u�q��!c�p+9�*f-Ģl��\�E������$ө�-��i@iP���]1D�Fmax�Ȝ�Dy+�k����x,�}�XE���q��� g�Ջ?����X�t���1�|y5���ł�.��틖�+�9��^�_�*.�Y����SeQ�6��~+O�<�g�~JCl��p2�b�gϞ��}F5*�V�t@��Jڅ�{�˹o�J�Hg��I$�5��\��)\5�� �ҕ38���U�0:�;��6��ZIA���H*Ȗ<�2��4t��M��u��b~�}-�������9� ���fuf�+u�-\�1
�>vKv�kҔc�(T�d�'�ư֢(H�����!��wxBI�#Ԃ�x΁R�Ș���ߨ=����������b�@�99X�2�fcPS&������t�I"���k�آ"$��[,��ָ����я>C�[�[@A"Pg�x0���E���%�_��E���{;��S�A�*��M	���O����Z���t�D$�jE-HF��1�Xq�թ~�R�u��z�=�b�
Z>Pk��A���"?�;���ۣs}_k��#��_#pՖޞ��O+u��zԂ]��0�)4r�s�j������H�ߖ�n޳�%c�<@6�eM�M��wI�2���?b�jP9�x�`�Y�z��/��<��V���c�!�����_ g�rr�����Ԩ��׹*�:$�7j?�(�P�|���j4�/	M���܇
��{�Y��P��������A�Q�v��B|��e5���g��Vj{W���n�z��I-����T�jS�ޖtV6ert$�ʆ<����?�?�ڑ�ڶ��x���� �l�սwMqt�n��R������Z�{d-`5=2:=�z`�u=b�F?����!����O58��H�~5�O�������Ǭqa���P����a�T�1�)���# y���e�8Ƴg�*��K�G�T5�w[�! U6V�����ώ���s���ӵ��5�հ�S�C�����p����-[VY��۹Q[G���DZ���b�HM�: !Q�>o;�*H�G���m{ �j^#PPc�S�2��Q�̑t-:�.���r�s�k�!���%UصP�L��(��E�|P�(xQ�Ib`�}ɸ�[����5���ҫ :��:��$=�.�H9扚�n��$)G㱈��h�5���_��Vs�����;b���Z���ۼ�%||�������DM��7�	T�ME��?�VL�tˇ]4�뒃?���
1P�M�)��x/��G�|#�]�OD��q��7M��X��y��E�R�._��Q��ӥC̔32��-�OS}�p0�(��3# �����XL��Eޔ�Yz��{6�uu�2�%��G�ƪ��N��=J��LJ�馸��)=cT���ģ�t�x��;������/�'B�%vs �9���-�Y-���O�t#D!��/�������䓧����#�A����*�[�)(�c=��y|rB�q^]r�W��`���7��Cq) �����ݣVa`0' W���\M�j�$XT-(w.����ሩ�7��g�}:��n��,��������<�3��k��,?�K�S�g�vq�|.�q|��鶴�����ێsat�z(��-�w�Ǒ��bʺ�jQ�t ���ã�P���2Pb�s��Ǧ��up��z���%":Y�0*�J)_�Nʔ�~��lU[m�7� b��*�,u���%�����pYi���8�w�>�d�#���n^��v�E�έp�c��p�QwP��Sq��@Ҕi�t�O�Y EՔ��H�m�������2�������KV5�.չ[����M\���[��J8�b?�N�Uиq�*z3�?��&�)e2R'r��+�'z�j"��P^���{���t��p�i���t���k=����@�Gj�W��x�,X��)5��:N��F�ɀ�ڍιKfV~�9�?~�#���	�(j��tN��Pl��I|��װ*�b ��UY��P=�\��s�`E��Yi+2jK%Ӯ|��B�<ҟ{�v���2�����2�(0P�������F���u�mu���+HѱDע�Ԑ�ԋ
ſ#6�;�P�s�6��L.���}�G���W�x�-/�zN�Է�ߗ�����u�ޑ�'�˕��@`@�N�� �`�f* ����4�N�Ǽg�F�¤�z��D�� �tL�@,�fCm��py�L�*��:_GY�#�kD���oV��;��k���B��	4LD Y8�Ȣ��/�\�,�Q�B����X>y�o�Z�j=�yz�����)���
\��_������F�Q��6WOm����6L������1S4,��-;�!g����g�
g��o�(si�9���E�˳ᜳ� E����M	�>??u���Y�y�P'�>hP�]-�as`�oaN�_,Q흆쵺&:�J���\q������my���ߐc������S ��e�~����T��c�}�+�����B�<��ڙ
��6E�R����
��U�k�;����jy���A5�ς*��͵�=4/d=\������G��ࣳ��e���s�|���@]�*�!i���H�V���ߛB�4aQ�T,���i~Ʀ�2i���;s�P8̎�������|�\��~.���&m}^�X��"th���ހ��
�5F`��ԙ�;�KLNk�N#��sS��-��"�P�Bq\ޖ#�]l���d�Z� F�/�6�;�=�"!P�@��Mu�Q����s����Ƥ0_*��}�V�ή�h#31�&�ًx�TNYμ�vM)|~����QwQ� �E�����_�\.������������~��8�F���n����p8R������~Tċ����_ċOk�Z%�ь�Xx��֫s2��n�O=�A��5eҞ<���#��r��q0���|�����o����/A	�BH��ܼ���
Ń1q�)���}����p���-�ax��jG�ֈ1� �f4�l慄�)L7�E4Ǭ��v�h�����FMw/��0bQ��t�W]�+��mи��ԎH��</�z�U�*[�̵^�U�U�l1��u9�qD��dt������Ɍ��ᾜ��Z�	��pk,@�%Ѩ��B%�QncNV�h5��/)��c��?�^R\�4l4�JGYKD�E���$F�ʒ��	w�"�j�݋Mc��-���ɴ��<���z,mΫ������KS�?�����C�U�FIW����{�ד�/�[ܳ}V��,�?Ǣk.��%�63�|~��H�,�^q(�dl�G�X�y��9;�w2l�Ť�0�A�z-��`��hu���l��ݔN�	:��8����Q���ϓ�XӖ!I���|~�d�yZ�r�^?8����Yr
��F ���_Q���b~&�'{29y+��������99����.�sfC���$�c:H��`��\����L���|��U7�o����4F�{IN�Һ��������MV�wy˟6�i'��b"ǧ��*��ؖ��-.r�����l%9���s�������̓A߱�?�`M��]��_�T~���L��pr���"���l�l$g�FfG����ŉ�wɡ�Y��і<;Nr��D����d�b�$. 
����� %��z��g�v��azs�&#DD��J;$=� �YtXICf�f��a�;ۗ=���J�~�d2\��	v��^?�گ4�0����R�߿���8<���B}�2x�*ˇ��O,(9'�7>���E���Ç���n�y����	���y���ݻ7j��Vl�7\�}��}�{9!V��+�����p鉏���_�i-Y8k3E� ̉6Th��O�t����n�.��󰸷F���7f�7U�,9���鄆�7�Ŧ�dX��ɽ<:k>���۷�uu݁�eec6 �5��[��-�$\7��֞:��b&GG�$�x��{y��]�?�t�fF���(a��6C�7� !|�$.
'����֧jB���V��dێ�xwF�c���2Ě66�=dD�:+�_�s���&70a��la8�e�ݕ`���d��X��׻tOr�N�gܔIT�!T�չ���L����~�ͯ:��r��g�Y���>F�[�S�/�!ł�ޱz��v(g���-u<$wk��az���m6sa�5.JQo�%�;�z�jΜB���[��}O<�X>|��������䁿�gO_��\�a �Gn��X��ft�i�D���DJ��=jl\��VI�v~>��߿��;����O��y �>|���Hk���2	��3ql�3�1���dz!��)���S۫+�(�IQ����=6nB�9��>� �~���m99�H�|�4{��}����ln��A�~���xC�Pɢ�.Di�A��TR/<�L�yo� u�w�N��*=��w��Q9"ѝy�;���92W��� ����bu|\�'A���^���j���p�zɾ��Y�{F$�E��p3_���b�"��<�Ȉ!S�i2�f��Q_G���	�4����هk�����X�1R	dJ��5*ؾ����	+@=қC##��s߫��+<tRK����<�`��Hp��B��v=�]�|��/��-���ttKϲ�j/�e�)��L9v�/�f�-ODະP�dt��b&V�dA��s8��i�n�t�i�N���p\��Vr פ� ���8�i���"m$��*��WdH������q=�x�I2ʇ�I� vwO.��|����٭z�M���R�WP@���t��ͦl�{@�j;�!����B̷2O��$}��gg�?�Z6��$OvhxOЇfuC��~(��-f�Az��|�oݕ�r�0Fߟ��[ې��ǲ�-�A����'�mrJ��!rpq�~���&�h:�i�mr@�ek�)+�xo<���h\�䲍lR�|k�q���HNZ�	�����ۙ�|)��=pz�F���6��L�$Sf �+cN.Wd��V�?�wG铧+w��5��3:��
���6`;�qS�j���t�i�h%�N�R+�ZT�^K���T�:`��WY5�m�����n�¿"���{�̀�| "�	A����d�n����MALв/�L.�M�VXB��?4,n/YK�x2fC�O>���lJ�}42|�bv�D��-:;��y�V��X�ȵ�U�CT���p&n��M�����)oU2��X0�x��'�09�.֯_�J����T��^�W��E��em�db�Z�D����gd�Bu��Dq=[���#kt��z�!���ו�#V�$}ԅ�^�!�j�^.H'l���u���a����^��7�����
���,��������իrZIt�Z��Fl��0�4�:�dr��8ƌ�a���,VW�<CS���kCt��XY���͝���0�ʆ9Q�w�F�=%�ڇ^8f?V��G�^����Z5�ꕵ]���lnK�N6¯1��A�~O�Q�kW�M����'�3�����X@>Q%m)�|󘱑;/:�s)E⍎���Tg������E]�Z�7XĊ��� �w�A/����������`�z@��˗��??���}�<��Y�vR�2,�*�;#��͎^�8�$R�.���l���I(�r�:��� '� ���>2�=��0����DY�[�v��pA��	[�[���`M�ݻ�b��$77�AB���㏨T PL�1��i�rG�:�Q5)�!���Pgs��d��p@,Vr̽f�<
"̄��A4�Kg|�F�y�!8��fI���9!�
�����c\�9R��n)��_�,w��u�$�8����1�v@�԰2���E��qԃL Ƃ���Ɂ��*n��:(��t7:�N�Bc��LY��43�X7�E70�5mX��פ��d�;��Fï��-���h.]>�˨3a����j�\�S�:I����841�.qc�U���4"訆h����4JB���"��j�M#t�ȕcE�����Uvb�[� w��F�م)!Ϟ��\�ܰ,r��� �i�>D\n�	5M{z����Ø���-wAi2��k�w�.'��x��@}� �M���7���}:���4쫃��E#���W�$%{#k�(سٱ\��99��jT��|tK.�����I2��Iά޺/+��6���<d�FA�u��_�x(��#YLΒr����Z��H���6d>X�Y�&��3���R��[���Q��G8f#��w���ޛ_�(	RP�F�Q
t�w�?]_MN]��6�1�!�v△�  ��IDAT��6�dԯ%Ù3�)�e�d�8ov����t̉��X���	g��Wgs�;E��Z��q�9�#�/,�Mc~:	,Z��Pnl�����ٙ|6gS���;r�̛��Zyi 7����FZ����{��!Y��9��Ҳ�a �i>�}m��W֕�Ѣ�܅�A�%�AR0�Y�_�+H�����3��.�xq,��oY���p|r$I�@���R�uD���A��ӠGqԚ�?��;w�}uu��7�*�����{%�y��
54BAZX����EaX�LX����	�����\���ߗ_�����S���_��_��`-X;c18��s��9�`F�u�х�A=f�`�H�2i�$�
(�����[�~f���)��	���(�-tP^�!��%m�/����M�`S���ZQ���v�vѩ-�O���y�}�V�NN�|�����tj�%��h��X�
:]���WXUgN��!�&�����Oe���Z��9�Q����Ɓ�@zks���0i{�9�r��1޺�������|}Ȩ�b�c�}�� ��h$S0V�=}�<��[��9���Pgُg�נn��m;�Rd�:���J��N�\�d�}?w�8��)#�}_����Ֆ@�׃K����)��_�y������w��Ğs�ڐ4Jy��&�[7eg�|����=���{.߿|�hr2�T��8奙����Ç����s���x��=������{��0�@���rvr����ٷ� 1=��سg m���3��W_ɓ�?�G����lF�� 0���>z����_�͛�dSZ,.ҹ�Pr"�g���↜�$e�&Ő���5v�]e����I$�Z����#ee��`:>�H��D:��V�� F-SԳk�`��o�,�w��|6UJA
ϡu<%�i_�Q0e��oF���7��a
Aq��RZڸ'�e<<cSz>�)�L�
�p�@����(��zژ�k�8ˋ��9\\�[��(��i=�`���k�����3��rz
��1
�B1��9�h��qAdwo����5͎�.��,Ugv`���l�Z-Ձ��v6���	K��Mi�h�k��M��i���at�.N��g 9�A�kn-
��tV4����P��VR�f}4Ȃh�F�bF��<�!��S��H�Tx-uO`�=28��Pzp�d�Aax��%K4�VBjܦ2������ɬFia�a� ��sM���*��x�������v�O6���$c*'�3s 3[_cO�Y@S����f:^�C�(��!��Hk($��܇��Mky�=F+[2Z����dϑQH������C�PZ�Sjhny'��2%NΒ�9h�`����Q�ލӹ�<~���B�l��5�мX�#�װc���ɡ�%�x[����t��4gr��y�?{(�e-�l�H�'�%��dp�;2`s�Vøo���Ck��|��/2[�u���:B�eӤ�m	���X0(���?0`��ơ�yc0�NI<bN!X#�<s��2 ca��������b�պ+X��t��swL4`��o��F��_�K>���ƍBw����G~���X�<&��;�,�\��	3�/��Pr��m�q>��yҁ�����=!%��掼|��R�^N��C	6y��Lma�ÿ�[*@i_�5sYR�����3��A*�W�^Ѹ���M��3�k��t��Q.2nN�K]���\!Y�� �i��fu,"�@7�Ve�ʈf��s=�uW/�w�;M�}8��:S���5r֑��~t��YXB�Z��0�>-s����9��*�Y�i'�Q2�L+�;R�ӏ�Vߢz�Leg7�\B9�h�&V�ƂZL*n�f�:���GjPZ�S�Y[y9h����/�Ԕ�GS2�[M�ã_�݆�8c��B��-���{���ڭڼv?�*�7m����&��ح7E�z��u���AH�щњ�XϮ����xWڞ����&�{�3����]�r͵����3V�� ���ێ��Į%;)�ZF`��~<ސ��?��w%�����ի��x���o����k�'��z6l���Tn�{k�_1_�^S��"��h25��L^�x��W�������$�/���[��_��(~g59�$�'r|tLa�ZҮ&����Ha5h��o6~��fR7���c�8���_�?���JNȇ��/�̎��|��8�qrF	��=��4L'��A"��a��{5�#m>��J�ݪ�JE1�(wy���@��������L�c�ڇ֢43�n[ ����Ҍ�SKS��1Ns�W4��C�,�@�Ѧ˙�!��&�ڜi�ݖ�����xzѴ/$�1g�hM(�s�/�F�۩�	����:K�B�{�V��1�N� F6�RI�4�sҸ���l'�~�es�3t�G`�R���±irCT��fh��H�_h$mA&����rp���C��^� ����?�oĶ4����"w͈����� ���.)����Ӛ��Q�33ʘ%�q�a�S�BVj�b��JF���D��V�ţA��*��FZ�s�9@g`6�j�@���Us R���ډ�	��X �9w����B��V3�8���4uhPQ7�L�8������v�ر�<��(��)'��ddU5g_�tb��4 9�r٬��/�-�>I�M�9��&�v�$9��$u؟��� ��9��%��������X�#�dd&����{���L;�� �7C��u?]X�:�f�4�qh��.���<%;]��\��UZ��;2�.�D�!{�r���Ӝ�!��i:�e�4�b$���+�#� �%��,�M޹���ø��;t*;����l��������	aT��j��[u�EF&	��Q��G6 M�u�-F�r��8C�#7,g�U��ޣo`��I	��ײ��v0C����_ʟ���<��|��c�''G���-��W�.�kҸ�%���]�怮�AGt#n�N��}�\@��x_.&r���}��◿�������F]�27ڞ0G�F�a����w�T�R��k>/��\���Ou/�ƫS�6֦fw<��5��5�icAG+�Մ��0�skL�*��'��!�+�Q]���B�A���n^^�r��nu��I�G�sE�5%B�J��L�1Z�hN�Sk��#�SԞ��c?�ٻ�w�)���L[38����a���i3�V�q=��8��֜����HtgD�"S��uO�,c�.���;^l��pL����Pȧ��|��n}r�֣_)ܹɘǨ�H�!�V��V��������pb䙎�]�j��Q��bvB�!�ъ�#׻W�����M���a
Y1K�<��hZ��[�E
tib���j����>�Z.d��T���*VEZJ��r�=6�]�QO@�o��� ƴ��)�;7�ч��Q�@n�|�6)"0��z�V޼=���dj�Hp����ӷ�
�||[���u"��Ux���$W�L3`/_�#���'`�ڤ�==KF��I2�n%�9�O��H��1����$�aݾy7}�F9��n��@9�����������g� �۷��ӗ��������-�]��B0v0��޻{��\��O��lJkk��|r9�1����4��p��7�<1��N���|67!X"�H;� Ц�Q�!Ðl++���7�s4��҃qz��&�Y�By_$GC��+J=W�)�{�ѳ@r�Y�N��"��l��*�{g�����gxN�����v���$9~g}mE�J&áC�98�t��0��L��8�Dd��9����y]h-��)G�C�4L�=�k����Q�s���=)�@Qҵ����WH-�.�	F�'�9p�xM�0�мe-�C9�[c(J�%lr��W�[�B#g��S��J�l"��Q0��fʼE��)��Xg�;[�?\���j8f�L#�i�נ�1��"b&�	��.:$��I[�o�G(l�7�����dSqκt��	����
^X��i�P:�F7�;s�J(U�x���
P��&��f�	i42PE[d�1
V��,������Zi��y�io���{H��~�	5���Gq�����	���� d��2��0NƾfTF��T����F�pv 7$�'�yb����g!�f�1�tvܓ `\�~�#%9Hs0B�<u��k#��p<E��.gq�N�̎�l��Sd$/;R���j���?�1��7L#��>'!�i��'��MS+�6B���`���iuF�$�i�>[�;`���qaȹ�x�Z).=�5d��<�Ԫ:���}����ծ��?Og���B��ߖ?|B�;����|��7rp��~S?��O�3п�����=�0La0޹}OV�a�3�I������ɓ�/~�i����|'���W�����8x�8�LF��x݁X�:���%�����s�*=?Ji�KX�����Z�alS&�s����ό�?xN�6\1�cl�*��q�^<á�d+������Ef=Y��N�ߋ�1r1 �cA��F�}�w��]�{F�\mnJn4��C�@d�P�u������l]����P3��ls�����{��Â9�5�A�ƞ��a�V�떭>���쑲�>(�w�d^�_�t��9w�?��G?���{�hZ�3�BWfCL����җb�_]iˎH���O�Hv��/��h�
"m|�1����fw��^ZWQ~TS�ɎH��E<����F�T��V���92�	� �:_B��e	��P����N�B���Ak��P�!�A�[]IoW�Ks��q��ⴸ��_�U�(, U[[7���0	�Gr��B�vwO�������Ϙ>��1���9N�Q����Xe��?;���&�n�G���i1�P1�����1�]�������Is1����#��O���C:^���p||��
�;��r�&C�0	���p�9/�I��]2�r��}�}�6Ϗ46X�~��?���o�o��`�Fp�3P��b(7w�'�&~��g����l�l����9R�ә�� ���t:pJ,%�(1ѝ�ی��Q��
euxp����mf��rxx�b���o3���ڥxwx0���QRp0@)'J5�5�������12F��5a�1�0���� 	�b4�Ҍ�`\���Q��q���\�\�1��တ^O��er�'��O������ �iw�ڦs���7l��3�L-�\%����B�|B�V�s�ɨ�%�dT�81��:,t�e�#,��s�XZDgqN�!ω5�#�gT�����}�\��$>|��������|!01��<��@��D)#���D��qY4��c�k��Ⱥ�bmv��g���\2��rH���'6hFc���D�n4,��x���Og������,|f�f�Е�8�DUyche4��?��3�%������{F6���Ɉj�` 0��Q��j��]�P�\[�5j�Ao�i�B��d�kBĠ��n��!��j�T$�=�,l�r��.�����ʠ�k(�zȠ6�Y{����d�@�ٮX�1� �٣9#��]'��<d��?.�*���]�:YM�膚�Ck��f��}o'N]-�'�3�
�U�<D=DԚ@b3�k�b�T��yc��{p-T�6��V.t0؋ �p%х:�)�e1���sӀ���?�A@� �trt	��2� J��\?��u(�߃�� �Y�?�I���=o^�˗��e����f`�<=�g�Rd�q�7�x���#�|�P�2�n�������Vƣ�$��Y����[��_�F�����n�@����Xzu�b���M`���m�s�߯����+�*�����]/��rxa���i�ә��~Ƞ(�8dF,8`��lc����J�m�=�4�����R/�Ǧ�L����6^d6],�]���c}9es��jM�D�6t01�_R�f����2mr������D��j-kL�l�u2F�t�CQ����Ĵ�^KR�qt$��f�=��[oE����Y���GO~�-��3$�r�P
2u�4E.�������J�AS"=�ß;Ԫ�]���z��"�7C �n�h|ƶ Ȼ+�W�R}�8u\��ܣ%&��<�Ek�X�р��0�P��t�"րD�́6�C������	S��Ǉ,VEQ�,_/d��&1\�°|�_�>��E�����+^���!�ܻ<��L��2��L�l���=y�b��wo�Y�4���+�(�#���^xZ���r���������ZD �e]S����7��2����~���r��m����Y����~��.���r*�m�"����7�_Q �x��-��~�����7���ϗ��x&��;y��Sy�.9����cڌ�d�_��go���[4�p���=�GkE���"E��E���eo���#�J�Wq�X��ܾu��`]p�7�5ooo�c�
,�p|��"�ݍ�tϫnp�@?�"183o�j�r��t��t>�����b;1��;�&��0d'��L�p�qc�)r
R��������c T�4�g�����h!;���&	�cb���Pks 'i��1z5ZQ6��00,�Fq��u3˘yv�p�	�r�B��e��F_�S峙����)�����t<��܋P?d_F+̒�W�3���Q,D1?��3�g���f78x�[v�eeÚaded)��c���<�fY�O�f�"�Y�5����ŬXg��	X� W����F���+k�.3iS��#�Ҷ�&��⠖ȶ4�w��|O>2Ufv�a�8k�tw̄�!�������g�^}~:��n"���X�O\3�0ubʲ�?��,��d�z21��w��h�h|Tb�L�bAȠE��D��P�ld�V6�Yp=CAqt�|��>1��}�?�;�]Ĺ6�EM�l>j0F�BP����_d���"XQ%H�`�F2�(��$vXǬ1̶��(_��1ke��~6�T��Y�f�6�-`X��ozjM�����W��	�W;�Z�)��w"b֋|b��lzɀD� �qkP�lp�Ȫ_+v?ּ���A�A��A���s�ӟ�%�$������?ON�>e0��1�r����T��uS�++� ����Btp��7vX��o��[����o��w���B��U��:�O���NS�]�Ng+,·�um��\�2\~���C�;�g;��4��E�s}3�^��rv>��rB��w��!�>p�:� �3\���t�V���t.��h	��P��.î�sA>&-}�N C?A���pa���&�M��Q�'n�{��� 5@ M�J�U�f9�NH�,��
f��vE�਺~;aN:�A��a���tڸStO���|loo?���g_DztV�<M���T��#�j����
��d#sHCo X�#^q<L�ݢ{���wl��as@|����.{�]��7�S�{E���-�7l'C��B�(
��=�?�qa\������O@�փd �J��ׯe�`��U`щ�Nc���#	��O�e�x�VL^��sb+�޳���h7�Z��'̴�4��) A����NVG��>�4��M.�(�������X����\�O�Fj������B?)�	?���$���`9�^�Qh2ޞ=A��Ay������U��ֲ�`��t:��g%�k0|I�׃h����o��뗲�w���yu�F�����7`䟬Fi\޾=����ߧ��1�P) ��T2S�����Fi�i�F�ע���w�����qqo0z��X����ㅤ��X��c{�&�k{4UBg����v��ƋF��H�8�qά��]vQŽ�Qz]��Q�)#���ـ�J��>WY�N����f:�s��(.&�O����GA������h�Mw�����ta��^B��J��28�gg\��z�@w��(
p����0�`�P����������sGG�I�}�}p�?����?�	���w��"t��]�u�8�y��Y�����67���5D*K:�yK;�B)Q�#��	P6v�M�
��3���^��޾}ǱDQ*��
ؙREo�+;Yhsk�Y(�@Rt����H]�b�!.�d�7����L4���B)�AA���0�Pj[5���D�0�O�{%ϟ���K�5i&�E	����S�͝[F"zs,�<gs�1ˮ/z⧒�禺*P�hefr�N���.-贠
�4vS{#Pk)�x�E�"�J?�H�=�f(��,5�� �d�qD�q��_p��M4��_�M+��ɜ�*�+(]|ŷlب��-����QT�o�,f��s}#��Թ�I6ix���!�Y�΀��g�S�c��b���+�4"�Մ�s;4=�&��~��M>f�h�|%Y�jq��Aay"*�0�Pk������������)��S���?&�-�c�������ή�0�vzv� 0��RA^#J9����ä����?gp��/��w/Ғ	�����'H�{�ྣ^Y��B�=g�,��=8���s�P��A{��앜>��	�ˢvT�����k׊�r�	4�'��Q]�PZ�j��;��C�yv�3-xO����xB�:ve?�ܦ���昨�	�aЙ��І��Km|� �7���`�-�Wu��1J^������X8�������P
�J!X��ųvMʄj��9}2^ۤ� ����}!ރ��ƛDU���?��Ï?��_Y�f�4N��$��eGcY��e\�̛ҋ+����� ��I:!�ɱt�y�~��6A�e/�8�]�����P9!K���O#D��o��b$�9�%C��Ǐ7����K���ݻ����8Ad{}m�Q��$`NN�&c��������~Sߨ�|���TB|B�AE�?�Bey*�>���P�Å=`�B���֒!#F&�Ph�4�|��T=_-��BV�²��_����/��������d,O`�!�A�ctr!�~��ß��л�-�W�ś�7i��(=N�ߝ��) 0��X!�����md( H MAT���L�Sֽ >�Z��<Z�(2"Ϟ�K��+�no'cm��K3b�5�{<;�Mnllf<<��ebK�vƅ�w�u �΁�b�><�=���`4�(��j��(�F14��(sF-����|��(8ҝ5a/�"�a�9ed���:�5�x4j��H�1�C�i'�)2=�߼����`��wT�[;<�i�)��,��wN{j�5�&k�`���my��I���?��tH�ix=j/�W�����
R�[�׉uC�E.���ǔp.V�{�$���<~�X~򓟰Y������y�r�SH�,ۂ58���B���=i�+�)!`���e�cu���c�k��`BA�y:��_dw�8�~�Fvn�0��Z�-0�yzO�&�����u��F
���(�s\����Z�N��jr*O�ض����=(P��6�D{��3:)���w�G��c;�I8�o޼���~.��3����ӧ�'g���
��7d�H�� ��q˓�Q]�Oq��큰��(a�gM~]u�D��at��(��[�}:Ok��w9.���K)��Fs4$��
F.ACչ�fc����!1�������Z��y,��8��caa�.L��F�nl7>Ėe��v8���eE-���TQJ#�<��|��B��;�YQ��O� ����k�g � q�f���[�Ô#T��ת�q�,�QfN&U�B�Yd�d� �ϓ�L��[y�n7ɐ-RY��F�[�U�+�I }X�XQ=2�&;^[���>B����Mzm.{�rtp�l���z�`�\��P�zU�lX^�n���-�y����65�%H�����O���j��\oΗ�B�ǡ���s��4�ۅsM�� ᢣ!���Z�c��;4�,��E@	�'�ן�ά��t>e�t��4[��؁���"d,����3���&�ll*����D3� s�O��V�Vwk�c	E�@��|Q�R�kk!���]��!j�
�u�A�j�Mf��A'�l��'U�ハ>��:6�ޚ#E���z��,9W���^�2���	Z�!C�*l�9!���#{}��6��s �aH�X��8缋�����#���bv7�7EFw���pB�P
�JDE[[��&��`�рF�ba���ZR��,��"��ű�0�W�)�;,P��Tf����9�Q�$牴�ET�9z���ɠ�N�$Ԧv�Q^p��r�g�>勽i�2�pK�Vx��ȩ�z��&��+��4�(�D?^����!u8Z��������Z�70ч�������
u_���9N�E�E@0/�*#��s��3���լ9���j@z���g/���yK�:�C3,�d��W�ҰG$eH���j����¹b��5��q����Yt�E�����N\����s���y�%g��|Bc��@���:��!����Yw!ڨI���Z�(`a��'DI)<X�Y
ߕpr߼~��HCv�)�D�.y�����X�)~0����}���Fc��؍���&92h�
����ײ�N,���t���g�YXѡ:>83�F��y�J������Yr>�5� �ʝ;w��ƽ�8#pY�1Q���L!G(<F��?���d��G
�ƶ (�̴� ��#���s~���;�G� 'C����+��'Ϟ?����s�X��`4�2ُ�
�Dd��4B_��Ԭ� ��OAM�bd_P	xꋐ;8�f`�р����7���ڭ�W�=�:�$�i�k4X�y..f������9�,���E�#:@!�a�7(oQ9@�����%�N��g�-���K��/�	�s�=����|�K��d�g��HV/D&r��a0n
�2Y��uE$�'1��%j~�����7���;V�X����03�.1k����KM���Zi�~�M�N��o~3;3��x��M��A��}ߝ�,���/�|=�d=g�+� <0|�Qˊr�+�I��:���'�kK�~�����r�I�*X�� *��Ov�O���}��C�Y����̉�S�vlz�q�DO�F�g3h���O�o�9�q��?k���꼇g�JV�b+e_�F�Ѱ�GT�*�w����n$�7��?ܙ�9����֣��+����K�/�#�;f��a���Q��x��d0S��+S��[�P`��1��u�ac@�`4�#��ӫGc��ݧXVD��%�dPZ��Co��%��>i�^W�$�p�s�\�l��Ko^|l��q��MgʚIdG\P���
>�~O��ߺ���O�i)󴼐�8��^Q������/��%����:!%ӑ�]�I(�Ⱦ����)<�^N��-���;3����;<ZT8`�v�=;���w��H�s�1�bfzʈ¦1v�<��-��ba���51#t���Ѱ0-@D�	����Uc\�0��Q��T
��� �8)���x���@è�kF�v�j��B|�V�� �T3��L\9V��3X�1��=�;��UYd�����s,ؗd�&
lxP_L:ְ��eaZ�g�B��X��Ѹ�g����XKP�^7K}����Ȯ� �c:T0s�aЉ(�U�PN�f�./���N%�fm�<��l�g�K��8�#���^%`�:?�ev`7�.9L(4W�#8_�X<�LN���OJ���
��Ŧ����hxϬX�3v�`�o�:L|s$�ݴg4���؄q*%���c<&��J	���s�<�b�L�r�C?��f//f�g-�Ex�z,83�*m&����vA�={.o��4�4��sC'��120���I(��' ������(�{���7�lp ���+�ej�K1���i���1!P�C,�n:tȔA�ˏkB4�"�/�Í #��Ұ���BP'�4��[��b���׺2-<�\�$.ƃ�̌�Պ�!Ϣ�sȨ���[��n�l$����N�㵷�/;�n�Nrn���陜�8����*kAP����� ����`��O�}Y ����|h��E��b�S���P�=���"�����9�]�
�.�P�D��qQG��5�F+ZoL?u��C�mqG8�#������q�c��+�����3V���J��Z�i�Er� ���]�ɦ�z}�"[�HYf����
ˣ�IA�]߹>���-�U=нy�o�8O�(V�!d����ha��a�?V��i�k;H�XWc�F�Gڀ�u%ъ�Cg��H<�7�PhPz����_ц�؛�<J�.�+�ѐA5�@� .�-{���PO)lT��qqF�Ǻ>���#���p9kg�˫���
RG��������N~�WsP��WJq.�a��]�^v�tߪ��k޳,��4�_��JT���U� W*��Պ6{D�Fk/B>�	P�P�f�x]�/��WvR�@VC}�UA�*@�dO���-c�E�������{3�����1vy]T�~�l�9�x��c�9��f
�}_�[,���"�v���(�3^��-�O>���?��W/�ݦ+�*@��K�N�%\mh_���[�х\�.]X��o%��${Y�����Mc���WR�q駓����|�:��9_LiL�_w2� ,�E��#-��QD`a̠�b�O
�P����Ͱ�q:�D� �r�A�7���[I�JI����p>J�+y�ؼKt�4�y����L���_��`i��ٌ��0V9�s1e�� �@	reZ�u.)��9��-����ڃHB��������tu]+�/��'_iX����j5ђ�u���5Jl�WD�r]*Ay��޳�����DT>6"�a�\u(��(V�a-�!���:�*�\�9�F�}f;��	6��ـ��� ZF:3>�)?�^:;c��F#��\aH���_���1�I<��A�+&��N���iV����t�fٕ�p���y�\��Zw��0��]�#��8��:<<�>���B�Q��	@��	3
0�jW��s�>9�2;�.�S�e��JLx��q�O��?����T���������	~����-|#K�,Cc
��a���Q�9�#s��L�8�A�I�||��Ĳ4��\*�~s��m.��`�#E~�(dՂ�Gb���T�(��/�Vd6Giߴ�����5f?:kS���{zF����*��ݽ���;B x��4��Df��66�n�9��p���)0 ���,9��H����BS	�T6���e�;�AT3����U���WK����l��~���VS��B� %�,�ʴb���)mP}���%RP��Z#萣�}9Oze!`���M�/�x��t�r���z�7*�d�g�c�eW�|{�z\7g;+�C/� �TQ�p_TsYi����FȞ�]��b��u4�d�Ϥui����q����>@Z�;n��8�����4����A��f��ҩ;憙C�@N�C�fʇ-2�g�w�ޅ�j�i/�f1�����Q���-3������WcY��.;�ݥ�QoR\dg+��=|�z��S��ڜ��T������A��C��z��A˯f|��E7fxk6�U��C��h� Cn����T�ϣ=5�l�e�μf6op&)�	�mJ&)p{�\o��b5DΪ�����)a}G�� dd�֛�5̙��qgĆ����C!�Y� �U��3�У�+�xG�`{!V6?��G�>�b��[�]uyS��YT����<2� �z��ת6c�M^��Cj���u�W�CDr��^P��o�,x����j�)VG��*ӑ��K'&:)띭7g�'i^��SFFQ�y��mBؿ ���x~�����5Ro����9ٸܔ��3~�^RMNX�f,L&�Z0d�-��܉�7Wڞ](��H9s��Q�v�χ�s�^�Y�	�y��g|�(����[W��]eSJA�T�����/�*�C��L�
��PfQ�K'�ndEW��B�"��UD�oW����g/��*Vi}`��T�Ā7Od�<�Lb�������E�3�`-m��:޳���,�+��>n�R�unc��iT(���u6��lЃ����.�(c����y���iD���j��v��s�ZSRR�̽i��-��iOv�
��0�5b��aY�o��N����я~L���]�Hs�9=e�t�ud�(�Wt͠���Q�$0Z�΀�_~ �������?���m:�`Ø ������`��53`/C!�ӧ�o;iC���9�/:?��qhJq�e_,��Z(��N�u��:p#O��d���
y2�"h6���b[���*�>G�m�fpp|���kc@�=���������!�pA=�`��~��P��k0q�^&�
ml��'�cA-2h�1פ�#U�Q�R�}X�Ų�<yz/[��3���(=G%�)�?���<=��E���%'�^�rv��c�DI�<ƻiL�{p�N/V��A���y2 �G�d��Aֻ�K�?ꌄ�����	�ޣ�`X48PQá�u!ձ�e�H!�Q��j]_��D>L@�*�Y�Y���;�
6� ��B p�l1�Q����{���*�uB����q�����
l�z۳�zޚk�Y�:�3��L ��q$����|�Y�R� nX-[߾3����;f�-���z�vP}��"�BT�$ ~<��$׀d����kԿ��N�����6��k*=�R���`���V�k|��3xj��ߜ��9���LP�j�i�,��ʂƹ^�J	Hؔ3~���f���U�:��p$Ϲ�ipHZk����*��hEz���Cu6��T�A���{G3�9b���'���,0��Q$c���'�}���es��BhĨ��M_�@�axP���N@=@�e�������܀qj_}a������E�W�_�%���7E鶎�%ŇL����#�� �I#d9n����	`�\`���n���G���Ɂ3BHpr�6=�b�M���%!%=�C��Y��`�ץt������Ͻj�N�c��ٌ
�`�1�"b^q.��^��M���2l"C lj�c�nj�ėjȝ��P� $��k���m�������Z�qX6ق�����޿��xp8[�n�ԋ.��YSh��\��u�Q��_�A"%�嫵v�9:�ћ�)GYp"L|~a�r!)0�A�4��Y��MM�sal/�-m����ˮkᙌbđ��q���mmd'��+��Y#D��y�<�
��H&�y�7����X^�~%/_�LN�|*���/���G-E8N�?o��j��P,R�.�WH�;(G
��Q��H��[�X[�"��յ����@ ��Y1&3�D5̮a�]\�:x[�J��h�����a�F�)�4��8�
�2t����-*�h���ZcX��qE��&S�2>��q����i[��k����_� %� $2k�>P�L���M�٪H�K�4`tz�ͣ[*N:@�O�A���}���%Q���G�W٦�5�T�����}�Cu��d�R�kS�\�ކL1�@Y�w|'��Q��X�K�gY�-�����L�e��?��tխֆ��C3�v-u4���re ���[?K�c(VƠ��}7�l������/u�YŘ����,)���?��\G�j��3#>�㠰)���ve~�|�JѰ.��k�kL]G��OC5�ٟJ]�1�b����u�q˦�J��� �D�����T�kFk���:R_��Tǲ�s�1�?a^^n�Ԑ���X����z~��&��E��>㊩��]9��V?�5 l2�\�<�o`���YG�4ϔx�d��Ǫ�����ߊ�Tj%B%�"����w$Q�{�:������Nh����0(��A[�줦`(^�]�ęxT�r��!��,8cS�36#���T��Ä���g?���'?���������Xdl�������/�X��&\�>�g�y9~�n���������ĕ�$��3��}��<�.:d��躩�_����;;�d�A�@(���{��<����,LF4�;�RG��gcomoS� �
��,�Wx�z�v��c�l�]G���%㾗f��#�����r�y2�z_�5K��.�Z�����B�DʚpëT�\����5p���XaCљڃ�U�9�+�E�a��V���rq���N�iT�x�:�@f0Fw���C03[��+��Ya����.�n*����~7���A~��6�~Z���iD؍X���/m��"PrT���V���!��b6��q7�#� �F*��7 C�Z�p�'r#n�������o��Z>��������.G�$vh����La��Z0Ppz|�Z!/�E��٘���s����o��qrD>z�?{���Lۈ����CeӲ}ύ�GR1.��i~��aՖ��{�z��6XR�13:u>�1W�h�����&K<�o�(Z��ۢ�hJ�붔E�j��?Z��y��:�[���s�8�Iфy��Ǟ Q�.+CdLf,ލ�3��I��3�z�U�"��ec�G ��+=U���{Sa��{��Ӗ3�~�Μ�h�|8���ƛ�U�5�.�����/�(<FcW�l�v
�h��� 7W�M&O���l����眛��j��{�'�+�Pl�&�d�g(�A�F��0�'��l�I5�nhHw��im@dk�=�B�D��|]�d���[,g�q�nCi��h���߶�8���hڠWL9>'<���V3�]�y���ʊ�rz�@�_��^������ߝ�h��U�-���*���ۼ���tL7�=X��#T����\�����q�t�cW���Y��ۃ(�a����lE{w(�bK�A�{� ��U�9]��ɴƖ���Jσ����~�6"�ؘLf" 6�a����7�F ���Ѹ]��p_�0K�F%jW�����t��_�6`Y[�� ���Z
���O?��W-*�Ä�./��:�,�4�����z�٥���Rusz�j3gA�l��}=���i�!zde����9*��a1b�����6K�ƍ-9=?b! 
[�8T�h��+P����x��b�u�������H��A8&�׳�3��i������l)��tg[��ܔ�t'1oj_t�z��&���p����UH��Y��!��Uk7>gaiTs��Vz�JYz���^��y����Y�縤�{j��8���x�(zN2�V�����:�2�K��R�Q9�ث=�h��~�Ӈ��
Y�4էB>#�&\�%b�05~\q���R�>�)�����O=8Uƫ2
J��EID#{�B��{#h� �6��){c#	��)�:�z��
'��/���Ϟ�b�G��wϞ�4)rPZBp#h��;�޽�^���T�Q��I��ue�tV�d�<w{s�� �%hwFG�����09:�![XƐ��nl�3���`,%"��o�W����r��(4�Q3i�l��c".�?�ñU����x�	gc�}(bS�@���R~*)7��(�/4�t��!|��=w�9���;9W���JH2��|A�,����{�@��=S�Y��6�]B��_���������}�c�Sb�8§���r#�
���BuA'u!ڍ�Q�cdF�ك�mr�$z����Q�0Mɐ����Bq@�>X�ޔ�wΚ.�A����E���� �;v���͓_iUlE���rv����؝9���[�Z�	?<��NKَu�f/��F3W�A�k��r��|�36׀�Q׶�A3�'��]_�)�oc���WD�1��|�cc�>�"=x\޿��}5�A公C����Q&;�3�V����m����@�T�Ѿ��d=�V���;��Y?V0��j������'��-���!O>y\f>@�{yiy�K'�
�m�t<^&����[��-�u���d{�Ze�e��̿�E����-Y�+Z��f��&	B�t]c}w����ƣ�C�l,�5��j�Q:2��,�h��
��6h@d'����?��b"�b�Z�
8��a��< ����5�+�Z�-/�z0��KEI�W�kQ*[��T�4���
Ma���9���+�>o��cFjum5*7�G|S^�����k�'�onn��*ї �`W��@����;����"�Fn��NYV�,L���
�UHq��87�O�]�x,;��{�Ǧ����<�aI�B�Z��0��M��r>B/ّ?`���U�o��+|���?s��y�ǩ�S����&+78;�dA�q%�1���+v/�=��[s�'D��o�_�W�ʓQ��2�{�Z����u(C�7&3�����k#�/#˾v��gQ���!�7\hTu�ȥ�ߐmMǂ=M���h4jm<&�ُo��V���߹�>��SYK�?�q/P��h[(�Cd3^�z%Gڭ��AUŭxf�����ք�Я��);8>d!5�5�7�&����!��L���ַ�=���hf��R#H�p�]6�����"7��փ
9�*���v|w�B�F���QTw&��,��UF�3Q��֖fz<�{�Z֣;
�Z wV���8b�O�Bd޴%R��l �{(���Q��6�����dm��l�ƣ�۬�b��櫖%E��gY�Dz��_�{m��O�Ő�'O�uK^*���Yv�Q���������o�۵(���j.B�a)k.gh]��hY۰�Muif2�=2���!��~0��� ����Fr�F���2~��	�,⊓C�VEi4!g�4b&}\�^�xi܃�g�wRn۔��C�{{�n\>G�~͔������u�}�^�j�u��Pڝ��x�k2[���X$��f�|����z5m�z���,�ܺ#=�H~��_ʏ�c�wn�A���C�
6t���������k�A&��3t���������!s�^��_���q7�[���=�z� ��?�  �ĝgg�
��<Z{k#T��d��5�<�Қ\���b&g'���r$X� �h�����/�.'V�芶S.v+�QB���cِ_�lԔ��B����`�ݢH�e��
'�R�WTJ�ܕ�6��D���G�����w��e69����(9c;x��ݽ˔������`�t/�k�F,`��C=��̇Z�����SQ!�
��W������J&H�*ʵ���N� >�j��Ʃ��E�-�*�nq2������w���H�H��|w�g~��	ˊ�m�ʹ�E�2+E�+Ю=��2�K�[�J�M�����ݫw �P�S<����E���5��U�t]/`�]J1Zc��}��<'n�[��'����zr�#�Me�-2k���~�{��C��XD(�A`$s���c: ����嫴oי���^`�"m�B��%C��u9�s&��ޱ�$pd{{�3���q���?��?q?�y�V�?�kF17�� ܸ���76�)�'x���{�����H1�ˣ)��0���U�3r��2�*I=�Q�9?�<V�3sas�KϞ���9��ru���	znH6.�W��^3]P�Հ/�/V��4��N�_�w�N̸��GR�m�������T��K�G�|T��un4���4�9됺�h�>(���zu�[��C^[U�;oK���>�~�z�ce�H�"�U?_'�j�Zg�l�)XS��xg��uNb7������R�ЪW�xu$g���H`}� f�l�%����5[S
�6�z�L/̀���~��̇>�#���и�_
�yN��R]Z���<�q�?~�tT=V���L�d����+���@��Fת�o��T�rk��t=�����f�h����~�DI,i�wl6>{�#;7o�'�|¬�h���~˞F���Mt�_����$#M:� 8=��ÃSj��n�V���D���*DO���n������^�x���e���8fɢ��^J�g���R�+o2�̷P��k���=���Y[�A2�a�!��(v��xmsm2;b�$.bn��h�9, xTRa�B�����WZ>����[�dW�Zg�O��=Ţ��p��B�hfm�f(כ/ jѰ�p �x����z������DFi�7��֪�mr�z�ŉt�����-��hc��ӆ��6�Q�OQ<,ZdG�	G�,;�c���.|�	;<�v@��䵃�B�v	�|T��*��c�����q�!���Ϥ.�`��1����kK��ʒ�/���(��խ,?��短�}�8*��ԩ[T.|��U!��_��J��� �?= 7����g�Z�
��Ov�}.}�V�WR��[o�����"�p�W����[9/�s���M��t�y�N�� �|j�]�%jy@�ô��s:D0q`o�����[���k�DS�ٜLK�g�F��g�����4(�����<.�@��ܽ-<��P+�8�tkh}{�r�c6]�&��LR����SJ�1;qy�<�ͬ��"3{δ;Ėi�,��Bwʲ���z����ޫ�����a$
�� ���,:�A}���]^�,H9Sz��	Q�����øl��u�^������s��b�����s�iv/���H:�����л13c�zІ�d0��t/���7e��-��m�zfѳWA�:���L�R���q�;�������]U_�q�N�"�@����(� H���[c$;[�m�ͯ��A�cҿC��n[���T(�R��\���6x՝�ϸ�#�����"*<��a�AS=�~�m�)0�jc�h���N��k��5�H����O�,O��ޢ�I�L��$���c���|�jc�傒�����O[����+��x�l�Q���t�/
p�q7������r��m�yk���Y ���؟ͤ�s��z�ލ�On�q�ِ����`C
�*Jۘ3�kA�_vK3,����,rX�:`(��!p<�R�%:�,��͡�^���������V��$�����̸rtp.��ް�K��x���(V���@�4�t�26�\ha��$����e��^̡�p� �a���]�{�~�V�o\W�g�xY��V��U����@��<-�s�hӢB�gx��p��X���|�6���A��8�G'Cku��S��ݪ=�60i�� � ���s�3������X��ρ9!�ب89KQ�UY�����Q��p��n䨹�����ޮ�׼�#�9�-�km�X	��WmJ���{3c�>H��b�b���������{�� s�:+�ҭ��ի�W�p����j���س��|�ΆV3w�o�#X�[�ƴ��h��he����Ύ�] ��$�������:i?�I�ؐ��<�퇫���ֶ�y���ȋ�� �}s�&��w�~� �?�P>��s!~��O���gr���iϿ~�*Ɇ����1�?��R��CQ����Ö�;hȇ��`�Y���O_�z�
J=�Z;�(o��%eΧ�z),}�b�ay#U��EV}O��sz-�]�13�Do�ȏD�zt�o�������{f���}�����e�y�`ЌN�ѣ���3���w�=�ׯsDʇ�H|f�����?�y�7��4�4׾3M7��y��2���~�-�������ÃD�^����u�r�[N���Yʩ�
�j=.���#k���i�=f@��X<ڗ�EGJ(a�B,�;���Zi�A�Ȩmxl�jPk�ِzס�e�-)�<(�}�^ӹ��5��e}/:~��J>v�/.���`j�ڇ�����N�,�c���l�[:L�:����������}� �@���s@Bu��	_�(ܢ���w�E颃�o��c��d�=���HӢ�@8/�r?L�Y���D�B�ɠ�I���)a�hf�6Y���>e��ӓ�<k.X�W��(�Xq�zP��}��m=$|�a����D�G���N��m��)P�����5r���g˹�¬K7"S���\��ч7���g����wHԅ�0j�����fi ����GEBb٭���G"��[��+/U���z��_��/���փ�;Nu]˛:�V��K���;��"�767e��N�\�m+��sq�I �&
1ah�(\�1X�d�9�A�]�*0xFC�5W�2�K).�6f�`u:�z��(�+_p|T�G�lVɭ�>�i�_s�k��Ã-u���Wg~e�]�x����{=@Vu4�d?�C�@_���L8����u!��9'����5�}Y����gB9}_�,]ǵ�j���7�����C�`��u�텢ys�u��5{�p"-����-���X6�>���ez����e��Ӈ���ܧ��>	�����G��>c������Ǐ~���s����(��}$_��Q"�G`���PЎ���I��鸫C��@����K:�t����������+�!�����ѣ\�aʧ�ڝ��U�,�
�jhKS�[o��'?Z�A�b�#�����$_�R�B���C`ݹ{D�%V ��Bg�����`ٚg���OD��B͍)�ͦ��^S��R?�R����ZÍm2*�
�}z�����꺂���g`��N{=h�p�
d}�XnÕ�	�뭵f�������K����[�X�~;T�/��|�˟��.&jG�Gu4���a�hLkr�bҡ2gCk8��H�B���v��ش���O���c;�πٓ��V �,qDY�X���.8�@�N��2,�W�ñ0A5��5F�e��s'����5NC>~��������p�|>F���ן�^��޻�������g>�����L��p����[���C��M!����?���l%����ɓ��,�#��yr66��˗������m�`�`+<"�:2�h� D
����]9N����6�$7�y��x�P|�c�#Y��Y4��Ah�s�����b99F����[�P�ה�A�r���F'�q��k��jy�z!g�''�}ODW�c��9\��|�����pñ_,*G�-���p|l���@'<�*�Λ��T�u�V��k6����P���R�I����.��s�ɂ!o㿥or6Doh�4[�bBQ��S�Γ����t1 �n�ml��
9�OÀ�؇ë�\I����&C�k'&]��`�a؀E�X�87�,����^$n���	�O5�=��Z�9�����!#E1��s%b�[�=]wEn��'���z�}%�g=Ց�e���9���i��|��ح������*���C�y�*{�R������˩a/��z����u�m���0���=�K/��v	�]�)����C1\zc���r��G&��ळ���2�8a/�_�o}~y!+�4	�	�ٺu�l�}�c�^{��#r��'[�����8'�ڍ��� nݺ�ݺ�B����Mt{���E^VW7HG����9�L��Nv]�r-�{�w�E|�֎^��G��bjc��f}��O��`!+(O��E�N��5ў�X�[dӯ�	�5������h	�1���"��z�k:�H���=�qI�gz�e˕De�ܾ.��k�`v�b�������Sr���v��4�a�'��x샢}KЁ��Nؘ1g9�������v�ד�1��eY���>�-F�g�2�"�s��5�k��9��yXz^. X���ND�e0HvȰI=��h�DVډ��Hzxm(�$vO��l0��"}����INIXD��%sh��� 5����k� J��^o����m�v~�j|)\�3�Dat��Ө���Ֆ�W^QB����o�P�ѷ�\����;�T��ҍ^���f��y~�>o��?^��6WaI��f���-gwZ�fuZB��˚�����G%'�ٹ)?����_������{999���S�߿����_�(,6]��B�53��p��З�2���XO�9c�2�`A�㱺��l��]&�4�3�TB�7��od1��,��Q���l;G��g΂5t�d�� R=3e���]��s]�:<�qq:[�HO0��ޟ��]���Sfw�S���1��9��Og��;��GZɽ�,�#��pY��y���䌢êz�Χ͋*V7��/��{�R�[ND�)���E���cM�G��R��tvL�9^_MNƊl%/y�����U�՗��xq�[���Dǭ����������.�D����<k�ADK�XV��7:܊Hp��?5�oyz��B�����9����P�w�Sn���첦�iY������qC5�����Qjɧ�6��\�W�d}�+O�1��p�J�d��Y@g!��z�b����&{��Ro�WV��W<Y���ǥwۮL깫�`�`��ǡ��J�hA3�⭣ev��^�����Z6�[YY�^IL����*�K�8`oۖ�=gSy��'��I��e*��x�B6�Sq��Rb��}���h�_ V�J��
�BgSf�
�Bp���� 2�M�5+2I�`�(�f�bo�=V��+S��]/��d�����	�$Ǖ&�<"��Ϯ>��M Ar5���I�I�\f�ٚɴ3�3\^ 	h�Q]wU��z�;�=��1CSٙ�������{k˔xtZ�u�ܤ��P*0)U��J�(q�"�]B�!���N��%tt9Ѿ�����ٚ���$�yJe�ԍD��Ŕ�r ]�%x�i�ULQ�й�b~ޱ��|���S�6B�yEJ��\�Q`��ȉ���O��N���a��>J�FH���
Mh�s�0>�V�zeȇU4J��[�V��Y�P�[M�F����(xg�C{��uNG��ת VWt��(MQ�U�9�y�G��7����3���]����F�.���aŲy�z�O_^��^��|F�e�;���)�y�����|����HH��9؟Uku��~�1#�r�*S�t��"Ѭ�M����h&]�!�_���G1�ֳ��⩲���&J��u�{�Y����؇��ϋc�k�$�c��):�I��.����ҽ�!���V�j��>y|B�~�!-�g�����}��o���\"ԨAz,Rz��'ʿ���ttxH��t֖�BlO��P'�@��K�B���y}I�E�
������O��ü'HB�r=�n�"��3D+r�N��
BM�w^��{N;pۖ�7E�-�A��}d��8yd� ;��C�Mz��`0�	�	�� �����l��,UH���&��	])� Fq�+D���m����Iy�KU��#D��ݙ��~Q�~�<���5�!`3�<r�N�1�b���(r����BNhBc�iG"4*�h^�.���n�#���U�U��]-zB�Ұ%:ntE����Aa��5NaB,_�T�K�
oWg����u�S��~��[�S)%�EjXH��dC�J���u�x���ǿ������t��ƽ1U�=_�������d[|�"������e��Rq#���d�����wy����}�t<Gݽ�AyFT!�a �M���D7ZO����+����J��.VK��oHV�N���J��)陂f�{|l%��+z���ۀ�a��xL/_�(t��r7����x��醾dCeK"��n� ��
"�߈�nm�vs)X�B�÷�;�g����k�?=� +]��g�D�^+~#����� �*�Zi��ލB9;It!�9SUE9����n2��+����Q=`|�[�}H's|��ƚ�m���=���/��N�|)���#�h��T,LLå6����j���%"怣i�:�Iz29��͠��Y=��%��X��W�
O��Q�O5�)���4�ג�l�uCQҸ�P�����XK�>�1?]oH)���D�ܓHAZ�X�Y�_Ѡnhg�{���>9����ı��N�x�ҧ{-m�hn�7�=���ç��"����M�R��G��7�ݳ�X��P�$�%��^����ʩ	v!�{�5-�����/�eDu�>G�b������Փ\nv�Z�M>&G����0�)���M�z$C�����fk��f�tW:ܲ��~͒梉c��Wo�LX�t���m�P����j��������ӢY��?�L��@d�!��O?�gO����������m{[�:�LW�/�!76h����k���L0���R��FGOs��L\��8��n)%,M�Ӕ�`6Y�&��
�lO^}߭�OA(�7P����Cj����A�x'޵������r��m��@_��
(/��DX7�����~��!9\Z,�a���Ujl�<L�>.��������U��O|�H��[���j�~��TtP`)�z�J�J���Da��Hl1qa��Lf�V������>�ݽ=f����b5��M�6�;�x�l�����_��� ���]���a��YG��d�V��SXBM)�2yyaQL���{� v��_e���5�%)��Ν�/N�e�y�}�Qz�Ibޔ�K�5�l]x����Ck��:�L�z�*;ƙΕ��)��^d�����������ݍ��-����z��pE,��$����p*�CW#������Vb5O�g2��/��s��a�[�>�h7έ�FEKKQ*|��C���FZp�:�unĺ��\U&��M�D���D��7KA�ZX?�"G>�E�XF
�0�+�#R��Fyp78��hS@�DV`��g/�GT�^+�N��F���1�
a���߻�)�+�t�^ƕ5N�~P�e�BH��-��>�+Cg�����5�ȇ++I��:�Z���P�M�� �<)+�k��(��D��;�-ee:OIYg֙����ZJ�2cBo_�s�%�,�*�\��k1�h04��VR��Qk:j*P=�pI-	���uN!�S+8s4�����١�MR��b����n��9L���C/���q-��FJQ���^�%���بV���6�K��^�l|C�Q�6�:T�6������}�rwcz-|w��s����ŀ�s2�����6��ܟ.�qA@R�ug�>b��yꚧ�)&^�^1z�Z��m>}��Af��E��딱a:�OM�CO�B�{���D��>���"�w�W�J�����rq���u}D��+������8[5�:�����a�m�[�N7�ͭ>�W_��6Y.`M���f=L����f��oǇ���܁sAM�F+8�Yvl�w7^)'m���u_)��1\y��<�}�*U��L�ge5U�N�N�.�S����r�=��7��m|�B#oq��0�A�MW��҄_�1��e���2� E�3�Τ�}�G��c�xi��E�E�����ݬfO�.̻���G��͒;�T�Q�Hgn>�eA��3��	.d��nb�o�;Cԁb_i��t2�t*1���8<<��GO�s(1���"lA���w�]�ů..� �Q����[��nn�#����4��ǋ���G�h_ {w���ts՘	�E��Ҭ�m*�+��	�q(>/#����纷���/���gݿ���5�N�f����F��22�Z�M���O56Tt����h��lp��U�ۋ�-��׶3O	�u��D0J㿌<���
��k]�s�u�*���7���)�j2��O��!���9���K`��A��B�V�Hk�a�<��5Wz�z�H�"�%��@d�=1&��(���h��2D�������*^#i<��l�:�VDR�x��{��Ҟ@��w����hV��6w7e��֡��D���q��f���<�\`��b_'�\�P�a,�sD����P2�%��idro{��Q�AK�`��︜e�J�Lc�gM��P��6+��΂̇��q�A˚$2=<���<��j�r�&#VK�+ӄ�)���}td�T����t�<�)������=�t�ɤ�h\]�i�H]Q�����V�H|�3�D�76�Sn��G�x+pM|ե�OU\��;i���Q6�+��i9��6&�Z�w/���D�)6T�!��T�f��yC��S�\��'mMw�>�h�`���Xf^H/�*V(�k80>�<�̨���M��m���Ğm���TPW������u����np�V�K*�W�A�}Ƣ�*�!]@�BȒ�zżN/��d��c���;b���=�O貸��Σ�C��G�@����+����Y���!S+�2�;���.�|��	�Qc���k�Ξ������ �<}�Xta�~�E����>���r�؃w-U��D��٥���	u�_�X&�i�����R�&��'�Ou�h��!zOM:��b��25��#�iz&O��"���|_w׬�,Q�y�&��!�rS��x�����tL{���5��{X�̵J�(�7��m%��r~�w]53P!ߊ�m�ed$vϖ&��S=�0)��#���1,4�$�9I'�<�6!+�D&��O��\q�3rא&�B���֞(��ȧ�r y��۷r]��a�C*wwcA�8<ܦ��M����@
��Ӊԇ?:�愇GGR�
e��'f�[�#h�AJ} �B'�>���74��.���];�>I�_�D�뽦�w� 3��DEB��{�Q{h4?UD���o����!�Jܿ�0fZltOa����S�Z�n�:W�扤L�������Pl����X��O���,�#�2������f �ӭD?�V{o����~M�ŷNsEظ���_3�5@�)�3�*�0Y�$C��{�)���ľ�ww���x3��� A�Z����~C�|1%{FIm�tjh�t���[h�hhccK��`������ǃBť8,�p��p8���x��m���'�RbƤ ��\�|Qů��֩�>Ɇ�;3D:�ė3+��q�e���� �	��z��#h��Y�z7qd1ߚ}�a9�bx��ˆ�jD��%�T[�Ȑ��n�}Ƣ�v����nc���O����LViG�nN���(E��↎��<��V꥖�Ƣo�C����^P�O�ה*�zo�*4�G.�d�kQ�ĸ��;�����U��(�����x��'}%�R(��]��>nc���A��|�npD5:5 jU;e~8e�aL�0�a�����[�R�T�O)�����	��.�G�u�{�@��5��t9c�~4_��g>�:�'l���Z,��(�"ڧ�b�Ʒs�x�8` A�̢�6y��Li��3�'�E�,��$�RE�z��V2F��#�%֚J*���]���R�N�XZӍ�V.����� �����{?�c=eoM).�v'̮L��?/��Fل��F�\����wRσ�y�<�F ���~/�76hƆΫ��$����g+~�h>��{��{pȴxF��-WsI��4�Jce�g�j��%/q J���^9�����&C5�#P���cWM�G��E&�;/�HA��=Q72�>�񜶶�%VR��x����l���+l��
�3���:D(P�ʶd:�ޔ�CG�������y:���`�{%��Nh����6�:D�[<qz���J�m�q�ڳ.VH�2��<j�zQ�R�q{w&�0#������i;l�39��F5�M4�d�5/Iz���]�숕�g��4R6Vo�ؑ��d����'��]�Ѽ�f�$%.CT�J:\"Ē�b.�>��q%�{�U1���6������HE���c]iWҽG)c|��h��4H���/����F�#3D�IFg��TQS���Ui�� ɥHH�TE��z��3��v?��x��P���~m4�Y��.��~8P^���1 ������B��,���EN{D�G� ��Vr����y���I��t����p�z<O�\�p��+V��rU��A��t̆"  4o��8��2��V�Ib�1��n�i+��-�V
�CC�d(��S����בR��׹�{����ׂ�E)��p�F�]QL�<t֦�_��O�
��?G��E��_WW�tyq-k0�q9���=5�d-VQ�޵y��w�^�D>��v�Z�)q�$�񄂞�"����n*��e����֝�u*��HӔb�)� +ڒ�Pi�eH�<����-�h_Q���D������J�]a7^�y�MÐG/�ƌ�Je�ƶ��w�(k+Gky�`TZʆ-�U�렉�|����$Q����k�+<�9�̂&^�qtM��N
��RĴ�u;�Mh��������[����h�����4�/�qoB�m�i�4��`����U��>0�
Q%�[�z������'>�Ӎ>�|uN��W<wy��b�7PB1�^-0�M�2�+�QQ���^���5��7#�U�I�tʹ�c��������V�p��V[�s)����Ƒ��{�C�o3D��f��lQ��6��u�-�u�c>�����tGS�^ׅ���p�Kmz<�rʪ]��ե8�">��[����Z�1�
˛f@s��7��ͦ��4�H��9"l[;R�w||BO��i>C�+��%T���1ybQҤ���j��Q{�������A��L�z"�#*�:���-dxLz�w��u��;H���c�=� K��Kd�=.؀�\E�c��&h��><�T,y�.�A��B\�F�X�~Ȧt�-4\�Y'h���'�C�!��!�ֈI������� ��it�\2��F�n��d��r�6��N�+w�ap'};���L����R��Z�?ɯA�w�6��qn��К�u�D~��T���-u?>��#&���ј�s�3�yt����#�	ȍO0lU\�L�ۚ���r���
ӎ�Q`:_�r��^*z�#�{�V��ֻΖ@2F|�q�.9��6J����ż�(ܷ���9�f��D��D�{))�Z]�Ny.~0C�]�d%�:.��=b9���e3��%�9�C�����1�c�(k�|�+��R"�m��>����b̥
��������>5V3@VtJ^8e�f�/G�M�;�����#�j�G�r.�^)��lE��J�������h�w!h$U"�p+��:Nx#k��t.(o�G�U!�5���H���aŢF���8�>��ho��� ܥWo�$M"��m)K�h3�|���7&�XK\L�f:3��5������?�.��rv�V
�̪��-D�7���uD=���*��RV�H��?II���G��jm8��L�,����r�%H"�*�*����|�^��;�=��a�b���Rs���xfox(.)�Gk����]�=w-�ǜ��$�o�df�T��c ��R�ŞA:#"��wD�H��ʕ�`��|l=D��d�xbӈ�k�������8Ds\tP����{�G����y�'�
ɼ�S&J��S�Iԣ^�ш����o� �Q?�i�^���DS
+Q$'Wgt't�;�''�t�H�x/3_X]�jh���ֶ)�\zˊv7Y��/�`,��늮�/x��$�`��q��|`�hz��Hҧa`���1$�.�K`� �i�p���U��� ������-x#`���'���?N��")Y�h
�^�&�����Zӝt=~*�x]n��{�ƭ������Ȳ1K�w��Pו�!�f�t���xk�
2�p��J�׭��uɆ����:Ŗ,T��N��H��A����.d]P3��v�n�c��㧬�!%�OV���k�eR�((Q�d�+��Ju����u�F!�!�[+���(ϯ���yD�*ư�p@����6f��,��}`���+q��� �t��G�Y�+��KC	���y�]�l��>C>��*�\�y�
B� ����6(�7��%!�
R�F|�0���-�h�Y�B `s��ӈ���_#���_	��z�0)��Oy���~3Q5f��&�z��&�H�t�D��{q~&Q��2�	<o���z�� �-�3����c���!��O?�рA��sab���|szMR��j�kn�'F���(�T��#%*3!��Ua��,���G��v�E|��<<�(�4tN���l���LR��m9�wI�|�d��&M���[��+L�	y�!�����LA�@�+���銡~,�b�r�,G5~e�P��R����:����M�JB��)����t�f�Z4r�M#>�Yni�F�|�p|ʶ&jU���,�nQ��7���JmT��������#�L�٨��롎�ϼm �l�L��[[{�.���[=�x,Q�+z���Z�\���5�y����㰏i��[0��V4�!x�d�?�~&J��xʿCN�1�o�c:��n�c�6��ʢ 2������dBr>X�q���P�y��4y��V��;޾8e��{����{������(T=O=�j�H_@�|2�I�K�ӟE<� ���2��R��=@��)�J��+�yԦs��Ш�.;���nOj)������hE�6��iۼ��k{�4�4�{J
�(�\);���UR�ʕD
�H�YI�U0,@/}K!l���h:���~
+����{ʽ���ϳЦ������z0��Q���Ah�)c�� cO���ے�b��L��h����oZ���k��<D�[MX��R���aoN;uCl��뒍�%-�K�c��/iP���O��on��┮Y�>:�cy��x�R����`�/V����2�`eh��(T���π`�!���-=�����>]^�J��Ύz�a=?���d�<��֭'�8&� �b<��W��F�h1��sJ7�,��4*E��[k:fkm��r�(���#��z:2��6��Ӡ6DJY��rw���^�r�44�N�7=����-����	�'�����n���b���I�{��+� ^��x"�4c#rowO2]}U�%K �� wu%iWS60Q`}uu#�V�oom�����h�J���Z�H�ri�L�%.�*��rݒI�R	�/�6�]ۚq-�@��:��t�J�U�nHzM��"�x�RxI�����e�}��������P�h�)>�4��H���J�4�c+pʂ�����`h�6�B���{s��3�Xl���/��!J�ݬԣ&�V./.i6�hBBC�����
$�>���
tFBl(�o�Bj@0O?���wLp��AZa��DAli�$-ْ{M[;}��s�>~r,���`+��_���}�_,�#�[+��8Pr��{����%|���gﶷ�K�l���
��C��ߖ5 �9�=�VaD���9uz��3GB�OcR	I��O���9+��a�����g�^z'��c������w���1�Wc�
��5L�_��`�u/}�޺qF�r�ϵ������w�lnR��J���kT�G���*_M����W�8dm�s���\��d �	���z��^�KL|��)S��,�����l�^��`Gq��{(Tu�&G��t&����ښL�F�3��;�)�|yƂi.�	C�0 ���,���ޞ�DqC�����4���_�����0�As�;���ekᥙ���b�:��8Z(H|?8�����ܱ����b�5���\�>�����V�/������`C��4�2������Qg����5OkB,&u�8��GR����}�y��~�;i�xs{c�go_k9�b�-�Z+�ʍ,�G:*�{����	YiL^�
y�f	���7�Tn�r�����h5mgn\p��2���Q�<�J��<~�tt��Hi�R�P���{�Dk��{C��H��d�h8�H���C�gD��5�U/l_����,4�������V�Jm��QO+�66Y)Ы5Y�k
CŌ���"�\
�n���I=31du�7|%zņG�l{�㼢juC=6H�7{������Z/h>`ë��L k�B�5�=7���5���&����Q�(67gCk�`�۬�VY�1��}�z�1�~�}�lqL��>}��t��X�G{�MTHVHE���tD�09 �@�%��j6��_p���p\6�6b�����%�~uF�gWt~q+P��S�L��+㿍F���lb�!��ƷG��x~0GR��?i��C�2�*k|]c�>!���j����#�8:�A�����3�HBf����+� !'��,������J�P	n���j��l 4Hx�|���������$��e{g�:��"���Η�҄Q~
#q�#�4��e��i�DI�t��@(���ip�,�OZM-�a#ue���
C��z	_�K
B�Fv[��#�@~�'?!E��Qv�r�jg��Պ|���=���	������0�=^�x׊��(���6Ҵ���>� '�R��ѡ�P���L4��+e��!C�?{vB}���������t�����U�^�0���,J��M�����?��Ϟ�wB
`b%�<(�c+���)?����䃯P����<�`!���5���|����ϥù6��L���3���R�6F#)d�g0��7����O���}}}I������b���5$w����}����=�εx���n� i]iV"M�+!Twzh���jȟ��;��C��������&H�r�C�F��(�S��8O_iM`g������ �ﺌ/�6{L�=���y���B�h.���*).��C�|����a�萮Ay<~��Oo��t����:����QS��RE'����\��2�(�K�<cU�5�`Z�{<·��Z�|m�4Q��D�Ӷ�U�T�킥�T�T�qFK���E�б|A��㟥�ƣ�]��ۖ0�l6������X
��66�%MR��U����B��vDL��lXI�><j�<�ZWZ<���-6:�|SV��$�t)d_�����	�7�{!Els�^�^��-]݌�~D�92'rvoQ��r��h�nd�C�ū��)�f�j?����,H!P>96��W��BT�ROg�5+M�J�"�$@�B�=���:�+�(�0�!�[(�Z-Jm��hQ��u]��"F�B��*�bmzs�ᄍo�a�m<���h�"`��^cʃ�b%O�D����=��z�M�I��#��������dk= H�P⍇#�����FJ���;DgK}#��0�h��rZXT�����(��(Ep̐�f{�Kg:s�OI���9@��D���-5��4i*�6h��q����cE���f����b�C�jw����)�:��潽},t;�B�٣� �*�@���ԉ�LΛ|��z�ч����� 5@�c��Բ&��Tꠠ�����Ɋ�Q�5#I]����n*����'����SP�36:���o鷿���7�����[(n��P@�hud��ve�'�OO�8eg�=�Ș�{#�\6�}��I�D��kt���/J� ����g��|�h�IH�D�_jK�T��'��RKdi�қ������8�uz������9�� ��@M�vY7gcD�����X2��>�z�Fsk	�D�4J���F�&C��r������B��!&}D�v�_j�(i^��?�9[�K9o4�DT7 z�*�l���[U�cj�/�!�����U���eX��ޞ�J���nN{��J$�Nk����=x�VZ	Ӫ��N*�q�P�/Tn�8�*.IG!�7�So�[%�����ɟ�`�f|}��ݿ�}��g�����/8o��31
�$���<�
�Ϟ�/���>��3:y����@�A�������)��/�ҟ��-����@`��{���s��>��>��������_������8���=����;a%����k %+�w��ӧs���䓏������� @�@��2�У�G���z{vI���n/����\��y��U�L��H�G���\1����8��nY��<-dHF���uKUr��
�R�R���U��$&�B��;S���4��|�R1�G��ڞvo^�Y\J�l)� ��AO��R@���)釪���U�l���h��W�-�0����j�e���!�Pq\�ЈR-jY��@�0��#�ꍵ�Q>�i���R���9���İ�^��"������+({�g��C��t=���B�| ڬ ����OK�S;; h�H�Bzs�E�c�V��%�v�F��<��*����U���1mon��c8 ��>��{Eo�V�a�=�_����"������|;�Ւ��$@H��WG:��I���}2>�&<������76>vqy!0��'����ت5C������Rau�{ɕ�P<��E%(�������z��VШ��)��f�T�}�����+UE��'J+��)Nӭ�LH��n�qfJ��n���=����ĻB �G?((�'"
L%��Q��5+lmFЭ���'j� �E�ZƤ{RҸj�<Y��4�l������*Y)�
ug�:Y���hEe�����m)\&dɟ|�'{�!�!���x@�	l|��KZ]���~k���V`E���{���7����쎕��t��������-����W[_��a�XJ=+��n��Sw�J�5Xl������~�/�D����ƑD��^��5k��1/_\�9��`��}D��^�:�W�����nX�^���pw_0@�{t�O���������6�O���O�	 u9�}EK���Q�sY���~�Sʵ�26'E���C�M�H'���4c�b>��R�o������q胔��~%�C����������>���E�~�:6��3�ᦖ��Һ���+�C ��F�:��'�J߲���{C3�V!*2�
�\Y
�8�@�����U��� QH��V����At'F��ޠ�E��fδ���|164����z�F�E��D%#�S���R��HSܠ�(�s�)�)mi�����-I��d�3���4�yC��l���Cm��=B�`�#C��QZx��
�������Rb�<D)�^Z�f�Q	8j a�t+�Ũ�.����b#��:~�G~�~��O��x��/ާ?���<	�hs��Le!�D�,��E��W_�W���>��3VvD��&�3m	��Pxtt@�|���=f*������7�h!:(2ÿ�w_�/�%���/��pO�Ge�b�Z����<"+�r�Ӵ�cE���B�y���������G���¹�*��8:����X"��}���_� ��VP߈0o�$�Z*����pve?X�u���Z�/��ꄵ�L�N3B]�����U"ǹ�"w�P��)OnF�}g�o������rṠ^1�9��ʒ�c�oXS�V�8ɗ��ϝR�H�.ѕ{�#f�c�<9"h�fk��d:����D��*�Y1D�a&�M��$��D=�̜�k۶Ի1�����aU���61���T�QB�F��=T�:�ꪕA�*SuC�����ڢ#=Iu@�fE�j>P+&���'���d!��;���i,PD�k�H�����0|e����@����/�^�z!�c0��>F}HUזfv'p�@�C�*�6幒�J�U����K���C�jt�0�����/~��-q��V����Qk4,V�hp%�(\�Up�(2Y�c��v8PF�[?�O�8�T��f޺����ь�F���H�"��O�	�{�6_����^$e'Ƌ;@� <ݻ;cH��$jP�� ��0ۯ�O�$�'�<hъ_�f�%��=��qNq�UVTzA�䅍�1Kɉ���d����ºV4�*��v �Tk�p��Jz�J�#�9�i�)�`)\W�C��2Z3|�ߨY�	�Ĭ&�T�#^�S=�����R��U���P���ڦ��y�^�X'w٫�V�î����=mmoI�A%�������B��|ߪ���.W3��.0e�����C����k=Ҍ�Û��i��ew����#VF�y�c}�ԯ��vc����F�6�ЗЏH�"j�����=}�������{�T7�(���s%]�	�"��	s��T�'Izma�d:�Q��P9���~S}�5��&����Ky��q�=������h?�c���E�t�uV���jgt�5�����	��e1�Y������/�(��@_��h��Ɔ�� d���Q=�E� c�Ӑ�������X
�D�+����*�hz'�$��a�@Su�y��w-S��W�y�ho<yFO�>�����^�|��z+ȩ0��nRx �d�Q}�E?��}:|t�QK߿��N�2�_��T����b���t���_琞>>���M���6��^9�˳g���ֻ��p�y}��� -8Gt���3>p!�o�����<gDx�����&���5s��Cs���-^�G�׬|�����T�� �h{�X�Np��z��{�V����oC��?��;<���4��m��(��yt�(�������������B/|� r�u�e���]�����l�$l�jƬ������'O��/����_�)���H<�/_���*�C8#�����hS�l�^���*DE�a����ۛ3z{v.( �$~��4�xDJ���'O��G�|D�NN�S3�_:�ժ��@/�R�B0��y�!��ŋm�\R8�D���Ͻ���"�ʩ�6)-�mL�kqpR�D�VM4a��ybVR��6.��U2��FI�df�h�)*�, �Po�t���zM=��jU��=ti>����yw�E��i�m9?�&txi��wr����nP��Ei�m�
ìr�rt�ƌ�!���	V�_Fe�`,g��?S�)����yq^X�mq�&�Z�\h{���%@��fv�Bn�%J1�ϹB!�Y�!�#m����"�[h��M��G�o���^�Bp�G���(�!���hC���T�KDCU�3@��9z"�Ag��E�˅�w��<w0ޱ�i��絡��k�Bʆ<�>7�%qG*�=��w����O7�������S��@�^_^ɚ�������S�����L5�t�k?r�5���c̉�:�	CCC� 4�S�&��A&OZG���Z6/6�����
���Ɨ+k�^�q�y]J'��CЊ�,�d7	$��OAXk�AK�S���Tb�I����!K��O��*����#-ԇс��%�JqL�68�*쭦�"�ġtpeԣ{�~���s.�b ?��_�i5��N�=<��)7�]��i��Q+�L�(�!�]�����-���Ƞ����%��G�D�%�d��׼{�fb��0>?�����TҦ�$�n����[OW��y��؂�����7tvvAGG�Y�8d#g��y9�����#q:H���%�q,�j��}��g��Ͽ�/��9���_�|L��3�[^�8��d)��!���*��Z��(�x�W
�ܑ׾ɜ�
��t�(�
}e*��zO��l�w"T�F�^���.�}�sѽc���88?P�u�їh���F2?��-�NR�;��l��� a���6z���;Z��&Ӂ�-8�"�I�L��{;4��ev��%�����YHW���e��|��lp^��+��&͉�|x����>~N���/�����_�?����?I:
흹k�d)���������/>�����ڐԿ�?���L�h65}��s������=���!�x�Q�^3f=vzwI/�ߧ���b��	����=AG䃐��h����N�ȐN p���F$D�b*SB��0�SO,�������/�X?��t}��fҸ���X�Xo�R��5�����b0�����P� ���DV<���"y8��g��/�����_�׿�\Bd/��~��od������
�󄍉'OO�������l\2�:��:������?�g�}"].��^��N�����D �\B�<G�|�'���|���nn�%O���H� "��ŕ 'ld�0���Ì�'�'?����9}��G|�'t���������9ݱ�����gH@V$�ff��S/�^�����TnOm�|�P�RV\Q~�����(K�T�T�D�Ȑ��d��:$o��ȸ���
œ���7��S�X'��a�Ʃҙn��6���'WX,��F\�x������ٸ����+W"���)&�èU!��q�����-��Ռ�`�V�m��sd�)�h�M���Œ"~4ͧ�.�e1^r�D�G1�3�1㠤C����cBG|KM��襷p�@�V�a�d��zՓ���ݤqci���D�v)5#��سu_�?�
�r\���چ��'55�Y{�)�`��mJ�#&��9�C�+���B��I)��w)�KE�x<�a��מhJ;��Ps���Bە*�U6n�7F,�1���|�G�~T�T1�(�>����P�WOˬ2���H�rI�`����R��Q�tKn����6��[W��͠k�q�Bm9��m�~��'��3Z�iJ�!���lܪ�{m�[�\7
��P��E��8Q�+.���8�n-~��&��b�h�8Y$�+�D����Z�>W��"V7�@20���C`�#Ln)N/���R�r��f����� �
(�z� @���"�ϻnC�3����;ԴŊ����s:={�J�.�z#I�\4����y06�%�ҾWh��Չ�p�x�o��LV�nY�yNO�����Ѽ�ӳ�c=��~��^�����S֡��.k��ZH���lL��J�_M�\�������(�(�;{�!_Л7�j3�"�IQt�p�D��9�k%BEJ�M�]#�B�d1�Ԅ6SA�����{?I�rz-p���RF�>""vś��������t��*�eNn��"*v�� ��wȊ}�������w���]��A�F�$�Ĩ�y�\6����B��pn�L8��������ɴ8A��L�uŐtݭҚ�Z2tVR cx{_f|!5�S���7�s�I&D�j�_�����'O����A�&8��R׌{V��JۇT�i�c���w�çL3+���L�g|<�����J��/�lp�z��	�<���~��/#]�����&=v(ɔ����Fx6�L�\����KD,:��TK����(*z~Y#�b�c��� 8��|�����������~�����+-"A;#W�����ÕAt�褙W?��p'�ѫק�ɧ�hO�'� ��՟(3���93�/Xi�Q�2�o�;�����߾X;0u0X�0<���s��W?�g����6=}zH/_қ�l�ң�C����`������=����_$4�n����{Ϥ���'��څ�tz������������g��}H�l��}�ϼ�ts����	���؀������ ����?�!uNW�>oI�PFCH�6�u�x���%�&&eF�,y�c��\�AG�'Z�A��������#Rn`��4�r�MH�r�o��u���eA�a>���2���δM��RI��۲!���0�4W�WR%(OF�7�m�'羥��t�5����y~��6z�K�-�yB�]���<�D](��2e-׬�wZi��(�pe˄GB���>
�7]?y*���*���U��kK
�dYwm�fX�"����k3��6����V���H��h5*�(�L��i��{-HV��)���%,wK�*W�"r�W��F�G	3�_�7�4����ׇG�4U ��/W� �
Q�h��Rc�U�IgC�y�B��!���-��8M{�������]��9��w�,<�Qa �'�{ȩ������-���5D�=J��C%}�������i���TSa��P���o�r���>jp�H�d��Z� ��͛_�� {��V}�	u��V��ߙ�����0�Z��Ri�S;in�6�u�N� �)�Gq삕��<6@V���ik��F`p��v�X��'cB}E�^дZ�фZ*�8�㓄��X�|��@�4�������0�!�0���3�)�d5^w�t&D+=6���$����G����������1�ٟ��3�����跿�+~oy<��\-0�57�4:ٗB��>"00������)�����d�������G����G��w#�:��,�Q���/��
F�t�Fj�����SG�T 9f���|a8�����i���=͠0�qݡ��m){�!�s����V���wr>�g*��G����4�/�N iG�{A�:�#(�KA6\6�(̷�SV�o�z=4����+�����&�-6��W�קM62�w���C@���Ό"�P�$Nu�H�����˷w��(xD�?a��..�F�.�!��p�&ӱ��Q�PD1�s���^a��ɓ#>~&�t�`��� ��j5���@�9밻�<ac	���Z���h �|��{��5�yyL�|�亢�C��lH�9 ��+���af���8�i���k�J�E5�{@hZZWZ�[�؀�j*�����zX����rĢ�����@��w��a�ۦ�����-���c8�#A�@=����X���Db<cA�X�I�iRU����}k͉b}�9,�G�M��( ���/����������Z�1���!gg������<��6Q�G�L(H=�����LT{b̀������/������K��	<=���w�}O�g�������?�g?����'��o��ڤ�����tw�d�q�1q͙�x�MO�l|��W/o���ea	�����b�]�V::&�^w���z��.a�r�j�.�@*\������v;���t��X|�ft�|7J�动�w�Bѥ�:Mq�ŗe��s�0(����#�F��B#oȌS>K�ZjE
�ct���{���P�8����=�_/)�*���K������U>�D����;���P�Px}��:O����%���L���|�y�|ӵ=�΋�m�v-�T���ŷ>�j0�e+U�ZK0!z��]M�
jpJkҨ]�EǘvU�S۽G3*L(Rc�`��]���w�],���g��`Si4����\!�`oɫg,�����U��<��-��H����"�йk�;<�j��#&����QxQ��̟P{((ƙ�������̳�*�RDCFj=ZUtQ4��	�'�W��hb�i�Ȁ>�LY�������$
��|K�������Hm)P1A�ȷ�fD�Z�*�/~EDl9��A4p.�p�j��D���9�$���:�Qw^�PH�����d��6��Q}J+N�]��j��� ����oX!b}��	j�S�Bɧ�E���-�qDE _�F�A����u����Φx��&�bab#S귖j �4�\~;���<ZR��ȭ?�X�A�wr"	mӗn���r3�"�-5^H�>8�a�D	s��w�I��?�X�?����ɺ���=��C��KY��q�hW���H��e5��Soh��u.
nK^3�N=g�����3g6d���6�T��X��B�N�JN�~�yK� ����J��Z3�҇KnibWǑ� ~�F�^�%p�K82*�]Cr�oWW�Z���o���.ίXO����H���u�|����w��}6��g�q_M0Pw�wiwg"F&��{lĠ�@"1��Qh�T������!��W���?���������@��_$kxԦ�Ѷ-�q�MϦw��A������e+�aH�oV��4��\i#����cq@�iR(���&�ʬ�V�[�brE/����K��׿�����cz����/���/����c� :�r�zzR�/�{��e.y�5�.s�aY��g-���^�]E^�=�bĈf]%ͨ/�5�"�x�a���]W��^G*r-����0�Q�0�K���Ŕ7�Hrc4���̈́�#r]C�9K<�Ɲ!���+zs
���`��Sfv���C	��(+f�;;2� D_��B4fv��Tʫo1� ]y}"��[����)D�z�0���c�U��_�0��	��w߽eKEߐ|Z���4���pg6�hē�"��C �"ݴ�}�w�	�3)��8��1 e��n���p;J�3g0Ʈ�$�]�l!�a뒋(!����R���6B���O���s�t?�{�[F����p�kI��*�M�S�By�Ź���:�<iqm>���߇������<%��,zbi��6�����.�s}���K5vVH���Uz�ӽ���ȫ��d��[�<�i���01o�z���DV�k	Q~U	�
�Z��nȷ��3�����e�w�ɥ!��=�J�8y�<���1�O-@���(��+ ���p��k1$iz��9�x��W�#�G:�h�S�r	�+���o�"�*�5��w(Ą�F^���qo�:3�����ZI��:^z��;c��\�_�k�x��P�t��<u�&��>�f\���D.P��5m��r��W�*]2�)z�P���Z~9�m�Z�Ƙқ��f���%ۮ���Q����09!3��AT�Kw
؜�@�n��������͆�l�bE�6h� ��x^X	�����|K#�u�-�����������D�{�bEn@��[Qʏ��بAR�
��(�(�~8�(��'�����ոc�^�w���4���$���ѧ�}?��~��pA7������}������-��z��3�aC���6�F�a�z�T�sZ�e#�Դ]�#�H*�%G`L��ьJqy�e^��f��ud��S��dQ23޳qP�Ti�*�:��HQ�B�O�.$ɸo�
��6%A���c�X2��n��}�����s�t5���z=����R�v{}��+ cYi�~���3H���۠�ۙ�Dݱnwtң�m�-o���.�,���	��W�a�܅ ��l�'@�?�����}MG�'���.���5�˅D^Po�z��F	 �!x��8�7��Ǐ�	�/^|+}褰�]<^ �^ߜ�/���+��l[Di��P�M���߰~����[�<{M�=���#顅z����B�������}��{tu}+�d+�L���d	I(Da�N���t��3�,�b�:��>��Ŕn�P��C'|s�� �(!��#�����b�-B<@� )2]� �$h()}f
� ��%2 d*l*�2E��O���e֥4F�ɟ
��\o�06`��}s;�	�*kL��<!��с\Kx  hр?0v��%��z̄Ɵ����~H+[�a�p�p���ĳ���kz��s3�|�� P�������PP���
��V�6�a�(��;��-��}�+ӝ�I��
�z�ɴ���&�D��u��>3�����i̢�I����|�Šc����jW�f�q'�q���6���{�P(I>�b��X���sv�r���n9�{A��.���~p������B㷳���
�=�����SM1�1�s�~������9&�Ey��ↃT$���%��dTA;~���vٟ���vz��,׸���.���&�R�̮�3�绠�Rq~`��������7��^F��&Zb�Ξ�J���1D���ߵ��D�����v�XS<�n�'�4,O�2'B'%'�{邺D��kTvl���]C�`y�es����4��xۥѪ�s�|+;������I�&����}�>/��7Mf�kk�T%������)O�$�֎��WA{�Q�0�a6���B]K��J��[$[_�����]�[�����E�M,�i�A-�fFЪ�9�t��4)ku���>�S�X3��u�r_���`�kl
Ws� �u �0@�ځ��f}��+qf��]��3��>��I�U��oU�X���d�����F�Y��Г�s������d��:G{Q t��tvG��aM��w���+����Ō�xԫ1-�Kɴ��Ï${cc4`��V<��_Q��)�E#h?�lO{d���b�|�d���^��t�����g��%S���M��W�M*x��K���R�T�1o�
Zg��*�Wi�QQ[�L\h����~�w�#M���G6���kz��A9:!������y�H�N�-� @�G8���ί����?i��{��Wj9c�G�R|���
�u�j�,KdU۬;֒�st�M�Q�C֩�^�g�V�+��]:��g��NS��xK�X'G�����G���D���N�)�B�Q/�:7ҵ拉��hDl|l�l�gR��G�L�?��(;?�}��������Ɍ�X7^��n�S�e���#s��TO���5j���6PAC�!�C�IQ��ѢD>������6b�H~a/��?���	)��O��W_A�?xO6��nN����l���B-wc�0�&���X���#9��@Ӯla��k��C%ƃ6=�~w#���d��!+�X��X_��葞!Q�є)Q��n�:9G0<��IckkO�0=˅��'���I
��(��x��=����)�9?�HrR/.&L���e|0L4Dd���X˽��f�c�����Փ$��zJR�cӦ/�B���5�R�O��7p��A9qC�v�-�)�V��)��#K��;JU,�5�)3��%�q����I�)<뚁p�N"S�}qͤ��{'	*�Ν�.1����$AQ\����WʽH[��ݓu�]��:��TΥz�B�	������߽3�><x��B���d/1��Gi�0<`|��>/r�In���� ��d���lf�,�\6��ǞkWl�7\d7��љZ�)1�C&�H�zDӶ�ntط�"�#��[K

������*�&an����@�CyT��n��A�r"�=����w��>CV��7�s��YYڨ�Bp#�cd�9�>�A�#�ߪ�=i���[�ni�T�\GK)��
_�APKL�ƃ�-�z(�c9�|� s�h&��ıL�F��Wli�A�O�/�"[�������j�Ҋ������-Ƈ 5�T��$�7��:*�6.-�hm�;�|�!R�Z����FE�K��}>�e!�D+�6�~ݧM��U3�� Cc�,$�9\JN=Q��;����hc*i$�I$�յv��Ng��Ǐiss��_��ǐYV����
}�d��{w$hWH�B��?n����}�Z�o6��7�SA��uМ'��qv~J?������u�xY_Z��ueC��M��sz��P����}I�|��CQ˙"�[�5ə�/#��m}ܢ'�|uye�[� �ⲙ/���Pn�t�Ƀ�:��@��4��_�����f�l��l�9{�z�"V�	v���ϽF��=d��R��/y��=��|�3Q�����g]�/l���u�'�+G�$@��K��z���p@��ZJ�U�+�{�^.�L�|nK�2}�2]�tͱ�l��.��:�� h�;��<�߇��[��ghY��������ᥤW���@��i��R:�#��,���;VY��Qԁ���K����C�¾,�޻��"�0��|�~�Aw�[��S-qd�
7G[��Z1cҡS�H�����������_�{O�����-���]ztr$a����/�fk�C����/(V���C������R�QZl&�߸�)<(��O@+��0J(�+R�Äl�DE*!0LT;_���i��M:3H�I�L�n��
�G�x������ٸ�Ƶ���F�T���9
����6�4T�J�TU�r-�޶�[8Fl��`�LX8��-�?$1Ԃ, ΃�P�[���Z�ں]g�ӼO	鷵d֪(�֘R���k:
��G�+��
s"�!����^�h�KA_�,ɀ��rd�O���l��s��}F��˺�8�$�gPI+�{���p��w�p�w���TMt�Dg��5I���  I�1}�*����������5�0Nc�=*���'��D/�v���]�ga��r~ZJ4SHɵ���7+��c���]���b���GS�M��z�U׊��VJcB��LF��B��uQ�:��o�!�>�~���&��DT#M�P�q7���ɓ���4�j�W�����D�S�-N+S�$�9QʩVe
����������3i�d^_k�i]�[�Z����
�i\i�Щ�C�Xi��C�i����=�c�зi���h�Y�l]��L�طf�{eTe^ ���Mۨc	�*��l��O��Pm$t�n[G��[�6���ݕ��<���d�s�Uk���V>ᑼR�좊E�876�l8��N�
S��+�g��guT��&�Ca��o�>��Y�*�RVz�!����%��C9��ЌX���������s1��	�����C!&ĺ�@$K����� ���5��Q#+p�~�&�0tnn����-�c�P����xyy.@=P �wv�y}u%YЙz�6�Ոv6O$�G@E!J�}7��>�S�O�Ջ\�̹2���a(>׌�R�gc �@�^��)?X�ρ����L{������>�w�.�\�]�	>����]^K	�����=�o}^��M�̈^D�T�T�: "�X3�vw��m��Ѥ�Mw60wh���5 J��՘�w�6z�L��O�;Zε�B�VX
R�p>���6 ���ь~RS�O8����O��Đ�wڠ��k��b�#pss���Jң�vw�/?���;�{��֠�+6bxm�!�����r���ެ����M_xj��3�%�M�O؀ۖLԵ�N�b�ҹj���Wyڪ.pO���*٘�G�a�$G���\�'ߡ/������1*NN�e��=;t�1�Q���`��?�Ew���(V�|s�
���3���t�	��B��
j0�
!M�Y���%'�H=�H� �E�C��S�d��g�" E��� �@�O<[`0-��WB0/~|)��b��b��+� Y�w���N�?�eي������b @�E�� *�V�;G<�ȝ�i	P�Ѯ03��Y�����M�̀��R�`
��++Ld��@�&Y�����ٓ�£-�����XW��\��]�Ԭ5���<�t�5e��mXAe���tUѢ�َ��c�{]^�_|�F���6S�0��y���E�1�9�^/OԻSkJ�`tb�V�mi`�<t���k��X�uKc"��!.I�@�/��Ԍ��QZN��~�$�T�T�)*�0��TR�{�\	�w�n̤g1�v�X�K�&3@�Y7��0D�ex�3��,	`m���J�D�E5���!����;I Cks���g�V�iS�P�Bz/�w�5�O%/ɼ���ء����2CԽ�o�F��aK-�:�*�5�,�Lis�҅$u( #��@���iQ��r/��7VHNY�sZJ����w�"1�͓��t����qSYҽ�&��Gw���Ɛ�5�n�JJ��`�Ӊ��&o�\�e$/���aY�a+�KP�QK#��|���J��߈|`��8���t��"�yT�qߐ�a�hA�Gu�x����!+]��:8_jc^^�	�8oϮe�FH-�y ���P�^Ȏ/�A�g8#���pbN&��\4�B�	�r%��W���ϯo������A����!�5�a�{`7U�H�)�^aY�0����^.EG)�(��օ�)�}��k�=(�7$�su�U�^	:�^U1�*Y����Y� 
^T�ŚM:N�O�7���;�0sd��7�ϝA��H忾�IT�?�^_�R>#(��3"7��Ac�6�P�%~W��Ơt�4�f1e�yʴpL�2��SV����~+H�K�[}���!��TR"wwL��sS6��F�G?��C�]0�PK}a�ټ���6����^���_��`��?����/y����=�b:�קo��e��Éc�u*�	����u+���єm��k �nI}��:�1}u����D[f W�W)J��Z�0B�ģT&�{�2�o�	7ڀg����F�Q���A���k�7�����}��.�zqA��;����/0�000X"����p�Sz����1!��
;o�VB[�k��mk��e�������d!l;�hږt��ka^�lPaP��Bx�ڂ�1E!���J<f(d�fŹno�|.��(U�Z�1����%d���v��U�R�JN砅���ZQN���¢ܦ�a�M�-�����TȌ���:+!;��tt(�v�}5����zD�B��О���71���	Ŏ�{=/(1��|oi�V6,�sO�+N�z�C������K�k�I!D��2��α6'�>|^Jcc}��뻰�b(kM�q�ί�p~ySks'�ϊ���ürj�?0�eZa1c���h��ߵ��R�����:/¿n�tg����Rsڜo�u{�5ca������2%�?5Gh�j� �����f��e �@�o��e�!�,��A�}�F����1χ���y_��O�(��<���OV��ȯyR)�o%Ȅ$�E8�[qa7rl���W��_ƍZO�T��X'�������V%t� �#�VUWvi��F�S*?�{0<��.�]����zK!���ˮ����"�'�vK��f�HC4��2��Y3�$��j��nD�u/$�[���]��T�  ��vF���,�r�S�41�ݮCtg4�T��F�lH�Gc��f+��yz~I[���S�k�f����Ye����Rt��R����LY��(��
h��򎎏O�����@���-�9���6�M��Z���':��F �jk5�
�3�+b�i�K�#�Z���S��ŧ�󊺵$7��ճ@_�b7l�ءW���Ά��G[ˆ��^�Wd����,�]�:G�ܛgCD�!����@��F�U+u��I��6� �Q�BdD\J�����Pzw���)�k��ݍ���9��������&�<����������T��}6�Y7s��}��3�ݯ���7�=�*�䡗ƫW�ـ�h�Eg�m����F]�9}I���0��I#��>}��n�l�_������x���菏w%2�: *TU����eFp c���B�ݻ�-��w&����f�M��$31�AG�1k�(����Nۚ�T�J��ʻ�	}��J�%z]��I^��Ζ(��~_kE�l(|��tuy#���,��s���a+k*HP�%~t/'���K���M1@�C7@�V�xa�q���	�k��	�}?`��F�R���6�XqN�[[��v����ż��@�� G���'xV�吓z�0b�y��䎭�(��Xě۩0ɉ�� �e���5���7�	��y�3y��V�ų�F��3�B��Q�BP>��;�H�⒭��IW�ae�Ԏ,�j��eS��B�#�k�|��Q=�6�c^nW����}�{o�GH�O��3\S
J���S0�G�d����s��_�.�?&�oK�����ׁ�폐(3%m��.Tg�F�Ҩl����������H��#Rg��j�h� r���G�.�޻w�{�����=wG@7�@7Z��J��Ͼ��#<��1�M����"C�0��g�ew������uc�4�DE�M<�}��d=���U�N�u߯��F���j{�\<ճ�g�v|�o�k����]nfOC�jV5^8���C�]dz���*��t�Z("`y���isl٦ai��lm!,*����xe���UP�B�lȋ��@*éH�q{�Htr�&O7������@S�����O�K+2(�>8D�#��%�ONUv�f��ęA���s�٘��0�n�L]���u<:��-�ik�f7|[�� �jVBf?�[6���p��=����z�I���EC��(�S:�^$��{&�2��$%�` ���	!k]_���j��͡X2Q_�`[��p����l�mit�VΔ�~GJ����h���L=�a��׳��:w�R��C���d�ۑ�d,-\� ^��xD�}�S�H7o�2Ht���A�`��6D��&�57���h����B�-���A)�zw8)��t�K5�>]�)���p¢#��
��դ�� %��|E�ӧT~1B�k�¹�����>]lsl�WI�+� �>Wun�X^��')�}z_����m4�lRod��xt��';������[[�Z8�b=t��u�GֽAM�6(2Ǭ�У�݁|���W�����eG��^�a5]z�r���A��G���H����F��Ͽ�B���y��c����B�kZ9eS�;���n���o�wn��urtt�ǜ�?\�ku`��l[y>WY�{��4�����Udj=�8֟',� �A�>�u��p��bȱ�i�Dc�9S�+�ga���r.4�������S4�&5�3p>PT�����;G�����>���Q�3�>���Z�D����&TB�?�kUЉA'�n�ɴ[�5lD86��B|��1���]A��d�����1���D�b���	�+�g�ZA�+Ԗ�fZ�B�A!�GhFC�VOup�tt`��=9��u36��g���\Ϭ��z�Hu��n�B��~,�u�Y���ܬp2�H����j�mk�6����E��!sM�s\Q�]+����i`���z_q���1ӗ��7��l����(]9"5I��x9n��㦥���f>G;7�L��۵Jz�R�NHr��:������D���o��վ���G&VԿ�A)������ڻ��S�4����/�Y^��S��KT9��{�u5hayW�*��鈔�b�:�꽗��:Y\�).:"a��LL6~�d�]]����E8����g����~63vrz"�ߥ���ޖ�x�@6!W`
"��m�<T�\�uW1�%vR\]-��L��I��z���Ă��3>1H|̂ā����H]�@�Ģ���0fB��Z)�Å�o	���	�v: +F�ۍ�F��Z��Up0�7���aͲ1��Ys28Ak	E�ʶt�$���H'"L{��!�,Pn
�(�~-�N��~5�P!C��K���j�U�z��:�%�G��20�^e=��m�⌘c� �/��c��R�|[qB�����!�u��e��@eW,��X��6[���gj��A=uK9?���P�����ّ���xr;��(R�(6�t�"$n>����Ai���Z��������~�1�Ρ��6�GF߱���Hm8�]PY��A�_uj������dChĉQyGG��啾��Ǖ�dà/?���]d1ĳ�����{{>����2��L�֮J�*ؖ���C�x�OV3;Jw&�v��I��z�;�lr$�~��͂a�`J�M4K8���CR�u`��5�ؾ(8@�º{/3b#�6�G�H��"l��4v���P��'��/�s�{i掌T��G3��:����n�`����h<��~:�Ócy��1���[q��p";[�l6�T��������|�p*�tdoG�ߓ�|�ȑ���b6!�����'�!�֥e�H��Nv�{m-�-v�Ւ��}u������9:�����B� �96;�i��n���O<V�,v�^.d4|d��^E:}9>:Ձ�G�@n��bG�Ǐ������8WK�9�@����>����5���8�,�,<G4�#�2,B��RZ=���t`�3�d������R���'V�IA��f��xz��ޅ*+��$٬p��w{��F���� SX�n�i2����d��H_��n��{I\�|5���b̢qS���`j�V{ݕ��!7_��0�Y��]���Rp��dv�G����;�w�6|�+p��3��x���L�3J�T���HY2R�ҹ� O̗x��A��(�b���|��F��|��ڷ�A}�����v��3���{]3o;�ϟl�w���nnB���NW�}4
��T�&j�]�<a,��Z�h��ه>W�#��W��z5UJ�v���O6B��������-M�LZ���f,è�����T��x���ƈ��:��}�w�B g
��d**�Q�o>b��Gw��;Ll��y�����%�#��:�G��'FEej�T��׮�_|vm�Y���4�+�zDAeR�70]邛@#=_!+f*�_���JVKbɠ<mS�I����#�WJ.D��P��H�y	���^0�W�`�y��[�ja�cA��c�E�6���	�G��X�c���d-ْ�\��i2ue_޾��Q��t���}`�ttpS5�ǽ���E���0�������e������Z9KM�m�[��g%�ٚ�Є����3�^�WWn�aD�F�06u�H�Am�\��i[o�:�ܟ��̶�:�,��������厴[}��#�h�[808t�֟񺼸P[k���������}��JwDf�8AFQ�9���jB*�eh2���sU���Iۜ��R"�¾��:n���^%��p|tD*����R��TC��b��<:ɠVٔ�U	=�����ͮ�C#�@��ǜqcKuF�Rfԣ~	}W��3����7�A�o0�҅yv1�Su~GC�gwq6$��o���歛2[����:�ݭ��d��g#��93w(f��Xmޥ:����:}ur]؊?���t۷�9�B����7ؑ��ޕO>����'*�����V60�"�A�'M��`�#�۸��ќ�๭&K]:�Ūɢv�?��ڍ�ފK��`��<b��-W��W�L�s`�2v�/ex1��P���5�A�h�tp�96k*�H�"�F<��߈�zZ��&}�_��|08P�`�X��FzF{�P���/&�%�g@�7]�u�ل��-������&�e��W��Z/Xȅq`s%=�piA�.W�ׅBF�à�����C����z*�fcY��R��e�L�]u:���f�s����E��U�(k��� �o��Pr�GAt��Jz��XRn���v�������]���F�[�����#���s�=o����Ee�����^%�4=�o��Yְ����L��Wui�#�%�g��fu��䯜��9��Ϗ_036Ʈ�!��_W�\��u���]����j-��-Ւ)��n���sߋX���m��񊆒Ht�*=Z�U�)��g��\:N�}3{X�aՎK=�.9ƞ�Դ�=��;=W�l������Խ��HA��|>c�0V|�v[�!�1;W���\�(� ]�-8��<������7G���f�'�Y3��*j��to�=�l���a��"xW���B���.ֱ0"�\�Ӷ�P(n+ʳ��/�B;;�β��{�'WB�h�X�gp$��x�m}�����`A��٣_�Cb��grY��8:���ኲ�ّ�����t�<��Ll
�!���h�`��@�����W�$�@����j4Y�Qc(�^����m @G��Q����&��R,��V/��^w��׳�����@�Sw�v�]Fj���v"�k��d�3	0?@\@��z+ud����X��͡|�˦z}u"�x���[]�F�}ö���ON�i�/�y}d�[֢������`jX�U]��RB��5[���5p.���d����b ��"��Ϧ
?�5���kVY^��vZ�et�Yٜm����- b�Rm�@��+^�������0�Y��5�������5)	Ĳ��.����5��/P��p��=��h왇ƀ��ߓ;wo��́��7��/�u�am�D�|�Z�����թ��+�D$�'m=�:4	|��<��:·�ѣm��O?�@·�e2?%�*��r1��@Y[7R�[-�� !tv2�ѹe�p`�z8ѵ��d<��ǲ�խ�^����笠_��_�o|G3��颾Qf��1Ͼ ͂-���}R��Јj6a�=���]��ΉOD�t$]�2����Aot	�@D�`�e�9��	���
��d`@�s�I�����X�O\e�-�Nj6XTT䁫�8��&�� �����~�>*��u.�w���V�6bˊ�:}u^
twg��̕:��5'Dq�TϹ�n��S�i9[�m*�n�:<�ܴq��UZ��KL��l��d�K>{U�T�#M�F���M)K��r�׾�l�-Hd͸�(�6����&�p�z1�§��S��A"0��q��ٔ��4�9�R�Y)x��pj�@0��"F�lT�����۳����H�p�|6�C��s�Cm�������+V�d�C����ߺqZ�s�`�� e4-�)SR�2FehƑŁ�:�2�:Gkl���qu�j
3��/����j0�������xl�QK�=K���^�]�aH)j�@�>��PǠ˒P�әI�2&PRk4����>0��.����cd���V�ԇ9��#�J�l6=�h���8RU!v�+���R����%U��p�,�gJ�Wa��.Q���x�LD9�{���T��UVfF�[��q�z���t���aP �ʄu%`ً*܋�ϓ�(����1p�&�Q@��>��A��Y|��r���	4�t�|��'{��=��d�B�_M2�&�a����Lb��ZI/�1O߼��{n�d{����x�6v��[��`�5,Z�nGm�2�L��gc*����!�&����b�ȵ��'�|�9��tyy���,Ś]%s�1��6�nܒ~w��6(��=]�ʑ\�"��"�Iv�v���5���	�d(m������5�M�$�ls�%9���F��d-,�.\��>,� z�n�o�c�	Ï:�.�S����ʺ����U�j4��sE���� �k��	�aÒ��JdnA�)�|�a���C%��Y��
ނ.�L�pIV�^C����F�|��c9::�^��.�����޽[��g�����J���?���?�����{y�t$�)j�Z2�N��P,��@/�������ݯ����>��ɟ����������>�v/�o����.m_ � 3�ݾɡ��H��6��'a� H�ke�`�bh$0�"A�d].G	}>�%�������w|5}²�LS-+���������Z����5F+zP�a���o��|��A� Y�f��D-�oY���˖
�Ÿ��c���q��-.|�MP��Y��nw�5"�FM�cs`�/���{;�S�$b�i�dA�P�,R���/�)$(bD��� ����%w�ݕ�����Nˊ��Ug���;�p��!p��cU�sO���-�~�~�+}��0�Vn�9K�T��K@NX}Bj5���Wz��ݚc��>�Z_�{�$/��H�_�J�8��m��%��]w�J]�~]��/��:IW��*$�����s����?1�\` ����t���b����z;y�oS��|%���s�n �{��������26�7���C����_��J�>�t�����9H�~Y��u�ы��Ꞣ�kF��\
��6+�ZL�Ki0W��R�r���ײ�F�����sWcS;o�ȯ���aYLk��d�X�0��c.�`��Oeww'�r�t��:��Il��0�^:i.D��3��#��q���A�����=��e��h��U�}�z���a�*H�kM*�9RE#�}b��X�Oj#�<�3�Uݓ�<F'҇ ��K�bΓ�W�*���]N�^Tk�K�W���F�"�+�팙d.
}�cˎ�p61,l�|kȸ��c��8+��e{�(K^q?��+	��n�2��M�zܬ��B��x�B�]�/�S9���ó3�#�A�zQ��f�J���������5��� ���L�vk�_+�B�g��'r������M�w������a�}0"nA�f:���f�I2`U��7��wYf��~��? �f��[�=r��I�+D�[mY��5w���4�̬x~���24.��;):"��k�Ϙ%����£�Y��Λ�7���Gt�<��qv�,.�A踸)�8]q!�(a�]�;��Ro'K/��I�4��_o�}yN!uQ��:�REG<�we�W��"</v��$S 	��3�4@�x��v7�ߺmX�9;� 4��O>��MJ�WoN�: O�`�i�*���24CuR./��>;[�]�ypW�����/䧟^^��r޹#7nu���[�w�^oAj��A���PP���WC'�8��޹~N�Ѐ���$�G�Ȋ���������a5j�̱�{�~He�-��E#��łJ�K��.��9�Z�/���?|�n��ճ����S�O�̂�#�,�q��Xsv]��[��ݡ�@(����^G���r��Ba����ܻwO.ϧ*�1b����N�s9<��1<��j_���Ŝ0)F_"��l84YY�Xr��0�����Z=:c�8}��'���q�@NN���G��f�w��������"�1�rzv��{������Q*._.ְ�S|fiwEC0j�����%�!n����l���uꙂMS*�:���:�~n/���ک���o������#�#�e����`�j��p\��A�g�f�5
��"6�6V��'�4�Bqj���p�FR�Q!��H�C���&�sR��AME��H�9�-�ʠ��!�I�����A����.��h�Dt�D'/�o����������je�%��te����q�ίY.|���]2�x_�MTZ�KjN��*�zs��m��H�l�Z������<�Wx/Ю��k�TF�P��П	�>����e��T���P}g������DF��(88O�ׇ9�G��¨a�d<k���h���3TX�g���Y9�垊���G��,q
� �ul�f���Ճ:����0��v�Y�%n�.B���\&m�tf�؛x��W���~W�����,+٬ʌ.�ca�HN�w]�|Tf�(��Cfst����k$p�4�k�5�b嚍�9~�L�k��g!�Q9x��Į�����H^�~��]��������F����E�*aRdn�����z�M�H�060�,�������"d������u��8�]�-���H���^�[���Q@��`�Ǣٰ�d9��h�3�݄��yP��GC�t�����#����5do�@m��8OQW�6��sB���m�j_�^,,�@�tX�md.��r_���f��M�(������k��~�N9�0g���N̋*X���_��\�-�� @d��vV��O��ʱ�)����Nl�p�O�8�l�ڸ�,t�U�a�+Qd��d��ƃwߓ%���zy,��\G����9�w�gަ��Z�z1Ի��������M:+��H.���ŗ߲���nK���Zn�ݖ�;e89�f�+B�`KÆ�89#�2r%έ^���r"�ǯ����g���V�gK}�m�׏����:$�q1X�+!c%yh��(@kM
/��˞O���.���v�q��|v:�/���Q[����R�Ou��ķ1��W%$e]\�`��׶���ɣߗ�}w�I����ν��o����Sy���5���P���sL'g�tT���c�bQ-�`�jS�:1�m3G]�C�)P�b�����D=��|����Ν��Kw��'%_�ە��7���T?7�'ZС�?�!w�ޓ�w�S�O�_ɫWHw��9�E�htX.Ҫ�yZ�XJ�r��s��R��e�[>x�U�t��1��{;�U#���tF�)qD����6�_9�zG&��cگ� �)��l���}7�5���A��G��Ɨ�g�X��{0�����w�(��l){��&�N�9̕�J��	��'o�fR�Ш,F���Ru�O"�������p�>5�]�[\S񭲃zTX⤢莾A�c��� ~6�c*1F�}��_��ɗ� d����|BUZT�$,���b�F�o��x�ƚ�חcj�M�{�f�8t���(^P�4�K�3�Cղ�n-��ni�s�H�k)e�d���r׼�<�P61k	�p�R�g~�����ݽ]� 4E�En���N ��6+���.0�H�=^3FՑ�&f��"k-����%R���ݰ�b��ƙ��:����:E��]2?.8Uy�6J{:ܗK�|��qV7�,d�]������lfp�TVE�[NYt�fb�$B����@vּĶ3��g+�S^��î	�cM�WB��5�*\�]�B\�o�q���s���_�H9 �F�Ƣ��FhK�0	u16���❜]1�d6��Z�Pp\�`d�
cB�n4d%4zD&6>�s�t<��9{զ8:9����̀`J�.ψt����0��dʽ �*���ޒN�O'��l$����Y�dv���q�nw�v�=�nݼ�ۀ���h�����0#3�0ꌌ��0.��P���n��/e*��`������\V6f}P�Z�u�1�hV[�c\#$�8�c�[�̅�tf����X��za�k�I;�*��%��ɵ2ȴa���5B}�p|d��t|kY�x��ٹ�@R�l�"�'��)�<���3��W���͚1P@1��Gg�V����6z2+���u�I��lx���C]�O��i��z�ܵ�hu?��Kٿ3���Hg;WY��%�fߓ~�`v�v��Vh�g����Ϛz��ȡ:��}�g�vL4��s��8���
�ޘ�����"ynޱ	���ٵ,[X�	�`p��؜���|�s��Pm�Hq���O�(��!7�DO�yx ���O��]d?:���`!�geɚ'7o胍ԃC��]���E���.^��;�u(�ˡ
���~y$�o�:3�-�%7x�]nLZ�p4��<��˫����Ҕ�����������g�_�.�x2�cq��=y��{L����>�xqgw�B ���|���:G���g/���6�dj��z|�f�T牢U�������Hӵ�<�+�����?��{M�)D�����p���'�IV
�T!:I��8K�3�R��\�"�Yº�6�������1O��Y,�B�w"�<�lWV�A��L���N�� �Y4l�b�����T����K�q��M��ņ���8Ma����y�b�ѕ��mjl��z�������c��8Wu�(��e�'>���c�z)�ӬAYM����
�����ux��hA/(�
�K�Ϲ�
�k
#Xd܉�:v.Y����z�'�G~��pD��g�������X1�d�X�lZ�`��H4�$��IW�۶BjD�?{���O<�J)'j]��4���f���]�΀w��ޠO������0� �B54t0��) �g
�ˮ����p�5u3���q[3��ƾ}��{4�mi��A��
t*�"�'�K"��'�%���Odk�=���ra#VP_%�t���d6���aY,�/2:�v"�.>��+"��Ί�8e�We��g�t3�E�d���P�N'F�����^�t�2�?:���{���p��`g�"Fٚ{�P��/� �d�9��G ����r9ҵڝJ��a$�3
���Un���XF;�AT�g��6t���������L������/�LpH YDXWX˳�u��u�������ߦ�ـ�P�K}45�^�͆Ñ^��ZZKo�ؗw�{(���V-��9���,gS�8���n�"Y-��} ��r�'z1,�"4�f�5��z�{�w�`��1��&����XD�a3�ytB��eAft8�&�f�Q�5��ۺ��s�M�j'��^��<f�l�?�H��lI*�a�_�9�����3��dB,wm)7|�����{1)�B��A� �Їp�|��
�&b����Պ���z�A<����9�y!;j�s�u.єp�-�ytr$���S�VK�r��ޓ�XN>�ό�t>�j��L��ZY֢Q�La<>���c��#ȿ D�o���:2R�����¨���l0[@��T���`x��D�Y6�1bD� ��
S�?[����eg)���z5�1
ƕn>�Et~z._��sb�n�ږƸ�7�_Z��n���9�/"{{�]Ámu�'T�-&���=��v���W��?���/��a!�BO�h��:&���y�����(����ڡ��G�ztn|����
���ܺ}��U����k6E�+N;>>���<���������͛#FHe��튱]z�q�ŨO)�*�s�(!"��T�Sr�����o^:u�j���<0�����O#ko�ګ��
GkNE�-D1��'���Cdn��*�l.���f�^� Ś�5�:��Bx��#+6ٜ
̎�a�� r�@B����B�(vP6ba(W��h�	�2�k�Sdִ���硷M�)�bi�0J�k(�r!�@�м�u,y֨F�3��
�i��v�,#�Yp(|��^f�χl*
!3�Q79��f4+f��	5��<�ǐ�,Ӽ����`�)����@&�l��_�_���#���`"Q��)s�u�;t��ϬfC+�s�fu���!�d����!c
"�Ȫ�k�#��c�Mk��4B�2+���\�+�yKܺ�]#q�~"�4:�	
:G�&���@0R�f���b4�a���ND�QѹAԖ�(��ƌ��,�:�
�;���e�y�T�1z�"i1�wUxs��� �����P?b_ ʯ�X����0HQ)��R�EW��-b�1f��_Ĳ_q�]5�yr�'K��"���,�5XΕ��M�)�[5$����ݕ�H��y\�R�yN� (�~�`���n
u1>�����uĕ����܅��e=����7rØ�$A������,\���^�=;�Ӆ����S[��u�M kv�e:c��S�	Y��4�&i"��Ư:	��B�9���Ky��:9C"9PB�����+E��(`}�z)�{�Hӛ1
��m�
�B[�H�ْ(@��-�{��|��	�6z�18RX�²d�mY�g�[��� d�~���I>�ˌu,.΂2�l�M���ԍ��!u�#6�EOHP�E����I�.�����|iA	�A(���p@ ��j�� �����<���:`�^5>?ۇ,�� F������ش����C�\�3����SOx?����>�Z���4{:.�"�&�r�I�D��kD��]������l���7�,�PO��S-���7���;��7�,�>���\`$Z`:\�97K���|���֍��S{=oV�G���t(�c��ُ�!��Nf�7��@�е2,P<�S�����L��(�f�R��FaTn|�˕�MV��)�`Ԡ1P�i�_^,��Oku$.��/��tP������U��퓮.�d��(�B�xï���Wrzz�.��zF����ߨ#4�7�f2�\��"b�׫�CcF�3���s=�������5���>���:��Ր�Cu,VO��d&/^����ȝ{w�giQ���,�����|����?~%�'#n�_0ʄ�����?\#H�B���)�ɼ+VUD.F	��J?�j['1���7�\��j�R	��T��w�ڜ��"���
O��/Fm�i��D�1�d4}M���<�N[vw���� �H�d=��5�����)%�3��tFnBb�/�u�AP��Z2z�p�߱��!'�5��{S2Su�3[rc��7�����!�g|�J�c�ꔠ�&��3`F{�g�,B��,؄!i)Q8�D���PQ�40�� :���5��,B�S�'!�����k�F�� M���p� ' �v��.7c7V�C�B&l|�& ��������{s��,�D��~>svj��@� O��:6C4ri,1P����.� I%n�P��H�
�F0��!�V���4�M*�#<���M���R��Fc�@�R&� ����W��{��(��>��M�?��N���yֽ���������C�}2���6o�>{Ƃ��lV�C
��\l�3ZG7Ȏ	�ɅY(�F!�%Fז�[�'�_�	GJ$	8H�0�o�A����(��J�%K~�>��FD�ax��ؐ#��R~s��_���	ؘ	����=qd�����h4J4l���F��x�p�(��5����n8�a�H���`
h���].39:��*�!��FM[V�1�1�3jS��'�BŲ��a�r�M�U􈙟�T~�)�W���U�w ���g�Jl:HcYl�Q��:��@PT��T6�+�W��m�����'�/�	r�9���{ �_Y��f[8ֻ,'\Fd���R��d�2G�:�i`�D't���C��@D`2lg{_���FȖ�zE�]��U���ܧ���9�duRf�|��J�̙,jU�r�t�Ċ�p�X3Ǿз+˺-�!#j;�+��j�<!+��l$)��Q��w=u�x2�t ^���S$���������q�|\���Q꺍��p$� >ʒڞ{�f޸��CقE5
�8�Y����ˉ|�v��p�z�/?~�F��.-{���A�j���_��\h�9��Y0g�uazlO�1�g�֞M��N<{�Jv���ܼ�/���#���]�Ѧ\�Bv5OГ9�`�)��:�{[�{oW}���;���K[��:��tU��|���I�K�T�z�0���n�R�i����<f��Ѝq�n����=Pݵn�3�ə?V���`�5�.���z1����>̂�zQ���Ύ����i}(��*���LPQ�wcG��H�9%ލ��z�-y-/�����!M��tp&�K+8�5'�`i��?���ѵ���Dfğ������Ά�l���kls��f��A9}-ÑzrOߨ����B����bJ��ݹ*�ׯ����A�*���~�Я�q�`O�K�R�!�B�80l�dͻ��t?\��[�����m�T
^�f��]:eɘ�7��W��6��<�Z��G-�7�e�a(�~+kd�:Mٹ�'=�@�?�+�S�+�6�M��/����"4ôOAC�/6<X&p0���aHommS�Ø��ǧ����tc�(��OJɷ���} ��>����v���8G�'�=1ꫛ�pF1�!<%�%�� /t�}s�!ܿq����Q<���h�k����gr���pf��+����\�ݽ=��{�=d���`k{�)sNb0���D���35:�4T�ᘌG�ƾ�QB��w�,����>�,82�A��H�\Tc�A�˭���;��FG���$p���>eR�cu2v����w8������w��{x8VGo
�耎J�9(AȎ�l{�(�#�}����Pg�L��r9J�Ũi}�$����<���w�����~��.�����v�2��IFN
cc��9U+�8͆���"ۍ4�����F_Z��%�3�o�  ��IDAT�h���m�<�횧����l�����)3�ESBV���JC-�H���22��.�{�r�<BSY��L��i��=�����J^�]W9 �\��啞���I��*G�4���Q����I� �$��J�g|�h�c9Ժ���FE���b��I˙�`�q
�B�����ܠK�{�@Bgp:���t���l/�����3��i�z�6 ��<����>iv����y4B�c�z�%\8h���p>�#r���r�raipмA֡�/^r/�>�����cy��PnݺE�����t!�Ւ	5F��`W�ߒ�w��-}A�<�X�mtF�w�����X_uƦh��)�7]�N��(�V�T�� L��&�hfo`�0&kc$� d�}���i;������s��b ��mZmZ����! M^�k/`�3]M_�U���VX��J�7���^K�C)<<����q�mcNIVo�e?W���/�ׇ���8���ń�=j���ud�2����j$�+JF:Nj���v`ݙ���$����ض����eoo 7o�ҽ�H�;Hvzi#S��9_M�`��έ��w��|���<|�/�n���,�y���{�����=��~�:�G��L��m������Nk���ިn4� ����4� 8���w�m�|�j`�6JQ_Y�ҚӐ"���x�z�H��UH,.���%o4`��ُz��lm���s��A��R|����1;̂ �s|�d�st�E�0D���Cv��K5�fLњna8����14ҿi�9�K�nU��~/�:�,&� ^Jopʆ����c������=`Ty�+�1x�j�p(0J�r�Q�L���WH����Π2>⭣�*�_��[�������s�p�Mqn�7ٺ�S\㌥.���.$����Kj_"��E�@ܱ�
������ǟ}*��+}���������/[t�ź"+�
���@ț���̚1àF����yx_^�z)��KF��m:���?� �Ź��\���u�ep�����7���?������6����%;�����h;kM\F%|pp�N"�P]gjT�)�����~l����Ãl&������]׺���ϖ���rV�
c��=�짟�R~󛿑;wn0���thJ�4�d:��*=+:���S����ZP�ExO�?`��=��ҵ
��:�b�0 �h�i[�iDsF��8t�,� u��b����X��F�zW�	��:�(����e� �d���䚌FB�O�C 0W �O.���P>��+��T�j�A�_h^v���9"��kJ��qS�F<+xJWc^m0[�/fzt�m��Z{U�j0�U��ͻF�V���!�m�M����_�k���,�����c���ց�D Ad�]�;��Q��� z8��(/f��"h�*�g�A��*� L�dQ�8�s��TNP���l2��ȥ���n�������������+GG2��T��C]�Jn��E�_���O^��t�m���s9C�U�^d�CRPd�	b�#Er0#ʀhq��4R�E�P���fh�(8GB��̡��[|�p�>��;+i�EZ����d0����ϙ�Y��u/�}�Н�X����8�v�?
{=Y
���(-f5�nP��d�������ˀ�7�|KGeM8��i�u=z_=z$7o����^���BiXM�/3z׭���7��1�uƹ���Q!�}-1�7�jP��ͯØ�LY:��E��:%���=�:� ����o۝>�Q| ���Z�m�w;Zu+ip ݟR�[5>�,�l�����g2�(�qW�G�t���+6]��WǔT޴�#z��e�q^��"���M�����^@����B��D~z�Z�n�1�/fk����>\
�8Ԁ�>���?�1����<���A}#���Ag��k<���-�X������k7��wX2ۢ�آ<GPw����}�J�&5��?��W�ۃ�_��7� ߽�/������?0Nw/��Gd%��!3%26�C-Ƃz^�r�Չd����jiX�z�XH�{�x�1�E��[�?x�N���77�aD:�2�Cgc����&���o�����Sn�����`t �8���tTP�f��� �68+��o�L�:n���<��fH�7��Z��6ԥ�?]��_#{C���>	��pm6��(����i�1v�9�� �;����H\s���i�ӿ��q��U�}�o�� �F\y�}����|QFV*GdM�«c�B������@>��/�o�7����Y������xu�_���祝����s?�S]w���=0��d8��XH���5X�B�>��N��^���co�.d��j�����t�B167 [��Nt��˻��c������prn����͹� ����X�8��Ҡ���`=��V7t>�Y�A�����ǿ C�u[M4�'����w�e	��
(ژތy��0ILgP|�H��#�yk�7����~�����'��n�06�:&5�e�8��Z��̽�]9=>���U>r�/`jȬ�<`������kf:��������4�E�g�T�'�g�!B����B�����23�	���N�ё�D���t�ؼ�T�����G�U��u��l&��ݢ#�y�.XSx��G����iu�����~���v?��dM��%!R(��1<��D��`z�Yu*��0&��~��P�Xպ��?=ƾ�	{��ɈNN@�"�ױ�󇺏�!��F���6��),���j�dp�'���Ġ�
�=���W0b�.t;7��Wa>rF�i�pXrfB1���+�U
÷^�-�7�x}�m|6LWZ�	�g.�u�3a,���Ɵ}��u�{�Nï�.96�t�qM�wQ��	��.�ʝG��a܌%���(� M^�q�jr��j���ɥ\.3��G����n:�1�;t�����F[���-�k�}�[=��u�*��͐��4A���=�]�FƲA���.�%���=�&�&9G�	8�{��5���2����9��7�X ����Ç���{�׿�L>��r��y������U
�r<�:֗��5���ޗ�Fq���v��h}x�UD©�҈�m�tNVa���h7D�re܃�1�C�:���:�Rw	yk�f�z�u�{��I����O�x�b��3��$e!�F� ��?V?��s���Ǿ��.������DS,�O���5�ַ��4(͠�Ѩ���}���fmśWGj�>��|��K�8��D�o�<��y��o8��O^��^2?��p��TΏ/e��uK��.��6<��g?�$�����ގd}����%
�����ր����x���Ԉ�lW�����5tS���P�W#��H��vWn�ڕ�߿'�|�*�=F� y(؈�hzqr@���Z��!A�`}�,��^3������Q�G��xu�cC��P_�/�wx�Ũ"U�0$	�g��'SP8�/&���K5�����Z������tm��9��u�iڲ�t���.�<�e��`�Ta�7�AmB���H�����H�X9u;� %�j��]il�Rm�jo� W���OUwY▯�ޖI�a�mV��g�>(�nT��NJI�U����|0>���ln�[�)�����?��?��(���7��~��5� �l��n˂�w'�4�` i�춛$^�φ��gz��~nB�7�}���z����A�|�XN��G�	��3'j@={�����Zȗ_��P PBn����Bt�?��":v�Y5	m*LTu�t�1F0������Q����	`�1��cX�=zĽ=����,���m�sF����k
�D!�|�=����<���"(_0��;�M�l�{��=ʖ�%��x�q�0Y�t;Xf W�|�@�B69ZX�c:���?=	
2#&���߆B����&fH	���ʋ�O����ud8���?>��1��z���Su&&2п�y�>{vAxQ]�Q`��db%�u�`.�6?��K���{Ox#<���_��f8Ԃb���-Y�]*��<���+;�J܇��Rf<��D4,3Q�>)�B`�A=�F�ud�[��F#<o��7�t��,B�12'F6`�)�]X^�8D�Wo8�u䋏��$bXS��*#Q�����Dd	��Xd�TR�>�AAB�uH�q��}	I�O#=:}uyfF�/ﲄ�^�+�����s�����*���P���UΑe̪1�?�ٝ��V/Sv�����5H��H��WLYV��Ӈ+�fP���K�#���$�X�L������R��5k�QK�d	�ra�d �i6:4V$A��X� ��Κ2{!�(�5�DT��T�e1U}K��!zo`Epho������&;@X�Uw�b�����=q�\G�~����:[|`c�k�찧vwwi�ݽG>��c�{�e�g���$%mx��/�%���������嗼]2��3����x�{$��X�A����(��r����<�'k%6�@���X1�B�ӭ�M1v}Χj-At�`�dϸ��q<6��ʦ
u+e�G%c*��Ik��ڸVc��HrT��Y�`��Gb��������0j��ٚ��7�9
տ�˾</��/��ӋW �~=�ӓ1�P�g�5�Vî�����١����r��v����<������34?�#h��x���|�t������o8���$- �<�8V������o` �����������������Y �/1��"!����ͮn�\��� 'F�|<�fk����l�`qiCC�ъbJh�
����7!�V=uN������+.h����]Q�!�	�����z�t��T�0�����b4b���T�l����(�~�,F7��I�s� �]H��+�и9�� 5�3�0F�V�.6���,��IY�F��������&��].�I�����f^�5/�^��}l:D��]Vo��َ�&M�_��{���-�*�P�0�Ҡ	_1��؅�]���z8D��t=����淿�[w����/���`w��dI�y�U)��m��P؜E�v�
�СA��~p�]�(P\�@�u�4h>�FO=�:�v��G�������O?��ݕu�Q[��v8 �-���Vgb����������PT6[p�X@�F��,n'%`i��@D���w��
��A&� ��� ����4E-�p�@ Z�^&?�z"��w������
����>�?��X�)i���ŗܓ�c�	�Cqqqκ�-}^�/�`���������O�tzfBQy$&�)kCSC҄�y�bq�^���h.ڀab�C��;B@�Gc��Cl�GG��8b�Q��M�d�aL������l��������?��wnJW�c;���d���D��W�um�D�51�7v�D��B����8u���fΎ�(4g�23�b{���bg�ʁ���zk�	_�s���z���3A�ST���)� �s�G2����@%�6Q�BW͈J�I��\��f��2B>VT��9���Cs���_�=�B̎����q�=k�x����o��%��yLh�m��N�54�f2���`�gNR�18�8�0B\�X��[���cg��L"��t5I�z�\�h��f�$�G�<۟��: ;E �)�g��œ.�Z�6.����o)��b"K5��#:�� �m�`�u髀N2����#ka8b�Gjd!���Q���7��Sl�s@��.h��_F�ML�s����<�'����3��\��ѡ��$�h�\��fx�zG�X?#�+`��lCf�������]ʓ'_���'��o)�UJU��u_�^���su���[.Yõ���Փ�2���4�} �"�5��=;�`�0��9�9�[���r�m��E{�Ž��B�6ԃ��#�2�Z\#F���d_���(�;�������3�s<"�V��w�
�+���c뒣J��&!�dCS�bɡYC1���������-W�ʟ��pt���c�Dnj̳��鬈�xjK���-��/��ձ�?PR¨F��(dX&����O����|���r�֮l�N���&,�OO�Ν�rrrJ'BMKa��qx��e�۽e4o����(���(�ِ����slrMF/�@�4�l�8߲B!q��[���B��1�2��b���	/�p�����4�Su��CĂ�^m2��,�l����A�Ū����I�{#^(|\#�偙F,�DUT��v��g}�v�1V�#�c;/��Q���%)uM=�`��m�A�\5N\"0l��y��P\d&�����z;}���7���,��p�8FM�V7$���,2U�Sx���a�,�����w���o����ot-��o���/���y}��nŢ-D���=�S����`V�i�i�a���5i�^XM�42-Qd��
�>�/�b��nˢ����8g��˗�(�Fb�n�)�� 7��ˋ3��[�7	��
����8�	�Z����i0#����?p8n߽K�فFC�La�RR �˩0���]�Kn����r�B�X����`VT���kh��n�"��a='p_Ȗ�cFm�:��H�Z�ؘ�m4 U��:u�<��xe,�/B������t< �B����B�k��N>�� ���v'�:l�P� Jv~v.�
Ѿ:L^?��A����:~�do߽)7����sna�4��\Ula�"���C�{\*�c���vY�[L	��ydd�t@#C��B�B+|��1Jf@U@U�,�z �b���u=�
P��A n��MH)�H��Cas��T�Tp��v5�"E��z�;�
�@
�j��Pc��y0dB�������f�G�2[�H��vS���Қ�lW�g�\����*fB	r;��揺ʷ
F���a�_�qv��܎�?Io�-�y=�$���Z�T�Rt�
f|ү�^s�1�c��Hl&h߃�Uf�R��j��MFy33�h����?��s��ɛ�.�k<�rz>W�xL���'�AK׷~F��%�[�=���k��{H�$��Y�r~����`��p��5�*�ZƸ�^^�w���C���_Ⱦ� @n�ﱏ���������;��`�kJ���T��#ǧ`9��^eg��Q��}	���\/��	�����?ȿ��S�??fp��ޥ~��X���Y��笠"��X�TeЯ:��
����T�OG�1�y�����e^Cԓe��T�ck���0(ڡ?�QR�Ţt���Z=:�ហCPG�F�ї�o-�lP#�H����I�p��2:p	�%+�/���\y��!��1����lo�+!Sh� ���Q]1����kI�o�`��P���Cc>�r��X�:W�p���Jm���͂Pq�j��X"[������8'gj׷�6�s��*�(�Y+P��,b1�dxq���Ru���=�I/�G���FW��ќ�1��!�A~�38?=y����j�j.uQ4i�[�(���&�(*������,�,���\�[Kv�� ��E��bq.����7�F��c�^5��eE�(�����0t)E�'�4p���"�����ºC��ryn��6�1�cB�ߩ���rT xϹ�8��E�2"y�e"2���6��]�Qʷ���x��]�"��K�=uv6X��Ki��/�bT���}i-ԟ��̕�wgf�}eBWl`e�����E�)�+�{8/<�Vó������?�ݯ�_�'�����������O����T�?x_>��.;��c9������"v",2�M�f+�����i��4�K<xL�c�(HȚ�/"Ww��1u�C�gP"��\(�]3´���h,	�r��e1�r/��77Z��rJ�g	?���oh�5�=6�q\Z�#�J|��,t�曗���o-
�U0n��o���r��>��`�ú�p�:
��*���3낿�G�]�5�V僆~�12�X�d�h�m�x���s	g��V�&�q�u���@�Z��K֙��E��D�^��}�
�o����� Q���!.P��a�5Eس��gFo�_����%��-�ssdIФu<��Ҳ�(^G}���Pj��Աc �-���b]��6ދδK��(e�88� �|$$B���ʛ�G��az+f�J3qt�!$nk��Ǆ�?�s8�7o�b�HБK�sTW�Uz��!�mK�񜥢M,�+����%$)�vѱI|U���f��1�4C��b�p�t] ���B&Ρ>�jz�%h����E�ޗ^B�	ѩ soV�ee�E�QM*�Re�4�3���C�D.���sA�x�AH�D���<2��K��qE��%e�$2|�j.z���Mכ�����VSbh��ڢ�E��!d�(̭�bE7>@��"�l��q�o~�ְ��u�M�8)��fU��grt2���z}��P�`W����$(89;����|d��+O̜�w0�6���~�{���:���,�D�=F���u���|��jE�h����D�����W�vn�?����R'�z�o�r�aO�(g6����|�ѹTv��P>��k���o��x��c6�]7	)'ErZ����[�oyEg9�+J+8u`�c�������.����e>�}��a�'Ȉҝ����k��8��!���\�m�`�$d����C�}��P�nN�:f9���%F���,�J��{j�I�ŀtt�+Ϡn�l��F���D>�l���wTNZ������rC�0oz[4�TNu��_\�o4>U'�`�6���=��1!���v���� �L�A��Gfs���[ЭХM���<��vM�}S��fȼ,Y+>�8P�wd�����~)�����2�����������O?�V�Ń;{[Rp2P�	��Ď�Ù���ƔQ2��D�cSxϰ�,���b���9����_Rh�'���	�6��w�m'��>�ja�ԼcQV�*�{I8��ІW�d*�Q*���P�^e���O�ԣu���l�d�-�0b���ğ�
a]��J��M�9�m�ōR�5���kW��T׻��N�8�a�ٙ|S\{?��HPv��5��uA��sl�	�f!��e���X��1�M�����o��7r��M��<'�ҝ�����f�X���q���䓿����W���+�o���I+͕�l X)5) NV��0�Ca�v�HO��A��B�sr�R�7M$��S�1NGhd�X`�U�O>m8!�2 �!!Z��$���"�߁~i���ؔiiNM�[�0<�qE��or_���0����I�\3r�ը�� 8}&��f���A�0⁍ȇ��<we��GaаW���_��W�M�ԿV���F�m�ό=K�1�gD���a�	j]�[V��gPP!_G�qo��� �x���
���I�	����~��0�ҡ�G��Y�z��ܕ��f�,��r�Ֆlaz%���{��j (���"�&n���x�|�z�>`]©\���̤5�A�<��j�.�����E�Xzr�5<���@Pn� X���H�`�����Q���˂U~-~�f��A��<!�PXd_9��j}CR�� �f-X���������x9ro�6�'���@�W�/�@�s!�Ɇ���B|%���<�l`Ѩ�T��0�zI��F��r[=���k��p�Ri�F�\^:���q�m�&g��A_Y+an!��qh��i�a�)Ö&?�z�j؃�/��Q�α-`q��J"� i�,EA�˜�~���st�N�х�}u��]�B�6o����|H����K��A�f(	uH��|8�) X�̫1|�敌T~�z�B�/t�����.��0��|��@�+"p�Q��?�qO�����vi���圈�������᩼yu����y� ��$�YVl��}��;{&)o��k�ҕ��%S�vY��«<����@n���:Z@��S[��Ɉ�1;�]���e�,�*@�˻�O5*� ɝec��|=�,f4��g	�����X�b��\�k×2��̰��0♽�esVV�~W��ܗF_�"�8Q��U���2IL30a�����=��>}$���}����u0(PG �z�Ho�f�AkB������笎uE&�e
t*H`拥��R��l8�+���xg�/h_4��:j4l���}+_���9|ŵ}q~n��@�����������[=���dgo��ᐠ�����kS�m�3BP�!=Gń�p�h\��(eV�H��i��:��B�N�r�>640�P~X�l����W0X��s��h	"������	jY�ո̹P��)��57ת�����B�����B�Z��9.KF���B^���Xޚ�����j��?F�����dr��+Q����يĬPr����JaV?�ظ�����Ee�/��a!+��"`ɳ����t��
(m8��/�����ɓ�鳧������d>Y�W_�Q��s�?ؓO?�T��ٹ��O��d4{_7W���zԡXQ�raX%�#po���@���YWע����BslX��2:Pj�s�~� �D}��j|��'�ء eDt[��B������d��5�f'ϘM����qX����m�tN��C�,�I(`����/f8��.v�i�6��"sՋ����a*�0VQC���=���x�#��sy���즣�0x�@��;�#������b����]�um���6���A@s^��� ��R���`�J'�u��h�oݼE���wO���HΎM�5���<A��v�������}���.��?���z�ܔu�Z;2��́�����~/�8=���i��V\���b��d��E��zvyo"#�:�p4G7�"�1\{�N��<ᕅh��-���&������L��=6�g9�,x�,<��)k]6���Q���\�F~P�ނp$�2�nE�d�d>�?"��S�f�Ȍ�w#k��~,pJx��:���4I��GW�n�̔��9#.y~3�}�
�(M���6��#Pp}Y�+t*�ksE�0�����ܺJ�m��'���c�j#��$2�G�#��L�`ڥ�c�.�;`���6R�E����8� 3U�rݯ� M�G�W�?��ʪ��Y�hh3��[�9����j���z��1�5=Qv#/��!�(	D|Q'�^/P��osߵ[*/��2��0�������8�1���YP�OGC��D_�(� K�>�I����=�(��[uX[M�/X�F�t ���v)�=D:��R�(�%�X�y��Y���Z���� ���Fi�`j
o,C��}T��DQ'{�G#f�� �GѾ���aD�1���Z�n7�1��c�~Q���Z�ewr��b5"�.�7��@7w�,tO��<	�� ��}�Z"s/��Y�$�#���W�R���X�^s4����zi撯���9kj��~��?��_�V��*��owH^3��-��k4�	YF��:$sW����}�8�I��Fr�l���Q�����	�c���V �<�"�f���y-w��$Q L�ǡ�����o3�$�Ў^��{/��ݿ�X�`�2�(�n�X*X8�`������Â���)W��YX�E0�?V��Y�4ⳝ0���FP��n�M{Y�dM6�Ō����M�A�BF7իFD���.�+�T�3*]z�ya4�`HA�%��l�JO�6&wq%����#������tզ��9!o[���(�I�)��<y�%��������F���lf;��s�l��<E�\�stČ�x���ʄdT�u���~NB�k�}�7)"}���\\I�~w{W~��G��7)���w��j��{G���G���_۸�QK*\�pe֕�bD�L1��mBt&��ł�5i`���펢dց��|��;�����rzzʆW���H{A�����@� 66ט��0>VK��'�I#�zD5$D" P��dF�ftޛ�5����FP�=&9*O�f�4�{{7��~��3L�_��ǃ.!�hh����x�Bl.mu�:�ؑfm�Ll�7԰(�}��<��]Џ����L9G3:m��	���r.�s�"�|�q#,�����k{g�ٞ���u�@���rv~&ۻR�6YZ�|�l�� ����_��} �nݕW/߰���3������E�)9�ͪޣ��J��R��5aEJK�d����P_�2륱X/��'�^hd�@5���ƚ��e��WB���j���R� Y<�9!�͛r���q�K� yLW�{�{:֫T{�z~#��0�J=�Fyͨ�h�c����0��%���\Z�:�p:ZMd��`���ɚ�x2o>�£(Q� �RU��@���C}y��,0���UB����-K�P��� 1��9�>�;1�`2?`�_9�$0����I���2a���(�w��&$�3�L�]з�tX��`�'�Dt���֡�ϲ��i�ƒ0K��كL�T �z����pԢ�z�b5!�_�t��ˮesB�i˕Ϩ+%|$�:�%���狑���9�ȡ��J��xynut ���qc�ό�G�(�*W������wz�m���?�ȸ�EQe������z������1C݊ʔ�p�  �d�Y_������sDJ�!��rf8	ξ:�k4yt���a-[Ӹ�O�� y�L4�ȑY��~������W�`JƹS�� �}�f��s@�8C�V�+�J.�o�*(wc�(I~������feVJe\�/���/�K�򩍓����S�ԍi�		��ޮ:�@7�'���c2f�z� ��l���&�<Z=��\�ʀ���n��7�:���V˺�Ӊ7
d����?��A_�ps���9�vU��h
�瞭	N��޴ɑ��Ts��>3���2��X=�s����|XY��ó�WvE�2��d7Y$�������/Nw���T�܁������H�p77Sӧ����ox/7����y�����?���<�?6�/��&��b���'�����e��ʭ��c�/,uf{
'�:�ӧ�D�R�"��
<�tO�f��hJ+�����3���(-�tp� -��2:�WԥE��� 8� �v���J5Hc�G��	��k�&�(Tu�V��֊��<�sr����G�(�s��t���m!�M� �9�?�bU�5����,��b�\ì���W�zM3+�����hc6���$�e��d�1��1z3a�E�s�������7����������::�$��~��>������b�6%�����[��x	�qX؋��6�5�N�1,
��wt��@6N�Bw�< J��5!���ｸ8�gϞ2����(�C�)))�@4�a����"�C% ��Y]Ye�t�u��N2{G�k���M��l]]����^;�����O��O�<A7 ���@
��T�����`��OOD^W�	Đ�<>>���_�i#�6�?�q�A�ļ��n�b�׎{�"��Qʰ�0V�ܻ�B�>�M��!� �
��0�����uf:~�@>��p_>����pM7|�������=�M	Qh �b��.�g��_Or?�AM�'-&���Hs�Yc3a�� ժ�Q� ���p9)�U�}V/Tp���ȭp�����Jlw���9 �S�?��~;�mJurQ{d���&�lS��V�A��b�,DK�ՇJ ę��5�@�֕�=���ת����`�����-t��xF�ѥάe�soN��i?Py�xBY-e�<<�\/�� ��Y|*қ�N��S1~��b�Xp�]̈XM�|�F�{��U���X����Nͨ�8K2vI%����ҩ8C=�-P9�b��{Q��VKBЊ�E��1���sY��cj{��2��@�su���Ȗ��T�@G eޏ�[�9�;�K��"�+2 #���;-��!(&�F�'�+,T�`��p�67�d�{0������!�� ��`��Y����g�s�c�NE5a?"�+��Tc�+VT�C�+dn�.{�={� ��IO�<>��/���|��z�)�(֤�u���G8��{q���*J���snbs��<Ͻq�6�Z] �Ug|��Hڃ�r�F�@��2F �|��	~T55���.���gIE4P#]�|��b�;�l� ��A��wi�&�lW�n9/�@5��>ܮ���x���'��e {�`s��{�a��]-o�� c�0�&��$����l���1x 5ٖ*6�LmT<�<}M�{��<�x -K8�B�B��X ��;�n~
�=� 6�v�#��F��7��~>.��E��h��BS��@d�����Wu�cr�MfQ��.�(����	�1����r�a�����B5s&�଀w��a���h�XJW�6���5Ҕ���6e4d&"q����LL�J7���_sҸ�/	e�4+�mTt(��kF�	?KK�� �s��@��c��x��"�?����#�z~�1�d�������/t��H㛱�����D�n>yG݌3V�J9� �HB����n�������˃�XP�����hgR�P���v���X.X@�� ���KJ�x��
e�v'c����Y x��v;t���Bj���e�r�:���IMCRw=8��!C��޿٦3���yg{}s���'���*��C���9%X(c�;8�q��}c	���{��y#ؠ��i�u\����6�;:>�#����O?���MҜ�������7�V� �ٟ��-�-膣 z[Z�ʖ���~�� � N�1:m��nx*di�"�J���Y���XL��t f��5���˫�/XS���v[Sƥ9ۘ_P������|��/�o�	��s6[�ߟ�x!��� >�$@�)W9L^̗��6R�8���Q[3�A��1ߧ~�u���z������5�B�Ǆ�pz�5E���:�7��QC��K��ME�	}\D1!��^0a�{a����^�C�U�!�v:Utx�U��o��N�"��`M�f� ��d2	�����l��v5�*D�D-�G�� 6�Z���F# ѢDw��vK|�*�W=~f�"5
�L�-"R�+U�(׸&���5g��,�ʌN��bJ�6�N��1M��zѠ�شR,��?��s��(6�M\z�9���d^�r�(v$����x�|�y  *gv�]`�o�y��F�k����,f�h@�1�-М <�S�R灊唚ْE��zԼ�� �㫙8]sh.��`?n���R�Z��%�C���.�l��}!c���AX�?���Z��y�=*F��-�8�X#���[@���
ǥ�x8o�7�7�5?��А��t���toH}_\\1 ����+������ￗ���rrtC*O�ͽ=���W>\<�Q�P�e� >�f� P��і���w�.�S�9�l�@�e�TQ�R�[I=aD����`C��~��WZ����R�!b�<����lGMGh��5x������|��?����0(�>�l��{`+[���[+���k�b�0HW�W�4�Sr�Lt�ʂ$���J��q�k�)���������U�ѩ��6vX�h,��9��P�׀��d@��닷a�/�ၜ'&&"�� lNp~(�W)�^�0N*�P{MK�La�F��GR=�,�mL�������������|i���{%�̜a��
t&���H�J��&�&_�m�q�e��Q	��L$$*�s����ٓ I=A�
E���E}�a>D����֤i��C�P5���|3���oy�)��s����3?������Q@'
>X����&��Hޢt��m��"~Z���q��AD�[ �~DtA�9?�`Ԋhp���S�y2�*�(|/lb��	��DN�S����;\� 4k.Ʋ�
�����,HׇsG�\D���X�[�"�޶�Z���̈́#�b@���h����-q|t6����_C�c I C�zh�����`0�������gX�Q9�g88��k�X���r�58�ё�E~���;�j��jK�y��셍|]}�@�?�rl6U��A+l�prq�'?�$�ʄ��యM��έ
��| 5���޵�7}ݻ"%����j8�+H�� �#�����ؾJ�0tJWY�����{���C��/��/�| o�ˏ?<����ʟ��Y/��8??�"Փ�p��p?&���<��r�_��,DP?�:#� ��j�_�����|�L�c��fo�%��eF�Gn��t����E v��>On��(�Q�l��p=�ͨ"��~Oy�؎B�_�{p^�i�0y� ̾���g�7F�jZ E7S�/d�+Ѡ��Җ0���t0��T�X���z�A�`��������!�Y� �7�S�B��HϬ�S,����4�,ȧc�� �q�1M�d��}�[�O�񣚹G �����	��K���g��)M��=#�zM챤f�u�3�Wu()�k�Ze�y��38����
�u���g��]�k�J^aXlY]�&�=�ad�V����ܐ���3����?�蠖�� �3Sl���~T��3�ўw�Ȕy���{V����)��]�]�Ȩ����y�
6=��O�x]{�;�lj���1___&'��`Ϸ�[�N-3�}m	��x��l����'� ��ư�]�H��P�V[!O���
����Оf���-&�����؅oy5264�;_�{A��k@�(��b��Ӱ>H�/�u��:�B�4�J�T����u�>c˚�)�����$,��#=�F����^I��F��77�k���f����F��v����O�	�[�l�`t#G'oe0�|�MA��c-���$�=СZ� M�;,P�M"��b�e���\��K�Q�4V������~���1$��s*忨�y�.��0�����������������������)j�zp-�5��J�W��j#�X߸��M���6��@]�iV3���1��,U䍶U�[�V�i1"�ȗq1�c�@:ˊ����(>8!W=Q��3�#O�-��bEZ�;hz���Y45�����������Q���:��,GT��Ũ�F�5��O��/���}�}Ӌ�_�HV��f�HMO<��ISF�n@�.�=mb�)W,���sN�G�H�O���s-ԧC�1(:hp�$�B>�E��5x����l��Q8���ky��m  �rxt$�s�6��_���M�s�٭�mљ%��ϵ5��u��s�yb��L�G��HVl�Gp8ҦL��=�������m���쪋ș�o[K�TР�L9�� �򍕖��eT�BA$6>�=bi(�r�D9��_Q=�Y�����1��\�z�%y��!Wa5(F�M���A=Fq1܄�1A�+�l/:�����ޞ�|����߿/���Wt����I�E�޽���!�^)x<z�Hvvvx- 8O�=c�x�gl���S��!��� 8>��S����ʝ;w�~x�	��o��}�����7�grC�v�r��0���W@�b�A�������5"o*_.֗!j��Yk��咶?}]?��ډWI��kAkJ3ό��'3;��Z�{��0�>R����u �tT	C�?�@�/c]�����j&��̎��E��g�ϔcU���>s�
:P��b�N�F��	7c�7���q���yYY���ħ�C��k�>�;Zg{`\����S�����wm��Ge
Nr�\�f�[�5P�2-��.���m����BW��.S������tZؕ�8�t>p�L�I�����M��A��J��c������"[D (�¢Yy(աv ��ʔjE��xȠCUX� )Fbs{�S�i�9�H`Q�MAq�v��vдI�#q.�&U�B�.:����OH���W�G=�\�~җ��?1:� 
�;pl�,�������d����`Oi��yƢ���f��a/A_�E֤���uH�Yh�7|�_<�ς�{��]��?�ؑ�oF�G��HiǿE��?�e����t���i�"��]g�k�8����#N�����u:��kGᾂ���2 Ȥ0ETք�9�̃�:I�t��y���l�$_�.>W������vƥ:�ڠz��M>9�џ� ��xq?��y�{�H̴br��[c���3���_��L(�eZ+�Y^*q��������#�_���m)���X|E��/�l�t�Z��~�W`> Ȉ��`s�yڠVk�vԉK����N޾z��7�������i�@a��D]x�x��IM�}��S�(<�,����:P��*��߼Liѭ�4JQf���	&�7.o�Jbbr*��)2䂶Z�r�6�ڲ�����4�q:g?�G�T���,���a��\������ظ#թ�Z"��N+G����w��}�zf^�*޲(�m�__K�l,Rc�Ox`>2�����=�{�b�<5b겭�L�a�C����.=�Ps���ɨ�c�_��*���a�Y �;����m�k����$8���Y[^afc6�n�W%2��(�'�1W)T6�,�tPO4C�T`��:�ZT���4���Z����ŋ�� "�7jbT�!�ο�Z�=fmF�d��.��Pr���7������e���� 宽�)D\P�>5��k�aL�����X#���˷���5���W�a��	�Q���]�`]˵�980��F�@9�*�|7�&�c ����!�б2�:��ɯ(���8��@������� `$� �`/|':��Wpܕ<m���y�X��AG�^ ��]r}}��N���G�-�p��m 7C6{Df��^��Ɠ�-z[��֦����P���{a�B��Z�I��s�)�S��~Qm���L��V��u��k�9�l�m��P�����{���LO�{~�-¯kDM�F�b��7L�&#!��HU@c�D熙s�s�mQ�x��@��p���١WN �Me[�X�TЭ\���e��&Z�X��#�Od���S��R�+��������3:�U^;@U��>�8z3�X��gJQQm\������@�sf{qe��ܚ�j@��I�6_1�U�'�J�Ї�5؅Cyӿ�s�~]�P<�Ҳ�m��D�f���d��9�����U(:���v�]4��Ǜ�>�w����]��
�/wJ�}Y��)�` ��Z�p	QASX!���;�q�d��^p��w�ԃ�^��}�c���֪�5!uYr�Lh�����w�R�r���Aȥ�v��pQwe�(���<3���D�����e{s� j~1���$\�
�w�T\�%{�ӌ3�LI�����
9\Y�~�@CDńr0g����&l@Q��D%�'J�½E�m�ƭC���[E���~��3���"p�M���䍨��@@Vӷ`c%��Kw��H��.����*���c�L�� Ŀ�Ϗ� ���Ϧ ��=������{��:�YA�"NQ�N]CO#��9=+U�s)E{*u�?>�v.�ɦ�]�<��G�k[�g"����[��>����;r�:�G ��jr&ٖ�[�P�_GM��R�����~J�vچ������R�8	8zp��Xd1j����5�dp�t����r��x�Ѷb��4yH�.ѨOθ����@��=��d�pr֤x�SWq�����g�4o9�� <>8�]�����)�Hkh~�-Gg����~���[t��o��Q>��?�k�R�3pd'� ����r���r�\W&u��@�s@N�]8�����s���a~/8�_�V ����څDX7��;��,�~�Ʀ�m���K��y���M-�P�����phQ��H�*���P��-#��)��'�)����0�/<`� )���Jp�(�`�w8� �/;o(�7]��@�T��R	���)k1�`0�j�TT'#�P�o�&�^�򴽵�m+c�t6�fhX��Wx B`H�� 8���e����:ܣuU�"��u����q���)�A�<��:�������p��|�� �qrrB[���/�_�!cg�
�c�qC� �>���g������ۍp��mڷ�B�2*�8R2U
3�)@@"ϸo�8Q�uR�lLg:k�����y��)t�:��l 0���hV�����lx&F�*�V�i}>@墲�E���@�`-��'��2�f�rU�U�UAH�j~5��E��}�9LhCb�M-*�u�V\�L���{H�U��=���ldT�
� �,���)%W�@�2�T�[u͊E剱�ȴ����<>x��E�ծ�"U���2b�F���j�*�1˛�-�Ӭ&&vN��ʢ��5p�K��Rx%��{*�'����戳���2�Q����5��af�ͪ%���҂i�Z��g<�ql)�M*Q$���
��H���RA�T�e��rm �hl#���6��AV��\��V�����'�jksc�SL;vNǽ��ա�H+��r��g�u~~v,����<�2��6��53@���xZ�o�������7t�p͐��rᰍ ~׽m�i2�)|��:��Y�!���_
�����|��`������,�.cY�zV}0�"ִ�6-H� ���H��-���=
�Tf�m�>G��<�F��	��jβ�zͨ���)�1Bry8$u�]�'y"��F �H�0���W�~4�x�])�����W����z,�4#��w�5�vm�qk|�_�P���s_���]\r��y{(��+�߆C�We��v5h�ѥQ?Yϣ��^#^
�J)Q���ИP6#���# ڠ�����.Q\a.�e����C�g'ǇO��>v��2��R^0�y�.�wU�.c$E��牛�(?���Gn#*����e��pҠ| Ry��]�k*Cm�hW��ΤN����� ��Gf�!�4���r����*����uiT�t��}���Ԛz_�o{$?�O,ʽ�oQ*}�7�i}��㒒�`?sR�,ʙ�ķ�k@H#�CZI@�0p�+co���s�]��A_�$s](�T�;�	N�q�[rq~N��'K���� ���_���I����9����w��	#��2:�'�q�	s�������/r�//,�Q��P��,��Sy���<a�͂���Z͉5�TI[l�x S .q�R� �p��+������:&)'���.C�M�D[V-�&P�{;��(\S�����$c��,�����ܠ�e���� �.�� @T=7���U8.
Ǐ������)�6
vu�(b����Z�v��كF�c��
JV�� @\^bft+г�~��������Bpee��r���u���^Aa=<<�gO��I � &O�<a3Jd@����_�ѣ/euuCnz}�|����� ,aV	<�錍���H��Z�ȗ�U�n�/�>\\�������N�Fړ��},l��)g=�4�SІ]��Ң�-~�����R�E֢q���T���o�O��z�n(fyn_�?�<3�)�0�G�T���d�Q���ޒ5�F�Ԗ�g?)gN��f�ѩ4S�>�ǈ ��4�u���Nc�� �Vf�th� O�t����:e������7lv]c�c�ĲdZ4�AOũ
ʏ�w8�T>�����Լ(��A����cVM@ǫ��ff�	$t���i�}Z��[Z��4�1�݂�"3SAg�zwL�0��ix���y^e
pFq�V ˔�Ǻ��&z-����|X��E$�����k��k��hua���dr%�K�X�v����X_`-�$�����Y��XXC�`#����!��\�'��8��Vkޢ�����=�3�Ha�����!�sqy�@
�,�����,�h����oS<g~q��Q����R��:���M�[m�mAE�Xsq�O��2^;�k�l����`+�J��&�LZ��2�>���K�e���d1e� �J 2% J0�@X6�lb�AD�T��Y�תh\��K�L�JmH�tM�u�kc:b\�����Nˣ�O8�_D�ޫ$oN�3�>��n���@L������m6�W<Z-m��1� F<��:cU�f���Q�n�#G5���H�t�3�����www��tUR.�I|,]]�=��<{2�]�NY��R��>����策�b�"Q-:*��^���V�K,Rt�~����|��&ۘH������i�����#UD��jd�ej\#W9&��53B�.��h0�cAD������G9�����@��P�ⴚ�:��c~ԣ9��/���-���,2lMn*�Q���9M/�i^r}U���*?|�EN#�w�|�@�B#ya��Z`�ğ�	�T���}-�֮��ઊC��R+
-h>bÛE�~��'�$g��ġv��6��h���8���FpX;�n�-mס����dcm=ll4�4bSY`?�9n�X/�^�?E���� ĂI*[����&�_n���Ņ���������2"�Y2b-����|�}(�fu:,���Y�ѕ(Pa��[Y]Vഌ:�*!�Eʟ(�������2k>P�r> 
�b�͍5�7����U������^{p��>�A $gg�2���"�(}sxȈ���K^�?�(�p�w��`j>����9�����'h��ia��W�_��C35�
d��0�f�qA`�,\ �m̺t8Y�ˠ?�3���+��CRBh��H#�������ǿ~sh6&We��VP����gz�kRvg�~-�[���mV�1;`W����G4��:��s+��Hoe��9����g�����ѹ޲�m~��k__[�g����G�um�fG ��+2�X9e�;b�\ܘ+s����U�(F'Yd��D�$d̽O��;>�e2"p@@��e�Ţ�bMd��XWiǪ<��,�u�.c}�����sH�J?���ݜ��̂�Q,��3�)��[ک�۸0'Uk�6E�:�לPovT�ǎK��f{q��Ґ���`��݁�xb��@�� ��f6���ꄃA%CD��ؠ��Qﬢ�4�re)��������UC�p- �E� ��^�� y���\��W:�l�O����!�l^��Gh�#;��r��E��s���,+L p\���,@l��YS�JU:��}�)� �>������C�����үA�umȂ!P��\��,������6
��sxNT�2�]R]]>���Du2������ ��YS#�m�n,}n��pV1��ߑ���Hv����e=�r[�8�:����a�,,t�ZZT�i�#�Pkl��[�B@�yF�D����ydR�@*-������`��t@@W��*Q�����ތ�<�^�mc�! R�m���;T`��jV �*`��K��^��vM"��(��x�yT=4K��H��%f3gen�7y\d���;�/*]�"P�1�`��v)T�QePy��_�{����~�v�����߇!��8i���4�*�UE(7ǽJ(\lx�H���c�����$���HO@�̢�t�����Q���~x�K%�ZB��0�+��D P�����*u�t=%�9�ޥ���P�������1���4_}����7k$�( N�|��>���LF�� ������}�B�)i�����ٵy+��[��ʴ[na�r>rdE��Ӗ��5Հ�=G�9�S�z�+>:<"��N<�#�⻶678jX�77�8�ˤ��v�h��sѿ��u��(�љeC��eUYD(c&����p��(�)`��?m+�g�(��4.)���ݡ���@L�j$��+'�{ӿg����!���R긻�k�J�h�c�R�t �q#+���9�T�fY� �2f?z40�}���((�D:�)68��޼���~���3�hZ�(A6� )Z�9hl�
"ʊ�Ə�k�~�_hJ��w��&	zM��y6��>�<<!�����h{ @�p]�4�>� ��qOp��~�RB���\�ju~~)?��"̟��Y
�+��˱�GE��E3�9k"��a�i�7`�*��1D��4��l�E���@|���[D>v�V��0�c��~kg#��9�ERt�������C���k�ͫ
Q��m �>�H���3���.���>R���<��f;����X���:�b��q�B"��d�2���!4���� rV;^�9hxτ,,j���U}_D����0�5����L2����}ĞX�}"�,�t��J�\j�J��6�L��:�2����eQ|aj6F]s:%��J����r0a�'��E�P	��8�5V�����9��;�I@$5DU��(6~���[��N�p|t�fơTP{�i_$�,R(�+�F���W�	NZ�t����Kd��6}=Veog]��1V�3�>-���r��l���j � ��4x-'*+
{wt��Y.g��z-������`�����ƭ���w���<���-988�ŕ%�S;��
Z�ؐ�`�:�y9>�d�����9;���>}�{yq��:kʟ�UY��T��@��Ȳ�¦P�M>�O'��A��d�:���p�z��_�L2z�YĄ��Xۄ�(4�,T��,�*�s*��ւ���!��p8Ќ|A�VP��X�R�\��������kDq�It����x����Z��f7�^�=��}���Drk���Vh&7�0S�Bv�6�ʹ�g���.���	�Ff�Ef�����5ͲT��[�պ$z_�M�(GV�{$�)�*���ǡ�C��9m��fhW��/nǃ�\�E����%�I� ��6��f$^r��%*�9�Q�//.��׿����x��5S�]Fi�����m[?���~
����7D�����"�J_��ک7�6SS�Ӵ�adܤ�P�&�Nԑ1usKW�9�s�������<�&�;��'����m���}�w����]_�f������'3���Ht���IMq��i6_���{��h}:_5re�ͫ(Cgs.��⹨��� 
 ���������e5lZt[ʓ�̂�����/�V@��u��!D�z��^ñ�i�@�~31�|>�B:�I��9�� ^�Bӫׯ�)��S���!��$��PG���c��'V���A3M|
��>D���&����ٓ�t�О��*U�@�΋�6��9 D`���RǦ�Bve݂3�@!(� F9� �z�?k����?������J�� o߾e��O����oؓ`io��ɧ�:8��<ܽ˚�8<���/���rrz"�x��Ռ�~(x �`��+/{Ψ���"��X��P���8q38
 *�����p�=uT�
�p�Qs�jijN��̀�>
��cv��a�k0Ĺ�9F�⺙�E1Ոs4\�4�$Wp��Ɓ�uƂ��2Q��w�?��p�	�:��xS�=�Fip*[*��"5�3�N
�كE��` }6�{Qx�ή���,�;V!ej�?��G\�,�o+�a�x��(��JRj�j��6�4�몬`�0g������ ���z�l�:DV����9��ņ���v$�]��.{<}W�������WG��*�ɢ�F������
�4�Sz�w�`�(՞7�N��j�~�yD��V˴���_h��U� ���Ƹl��x�E���|��0�h4nzr�qrWu�
:@B7�QH�A��@yN��j��U��@p7��Ȫ�\�al����9??�d����Z��� ^�O?��\��pݠ����7J�z�(��su�c��Q��,/.�����}j��й�s�A��y�y���-��4&�I���!��(�m�[X6���!Wt<I��l�g��T�Z��䔍Bc��:�޴/���s`E� �^{s@ *h�I�ıkg��d�y�2�,�����s�gQ�VX�:�æ  �R�roþ�v���B�kp�X7���5�,׍h�ä�S6.8��5gh�)����e/���1�z��֌(5��)�,�Z<__��L0�k4�u9��N������h ��h�O��vډ
��2���@L���ө�����/��e�fJ��V����

�"֋l���:=���=S���M��xks�2�qC&7�݉�f ��Hn�i�x�E��Q�gϟ�o~�[��?�.��^T ����hx̲"(��F�����=�0'������P�A���=�XlY*аp#u��(]Qj�'�R#=
�|�b�s�k���83�����В^� i,��i�0�z�B;իd��������wZ�0E�\�g�GdD�ǜ��_�4��%,�<��#�ԝ���Ο�BC<��a�\��*��cpttH�����b��K�����1Ff���\�����Љ�������}���n�`�IQ_K�����ܺ���"����#�6�+ ���1�	��_^@�M�������Ă茪7����`����`�R6A_9^��&l��\����B�`���ᘷ���͵�C3�͍M1�#���-��8 %��?���^�@a�>-(�3�b~d��`1�����9���`�u��Y�`3~����h�*M_~��<}��@Ը�0��� ���F iW���K� #�����*lz[����ns� t��Fԟ�� B����b.���Ӡb^�n�i�������9��%�¹�AE^3!R� .Bo���q�l��&)���LiES��Y`%��Z�ZX���fus(-JE�:9-�̅�O@_8�������<:�Rb*7��k*_�_N�e�R�͌�8+^���W୵�����vmV ��]�Go�g6�� l�"�J��D��c�hRo�u�&n��#ś��y����5��\W�����-Zv����U�ѱ����A5%�Ժ\��Y�hYS�����!c���TI��>� j�v�
��y�u���q�2WU>��U�Xci����LJ:6�tR%R����\1�D��i$���A�;:�� ����Ѿ=c+�3!�`k�v��賻ᖍ����\��V$��/��upp���Z�6+8�WW�yI'߇���.Z����#��qVT��\��R���6o-aݡ�fH��0`r3���~[6d�}, ;�c@����D^�z��z$�=<���ҾTz\�m\����Z{��2f2���|Ľ8���x4�g#-Z�Xث��U�+g�l�'���>�3ۡ�A��*�:�Sm2$�봹�)�ނ�:�[S�����6�IjY�����1��w���{�M.��FM3R�(?:�����H�M×�!.`�M ���w��wM����O��6��{"b�eb"(:Gb�o�:�I2�g<��"��F���>�����-�`�/��Tk��z�E���j�*m>��O�����ހ����O�����������ٻ���!���&���d�!DzUZ+�s��S�E�6�����+���Y~������Ӭ��YY���
utR^����o޼!M
���7ÓR�#�R>���\7N�������Sb��OD���马"����fzf5��w��cڦ�k�_f�smD	�q3�!J�T��=^V���΢	�����1]��Ȼ�;�h���M�-�W�%�ӡ|֒�r�E#�=����(���j��Q��SF�)X�� p��d��t���2��oDsD����/ұda1j��@��N�KN2���<k���O�%7|��t`"	sl����y��6I(v�ϸ�Y8�;f��<6����<�O
�nB'���{k�炌����Ń�@ �2����A�
�+�7A��N#��_�~���rx2"Χ�[�.L��w~^3'(����PbQ�v� 3WZ���?<<���� ppn �`�~����f�(nG1�_����f�{��T ( �Ĺ�^�� ��h0a�Q�2Oe����,��@�o/���	�X����XN��W�E8����| ;Z3�r�Y#ܕ���9���ݶ���Y�=6�P��ZȌH.h_�sP�SI��t@e�N�6�&�'�vw¼�>�o���_ذ�ء�j=�b@g �c���B��`e^�g�2~'\�/����?��ȦPJ��[͓R˦�(:�����"~b�0EBUޕ⢢$�X�Wp��Rr��V����\5���
~J+�䕚
�:z�1J���1���TƈMHgۢ�6e�&I��X�� ?[��S�~N3��D3�5E�T�����^���,�0ob�+�n;w�M�9W�c�{�FcQ����Fbc_j�D+7�B2TZ��uT.�RiU�D2���f�QW��DD���}|8|K7 ��N&+�������1u��|�J�/-����U�髫Kr��=9��g���}*�ẑ�}��=�54�+`w�b�@˓�Oh�..��*�k���AWsD�\����2`n��o
�D5�9�"�p޿�{3 �a����6 ���yU�[-P�
�b�������������s�]�J�D�YP*/����ϊ��`(�h7�����3�z䥊Z�Y ��^;��BpvI	f=�X)x���Jn|��da�ծ��L+�W�-�n��	,����T0�Q��E��}�W4���C�㖱�S�'���ǌ�&q[�]�߄J�x0$5{�h�T���i�qP������舁96������`O����{��2Y�����"QqO� M�:v�������4g�*�����Ch/fFc����f�0���[�؜�6�
J39[j�|���(���/�˟���h�<�0�0��Ј4 �e�:�8�#�gO��������`D���A��B������̜��@�-;�{�6�):���㖗k�9�o��E�	��	��Len9��R3�쪴IN�n�(���]�;����X5�!�GW��;|�&ʟ�[õr.����w�E�U�+�P��#]�N���L����@��|s���
����.��lC��)Ypl��������Ce�O�6�G�_����M�6�3oM��J-�e���	q��9�*���e�މ�� �������|q=�ŋ�@���oo�����E[ZT5ҁJu��;}r1���*/"���ǹ��ƌ"��e��$$�����F�"�0f��ܜ�/�d}u98�ox�>�s�[1�F���a��L%�0[N@wZ^Z��Bq���#-�fv"���dVN�O�;99��Э0� ����wzv�B`<*J�"۱G{r�x�lv�~��|���w@���
� �'�u�h��h�n���x�z"�Ё��j�I�R���j��Mo�����VG�g������#�2����hT�A7�T.Xn�S��ۉ����"�0���	@�䪜�s[1�(l��de�C�*���6���g�#ε�wyM�6��欥J)QZW�G���z�MQB�P�rPo���4 �N-9�먅:��
����0�����(s�M�}X��+r<XF@#����|�J���V�y���:ޑ^I1s̚��W��2���ȧv�mNL�I���q1@�>Uۊ�́4Y�q�\j��N�ޗ��"	�X��8`%7�����ݺ�!��J���O[��_��,>��}��SFk���F@�>��;0�9����P�2�S�0.r����P&���@�ۃ�������7���<}���p<x�������kc��?��o� ��͍u�?y�S��f˰�T�˨�����z(�a������B G�����p.��< �%ع��&�gN.�/	�����p5����ZJoÁ��ieޤ:��e��aa�~׷E ���C�b!TE#�S��FO,:���2[������Y���J�Y�iV� ��i1�Rv��'�C�Z���ө�Xᤔ{g�sT��[l�p6�63�� E_�Jk��m�p���uL_���;�fF���%�d�h��\+.+��!��ͲǬ��U�.<�XG�������{���9���d:�6+�Z��1y {��j�@^�x����޻wG��Ʀ�����vw��_���z8���)�����jGG)���I���@1)"�(c��2ե㤒��4*7����f0؈�"�chA}M��,:.|B�Q]�Yᠪ�d�����s.S��q��)E�j��x�?;Qf�U�$f>?�+>&��<��O���Z���� r��C����<�wN6���}p���n�S^����m��V �"7" �/M~�d�@�"u :6�L+O_��Ŋ�3�iw_v�9:�$�.*
�&�Q<��$��Օ��'TOiD ��N)1"�m��� �Y��np���d���v᤮P�qX���� ŉ�_d�v\&uE�ҩ@dT�Ѥ�z����3N�	��U��U��1ib�\�U�x�U�y�ZV�^���A#>�%��y���E�����$(G���N�:�+(k躎���G������e` ����j%�E�*�)YPʱ��g������t��W���(Q~"����F0	GF�'����Tp�/�j�p��H� ���}y�P;�?�y��L���:z��-�,t"�&pT����M��Y�/��*E��x�Wg��H2��ֳ���i�2o����_���u[E�w��
#vl��&?��p��yvE��  }6%���] 1\7:B� pu a�m1�ZI &�5�f!��nw��VD�B59�iA���21%���� `����K̢��ç��o(��p�	��,&�Ċ4�.�IԱ�~P�6<5��ݕE�9�F���L]4�'����GDj�R���!�*�2�s%�FTg_��Vo���S�u�yn&XA�R��<b�l<�۶Z�D�q��E�k��z\�QU)��x�eU�V���	�tz�gv��� 9��-����\ �bT�B���H��g�(r��e�b�md]WWda~N�����N)�H�[3�IDgل�Da�ח�iz����Cl#���ޞ��.������M����s�i��ƭ��o�����Bhu!������f�CY^Y$���Ж�p>k�\��,N�,��uN������B;��Qh��,"�|��Rs :H,3֑yր�/���&����g-g�Uؒ`o��f�Ɗ#�阚���k��e<�D\>�X�u��z��	*y]Z�C)Xe���^f���e�h�`�~3��O_�v���]̈́��O� �̾qF!R6�5m�̈I����X��cn�.͌���a=�T����a����h�Z��q9�n�Bum�$��)ځ1���1����I�'��h�[m�G���+���"������e����o`�d�"�]��.-^W�j�~����w��_|�YD]���˃��3�R a#��L�+�S���]�*�.�D��bS���;���n��Xx
GB{Ԏ�J���|���y ||��7�k&�ݠ��ePt��6��]��*����46��H|s�}j}�QO>�ܛ}�����M��پ�}�k��"-�^�E>j�B�O�O4ƠΛL/���%U�5�sѾ����0N)T4��ފ����L��X�Kc:� �e���")�$�j8��\�z �ð8�˲��!�WP��sn�Y�E��.�h��BH�A�Ѱ��k�./��aQ���sDa�o��*W��f��=����)2��m���U�@4{[@�pQ]apL�0������ڻ	��M^�Ne�:
(P��6�� �`R�$j|���y6��E&��aT�cG��P��켴0O����_?UclE7�+DM@��&S� NH�B��K��� %�����=�7�S��t��a�������楬��i�]sY� :삺{�@u*\"� "������}�˯�}���'z1����%{{�������ѻN�����ap��õ*:RPVc�Se,�"��1ar�-��Yj�=�\j���"��u�Y����8]�xp��X���>�­�lnc��E.б5R�]FYnd���z0��a�`�-�,��H,�=�L���dȬZxN�@U�u��R��5�L���Ry<��#љ5�5M��Ȩ%��
�5�.	xh!��/�	rzs��e�煩+UY���(�z�it�-z�s*��6z%�_Eʧ O�yP)E��(t�p<o2����٨`��	�)4�j0���P"f5`+Ť}c�BՉDA���D���T�� ��e��K6�"]����T��3��-�d7`;��J9��&(h*�v��� |����������b-�d�ɄS���,�+l&�|I{� ��ŉ6���/���e���]\JfDN�C���&� �z�
_ �;B 0񋯿f����~�O��Ç���[k�^�I��ka>�ȎN��ޖ����v�wV�W�7u�8՜dd�17Pk�t�Ԓ��n���&Z��PqS3;��Q�X��6mō�
��$ٔ���o֧9��]��]���lnm&��!�����M5��K��λ2J);)��������s��͆A{���!2E k����WU��uM�h��g^�޺���`Zl>��͇�٥h���"��_�MjU*.*��B���R񂍽	{7��*�\�X<Pf��|���o�W }���fp#��4�aC�4(�@p�s�贒����;�~��K���}����_�YXK-�O�������ރG�ۗa�ac״�R�b���.�K9�A�I:UuѢ�9v�dҙh��n���`p�=�9�]�\���� T	�i�̩�!۵��͊�L������ �ͫ�GiF��;V+�D]�w�I#��|}�;��OD�ׇ ͔��;|����^D�����uy���NbV?a�7ri�zLR�ĽsR���|���o�r�`wsk�N7�t�y���5�V)-���l���,�a�^�q~����dG�ț7/�;c�R�Zg�+_4�������� E�-�'T�ʣJ�N��o��7)�Q�E�4�f�%O����t98Ϡ`iGl]S��Q������
�)Л4���bD)o��D��J[�N��2鳳� ���b�np���a]�縹�gA�|��`bQX����Y���-�nG��'w�~�w�G;��dAQ���(�����ԕ��l��ƺ�9C 4^�{�����.��o����7o^q���y/��vM�*+�+���9ܘц� �]q���~��R+�a��?�9a�GN:���_}+�}���|y�oq����g<�2 �ࣥ���]*�`b�?ךc�����Qi�0K�4n=S(T�}l&x-��@�i�� �ls�Cu��Cm�������H�#����!����xe��
�¸"���4魭(q�p�{̤ {&Vt���g�����S���Ŝ�Ek���sS���������#}JY��ȷ(��Q�b��Q~�k�4M���e[�@@���J���Z��8s�Jw���2�?�71��d����Y����z�e�>��!l6D��1t.K��4PF	z�2�8�����/��3�+)��P��9!V��T��y��-�j|����"6��C����\��ޘ�`�We���� �R��TP��M��J�|Ŝ $P7fU'�G��Xs�C
�S��A��k��s��T%�/��./ӑ¹n���j�Wk[���?ҙ�-�sp@�����`S
���z�X����d} Hj
�_{�h�]��yY��]"�
�)�4(5B�u�g?�Wl<��b��`�ׄ��K���C3�����mE;���O�)��j]K���� �<�i6UE��d��|��.:�NP5C��fP��Й���Fr��1$�kc�*5%�Ź"P������H^?o�C�̵�[�R�� 4����f����G�B���5,md��Y�w���{4��Pj��x<�Viv�!�?��_�&̓�i߳�"Yûk�l��}/�\Q�5����. 	�UZ�J4���]B �C���}k*�X�c�L��T�������������˽]Y#Y{���Q0��++k�0�؄GԾo�nl���0J}űc�����4n*�p�6�M�l؈&��p�Q�$Q{�sC�#�:   S��n;iw7�)�g�s�G4(�L����ܜH�D����3���?3i���E�M0�k�|f��ь��gQu��	T{S/��1s���w(��TiA���ޤ���k{�#2h���e��xev���W�S06��F@����66���*U�S��D�/������ږ��-�Z�f���)��������i�����p���Z]S�u�9�]����]^�*�pZ��6̚����jb����)�'���"��n��G���'�{w���{�c��#�������¢sD����m	)���>ٔ?�qB3�������|��rp�<��oO��'����'����,6���f+�40l
8Ѭ��ѱ6[�Fv��G�`ԓ��ox�R���ux-�� ����������`�qwZ��2��	U����&l61d� �b��cm.�j2�߼&�
u;�9/���'�!���ׯ�ʯ����T��	��0̵y*v�]�ʳ�O�Mr��n����=�riE��@S+���w��&�g�EM���|�������܂o��RxVaGATx%�Ơ�܄�����ٗ�-~)tܟ��5�����	N?�5�d$���`�����Q�2ΙFеhIJ.i2r���&BW��xd��$�ͺ ��Ri�ATu��b�_z�Ĳ��EU֙����.e�������=���@����lat�%^;�_Fw����u�L�ծ�� jc歇@�p�ĨS���X1���+�V��� ,:n����ƥ�X1}�E�<�R�:"�!4�VF��|V�^����=;�Q�&��<%�+��e�3���*R)(�*u��:]\T�+p'ew��O�wE��0�}g���- S�H�����~h�v��"8��dߐ&4	��� |�4��ڶ��״8>@��j-^��-`)Ɠ�Э�������^�	�r}uI <�=�7t� z�v�Y�v'WY��o9Fv���5kAp��	��fqF�B(b���9Z�r�ѭь�5T� ��2 "Hs��#)��-�h�[H��u|_N�ѿ�'�8gE�Zg�B�EJˊ�k�e �O��Нɾ��
�5�Te�Em"����feYOy]GQt�/}��<K[8�?ݬ������c��&`��t�h�`�����A2���RuG}*'x�,�Ja�v�y�&�W �w7�D��e��:Ea����d��6��� �OFƀ�{���/�-h�,Tϕ������ҷeZ���)��TeS�;���/@g� 6دW1�d����4+��"x�04p`&�S����co��	����#B��U#�XȬ�@��<l���+j�
C0<eC�����z�*�gkY��=�(NoH5ӛ g���c�tޜ�C�3N��a�Oo�c�O�x��zc�7��!J�oC7ӇIQոi~ĵ���i o{4]]`/�*[N���\�8귐o�S�K����អ���7�KKDi!���7
��B���J��e=l@�<z6�}��(��I]�.(���fvtIn���c�M������zAj��ҙx�|����я���f� (�di-0�e�碝�[�n�8#kiZ�g��B&N�����C�;|",�^�׀}Bڲ��iF��Ey��JOn����ol�S-
kcqi-8��h�V���L�#<�d4r��K�k+� M�Oa#�������6a ���%��8��Q�
�oy���=�&IE�׊Ri3�K4�hH��#8ΰ%�}l�v�I�J�2�a�&��#̒X;��P6�8�J���Sfup���5�����d��+_>�
��)�Gw��c�H��cy��1��`|qLf�*�<u�ǈTui�XJ#�&d���"���;�I	_���&PNi5�u��W
�G}f�X����;�B1g<��J�>���{���~���  �����L/T���Gf�
J,�M
��6�\-�y,��[�3ډZF��,Q$�a�Ն#�"ݎf#j2h��#����^��n�x�j��:�����1��:����e�(TLȔ	��RL(�2�.9�*_��ٵi.v�J�ZN����ƴݘ#��@��pS�X�C��^D"Sͣ�XG丷f1x(��{e�fv~�	6X��E�s4�&k��*�*M����т(1ޚ㭁?���zT���e��s��b!�1�J�BV�4��ά�v���*��ɸlD�*��^��'(i�/`Q{8g��hz���Q��0���V�ޠ������	�?��^���3����T�z��AЍ�`ï4����&���y;�9���K�v�3�)l���>3��7����� @G ��j4�Ih?O��E�@�{p�LKz��@�,�|8f��M(��z��`��nA�ɨfE�W;�R�Z�g:?m-�C�\�;}��5��@�*�t����=�72�<Nz�9�� �Q 7� w۵�k�Q��-��7��;�WM�w����N=�G��@a�2_W�JRD�O��!���~��fms��"q)Ө=��5��%h��f?��<��7.�WУʌ�"<>��(������{�~WڨpG6��"nm�ȟ��y-d[TJ�w�~��w���_P4�6_FFQ<k�!�GM_HaZ��ĸ��fX�0�
|ԥ�\$�fQ8�;��<KV�c@�hN�w�q@gi`%����Ζ�%���6Ӱ,4�"�~wc��*ީ�������m����|��t^��=�񇸡��U5��45�E���DfS'6���C�~����Tz��&��]�.a.�������vxCu"̓8&�,��X�_�L՚ ?ڙ�!��7����o�G��@����l��')�?��ٱ��3�6?�&�4�� ���[��&�W�E�o������]`�v ���bЎ�*��ق̫lb�������E���.�鱜���舼st�n��p��f ��8�ݽ}9�8��B���¢ܹs 됎<�g=���:{� z��ep�Ǡ�#��H�s��޷i� _�$��?��5/^<�2`�Dѝ�c��Ӂ��	� '�n��ұ�)]�uձ`C��һ���pZ�R9̭6�%������t�ƃ�\�$�"'3���Dp�QqoaA����}(�|&G��܄>
���n�fp_dY�Wo0�'v:?9bTэ�54�ޕ#��4�/�d2Չ��%fF�4�C=Q�w M�����&�2�c휌�����DMdG1O!4pyQ�>.��gg���Sޏ������w��Mb���}(0D�����d����B��	�x��]
~}�r��R3�v��V <��� S�5톣iE��\���w��F
B��uq�3m��]������-���T�xn��v��Ѡk���(U�Z6�F.�ABmN���2d���ΧmA|z�J��}��J{c���vo{�&�9��M��N��u{�;�n��qR��ڵ%T/"eGxnbJ9����po�T�DmF Dn��_	״�� a�nom�Y_����T�MT�w�pam�\ =�i�a-��Z��a]@����LȄ"u�m�\y��	�4�W���@����>c"++k�
������*dh�_��	��� Q\:��:@�qO˙���d�&�*� �GP�#Tьr�"̥`2��ՙN��T2Xu)�FTm��
����G����V ��-�����Rj����(�.q��<9�q-׮�g'f�����p>�I�d�`�']�c�k\W�FQ)r�A=�R�W����'�RD��O�����i/�O�8�����CU���i_�K�����!��Ʀ�^^s�<�����'j�nN�XF��H�6띣O=A�W}�&����R��x��yў�$�  �\�fO�1�3�p�Yu��A�q�PÉ��0�������vuu�HY�È0#UB���l���'jIDry'������V�m-I�� �IoܨVԑ�BVu0ǔ�����Po�����+6L*
�F�P|YID�GC.�n�E1�o�U��ܳ�����εx������<{�B�-��E������p����g@O<��������s�$�t�Eg�9��Y���#!���vC��i�]k��2cQ�y���ѹ|W��Z�˫���W���=��g2���lm��C� ��.���N�{xrL`M�X�ܸ��IUR��Dv$lX��ޠ�+s�ql���F��88��=�OX��da�0*7�ڑ�G� ň�"���fP� *�$� pwg�JQ7a�x��53&��k��O��2N������� z}}Kv���f�6�	�p\l��1!
҅A�ʜ�r��`샃=�g���_��_�Vtp�|��?Jg0�j��ɩ\0E���m�1t3Ǟ��c�L���,/�`u�S
F�2�$w�FW� @Ѡi�q�d�����nQԢ��0�C�'��uc?(��05=s�#<0�:�yF^�~��1��ǧ�/�|��� ��Y����.탍��\�K��FJ1����JtZ�LQ~�"�I\"Q��+(�-�����'X
*jhH��qK�p��&��@�(� X� z�]�v@ų/_���s���#��Pm�� 
�3px��΂�X��α�*��m= �I؈�(E��l,LT;͎�Ȧ��cG��D�@�Y�:��M�#���)t�5�$�l��َ���,�M��#���e�c���po�5�C�����U��$�x:��)�2Δ��0e���r�%��?\OQ��خu,b��[V���*DV�_�V�j�}����(���N���&��u/WvB}O��j=b�k���W}}WΚ������4b��N7 d�
:��Gg�%;�+r��%�ۛa]�X��Qqm���#=)u}�;���*؛sJ���t����|��y��pN8?�RP��9*���?1Ӏ�:�/�" ��=<d���Cq�	H1#�,G;؎�ਂ*
��r�G�{��^f����Z8�+u4�m����`S�0` �}|t�M�p�&lއ����-{`]����̍�@���M�4���lez+cE�w���\�����`W{�	k�DI��h��n���4@k�A6��������%�V>�ڨ�k殝h�kk���߮űF�����[�j�~����j����HGf�܍5�q^^��8��G���t�a�u��ph��@�k��~\2;
)��XG#Z�:(�Dp_�g�7m�f��T�pdI�N��Y�����4(�Fе�Ȇ�vF)�cPqw�w@��:1������p��D�sy
|��_�x�?����cؘ3Hob�@/��'#�VL¬�X�G���-arll�*�*��ə��9XU����p0X�d�־w����0��`f@l��&\+#�iܗ*����#��Ґ.�������y��C��m�3LG�7�=���nD�|dS�6er��-�r��,���{���ؤ,����mu�W�l|�n�MV�U �(���lF�[�&e��,*�f���Ip@���ɓ�O��u�� H?������|��C���
�ƇM�]bcB��pB�.>R���Si=5X�5��� �X��$
�������Q����p�x�Z��ـ-��,ln(D�2
6��+ҥ@���/���_}�����)-�T\�OY�l&�$|���Z� J��hoo�1 6O8@��J�Y*d2hXN)E��ѽ�����o��l��~�b���� ��	��F�&"(ء�9�E�c�5�LS��2 PT��ly)�k{A��f¨R��(������<��H�6�� z� p�2ߘK+��W!ԧ��9�
�>��Vf�[��^ʫoy?�t���U�, �a�y��_�/���Y���SY[ݐ�i]���K��RC5��3��$��J�Tƹ�p�.����Y�uq6Y>�9��|wA��KTl�Lz���>�e�(�ṟ�����~��{�`��lms?��9~{��[-.7yVd��k�k�9Vq ������!���@��2h����~x9&)�vw���*���z�Jmr�R#���s�<���Q�F�]�ﮣ��k5�
)`_ m����5ޫΐ䤔��iH=J�v����֐(H)S�D�oj@?�OHǲ0�2�ZK"i�}����J}V��h��<f��������X�J���XV�hf��� ���C̞Q���Z/ ���'I�g\#˝ �:�թ�IYbs:|]1�7����cu��_	>�V�#��Mտ~���7�X��tY�C�FפG^]���@����Oڛ(ɕW���Z;����lRE齙����l��}�3��h4E����n �P��{�/�q���	��L�,V�2�.q#<��?�����W_2�<jP� ������{��c,�ǌ�^A���t���X���?p} HJ@ǫ7o��?�}B	N�ڂ6z G��2���x��m��P� ��	Ȑ�_-"�=��BfT`P_��XQ^��T��+����%X�c��-k��.1��D0?B�<��,��ӷ�T�� �f�W	�]k8�϶��j*�|��L�@J�XZ)�g�kG<��< }F�Y��|CT
h�z����Q�x3����e$�OgG$��6}���=o,}��q��g�c���:���|��GPl&�t�3P�z��� �Z�QqYZ��5��͎�����۞�sڠٖ;�u�e*"ZZ�)��1�q�����7������x~Aө^��'��n�n������ͧӓ��A5��9���Bow+k��ҧ�,��uQ�B��t��1��fP��Z��v�D帥����qrF��E��g���c{��*W���s���Ȏ!jP3�� ��lq��se�6�s�|{��{����6�����(�c���*�Ҹ�/w����Y����7T��� G%x*�x���"2�)�JO!3S2S]jUh��Q����=z�ie�-2mr^eS
��*مJ��'ws��o�����G=�zԳ���ُDÊ�R�0f�i<O�"�h����F��E��@zr�6�I���GGʔ=pҼ�J�:y}"߿��u)=(K%�L�d=_�����g�( z�'�}����r(oN^�r����$'��ٗ�R�;;y��9Ϧ� N%��^m4Ea�
lp��O��Ζt@��.
�5Ӊ(ʊ�?b��X2+kF�1H�t�'��8�����{�*m���b�v�Iٛ�d�˗_�	�CQ�xt����"�߀����YY]G�4�I��t�����ȡ�
2O
&��څ93U�EJ���aJ�:��"�n�g�vL��;�kx�(�Da�l��슠o�.��r���Q��1�˟�����7�S�4������N�=}"�����Qn��d�X����b*�P̑Js��er0&�o/���x�&�����"�a<����>/��$��B^�	��46am���&�^��I�*�l!��񳏸�X� ���E_U3�	��y[�x��e�� 䤋��繰:�>�����=ұZ���P+b��r�� �ٶ̘m
��?1!�t'�TӁO]�P 0��b��*úFD	Q-.��2�ޓ �]v�X�y#�+*�R������~�h��{v����k�)�Ĳ�Jg��}���هJ�Cf��=�bI��5O
TΔH�[�-f�C��@w�c�V7�t�ͺϊ���o��Lm� ��e�g�fP��kc �M�}8?i��8f5�`/Y ��2X�K�?N��i����Ҵ��l�{�K��9K��u����ɂ�Ȗ�Yt���G֯�F��<~tL[�� ꖽ9VV_:�Cu�l;��B���DN��6��v5��Ҏ�&��h?�iI`Cآ����Y�զ��kt���4�G	X ,"�Lelg�^#���c��>z��vM�J�+��ި�R?u65G�H����I��Xu[�e>���N�I�������=9�o��v_��,(n�>���?�v˂e�h��`Jl��%1�be2s!����`�^�R���  [�bFS������_G�ml8g��ֲ�y����������6_���6!������e]�F�6`�X@�Z�*��mG�*|��#{��8�i�H�1�(�AIz�A��@J��[�[��Kx~X�)�a��f�@�J;��(ju=R(Qc
?|?�$l�lk����?�ǻ�x�x@~�o]%qc�T��7���(��h
�#J��T�O��G�S�D��t_�3劲p0�Hˣ�j���`>J�]�Eqq��qo.���)Q���N򄫌�c\L��ߗ؜T>���������Ma���_<��C_w�B�|����� �%�^L�\ћ���O�y=v�ʹ�V��i��9%��%'EoԮ�F���-x�cN�CF��:^!��Y��4�H�,�{�m1O�׿��g��y��>I�=F�ٝ����> X��7/x�L����v¦y�+Ǻ'w�SF�+F1�S�^P+���&vu����Y�`���_���9��A1�#6B<;��q��ǂ�'����3yt������Nr�gT�N��x�bn��E��7�_Ѡ=���w��z'��/���E�;ܬ^/N���������?SU�lD{�62_-�嫗���gr7Y�������^iF$�q�V�����9e4do�F���\쏞=I����,��S� ��W?z�������0�q��=��s?�����"ڏ����4��*�A��Y�;��O2z�}��e#������M����P+����aP�V�g��i�(m�H5#Fg�5P����X�꣧�pc���ɿ������'td@m�N�r�N�}�){���[?yIЩ5�^`"8���K���ҵN!��.�AX���D�	6b�<p�hx�fh�젫r?�%i��3@�0�Nv>O�m|��������~���#
`�4x����~�*P�@m\�gH2��M�e�to���uOvҳ�Z�w�7���ƶ��m��2�9�D�P�g�x���t�h	a�!5p�A�BQ|���J�q��������>�uTz`c� ���r�!�E��NL
��Ղ6oC��]���1�ܴY� ������z����S���W�A�-"�`�o��T�"��n<�Bx��w�J�[H]����!_���Z�[͜���z}~������^�j+��K���z1I�49C��tk4���x��P��R d��b�T��;6���|��Iz��5J � ��{��9�X���}{Ȍ
����o�:*\+�""t�p���,�����)�^3�� ձ�lEZS�
2���,���'�C�z�����ӱ�M��� �9�C�>�H�e��(���^��:�|�;�yq,ٻ�DZzJ�R������@��q�E�۶9ڵN*��)_ ������lH��Gc�4��h�m�!)�ϥ�M T�>g"H�{U�׃-�2�~��v0�:}W�i�����V�(�\���>Ĝ�	Ev�������h������~P4�dy��,G�Z!�K[p`��y@dd�� 8������
�Ҳɲh&��S,q���X $ ��� Hk�Wڨk`{(|����j����+Ɗ�L ţ�{���5��l.^�C:��|zz;����_�\�#��`rrP]�tt�>�*w:Z�&|i��A�rP2��1Z��<����$v�j̭9� ��
6lDu�P���̔�΋�Ep0�0��ܱC���hȨDk��X}�{�|x���e�	�1>0+�?[&/�X*A��y��t�eB(�%7�w�/k���76������<���&ټ�|:�Z�HYDFS���v?P��!(�Al"+Bw�4̝��}����Xj����H�v�gߎ�߾M���������s5�HG���]v̬eBӚ �
�,D�A�"�z�s���!3��gg��.��G�C���B� g1Ş����4�_��Ŕ��F�;��{�������_�����ͫ���VF��:������-¯���}FzZ�~�@r��7o�HA@ư�V7s�(Q�^]-�׿���������+m��	=�J�^���`d��*m���v]�?�^��g�$}�N�p\�Ӎ��pԣ��R<+f�(>&Pw��86���� ��V�;����Ŕ�����Y����t/����O�����M�� �R�&3��	iLch���Z���)���bVZ�]:�:9�s���嗿 ��L4������G y�!V^��ڈ������y�^{;��cs����e�ft����f���=�hy���cR�07��<6��;1:u��"V� zAD&!aS����=����'����^z�����  Su��X&i�]��r�Aa�qK˜}��$T���e�Ҷ�G�N��bF�>��P8�$���6��l�<ޡ��x��
�!�0�P����u�L-*6�m���^,��JWe��WU�)L���nM4ʇթ��/��֒;H��h�ȣ�Z{�E*��@�c��, ��Q��P�%��yT)���"o�(G�h�n�.�NG�K;8�(�M�\�J�s�ϩ Ȓ�r�^���XN���<H���y}��F�z.CD��dm2�� �8�c��� F��I�!�ǽ�}*Q�^��H����3
K ˇ��_����ŧ��� ���ޑ����1� ���:I6u �����2�X�k:x 7s֬]s��=>�L`_ �!��ܫ��7>y�Xv�/e5{#��;�C�]~t|(��:��	�{��ЀrŞVsQ>�F��{0<��V�2Y6 ����P�f��p�(6�o��J{��ɩ6vEC�䰢��o`��>�W2���
Mu)X��
߶��?�N��Z�(��Z����Z@�5D�Z0(k��������E �cil�u��-�u7����_�3u���J������/�X<ka���qf44G��!3�,l����p�>9�M�� ̬�n��`��4��=�u�;4��X4 � |�V
R����m�Hr��uD,0�z���̚�o���'�}��������o�h�}Ӆ0�=�o�3ڝ�e���͞t!�^�fO�ю�S�Bč�Kk�4�x<�z �q?D=�H�JS��.;i��jw(����O&'�4�I�gJ��������ۏ��d�wT���-��&2ϟ�<K�����>n�׎�a����A���?�������-�SNv1����G6X�Cl尌Ѵ��KاB d��$�]4	�0�5o����i����77r��Rv��soiX0 $�A`� �=O�x�h����+.RQiB�w4���?潠���-�Z�2��bmD*�v�j=p�Ɍ��;�e�PjQ��ԃ�T��z}�29�����wjH_Ԟ$�"D�
���r��I�$$Q�� �
c�ڪ��j����r͌�mr�[t�m��E�C�;:ڷ�����n:W���³���CէS
���y_*��A}:d} ��g�[J���Yȍ�v�l���.�3�"E��F�w�@���q2������bpDI!A5���@�������t�Z;a#R�Z�pn�����h/9!M�ǙD�_�2�. <�� @�:�G��ˢ���=�Y�����	7��:����ܼS�4&�k�6���=j^�U~��3*�Q��
Y�ێ�ce�Np�071瑹c��4��������=���oӹ�����O?��~�|��׼���礢`�g3\�>�f�u��q,�H6D�o.��c�C�J�%R�ǹ�=��ku1[��.9Ő�FJɺ�rI�n^ZD^�.�J	ّ����u��X�?� ��մ�N�=�@��
F���4ᶋ���K�f,�|�ҍpŘ��Ŭ68�� �z���������_�R��]�XѾ̋�����s<ԨsE�67Z�!�� HZ��r�����rسH�p�=�u>*_�X����׿#[�T�V���������G��O�ʳ����=�Ϳ�J���n �ю1����_���6s
����#;�����3V���5t���''<7(�;�x��H ���4���	{����}p���/SE�]�9��ؗfi^C�MQA�C��G�s�!�ZWꐡ�mz}C	�G��GO��^w3R�P�r{{E�Ԯ�&�u�ϩ��R����Wڙ������b{��8G��D�E�Ӥ-�_[kRY�5���Y�{F0�{�� XG��U*7n-K�C�#�e�u
_�N��?a�RzP`��5'o޼M{vd֞2� ɤqټ� �8���|�|���Qzl$ƍ���;��?��>T��Vi�J���b��@�nYW��z�N�yM\$�'����CVC����h�bN0,.�	CA;$zC_�,P�m*���l% S�GP=�X4���H�י݄/` �	d!O޾���˗/���	>��O���||��x��t8.�7��Ȯ��g�-�H"bk�Α��^iGd0�f��T���VN�Fj5�M�f���v\���^�)C@�ݬ�s,�[xşH��K7|EG�
uV?���`�I�Br�7&������q����{~����7�H�!qI=�|m��v��]"
x�Q�2:`Q�wҙ~��^�6ͭ�������V�b�����z�.GPl@�ۖ£9t8\&K5��r9*�7�E�29y��wƔv�L<R9JT/m|k���eTx�? �Di*�������g_���P�?���	��aq?x0��b�Ti/m|#�D�y��:�<)����5�O��]��_<O`d�*m��☡`�{{w�ByfA����s��+���tZ��A^�����9{#(��3v ݺ�dX�/Z_�@O�%�|P2xu+q��c!_�;K��Y�zP� �T����	798���>�zۼe���@5�I�agt?�þ�&S�pX��A�cJ0Vɜ�\��u:4���Ef�i�t��}د�дo�B*2NNʐ��b:��Zr�Aq�j�@�@�y�斀�;ՐI�q(���}����x	�m�5����I0��:]3��p�)����h��BO��b��¹B k����t�˫k��뫛,rvz�5��FF���]<����wx�����ޮ��p����ξ�K����T���Ь��(� �ɍ6��VZ��i�0m�ȵ��T{����*�c����L���ah�����lKSڬ�My֢�M�5�JD]gI�Z��˭l�X:�n�=�#��ux�HC��M\$��h�R�<n-K��Ѯ��O����)����@Fb�[��E?��EJG�p5�޴� Fb�l~�Ԇ�}X
�5 ��jE�d�;��S�@Һ�`c2�>�aZ�xz�#��_���Wo����,���~�Cy��1}��H+���Cؿi��P��`&��� ��g���׿6�1$�IZ���xԦ�6��瘯��	�x��.�2��W���N.M�z�����c��۴� �%�eJ�N`Oj9�,=y&?��L���wr��L�P�Ek͖O�>&�Ac׳	�e;|�Z�0���^�;"����h��{����m/�m��*�F��&lk�G�n0�֘�i~ O��q��!
�,T�J�t'�V��z����KUG���0����93�����{R�5�K㺎��
6K��E�F�o��I�K�A�S>�Ni�������}?����_6B���Q�'�f `���^��"�����q��u0G��` ȹZ�Z&U��X�Vc���P�J(��, �����\~򓟰�>�(�I�9V�qS�z�SW��{�㰤�h{F�a�����i��iV6S\�d:�K4������1d���gv �����U���8�5�ӫ�,�ǆ'|>�#��m2����1��Ő�<<<��˾)��x�Nz�'i�C�O!��N�n�����'��#�W�k�Ɯ	A3��GJ>�����	����ϼ�p䏿g�l�O��x��l��p�Β]�+H�Ηz�b��8��=��1`� ���'��� @��4����(,j���S1z����k�A^-V��3����L^�:K���g�p��n���F"�����i�lHB�b~��x�h�T)O��sC�GmL�mvV�n�}��i�3�:�G:�A�S�VP�0�S��ң=�:A�i:�C��a�k�s����j�f�^	�q3o�rt�	�hu�h�F�jJ��4d�ʅc�6�8�C8C�ϟ_ڄ��Z�mֲfk:U��ْY ��,>c�Xa�_�-�tj�&�V% ��ǓMc�3ez�cΧ�2͙ƥ#t�'�yM�F���V�!`Pm�dM֐�}�r�����������X�F�n�4a.b> ���k]OY��%��"��	`�P~�N� �K�t8�H��K�����i#�9���)���:<�]�M��CT<hq6��u4��a=�w��M���v 6߃9�pP�����G���z��׵�w�|�-�	|�.���\Aٛ�t~�2=@\3 ��M�ĝ]V�ܱR5)#�3�Zm4�.q�0�zPc�Y�MРࣱ��F{ҵ��Ae�ɪz2�=�>��F �U���d�
wa#A�A�I@���ժ@EZ�T7����oT��U�2��o\"��rM 8�^���*�}*����=������3��	�@/���cf�_���d9�!MU9���䯠!]�}����1���+m! �l'� -����@d���1�wa�!C`�U���̐t|�%��Nn��u41��k���oйvv�^^)�vr�~گ*��B������P׺�J��9Б����04�;Hkz?M�!��T7rۛ���N:sS<{���w�Ş�Y��Y�T�@]]ʛ��v�PgD�W=�"�R�Y���%vBmS6
�9����*4`�#/_����������n'L�ɦ���ܫ�1(#�S�b6z;ث�ԁ3��݇��z�Ǿ����Mc	н`���_� (��}A���0�aC{�hv��4c����{��D G%�W<m�|��.�:����Ήl������W?���i�z)�R�AC�,#�`�ұ֐��>���S����w|��&w�^��~����o�yЙum� \��<�i`M��#��`pa��� PX�������M�l���᮹i��j+8!�RWE�Tp�8z��{Z��Sݐ�lb�܈���)_mx��Y,�	�X���}������`��XD+�ܴ7�����`�>��������Åwn�{�uY=�����@�E�:����ϫ��+�c��@k|q?i�qct�l�R5X,��Mi1l�Ʊ�&FP_�5��CύyQ�4H�Nn.��ե�|~*�>�N<t��q�_�U6�^&l��g�� P~�Bnj��ns�0ɩ����*��I`����a`�Q� �a�S�G6��dx���MED>#sȊA���6<�|��q�HTC��s���k�~-��>�b����>�1��A�S�Zj��xޘ�������j�f8,����T�g��̈mtn�����b}}=�����o�E�qMp��U�fK�!ߩm�u��������8f��!�V�߫M<rU!�m��'�&pɍ�R��ל��z*7EּխR
Ti��}�B!��� /Bp��R�0BMGà8�S����ۜ�E���)z� �_%@�����IA�����6������cs"܌�`�N�j���߈h�"�U�	�Cr4�Q��+SK��|2�U��Ik�fņR��K��i�q
,�4U)�l
���\e��"@��0j�S���0�=�#
����y�umN�RѨ�X�<�U4���bצ�­��`��,j�=D?Wc�8������y��V�xC����k��`�q+>ÝV���H��
{9��)�m}w!Mr�c3�5� �3yptO�K�;D�ٍ\]^�۷/���� Q}	un&X@Nf��Wf�1��@�4kZ�甕fߟ���R�S���߻w������������f�5����[�^A�s8���
:���s��:l����`��ͱ�Vdq���B�	�/��I kz)P����}R�����Ǵ�>x��8
��{��t��P����?�p%ʽyk���׳��	@�Y����F��ӓs9G?��SH���g���E�E,��*Ip�렶���QkU��W�6T�ɱO�H ����$y�z�>
Bv���i�3�,%�]��}f�7�{Qg�k֟�V9ԛSd�c��q�����"��S�.��޴ ]1�+̉���M�!0]7��.���7�j��R}w�M�O���17��ϳ�)�32vZ���<�=�X~�ӟ�.��=a��͂��T�T<�~��lG'_�Ҽ�P��=O���?<���w���ݵ�!�Ņ�}��XFC'K0#3(�E�¡�V�P(e	:�h��<ʕF��P���D2�ZH�I8j�&�e�6,̑��h�6ת��>I�W�)�ࢪ��c�:��I	>4o���}q��@��@ޝ��28Ѻ]~8�ǎoN��}��z���;l�ݮa�l�����΍ًOln���
����s�c��xdT��e��F9i�$9����,�j΅�]_�E�u������5A�ӹ��_H���`�h"��tr�c*o�>���r�u���AUG1uvHd�ܐ�{J��\������qִ2d��Q�k��I_�Y�/�fl<�n�c���RgX�{??c���� \?
£�@`*X��V	h� 2��f�
p2W��e�>=:�nh)�,����"�Ռ ;�K	�n�v�7�Hu_���`NZ�z�¨�^�o^rq��!�X�Wo1���ܚ.���1���@e`����{oo�����:���f1@Vtt�����fx�k�@��"�hH��lp���['x�w��X�VlD.�a�49s�޷&(�	�ڀ~,�rswˮ���]:Đ���C���H���(�+
�T2�)����4
���5HW�s�) :��q������=E+�J Sֲ����\�H@9Bd�����`�: ��G�9��:*-ٴ�`��;�<�g��g@$�k��ήއ�!h}���m��}�{�mf������`��u�E]w����-�[�\'�0^(�;�QlE���-�j�k�9�.B;�3K�9ms@Aĥ�i�Ls/$����_rЫ�D��NvQ&W���Wr��T��8�����P�{��$�Ԕ=� �}�1W;�zu�B�p�Nό=�@(�J�F0��Ç\V�ٜJ����>b��@�����g
{�%�X�>��/��/}��Tww����^>��#9:��5�o�8�>�l�5#�}v~^�.���L���m(}��'	�O�}A���Q����tpx�>(�~��tM�������<'���^��U�嗻 ]]i�3�����؊���F��Ӥ&[�:��_�����#����qW�G C�WJA�)�A����\H�v
��3��Չ|���rzv���7����]6z�~[�K�w�^�q>Q,�H�,�����r@;��!��<)|6��ᱚ/���!�6�(=��j�(�@oZeh"KZ��@�v4WF�f�P߇�@��h{%�	`#�le�*��-|�P�(��
8`.�L,�zÞhڮ�ْ����G����_��/�����7	��lM욖Dk{��
N�d.��x�T�R�53'��ŋ�����=�U6-bM�y_#������d�T�M��@��}Frzz�F�&�n$����;�;����Ф��D��kF ��ݽo��Ɯ����i�I�lH���D��O[�Q�;��^`QFJh����6�z�[���W!3�s�~����6��n]�q�2T-H1���lG46�Pgi�Ъ�&��e5�"85�x�N����d,f�L��� �غE�4�zD�&��Q����s�-�D�����"��Pi}o4C���m��b[i�a7̕�W�s'ϑ�t|����Γ}�HF�B�z�������/�k�:�z4'��-Q'�r�������P� Y��*�����F&�ۅ�2�}����@E��<�8��曁�.��$��������h�	6�u.��,0��i�;<R� �V��Q��R�',xJl`�e4.�n�@L�}H�m�H�ǲ^��a���\�1����{��n2k�J�1%5��oL�T���M�h69��x�G�r鑢����5��ZC���h��F�X�=˂ C�` ��5ǫTaJ� �|�Tx�fM�^�u��G��Ω~��:}���}�� @�{o5� �i��	؜��^3i�������[��^�|CѺn�A�@U-IM�+��~M:�jY��~�TC���{&@5�xh���U�U���TɫۇR��Dq��?�P�4tY�'�s�j���'w�*���P���b!0��bLN~��G3C�n*��V�N���"�؋+9��@������6�l!����h��\��C��i��斅�p�����
�#~�ߞ���l9WG8Ԥ�' q�捜��PȢ��YPW����_��\#�b}!{����������ۿ�HՂí�N��4"����k#9T�3J�x�e��Ӈɏ�K:�(0���O��h
zcH�auXs�zAa�Φ74��Vr���k#pǇ�f�����Z�`e b~�f�u-K_�P.�J"���}��g�/?���d42�ہ5�W��=fH`��sϔĖ*0�˷߾�W�O�j�PrJό&P�l��C�����ђ��Xl}��+�u�
���,�Ґg��1�y'��'������Z��g'�y�/Ch���	ȏwj�����߈��[s�P�$��&�����}�a���Ǐ��\GF�>��l:�Ms����f�gF�  � ������e>�R!�����?����9��fL�c@����&�|e��T�d�(�j��ӂ <�82���0lP��@Q�:6Y�<����^����S���C��V�,�������&�KN4��g��\�A��	T��w&K����܇2�|{��xC�ƌ�Mv]3]#���W����Xu����A|�������E���?�s���;xm㚊_+9б H
[� _�JU�_M�7��q�Ho߮{��`�3P�,*u�Um{;P��R��I�eQD�u���!O�8 ��[T��Y�ݙ�
�y�N+a�R�к1��!����K�1'؂W��F�7a�*����x�<�%u���+��tk&�u :�ޮ����-�-�5��Z}�Fv\s���jm�U̯��y�Ȣe�ݣ��w�'�i�6?3�u����ϫX�����(�6��k@:\�u���Y�e��B^k�Z�Xi��g5����0��k�A�L�Q�fاN;��3
/���?ɡ�I�
�|�+s�n�ktOo-��ο����`Vt$f����e���u�Ǧ���-� ���J5���������oM�DA+#t+n��R�U��u�1[+��3��:%\3���#�Tɑ�-�~�����ƢG9zFM�f(YS%}�k�z�M��,�ij!�S�5*f��J3.-$6��U�J�rUU���$�JN|��$qz?q0,GT���B� .�[Y0�@�`�-��1>?<�c~��-D�S���A%�M�P�&��|����-���4���� �	}��V�4_�ٛSiX=��}�����19/�� �����M��Z(^p�L�W���R>7���d$��O�y�����)j���?�ͫ7�sg�������u�{�|���r`�9�y ({qy�ƅ�V�W��;�cP�A9�H��h ���t/u�[���{��[c 2��i�syЮ�L��i�^�rV�������/C�
Ƹ���7����fa�����̓��>����?�� @����I�{������o哏?���=�T<TYKI�e��Pxܹ�lp�qw������1���iSK��rT���!�U��Ἧ�����:?�q���-5��z�� �{��)�������u޼J����!��D�,UC�Z⸥��Z)h+��F��j�E=n��˛���U?��f�'��`�Vf��]0�e-2�G�����{�5ߔCN�=9y-�|�Y�m�1�����T/Y�M��T�B�iy�,뀛�¢2J�Z�BE]w
w���W���fѸc���!�¤��vU��qF�yjW��+F�ώS�40�\�[���;F�\��3˲2��T��l�$�b���b?3��x݀D�C�7���7���=���C7�����K�o|�t��Hy����D���ss�7�����g���Wn7��w�����iA�����'�Π���M,G�t�7R-Dur\���`)H�'[Ӳ6�?��	���\c�Go������r&�������5��c`�{���I��qo=�^K��q���;lG�;>��s�[�Y=t'�[�X}g�%�v�s]zۀ������q;~<vx1������=w_�O��>�6�|ݒ�{��Mk�u�@(^�a��L��J{��\�x퍥ȡ@B��ҧ0�{��׋�1A��<��b�������$���5�oU�9�c��<9��,�}�c
�,�h՛)�<���	�1�п�ސ@Gi+���4���R�Z�xUZ^K`+]�u_J#y��DNa-���:�^��/D�I9j�w����X{U���PEk���x9���8źM�\1����Db����5���O�U?;9Y����s����Ilٙ@H���"I�Z��©����?LT ��ބR@C��	�$�peY��t��c0L�>��J������i���{f��PzV�e���ԐG6ET�Ϥ�$�B�4�Rq�d{�tzU�k������P-�C
s���>��d)�_��o�~�1�w| ���__�H�Gm���ڏ_��2L�>ؿ/{�}9���<��V4�	�u���X��yr�N�!�	������L.�/���Grw;a3�ir�v����=9>>�#�Fk���8��hU�4��=;�g?�<�jT�R��4]$�2$X98ڧb�1�����/Pb���0����n�I8K�����t���BP�.f2�$�����lG�NZ��6��[&5��_�`fp%M[��5R����-�k�X�g;M��*���}���^���̀@@�Ɲ�!��Y�ˁq��(����[��1�,[-��@��X�UX��-�B1��_O-����ZR��_xc��?���W��U��U�u@�����bph�\Z,���nm?�֣+Z�Uk>
��Z�&g��_z��/UU~�jYA���Yv�)�t�v�~<K�V�y@?�&dNp<����km������՟���~��O��7����&���.lp?}����_(����<p]k�5��"Ǯ�O7iE�ȯL٪�Lk$&p \�N�Xw��+1��]k�\Ur��+��b�l��GU^ ���&L|�rG�~�F���!v���]
�調AO���3���|��L.P'�7{ꊃ�s��t:n�{�J�j�B�����㻫��5����aa(|��c)���3�J�ZZ$Z��(��c�̻kU�3f�5)����mT�������θ�{q{�U��x�Sd�<��y�����u��]qeQ�X�1}��tH�ڼ}�t7f!��yg��Q�{�����~/ �_�VV�=�`cX|�+����vQ>?�����3�ῃo����$ਃ2����^�Y��ި�L�Cw.~ĺ��5�kd2�L.�Vۈ#�t��*�)5�irF�D��ʔDs	X`Sӹ-F�+�z<�
0�g�4����T��(/'Wtv7����^�Z��o/�d���TiDň��D���%k#D����U��g��z4j�@J:������6T=^Kg���%�Re���d�l�Z�'3�VQ�n|�"�MU��o��#�Bb�F�S4 [���+�z �iA U�	��v�f=gc��sq�~��Z���� ����X&��S��3����NU��q\L$�4�['g9gւcY��D4.2:U�O�8\#��V��TJ�P������}B)�z(�v�:��h��Q�r�g�%��T��� I���LT�zP�`�����3����7���f��piû���膾^�ҴFùt������x@???��.;�62W�4.��)���@����r���`s������,� �W����}�iz�*l�&�3�l9�p�p=~�$��LJ3��� �E3��K�Z�����Ҥh��:���hԬ+��{�����!'�NXL��m�Tc_�+�s3��a[ܠǭ�nû�[���N�l�B욬��Wi��C���� ��N'���7�Gu�`F�q�>�,8=���39{{&w�� �5"0W�q�k� ˨���٠Y�:�u]��%ۡ�uۀ����?�[>»�탼��;�c�����ͪ��h"��g��Š{#h4�E����f\i@�<���m_���o�}}x�P�l5逹��}�F�8�^u>BP�H�UU�gZ?/�_�+��J�N"�������f���{�?���{T���@іkzc��b��8{0�#~���������S]�� �!l�zY׾iw`E�1���u:��3�5T~�]��5E!%�Iӂ�x���,zQ�+�qe3��b����f �����L6}��Y�8��|��޹b%w��T����z_Ϊ֤���^����<����q?�/�������λ�︛�n���8�����Pq�w����A:�p�sg܎t���]���U͇����/��s�6փ�;�������%eV���1ݾ���Qb1i|�I>C��aך�U�\t�Lw�R�~����Ɣ���B��׌u��؞�Ev����E�U��c~�;�R���[^]� �9i�k�6Y\��?��r�{��S]���J�s}W��2-Rk�TuϲWeۂ�YDb��m27�7y�#\�"9{5送��Mz?���JUd��J�G(�-V����C�:�=f���|f���'O�qg�bQ�_�6�g�2@H�^��[�2�4����6ݳ�P�t �1�M�l؊���q*+X�j��d�"�Zz���V��9 �7Ƈ��J݌ j���f1�*3$��JYsֺCua�\�Y�v�7���ƞ�3��/|կ���TUN#�:ަ*W�� ��D?��ӓN��祮���&��Lb���b�f�V��r6V��v�Y.h�� }=���g\��8�_�G�ʗ?����*9ο��Q��t߽�J4����٦tG:��>N������bJ%�U���!�z��6Fhqns�@�f�|(0�������Lҹ���J׎�	�C�n����2�2���-9���ImZB�a���!�fP�V+]ӈ跬����'�п��	�:_γS��)�>�Βӷ�ʠi݂Ƅ��XS �&�|zy+����8�ד?�-��0�c�|�*��҆��jG[�)t+��*�N�f���X��b��9��f�
 ����t�Ǌa#2�KR��1}@�\^�`o_�;{\Ahv�y�+�F��ۭs�[#l�x�{���*��Zn�gN�Q*��=NS(��=�"���%_j��t����C�H�B-�O6���\�GO�������jB��릱c;M��oCq?Z�m����d��ܣ��Vk�b\�@���X�<�)�X �ȓ^]]�%�ww��_��W?;���R���?J��Pw w�ܱ 5�_kjy���F�*�	���`4��9wdj�נ\�6�qޫn�M^�Z�ޚal�hC!IZo�. �Ic]��!���̋�( ��ܡڜD�*yT�fx7Y�N�`��4D{�t7���S���t>2ϛg�{�H��1Vz?���;/�0N��Ι�S_�3`R���f�����'�Q�����F7;�����N��R�m߅m��A$wj�������Cy��`tT��r͞mG�ϗY8��E�g����7��-z޸g�&�13�=yWw�]S�~��ɆA�^�y�1h�r�B�M��������u��(V�y�����/^d��[��8�{/7�n<r��*t�"�g��*l��{+k���T�,���/�����Ū�_���6a�d�)&��:�Se���u���\OXC	˛�	ճ>>�����®�p��XTdFP�>�ݕ�t�{����Å����q+.'%R�A$E�h}=�]���|�
���R�L�8���w�խ���9̢���u(�t�6�Y[_U}B �6k�Н��NRbK��_0�b�Z�Z�~�kQ��t"y堐��J�A�5�lP���g������.,x��܎�[tE��d�[��~��,�ӻ�qc`��E�[֧��{%�����jA~yr�勧��/~��� �s�Or���~���)��/L(!�6�|��k�yq��������Q�:����r��a���'���]ܱ0W��U�']-N�T�����*c���Y�g86�[5�ۓ`w�����o�� ��6��q��υN3h0�m� �rvKP��[��'9���O�E:Dr��ҺR��s�1�ݽ{S�k��� �I?GW�	\���?�@˻�����^������l��ص�!>V�G�m��|�Z���֮@�s���K�^p��>7%�c �` �ѣ�ev�ɛKnm�W���8���l�F�|Cͪ�P� ��*6��fYߘ���x�?��"��G�l�ʁ=��'wc�}�`�p�Jmo�O�c�x�!@G���S���ն�ٲ���S�Ҡ�{���������p?]T�{�Y�v(�j�HÀ��-6�e�{k��@S�i�b8�~����O���0�Ɋ`:A�xD^/d�apz}��LUz��Z$ �b$���.�r<)z{�r��.hWkS��k���e�f�S�{n`�(��!TG1!m���oO�F2�ĢR��g��P��bb���,����+��]�\o�G�y��=�|�ҙ٤A�b��Z:i�ր�Gc1�/F���;�ـ�[��������3�}�� �C^��$S�2�
�{/���[�е{����Y̯u�Y:�����l;����8�c�q�٘m^�;����W��}Q:CW��f�8čGm~G�����+��^�1��V^e��U�$��ׂgn?���Y�}�p��1��[6׏�S"��5�kt�����D6#YF��!�����J^��5Z�+��S��J��4�[���k�HMH
ě�X�Q�CY=�*��?�X�-��<#@��HZ�v�E�2�����jL����?$��`o�Q�W��gO�[dNz��;b��YaK�Fզno�>@���Ir$no'��C#Ε�8�x�|6�]�> c!���ʛW�^��� X|��{~{+��Q5S�8>�S�M9k��Sw�z��V���Y��}�vl]iѥR�U��5��)�	Y��t���@�h���I�X.g�]l���B�>���j�(�~f����AF�B%�}�t��5��0z}�epn`.������bM��r�l�ڸî��9(D�Nm<�	ĺ�z#7(jy��}������)i�doԗ�������w�M�i gՊ}"ल������}�7[���V�>��ו���T��l��}��zf�S�b*�ڷ� }�PR�kY��4-�#��6+��0J#129�5�+jd�Y[��i����
�K�cTc�G�`k:�p�z(�m��SeI*+�0�X�,h �j�'����xLq	�c.�V�\�� �.�V'[���6ۿ�~����/�������Ϊ�a�!����lK��2wMŠ�j�NWT��*���z����!���J�TƁ�3>q��g�����|#.@G��f�"��尾;k�� �_V��7ũN>�8��W���d�>�5��H���ι�HB@R�q0ռ�F�˨�٘����~5�c���9��6��vfZ�T��7�m�d���7tkH�Z�m�9�ܐ��;ؗo���{�:lЮF��~���O��i��=���kv�mV��R��x�д�yTr��eu/ �Q@���΢t��__�f�o(�Z~� ��M�V���v�T?6�LB�����'����N�W�^�
�eX�B�!��L�G�6�߶�
 ���6�uy���}�#���H�w��)�M��<SZ�"ߞ�]V%��J1P0�i�_y�@q��s�&d�_%5d��r,
z��~�]��ͥ���j�39��F������nP�����[���,h�wu�5#R�!l�>�q�'����.��\d�z�w�E�۵�Q�D��3l���X����tܫ��x��k����+J�%_�F�u|;���yt|n{VԳ�Q��J��{��n���|��k�uW�����y�9�l�Ċ�֍ E7'�
�C�P�)n�򪚲9C��q��RȠQ^��cӁ=�c��I��B�j<蟤Ʌ&��^��V�55�L3��d+���������[���r���������/�.ɱǸ]__�:l�j����-� 轀1�#��F��RH�/Me�7J@%�aS��:�XCn`	�A=�z*��Avr8懰����4�j��-����q��1@v��
����.�h�3�<𵦢#DVF�Il)�
���С:�Q�R̭h B���p� �p����+��G�89��*�v�G�CȲ"�=L{^o����,����G�B�4o��+�(< ���_���U� B��<�����1XD\;@F�z�����Q��)k��8��q�,8��`�{4j�����K��}6��7�^$��&ЭP� ��!ת�^�0�٣ƣ��
�`s�"��>H���e��2�]�h��B �m\�� @A���Z�4+ �b�le�s&=�
ҽKmf�:q@%3a3d�כ�jo<���#��+��/5h�_a���Ǣ����>Ѻ��h�@;pk�W=�����Ƣ�|8��چ"��+�2j�[mnZYf@��w�pY5�$7B�ŧ�:طZ�.��-6�2��I���Z'B��?gzݏP���~n�}���l7/�7F�hf7��CW-���n��4l)�%g���q)�m{�~)_�5A�aMy��7T��wyqaʮQȩj5P[`tV�J(m΁�3�4#l� �]�l���su6O�J/����J�B��Ҿ{����f���1�f� �b �ȿ�sW�7����/������������ޑ�}�����o��G�ӂ�L;�5����,<�̦i���M!µ�{$��7F ��D�8�R�t�{���#2�ǔ尗���B��P�)u�v�v�ی�T��L��~����ͪ'������A�1g�>'F�F�3����ѱ�d�R_T�����Κ/��x�q���\����s�*9����w�E����ɴ�֌�y�\b��l,���yh���|�(����?K�c��c����w,����ng'ύ�/��m��ѕ�#vNmak�s���F�����^�g(bV6s眅�U06lw|��������5���s����H`[u�q�ي�:r}�l9��X�����t�73��zvu�<o����@���ZԊ��w�g[�g�,��Ƽ�,�M���{��Qub��|��	��w��
@�㨸�Ė��G����4�ں`Wk��*�m��Z�3]7�t�>�Z��nC�vu��>��Mӓ98��pG��T"���qo��������ݶ��<9�3����}r�*9�+y�����d�?����P�񾺾 '@�0PN�����Bno��d
� \��Ta�"`뱩�^�1 �)���C!�LPd
-x�K6G� �t1�c����D���)��f+
�<��D��[�q8�P0�㏂N�et�#�#��,���X�r�m���sa2�-%�B���&|>`�j��B���7�̹��LM��=Tg�q��` h4�#p����?����G��oA <��h|��a���������2�Ģ�� ���V�5}�p�R`�1{���$�iy���.>��S�����UN�Y�Bɽ,(��k�#�b�tv��5���iF��ˍɭ�pD���P�<��*��*#Z�\cڠmc�Z�Q��H���g�f�^ГF���G��.,�02�o��F�Q�ʲP8�h����)���S�~I����F뻽����vC�߶},mދ:\d�x+�f�e��慮���*���G���dp�*J��Y+�~�+��D�/+gTB��S�B줵���rr����n�ߡUYM��@�y/�V�|�zh���mk��4H��r��on~��K�zP�*(��j���\N���
���=���C�����P����� _���}�VG������f(�RZqQ��d��٭(Kb9)��vbO8~��(�޿G��Ol������u5f��~2B��߲�$�=��K2V������eɮ�}�,L2D'X �2Z��fP��5��hؽ+�G���0�����,:|^_k� v��$����Z ���P���sy��;y��u2�؜R�����u�&����J�"]�PmK��(o�9�>��S�;*n/�Y�(�Ӧ��lU�B���%G �3�aj�x��c�-4_���q؅��@<�\8R�::I�*w6�֬G���,^�S�5�#����O׌�u[����6 1Ƿ X��N��ETc+�j�5�����!��놯4�N�q�~7��%/�3�<�j�<"�#(b���!��Ν�P\W9�sغ�j�b��=y�U̯����<*�h�8�;�����'n�����`O�M[ Ūe���_2���e����w1���/ؽ�gLF<:墈�m\���o�"?����h�9�y��"�����(2�R[zJR�B�9��j����F�b�Ĳ��H ��f���kc�/�b������k���ZO�f1������ϟ�J��|��S:w�sf9�=�����c�<?���3A���ǌ��% A��ޘ8@�wo�P?y�{{{zZO?zJ�U.|���3�0_h�io�ǚĝ�C6�c�`�HYkqv�rC������A%� gg�`�a&�/���Y#<(A�?��bz��#��
Kk��}��X���!�:�oo�`��������Ʉ��x~�;����I`:!�:K���Y�����z\�: �{�@ ���>�c�QU$̑�tlUd�г��{�4�+^7X	{	��f��|u����ܲ~��=�L���eڟǣ1��CL]q�K �*k���@f	~:~����k� �Z(�ms�	�ҟ�h�������k��h$9ST�Kdc�iYP��E��cgp����.�5���f�s`ߍI��#�Z d1b��]*eh��/lvSg�	��ڻ�|�5�B�ѽ?���pstQjߧ�gHa_�B�b^(����n�����ڪ�ɡn�1)��d�)�0�Y m臻�
�" 6V���d@��~�Q�
Gƶ7��M6�1��8`1���������X�6z�,
�����e�g
����)~v�ۺ�W}B���KW��j����w���b�:���cd ��@=Z=N�Id��f!���:�Ӷ���h�gd�!p ۻ&�HAu��H�����pϠ�^�`G�*h��C��r~jsڻ�Y:ǐ4�;$)$v�#ۣ�x|pw{{� �& �R�P��?���$8'ۥ[�@�$�	^" E�N�gUY7]�:���kaiTB�������m֔���h����M�[#��#M0lHt�EJ�t�t-P���������� Fysr&�7	)"�20�0eS*JJ��2}H��Y��Hs�<)%oޭ�i;�r����h���HrO�,LV�	"x륦��Ue���QF��q��e��6뮓��V��l��!�ϛ,�;��i�9�r�Eō!�w8���k���om��M�7F'��Mg,�� �=��{$�����X��;�t#��vƵ;����w�]���eZ����QU��y1���G�m)
��Ꮝ[0��6v�&�rc�|uf�־���g��ƀ:��Q%0��>}������;�A�w�5B/Y�$g��:������}s�l���fko�����y�Q��Fӌ�7�����=%Dk3��ڃ(cP-
)��
��A5ҵ���T��Dsr����\�:}V�Nt�����}s��溧κ�KMU��<�h�$�� �]}1M���^�!�BAI�Αi�c�Q�:�����BP ȍ.����Od1����i�[�?'���/dg4���}�m��3��
���?�t�=*%6�����o�d�`�=���y�+6��6���1M����~���� �'/W<(T;�21c�'8��X�>��	�~������u������4�5�����x ��#ӎh��,}�g�,"{�C ��B�����il5�U8���P7�C�d M)�h�������qm�m��0��ǿy���&bA	t�>y���Ц��ߗUrn�O�����}����i��!G6�u?il0��0����sƻÉe�f�  ?�IDAT8?=�&���5�c-22�bs�4w�5[�;j :SCe��={Ƞ/"���@�]9)ӖR�8Wz��c��?�1�;�#"�k-����1' �I����:NEsA����W��,��_�~���s]��|��-&��Q1Ԅ�J}�V�\��ΨG&@T[�-��Ԯ}��6�4;�9��'��1	Ӛ�����f�X��d b a#p�FG&X5h�J���4�Z3^bQ�l�����g�.�*�GEx�{mw}��DZ�����[1�+F�:�����Ʀ��C���l�ăO!�_�J��́C1�[�S��ܠ���uIfCٿH3r�׭�TZ����X݊=��Lך�� f�@�֪��|߼���ߟ����u5I�Z����6 ����03�������F��͘�1}idZa��n4P�Y͆��V����qo&8g��N'���};�H绣�	j�on����r/��#}`�������g_�^��'KF�勗��"�:��Tx:���4�3(K�Y72`ڥe�f����=
� ���X�%�`ХBm �Q�t���F;�����AQ7�^eѕ��WխX����!VGz�%�C6��hal9�X��Jq.ަ�U�|�zd�EK���2�O��&s Z���b��d�^)�*Q���L�u��+C��o$�1��� �BP5��Ǝ%���
���-^os�1�S�f Jum-�����Ӝy�"�n�k3^�HE����t|�4@T���tw�CGO�d���pbi`}x��.}�����ؚ��!+L6xJw�z�}n��t\,K�@˂ ��
$��c��ؼB����7��}�.E���P�]Dh�����Q����cu��v��/�6*! *V��0	�gJW�L�,Z��������~�
wu��'�%���NIVK�����TSb	 9-��yG\��2Z�sh(ẖJ~'��G��đ�����A��o��?j���s�Z�m�������~��:;�l�Å�z%���4ڟ��d)�j���pS%�����l`k�d3�!��Dõ "mF���/�����חW�x-fs�K@��$���&�{��
�Cu&p��n�/6K��P  ��_�#.��׬}i�\{f�$\�ʊ��f]���C=Ơ2g�)��x��V�6��#1ӋP��,y�,ǊYd��Pӂ�D��x��=�����`���bs�:(Z3�Fs`Xaa�m�����
��vm4	p@@�9p
V�k&A���Am��ޮ�1���-=��==N��-#=�QW�<d�S�ͪ���gP�?)[��~�޼Nc�y�DЋ��N�����@�=�N�ooh�p��#Y�P�b(���������f��eٰ��<w��a-�� �\�x�ؿ��ϥ
��G�m���j���Ț����|��n{zv���A3(���Q��>�6���6��"w��:�yHT*dá����&����_�F���e��G����O�{D�ۈ��f��x�Mk�(LжȐ�mX������D��9%\��
m1t��ںhN�gm׷c��j���WkC�5�	���u��Q�g�Iߛ���u��� ��mP�[j����z2�Yؑ��f
z=�k��ό��(��m�����z*�0��Z�>�Jk����_�NN/�e���� ��!�M�{�O֪>�{�=3xRѮ,y^�]� ��>z���C����c�F��������i�Sf3��� ߾Xhk'<z���$�����Wo^}����ڻ��2}���#�Wo�E~�Ziq������!�E�h	8�����*������4��桲�t/"C�zD#�(�1bF-��Mb3�ǜ�tC�����Eӈ��GZ+"�&��6��d0��+t^�dEW�(LὨ;Ag�H��/�:$U��(Лf�%ra���.��<���
0j*tq��L���f���IM�A�8 ���t	u5:
�6kB���*���&�M#��4����t�e�ↅ�7mc��J���	3��$���t�Ū����
g�h�^YJ�[�pLkGZ$yE��t�Wi*�0#5UeQP�C�j�SҰi���R��zwa}�+�R�ץ��w�iC�гV�TO��)���\u��[���A��>��� yGa�h���$1Z%6�O���>kuuHڨ�<W��C���[���h��"������Sw�j�V�7�ΥM��ezN�	l��Q����	��8���j��3- ^�����񸲬&�L��,���\�Ώ�!f!�ɧ�B�7�m�T

t�i���4FҢf+Kw�YoL��Ve#ښ���{�`� ����H�g��21N6�{�"Wֽ6*�5����^1��ǹ� X�&{J�i�T�Z4�c-BYY42Z3L�`� Xk��b/�H���I�3'};��땄=l2]�����.��9�*&�.��T�gG�l��(�ϙ뽶9�>wyy�E���5~{��<��Ğ_Xp#9t���z��2kRE \��ڂz\"��X��^�Z���tjj���t�wx����T9����N����]����_.W�L�٦I����-�\�s��8�vE��c�}5e��R�-��7h6U��~��{eϖ *,Ik�����&q	��=C3v���8���@�r�m��1C�̙�S���t]C"�H�dmJ���B��DPO��C�}���Y�CFvㅽ��q�Y�r����`	��#��C���>�
$�߈��kCDz�v#gfJat���/>�hYcmQ �sn���f�ofd��E'�V'��(�'�h�H�f��(��i�>κb�:銁����"��5�=��xHZ'�� �AN�g���ߣ�V,ox�9(��#<
B�h���=�Fp�`����3k�i<>���i�x�F�; ��U�xўĵ]z��Y�Ŋ�c�~��
�|�,{A��-�%]�����`T�/��Z2P�F��j���@i�nI�S�ڜ�3�%3E�ǚ�,���S�F���b� A���^�5P���Ͻ�=���f�gAY����s6�wb�
�,�dC0�	iӜ�����SY��{���B@�-��C�R4^e��tMv1S9j��J����&��π�tF���T=�Am܀�&C*Y9�`H/�]K�:О/��X>|�,wY��V}h�-�1����H���I��]^�����I7L��4�x�5�T5�q�L�􇢁7�(�d����ڈʺ6���Q�s�������Jϲ�'���N�~�da���@�9��  ��3��#�iA�_����xu�g	�h!�>4�F���-��ㄇ7B�ԀH�R���O0��9���䇃F(� ��h"B���v=&�J6�#�H�r�j�CP�5��1JE�Xu�4Mr�XW�g_�d�u]wn��̬*�@ A[8<��Q����:�s��$Md)�i�V�A$��P 
������}Vsnd;�d$���{��{�n�^{m�I���(�1l|��K���2�\�L
���t���H�5-�u
����)؂!��؉����E�EH��;�<�ɧD���Р�t	&�v&��v�pfX���E�?+r��g��}P�Z�C<_:��<���T��Q��|e�<м�|ނ���|��%�*sR�JaB�����TU� S�)���YH�a�?�CZp����Z_RGqҗz��>���a�:�\q���I�����~N*�bu-������D#Qɲ���۝��v�?�s�g;9�q���@�6�5Pժ��w>�~)�<���{�2���q��v�w��_�$h&m�UG��@�[Z!/��	"���'�7tfHT �w�?��	]�϶;I!	UB��y>�u�(��|ĳ�D��/�c�Q�)��QB.�J��젃΁Ȕp �8;��E��b\'�$�t�c� Μ]< ���}��/���Q��28fLm��s��A��o,ъ���p���k��eSsF�(V#�I������j�<]�%�Y�^�Q6<��sD5�i���)�n63�?���U2���T��oL�J��c�UlZ.y���[+qpB���@4QF�5�T9[^�����;�|�/Fg']!��X�U�j�����j������@�������ܥ-�^�������T�R�<�0�&�KMΖDs�2���
N���>���*�Y#�ܛ���(DI�������m�	�[��`F�� 6T��	�`@�	S��5U����$?��RJ9���MQ��q��x޻��� F6�L�넏3�[o ��H�tmR���B���U�<,�&�z�h��g���X�+�U�fW��d��FP.0��#ΛZ���3���DcP2`��1T�����$#Ɔd|��5�b���B§Y��������R"�̘�.( �ē)�L< �J�몞ᢺ^ +j�sE�p�t�]���~��s��9��`�.����v�`PR��R�S�h����`�H�/��ar<��\v�	Z&�H报�+l��� �`��dS�
	F�48��ĪM��g���*���a��w*�0�I�7	fX
9�`)���Q�s�A'�O��bV�J*��>��������v�3��É�V׈3�0�U���O1se^�Y0Ȧ~mPw��+�ťyQ۝�Fp�Xl ��/�GEEښ��2������Fx��7�����'��G���o���g�mB%�%���L��ϊ��l:y`p��}d�̂#����8TIg�\S}�@�W��P9��4q���,�ʈG��(k"�AY������������v�7�l�tgI~V G�jKߝ� PGY��xS���to4R�% ˯�Ԏ!M�e_�\8�(��Jz8W��`�<�AQu�$W��xJ+��W��?eÃ��${��ki�g��(�X�L9��A�K�2�1��w���&^�8\ۮ];���&�J(-��~0�C}h��tLW>l���w�4��A��� 5͞zTe�4D��^g���>qI�_Y�#M�ZMt0��1�L�P����"V�{�j��S�H��b����g�[&��h��Q��	9�5�n�"25&�|)k���0 ���P8Qh��U��u=��h�ʅ��\�L�WupІd����z%��$���+�5�mEm����+�=VC���H�)�j~� �45W�&�ˁ�ԀKڎ��&?W8��
㞛F��=�@�����/~0��<�ڒT��9�l��yv(#�c�����ND�t�[�-�C���R"(�ȅ�r�ya�܆2�A�&�K�(��@P�t��3j��bl�NzQ�ʖ9� 3q����{��ęb@��x�W��A�������J0@�=0��理�g���K$]+�?���zC_�8n-�,I�R�&g�DV� ��$�5TM�k�P ���%�f�{%0a`�D˪zh�*x~��it�*֕îJ(|ذ��J��_U9�L- 2�}ɜ>�QSevfr�!jA R�^G���U\SU�c����m. >��kµ㙀����`��cuj�쪯q�l���)�L
Y�O���8��)�,����A�|T�De�s�����Ӂ��sH�}Ue:�����`�
�0��k�5a�y�č����Rt�͗��Ș�$�+���~�π�<���H��#y�"��
��=v�!$�L�n��S���w�c�R���f
��i�J�,�%*��x�Dn�{&5��qt�$Y����:�w �Ô��:n!ד�O���>���D;�m�of5K�k�@������M��l�~��څ��e��읲�8�B<��S���"���{Y��W�;V���j�^���Bq�f%bD%�ܖ/1m�nC[WǸ*�+�A�����~%şi�\�JA�0}�M���~�]� x���vg;!��qL�4A�P�s�%��5Rŭ���`��~[I)���,�a��h]:��o��o	ޜ��Td����طc��^���@���cbY֢ݳg�v��v1�h;UK�|��n����<!����#�xߔ��|L������W��w7�D�}~���#8D:�b��+	@��ga��y�([�R�={�������w~��_����{E� i�TFGS'``Q����Ǳw�\�26�dҳ�q�9S�\�9�:��~���u�,5u����F�n�R��9�7`��h�������;
����#�)�$�I6�PX�F���j0��A��Q
��wL�*�U�w��g�n�C	�y8R�$e�ˣbh��4'h�U@���$��R	(0Jx��T©�S���C�dF��P
[JM�!6l��-s�gr�,��e46�dz&�� `���>p�x�T����7)!H��`�0"��	E�%U�R��M�p�,��g'�H�"/�Z��4w�4,M��$���B�|"_���~�����ߣ��,�#ò�����;��y�P��נ�3J�[W���x��q���p"uPr��r��%g� AG���;iP�_���NHAHA�w���?�ѕ�[=$�TGZy�Ղ~���_���z�v�� UFũ�}��ܰ��n*��,���v����O�҉v��X�p�uƱW�#��E�����D��J%b�%سȩUj_# )����D�P���d����d�+��q��vX��_�u�{f$�_ݾ/��;H-��l �'���|�3��{�D!��L���W=��-0��/t���r�xm|�Z��~oC�+��x�+J=u�wP���VJZ
!]�$��v�s5Qs��E��[��s��|_���I�������Ƅu���;'�����Y�:���J @	��^gXI^`�tDf �֏����#6z�P� ��Lp�����B�ApT��T�<�.�x�hIr��7$�J�z��|��!��pog�3�-�ׄu�m��a?��A���K�bJ��$֏����}����>�7��+���������k���{���L®a��o�0�Ğ�@4�z��,(9}���16��`j�kTQ �{�ac:�{�[�����J�9�A�p�0W�#� �;��CP{p��'u;ڑ�p!V��c�wQ(�Z)q�ꐋ�5�'SD3],��A׊�,|�!�g����ُ3��ZyO�:��#U>	$�2�������(�M�M�>n�8���!V����/�� ���Gl��@&b"J���@�!f�E�s��{�W��>' sV�p6�kpL�@J^��Ԩ�`U��pЛ�k�^cVO�h�GUi�X��~�I� �Ǔ�)���,`K��$����B=�[�D�M�*����-��?9m0�5zc�n6�F���@˜�hA&JM��ӾҐX�ڑ�r�M?� ����^�L�/=be`���}rw�% ���5�Z ��Ӂ{{�"�?)���A����(�Fⱉj���G��ZɄD;����������^*��Y8�s��@�7�x�T�똬@�������_�x��믿������7o���O����Ѩ��u�FB�eu�Ʃc!5��3�	�&���sE��j$���^�����!G��A�ΜƉA��`����~���_��o�����<�铸JBIeV�A����xou���\�E=jt��l*��@Sag�Y�BKQ��4�ZB������!��ѽ�*�~sҧ�
)e�(<�>&�I�=���+K��U���\d��b��;���^��>'����`~f�Ȉ�8ӥ.��]�};�bc%"I��vP���&��#htIW�1��!M�5�3F G&��fQO(�MX�;��1�֍�� �,3?~J}(��gO����y�O��Yt�5_�|4O+)�Xn�rU'�kp�����Lȉ��j��Yf�t$��E!dF�Ԉ-tN����j*��F�P�ݠ!�BF�C��;�����Ӛ!p@�鱒�����fä���S
�ěUC��=�Us�g&&řz�`������z�!�7Qc"�+7ۘ���G���=�G��$[��9�E��~9�HzRH˳��{^��G�A�F�sV4�Q����ڑ��aؤ��?�̓;������==���[U�pV%�@|T-�r�fc@(�zv� 
�ֵyp������D4�|��Th��fR=����0�(΁�n�i�䌠�(5�����F�/ +��Im�A
J����j!�ř��:oI�9;_+(0�{�j[��}�J*�B*JD�v[�W����B�����:mw ��YUDϫR�B�g�TS�5������fU�]͠��(;�T*U�W�Ӱ J��U��!p��~�3��DNG�Z�^}m�&���|U�/S����6���߻���2�,(kP��Վ�&i衦���t3�k�Z��/.�X��B�W���գ�����(��IW>w:����9�2��AR�P�������@G��6��� �����+$M.�S�}�a�j�� ��v�)+�$����CIJ��,~��6%��j�TS��
�)%�e����4bu�"U��f}��!/صܔ+U
S�r�Z0ț$���#�ox�"�J��[0�~	j��:�	�J�N�/5� �@�v�����x�n�,��"�J{E���v.W�_���D=g�mu��)xC)��z���x�jrnMM�s]�����l��I�Ģ�����{�%I�)&���p�N�MÞ�~l�^,��j�@R<��xM}�����@kpC~�p�]����h���>�>~������V����؇����y��{��������G2���������؊́x/S���TC���NA�lJ�6��=�+^Ԡ����kJĥ`z-l�; Bov���'��� "@	��\sv�~x<�ic�aZ22FQTIߛH���` i�{[��1<��,��"3__{]vT ��n��6P�>��+VL Z��v���ٳ����?~����������5J:*��2����5�+��L
4�T��(�g�2xj��q�3��yilH��u�؄E&D��&l������|������O��7��m[����w������=�g�~�a�AI�*h�S� ��%�vBΤ��o�8��ə�/I���� ��
<<��0�%8t	�J�*St�M7��׉��ŝ�%�9g>���i�J�T
��u�H�/ٍu�v�*��T�Q��|�ҍ٘�ڹ: �H���4@�	�T�D���i�i Hf��xi*_|�@�����;����s�4NZ�c5�Yrg"I�j�׻��V�JRt`���i�Y�G�(�*'�w�[n�@�`[� ��{D S)��L�$m�ޞ	+�d9����F@d�.�q��!pA�6͉n�Ό8$�D�#nR�b? U>�zdJ�z����R�(�OX�\ì��o�E�JC��fz_����4��Ys�h�>���I���9�5�F����~Z�e���`x�d����1�FY���X&�����݀;���D�J�\�I���d�R�mMRN����x���c~?��y��U��k�^�9���{u���rR�3�%&
:�t#�Pa1>���l$��"U4zO3�e���%�K����}�r�ӿ�<�Z�;x���q��?F�0��N�;��v� ����ǞƑ��+�����s9�r��H�Bp����s1���8�d�B����WG��|H�� Ei��Ipb|i�X�������d� M��x��{J�GkJ�K�JHAe���dA��w�gU��6|�N�'�ךY�ep��3Xݚը�a����v}����d�����R��-�L|r+��K%��� �+WY
SogWר���nF�%"��.x����I�B��o�gm+�T��a80x,
�G�c��%���� e�x9���U�H�6b�aG ӑ>Vqxc��?^���44��z�(���l�����o�#�uiJ+���o��*���> ���,u�KvmV�eP���f��`B��q8�E����� �W��Z�ܭ̫<{��J���:��)DPK�����y#�"���U6s3������FF{�Q�R���xͫx&����
��D���s�9D�l��(R�f��mB�f\���e�<�7,�ʇ6.2�7Hb_����Ha�����V�(fH4���˸�}��V�!����*r�+GW�OT���=;�!$	细��w�D�8�h��C���@��*����Hh:�`� �a�зq�.YI
� ɚĊЧ�2�I�K_H����X��x:�F��FS����]C��.ʠ��Yt����U�,[D��8�$(D
;�t��® �!� �dA�m$6�j����χ��~���)���?M>P
>>��_���}x�G��i� �j�@�Hm8m��
�χ���������3�K��ǌ�eƸ��kS�W����_�L��x�ʻO�~�w_|��_~��ovu��7ϟ?�X�'���O>�����n�x���O���'�������'u�lmS��B0O�t�k���$''�^˃ ��V	43�~E�M �x�I��|gV=$���� 8��am�W烹����H�r�D�M��P��#M�U�,e��jq�|�P>d��3ҒO��(t͙�FWZ�PJ*T��f��]D�J�"�~ +;L�^�*������Ӛ�.6x�d���~���6�p�a�r%�j�6Q���&f$-I�M=�%%��$Ĭ0u�:P����Ný�4�#ҳ�D��S�k`�'+�N������2���h1u"�^�u�ЮJK��`�{;�4U6��Iy�LS[�SU�N����ۊ��wrԝU��SD#[U��u��x�X����nu��Ս�Iz�TU)�Ӱ�Tj% x����LK�F���e����i�q��D�-D^|o����_Z��3���k�W����-��?L�����.��$�� ��gum:f�9�{	�n@��x7�a"������jX&:��DŽO�"�vA�(�la���>Go�k�>P�/q���7�	 �c���xG���$7h�n��� w1�F������&�&��
g6 `��s�9'�fU�g��*(�.��٢!x$Yu,��s�3��׋/�ߦ���Q�k�k�P9�	�*)		�&��֫���rz�A�Ѧ�_\Xx@}�71�]�g���[FSlh�po��פ@�/�?,(�{�z�4�NL8'��R3ep���y`��)��x��\���U�3t��0��^6�����9a=p֡�zj���$K�^L7/]q@��syv�%X$��^�9p��k�d�5��V(E�΃R�Eԁ4cPD`J|-; �!���U`Q�T%�S���^f}t&D!s�<��B�o�FX���%����<Ȍ���P��'Q[+Ҏp�
P��dn���nm>��8Sz ����9I�'����K6��+A��oI=K�U��5HQ�:s�Q���|���z��O�Zĩ�8�na'$����=����aI�KSW�A�tJ!� �(��6�k*�$�������p��Q_��?L�g���uh�OL��rVYP#?����9y��d��L������y�-/=�:,"C�����PԞ�9%�U�H���en%]�JJ��"@5CR�c�8��[�Mf��c�����w��?C��~�Y���|$��P���� =�l�N�,���?��I�B�]6�g��0շ,��y�b�H�������"UјK�j����2�U��x�����N�j.1'T���T�g�Hp^�r+�:�����8�Y��P�_��7�Tg⾹�8�W�U��%����_�꿼���?��x����y���4��]�D�E�o�t���$�;ʊ궟b��F��ԋ�o�����զ�WM�={�կ������}����<׶(��~���g_�cHDʰ������������?�����+1������O���w���yY�9@EVƬ�kg'Y��Px0����y�a���pss�4�)�<T�^���[:3����6�Z��P���S���S�/�9gV~�Ed���
^���@Մ�e��m�����c3�`��`�a���	�]�d��ٞZ�{-������O%n<�V P@�G�[��Usv�(f�lC?��Ջ���kGY�a����Z� $02n�ս
LL���BR��ܝ���@�G�B�}O���*PU�W���8e���5d����)0�g5kun^�>�
�ʗ�3S�H���?���8GDh��0�|�p@��J#� Q���8@�0�ԝ����*c|ޠOf�+'���Rp� H�
�FW��lg�nM.l���<c?vv@�	���L�㹗�
RZf��P�y�ݔ�)95���d>��CtxT(I��)Y��z���̔��g2�Hn���A`�a���(~$�V]�� �!5zrU9èW�s���ěN3�O�Jm֋�G�NY3�@� jNM�7���|��uNIVU@J^�5��=��G��ݐ*��Fbns[�3���6ژ��í�
�R��� �@%O��N���L���c�sRJ+R��9����� �����@��q���ELp�+V�:���@t�?��i�>$%�cIRܖS_���(����A �!Q %l��U��c��B��H�+ڣ8�#�L�]���S?�)��2\ ��0�8��A�i�t�����_��`F�/�A	���h������ͻ��3yyP�,���Ftc���B�="ч*g���F{yrb<ߋy��	U��F#fE��1T�N��4���6h#�E�8d9lO3p���pD[��|@����{��vEp�L&*��)7�r���#��Z�ip2j�����g ��^C\sSQ}g�Ph>�f�LN�'%3���m�>�]� ���ԍ�[�ݻ�;	BuHB�����$�$�Lo�T�X���zu��{��kH!�^��X�b9���,�bbE�"];�M�8`��{�>�׹r	?��.�92+���h!	L1� ��P��E"8���sm�?�sNf�^���b�K�A�\3!��b��*~�g�R'��sHc!)ν'���hà� З��3��H�_I�h�Vd�)W$*H�%�>�N����|�.���Q`"����z�6.u�x_P��s�/1�R0^bx�hW6�,q��{�h����I/
;��l����f��V�����:�G�K2��x2~���l��5'r��-6 X��Ps:e˃�I �#~�>�c.j�,����7��?_����|������w��5�)r�m �wpo�^\>7�fe��'�F�(�7\-2&���NBjj�6��7��ç_~��Ͼ�������?�E$`���<N����>��?�'�����;O�~��_{�'_}�I��<�&�f3Qe4w``��&����pgٽ��AK��^�I(|8(�VeE|H8v$ 0���h�
�~8bqu�Gk8ҳݖtL}���G��������`���rUE8m��C�r�$��X�B!�����&D�Qb!�A�qNF�5�Ƅ�	��z˯�.��M�Tb���GB��C�.��$Eij��hj� >�8�
ZB0UfE���0֙R���$�ݤ�[.P����0 �g!�?VRP=X�0��T�K���\M�Y�|������p=_��N�����r�h��d'c�}�Tm��0JT������G�t��i!ĳt�U�k@��t9�jtK���nSeR��J���
]���7)��򪻧���^^^�:�~��c})�J�w%z��u顏��j�
�BWp����������oo/�jJ){�iJ����Q�� ��_]� �M��,[�p�&�[��~�L�*p?� ��RU�p܇��K��\6��=��`aSpNX��k�}��X�r��{L�yv��1'M~�g�@2��j��������PTɀ�EE����Pa`�t� k�ݷ���,�8��4�idz{s>��3����\I6�u�O͹#��6R?Y�W�k����U�>��Z�)�%6c���88��'	x9���S�L����e����d���j�G�-t"Ii)��@�,����3��Te�ٹ�$��)�RUH�۞��Z���7K3����B :ae�+1	��l8�D����X����FTYW�<�ސ|_<8go	�Y�C¸���8�C!��=�/H~&So�8�o�Ps����in�hYw�X*4�	6��+�sLZW1��Pir���zW;T�ù;T���
�P�~R�ޏ��8�P���n\��3��z�B�yp� X����J�*�D�q�sjPn0J�L�A{Zsm�C��*����������&�VA~P4}B����St`�.���M8oE@9�@g볌j3@��7���a8~�;���
�����>�i�I�V��T%�uP��R#u�	��LcLgHU����l���ld�U4QKD�c�Ra�"{�VJQ�t�Jt-���^�[%�Qc��-h���ZU��k��
���,�]���+�@�I��8���4�F�Hc\4Ai��LIG��i���@�#��Z/v����H�F��r��p���Zc�D��ٖ�+f/��jդ/ip��dOp���=G^���)��V�^��,׹}[�=���<�9e�ŉ��B��*� �Y ��F�I�d9M��Ͷ��s�d����_�����������|����������������Q
��g̝�Tf\'@��4Y19�`N�(����������o�����}���/>�䣿N9�?��9�|\��������ݻ|�᫯����������=���5!O��Rp�E�f�ġFER�n�Ŭ�^�W�:�p�HQ��.���d��Q�1"	�$r8|@֮�%����j��Z� ϪZD�E[`r����N'�{��"ɥ��'�3�a���#����H�^��D&�`�,,r����0I׈��>�+ǰ��iU�ss;�EsI�Y��F���e�jsਁ4� �M�XN�'��Sk'�/�Ehnj������g�'�O�'O.2\(�π3(;l��;�������k�s�@�@�1���<��g�����`�\q���K��A�#u�9 ���!PT��5�
L�p?љ�rU'�ϵdJ+����eF�8��Ld포�DT��|�`�
:�{��r��l�����~"ʒv|�f��Ȁ�����"TL�=%� 	��7+&p�xpTk*ӔW�����@��.�|��rf#��I�)�ENUN����6�����PQx`�n��h��^�4�s���PR����=x���B ЗؗwBܝ�ñg�j��*'=L�������0�P�{�l��@q�W�	6  ��玊oo��Oz+CQ�<��~�`��=c
��9ONf'�Bݙ�?b0�$#9薓�KV�E��y^q���
������F�60��8+���dq��kM ����0Mk�{ %�|"eF*jxCN�f����+��䀻�-� ���x�H0��}t��:z�i���ob�[� �p ����D�,{��׺ڢ�Ju�E@?K=f���
r�*=%_I�4o�E��J=���0}���m�4���n׹G� 	��T� .��>T����}�y�����g|�?<W��;�:����kϳ�H�(���3:]L*Լ���(�S���E�FU��hb���F�Q�������E��ٷ��8w���5��c5��D�m��3�L�qoSde�	r�?��dF!d�}ݵ��,߷��ω҉ 1�0��i���2J0�90Z�F�2�}S=��$@>`�NF'�-+�5�CWL8��8�͜9���ǔRA�><��w��/��*�
��TX1�}r����(��5��V�H�u��$� �o�q$� ��~�m!�w �����o�'@�FJж�b��$�d�C�qMɷ�R,9f�􌢉��f��ܭL}����)0���}�%n��,W���""�?���ެ�l�낙		8e�� J�D�ʐ$�{����|q��˧��g��O��?<����Y׹D���    IEND�B`�PK
     ��ZH��X/  X/  /   images/78e6be4d-468b-4075-9957-5b4cf1a5366b.png�PNG

   IHDR   d   +   ��-�   	pHYs  �  ��+  /
IDATx�M|t]�u�~���^�h�%�Ҳeٲ��ǎm9�J&�̚�&+�x\�JfR�x�8��I�Il�vl9vb�*�(R"E�W�@������{����^	$����{�>{�{�?����{�m�����Vu�F��^:?����+�' h�Ww�i6\s�-�	:<��G�� f�nE�����Aw8����h%D���N�@9W@:��m�xl�c�|#�e����(�vv6 ����`�~�ޅcj�yLx-��4�ip�4���ǋ�� ��{
B�L�}�%�ϰP�[Cc]e�Ab��u�`au�S��3\��AV���V�KEl�r�9����J�s.�C{XܣNq�0��˶�N�_U ks�w�\��_~<�y�j�s������=�}�;{_��_�,�m�\*a������ۺѿk,Q��!�4�F�N����%TtuV=�4��'�h/�� 2E:�r5�,%�`bp �Ǉڰ��+���.]��������]�����C�a.���l��kiT:�B��m���5"K�õ��}����D.�Dkk7xi�K6��,�����.�˕P��`�hE��%��(�ܹY�26�W�Ќe�S�'؈@����L^4O�ht�D!c ���[o ��*��
t��G����PKC�����9X&�����7.�������گ���񠹩������ʥ"���W5]�����a��,>�#��oMH$��?���4n7�H#�u4u	xu�����z
���?}�ٕfJ�|�#A�OGE��ky�>����o���
�E�������~��j��PA�k=�x�����cq	�hf�\�7��I�*����Z���d�k�����7?����)��@.�F����+�nđ�]�X�˷��ь�c��wb|}�_�@2�kъn>�?�g�~��m0��1qg�H���'������f���<t��{���׽��F��.�-�N�(���y)�S��9_���_Bsc;w蠱��������īWR���_�!\bDa���f�h׮�A$l���lpܪ$U|Xq�hj��i{����g�RZ5H$]�ܚo���?�;v���Ml&�ğ|�k��`�0	Y�Kl��|���t�[�?c 7t���d���߭L�{nD��	�X�	����&�gG��EL$���H`�zz�����ճ9@��������g�����{3> xI�}��7���%b�L/���:F3cݽ�4����'h�R��=�{p��7�%�*ܤ���쫗����f �N�bg�N��Ee6��V(T�����6c��?y�fff)>�5�z7��W�D�Q�~�o���]BA�3�xh��b�Et-��YL����Q|�/A����߇bN6_�2k��=��u�t�|�{�Z0�]A�2|o̰l&I��h̅xǧ�����$�`���9�?��w���	��)BM�D2Qd�0�{������5Ģ^�b}inQ/�q��U�J$X�߃7���7F�w����8xv�5��^;	��\L1�p��`�2�>�������H|��u�x�&-�a�Ӹܜ!�r���
���!֫;X[[��� ��E�NI@�)�:B|��D`|��8��x"�'���&�y�>�w/�����9ъ��n�q7^��-,�6O�.��|M�GH�(��s�)d�S��!���U����xhRM���sE|���vB�k�k(������!����Tx��T��2�`��?t��#�����v�'�ƣgG��	Ȗ��m��A���c�@�W2(�ʸr�N�����
n��hd��G��r|�3�����Q�=��[G��(�HԈ�^Fs�\b�q�Oʖ|hlj��[70;;�B�?�\4B���~ⱏ�}�m{��?�v���;����tf��� bZ{�k�`�-�]=����R�W�x�Ã8-����Y$	�R��;b�Z�I�r蕊�VKd����Y�w
>��N!j�l�L*C�Q�6ȗ~
�d&I'j�73u|I��lT�`����!�̡�1�L�n���A�!�����7�o��~�dYķ�-�QϠS���_g�Ma��	.��ح;�:�0o�X�}��R[iF�*��0��H'�X�0
��*dpt�)�M!���XTe��I=���,μ�����8�b�"�]B(`c���/=��� 򄮷=����4#qm���Ja�,m�@	edL$:����������X��hh��t���BW,I���B�wk�CS�
�d�i��d�LT!X@�Nu5�K�r�8\/�0��-��>f�6�g?�M��m=�s{������x��;8��+�����˦7�ԉ��%x#l����A.��k��/�i_ ]$�k4@������K;Ig��N9�e�����9uj
�P�rfй������G�O,��w���@��>��ˈ�hdl �bm��ao�H&ᦸA�B e	¦�2�M���Jg�6k	t4�w�I|�_`}e��+
BY�X��6.�R&D��4b�5��}���2zE�4y;O����zWtY5쪐$�����5Z5��#�*�����{�TV/%���I8%Se���F�]���M���������d�t���rv�-^|�S�O$�W� ��D*�Ask+��ߐ�ڂ������ ��6�~�����y|��#��՘�%�z8E"�D�Z�<��=�_�@�FH�N���"���H	�m��F�0Y!�ym������'zB�p��"�h$�SeIZ������wu$K8v�O����a"P�\S�s�#t�8�(CS�K�����)B6\M�Q�F��UE*�jD�'����Ocvf��oay~�B9"��`�Zny4�L���t�Ϟ?���[�>n�6v��1��%|�C�cGv�����S�����s籶����������/��;X_^���C6��ܦ#,<�'QϺ��#an.����(QΧ����RYU+���:�}_+b�w0s�*А ��94z�hb�V��:7���J�I]����<�9~�Pq;%J�עpe��A��c���ԭ����Hg����f4L]e����h!��NQ��ȯ�����T]p�E_5�����\�̚;���|�K�+�U)�f�fZ�3S'�y��F���>����,2�ė���{�z'Lm����ӋKo^DCS#F�C6�ơp⥗��y1[-�B�R���S�F,.�7>�(~��8�V|~���	d6f��O�Z������i#��g[�ǺS�#KB<��NB���Fq�^-Ĭ3T�u�m
��Prl�w�UI[�e�j�.�;�	������mW��V-TA�T�@�~�K�Ш����J3p�E�a�ܝ^��"Lf�MM"�]�p��I<~�8����dpeU�u�bӨ2�"i����	�QĂШK��Q��ۂ�|��H0P��:�J�нs'B� vt�ӛ�
FT�vvv��'���D=k�]�12ԂC����$S$-������cA�Q(l�X�<���A�N8����a��A�e�\E�I98���V�1id��+�h�0��=�U1�:�{�J��̐
|�XjC[�)�E���IqW��U�<��H�)MzLiFl�6��3���|=��!�_i��KD���y��{7���q"�ĩU�v3S3� 48�_�0���Q�꛰����fG���~H���"��;(����$X{��u"��Ǚ3�����K�/�c�~�^����1SD����bɪ�I����]�8uq]5�4We	���8"�~����Ҥ,Q���ċY*���.�+��g�p
��~2�f��t
�4����"M�M�*�^byLI����^����\�� nMQ��=R��i.E�νf3�9�Я{���*K\�T��wHd�٩f�����YE]w�����ɚ�[:���}gg�J2A��/0�Ө�k���,U횛[Tk����2pw�3��9�i"4��sJĺ|��o�.��������ǽIF����(樴���F����K-�Ngc����RD��KEGg�a&/�ٖS�B�h�P�����	�b�J}k�Vv)8f��	�tD@�x��7 ��R"�b1�Tw���!D0��g������(��ڟS-:�z��/�Tq��I9�Q�����.:�Y�h�mۤ�������b)�;H|hPj4|Tyo{{:v��xf��;Q_߀{�>ass���ލ+W.����ds�n�SF/��ek�Ԕ�Qf�J/*K�EIoו@ljh������c�߂�o�E4�������lJ�����#3��	�D���_GT��(�Rd��,�.k��b]a�;ef�67�B|��1�t�z�
��+=*�"dY!�0�9U���t� aC5*c�����#���ҫ��ba�t��Z�Ʌ�D���x�j@J]�*�!��`�9��2kA���Ύ��O�ڬbL�)}��ưo�~��ݽ3�����9Ҹï���1�B�Hf#�� ����v��Uu
9==�9���� ��6�{���p��yzz���$q1����M�=�'�ebam�Z�$�����̒,)t��^ Gj��
1��+X�lR����.6�6��mx����@�z��(�^�@q�F�0����ku���1ᛛ(�2
>F�M�ڥa�S��ҩ�XU�s���ᕂ�U�.mC1 QVQ�R=_+��u���qYrI4�G��ފ��5x�:eBV�j;�b�R0Ub����",���!��������#_�c��u��!����_��t
ji�>rǎ=�����q��x��̒�����X\�G��,B�+,f���굹ZCV*5i���S	�S�ʅ(	)^�.��ѫ��h�7!5G���!�����;H�}XN���� ���fk�|�r):ӻ��c\?3��� �#�U���鵦��Fa�P%�:B��ڴ
���=X�#����k�Ȱ�ttv+C%SI���f��BI�C�v���b{��:ݎ�SZ$���#��a��L���I�n�6�����3L�(�]G贈�tH8���Q$i�}JV�6a����Ԍ��_�q�;Κ�@�kV|����C�U�JF��7p��L�-���+�"���716�w�{�N����y�_��0J˅�bm���Aj�k���#_�ⵛ�������oaF�h=�N
���q�5|�D�P+��W����YT�Xo�A�u-Έ|�a��?���Nn��g���޿���ۯ~_��p��|�_�	��'?�	����'�_�����7�?�=ܼq?=�F�B+��ǨꍨS�S$ư��Jt��_Y�d���ޮNCB�N�<A��ѮM�=���D������0�%���0KE[	y�7���7��܊=C�=�H�GZ FU�JѓtԘ֯�|�T�YZ\Rٲ���o��e2d%^K�hP��������Z2��F24o�s��yk���z'ٜ�����c%4���Fc�N�������j��j=���Wl���!L��v'��V���T<���M����E|��x�(�f{�ܾ5���:���g�������?|�m؈o)�C(��(����$��*U�.�*�PH�+(�BT=^��8w�"�= nRY#P�IgԙL__/nݺş�x�cd�o���lꤝ�D�ѕD�%8������ab�aJ1����)�4�6Q=�*�71��cǎ$X���Il��B[BdX��D
�d�i�ais��&��5ǌ�Z(�&QҖQ���@d=ٽx���|k?F'���aᵻK�e&��BB^թ��fBSm-QxX��z[qst
+i9��Ż�h�YŲ�{����;��,����C�c@��$���`ûѹ���b��ј����:Fo�3�4u,�F)�Yd~Eah�Ճcz0:v���4~��UH#��P�|_�GM0�S�mu,�ЧŢ�6�U2 �ߋqO
_|����p�}Y�õc\M5
ų�ߡÇ�g�]�o��^����k�>��afSy�lo��g�U�2������&���b}�߁ŕ��q��D��\����h�l��sױ����+v��aF_�FaZC���!!8��5��E����`!W�\2���Fv��8�,]�o~2����XA��Y �X�/�8�Q��+X^_c-l��l3T���7�g/]�X���� �a(����+�5�o�,)�I�Sgy�ӯ�����!�w�VA������i��~�?���&�>���53;�XK�f2.�ŀ�������FV/���J��/%�%�H1+��G.]���\���x�-}|]�x�����}�#G(��{K�X�Z#��0�ll�dr�Hl�H�3�l��d����%�%�Ҁ�ES]��;��G�@/����yDvt��zC!��kkq�շ��G?H͔�W��m֖f|�?¥��X�*��7���s�\�s��3�Q�l̃�^>��	��yp��k��[c@d	I%R�,�Û篓�g��Ԏ��4�J~U�SJH�z���<^<����G	M��_�f~ы�}=z��������ǎ]�����ֳ��e%^dlF�/�r��mܸ}�\�\[S�9��R�v"�ٙE,,-a�Τ�� �w��hi	F|3�䧔����#�����p�)FN�I�L��1D|�Eֶ���^�2�MfP0AoO;�O�M�'zXX����Ќ[�����,�z�P�5���1¢O�>����q�/<�
�W'�8s�Ml�/#!������k�cvq�onRP���Z\�cV-S �#OR���Il�khD�^G��PL�h#�����d�	��#T��à�˭N�H}�����渹��.˫I2��	fÐ�l1�m((���� [HˡCEġ��K�"-��]"d-Q��3}]s[_�e�d�پ�tr�T�Q��Onϧ�Y�;Bah&��m�jj���#T��t�<d6���F�|��dO+�9,1;���(]:�cz��\�ƽsS�$u!ս`v��`�y���IA&���d6d��2�}{������8�Fh�D3+^��ĤD�˔1��B{,B���a�4@WW���݇��V�{C�~��u��ȗd�8�>�����N��թ.y��\�%T{iq�k��s*19���7�F�~.fS�Q�,���C|^�Ir0%�O®$�2��{��K'���ϛT���8�F�&O׶,��QA����;S�o�������)Rm.L"�B|��냱����T�9L�l�¬��Vr�����U�\[�H}E;���2B�zUJ&�i?,�*�~��v��g�����w��]Y��}�D�y�07����}���ޚ�3O?���M��^���C&'g��\�o�Hll!��d`F�ILM����s�7����*�PvL�d_s��<	䮡���XsC�f�
G�`l��	D��K�tL7ɋ�Tp��nu��$e��}�bQ��N2��`�d����o
ֈ�!
�!\�8Ͽ(0��މ�j�=���$��:[�g�x����y̋���h��lfP4Peߞ�ŶI1G($M���`b^q�i�!C
�t�����i�Bg��ӵ<��>���A��O�|u���Cx������09�˗��9��\����YO���W�6w�I�1p�ߗ�Q�=�m�P1s���j�h�J<�c0�n*���[
Y�>q��#K6&�H֝m����y��;b=��_��khO$���}cU�Wl��QB�`l#/0
9-ӫ�srV����N`j�l
??�IW�}�`���y��A��]�0����Z�|�lޕ��仗W$}��3�+�qն�q#��(:q���,��X����a��Y\e���T��ƈ�6'c�!,�e�<�@evnA��E�@S�� �ݍ I�'��G)�9���Oa�zd7�jF���鴁O��Y̑t�ͳ�{��^rZ)�;c�Um�=L�WP$�K�2J*+�4H��OZ� ��c���oavy�?���~�܌珛n�N�H ��$E*A�~��xMeF8U)�>dɛS�M�����SSrEb�&6Dѳ��ؖ- 5x��Us�]�q�>C��%�qr��[��_�W�����Es�$�5�J������QM�mV�`�9z{�#�{x?��ȼ���mZ/���	���$�7!��$N�Q�SSm��˓et�0O�;�i��v�:�"KA(��D���_��L��`z|����V�w��O؟�Vu��u���Qu{}�R�oQ�kk[�x�
Ƨ��������O��GsgWׇ�ݑ�e��;y�ߘV*T���B��?�����}{�byn��e�1L���PS�@ghj�E����;8����"�c��p�C{�gZk�жjU�������US�%��k�*�c���0v?r�#m��A�j2�KH�F���Z�����"i3�[���C�~n��Pl�X����Y����6�=U��t�9�{��v�e���ۄ.�ڡ �ˉ��3HRf��fjYM�L�$��v&H�6ˀM����	�]4PĶ�5q�\%����}�5���/�jڣRϚ��L���]M�gzB��H�5��ԩ�MM���>���a|��_���g�g�El96��,�UN޼�	@a_��$p�n���{.�M~ST�3��ڦ�K�A�d�VR��'޺�� ^~�u�u<v�8�I�Ͼ�3f�k�&�NUl�!9U�v�%��V55o�)��p�W_P�-�u!���xuu�dː��WP�T��%����k�O$+��7o��V�B@��2z!�.l%����}�W�0-Pu����;���I���k5);�odI2�`̕S�:"�N���n�Y�.�=Ї��"�T�=��~�E���A�~���NI����YuX��¤yr4I�z���~m�Ʃ�Mx}r~�4g�F �G?�Q�u+`�P��C��:iT�	S�����e�*�h�jr,�֠)�-���9����8SW�d2�X\à~mMLz��mAfh9E��,�y�[;'մ���J�#^������|�d��pWn�a-�t$��}|�����be=�r�(���D�����Jږ �[8px/�\%�#5�����,>�k�U�:�e���n�`�9
��XNu([�7$��r�Q�s���\Rby<�R�0z˸3��
E�iQ�҈Je	3f=�^D�a�t!���E6=D��Ԧ��];[�hg�����PP9��ܩ	�|
���+5�kշ�p�z-�38ֺ{��"bb(�M˧OM G�����o�N�˹�Z��(S�x�ɇIL����دm��j�5�!�w�A� v���f�L������'�?�Ҷf�������2>���qwl��#Gѳ��|)�PF�[�Vn�� �֣qk�1�jF��éh��d�ɭ��JRJ�M���L�6���#���C���W�(��d
j"D��I�yt�Ɵk�lm��6��2��)�:%˳�,9�2���5Q�c����*�;��F:?<� ��
�� �^��:�N���5� �&�n�}�r��`�:>��g��NS���u�B�9Ћ5J{g=�n묝sSq:4����c�d�9��؍"�ˢ$��1=��G���8d�NL;X\����ӥ���k�q�e5=�)w%8e�U��Tj��UQ+�
0*�1��u�����������r��g��Vm(M��E�0sB�1�GM��^�r�c���#�Kn��)����Y�yHg}aюLAf6PI���l�G��m7�bp�!4D<��N�����ޕ�3)C��LJ�˓ �3�����/���l�vKJ\������/ߢ�iC'���+��_^�v�%�y�in��s�3x��>8����J��V#����%����ױ����M���� �����h�Lx<�~_P�������
F���8m����ƍI<��1��ѯR�(^��!u��W�W�O!_��1�qА��H�	y5 �QQ��
y�M����j^J�5�jj
�(����vY��������f0�׃������˸�/�-����?����}{�z�&I��^�1�lӤ^��A�'�G�ś��[F����\E����8��݇:�Jh����7����O~�WFz��(t��I&�]䅼�r��~u�hH>O5�5�bT��$��[=��W�c�{d���0uDK���؉�v+kH��u,��ѷ�~L/na�p�_zBB��Tk�ZX�5��[��4և0��S��%<��2���@��A��^��Q؀���鉢�lt�]�F��D�)ݲ*�q�!��4h�,�0r�8�BaG�|����dm-d�byq����'��zc��5"�n �\Dfk�6��Bj[�H�h���
v75��?xJ2XG�;������L���/�$��T���S'�ce�} ���J������|�MST�pSO���P�m��țz0G��g!.����G���c�~ܼq�~����&]��Q�
E�j7n�V�2G��w�l3��	nN�o��꽲�q<��r[eo�����.R�$���Q�C���)�A�_�ɴe�CB!�L�z��x���.Z��ۍq�,�[�h =#�XX��LȰ�О.~�������֥��ئ��� Ԫ����{(������3+�r��5d�������?�Ᏹ��lm�⾣ǪjX1$�FO]�1$]ת���	U�j���,�Ț�ʖ������h��¢�ň���$FG��!�g�<Qʒ(0��,K���]�hk���B���:��
���$����{�Ϋ�n�
�����h�#h]=m[}L@�2��W��Q}�ǱM��.#�������1��F���50�@���#p��,*�C]斩7T)3|�ݏݴ��}���x駯�Lfʝj}TO0�����$I��x����"�Xoa}^�dڌ������D���]bMZ�]M���85��V�V}�̱UKYZ-��7PC(V������9$W2���E-5}�-$72�~{���II�m5���r-K+[d%M��k���󞎘zش	s��<�T̬q�[��������(�-���e9J�Ȁ�Y+ʲ�LY跆F֖�;5lΟ��b�҅l��;�@̋fR�8��P��yA\�6�'���v�3��jFKTx�{����W�e&WD>[@�賣�E����8�̱��Z�����ځp4�j;�qRy����r��h�$5Z�4��N���^�4j"�9�/�֋�2��;=WA^��xў�j�IrY�����
�>�$]{���T�Q�Q����+(�*�$����F�x�d��ҡ��y�٣�Ac[j`���H����2f�F�)G�U�4"�k�}Ymu�'�>$��xc�@#�O��"��Ki��/����#DgޜDYoP����*z���@>'�u�[��^�_0�c֓�F����?�Ν���	o��0���*�^�/�!2WyZ�>	�M�Q��QU��skOw��G�4EF�ezPf�t��Md?�Ψtt�h�z�Veb�q)�r	���lI��%��Z�D��<��������{��$GEŠX�P*�� ����<��CE�B���%���W5�d(��>oΈ�J��	J@���3���7-��TXÏ�����/��g�x�n�\����:��NF�ky���U�u�ɓ�PF�1�6d�m�3'�[k�9C�e���݈g�}ssm�����y�mG�qyF�)�Q��e�4[Ȫ�E��0C��e�6���iAM�h^5�%PUR��75�o茸|Q�k��b�#�c���¶:$:+�*�t�Yf�Ꮳx��"ܸe�	y�4�Ϋ�v�ٕc��(�/�xO�.�I���ګf�,�=HG3��85�/IH��:@��'Ȥu/MBy�R����ZM?��2�9�Y}TC���5��������_�v���� a�E"������Z��1�    IEND�B`�PK
     ��Z���y �  � /   images/483af35d-09f4-402a-a8a9-75c28eb4643f.png�PNG

   IHDR   �     ��   	pHYs  �  ��+  ��IDATx��w�$Wu/���Nw��LΚi���	� �D�/&0�,��D��3H$s1&^[`I(�<#��h49ϙ�S�X᭵v��:G2����}���OG=]]a��+�V� Nm��SN1©�ԆS�pj;��v�Nm�6�b�S۩M�S�pj;��#��Nm��������X,vX��hoo���vj��h{I�������\���f`E$��d�O�q�����97��������yɶD&`b�Fmd��g�4�<bsv�:hY�p:�
�jV'1B��i"R�7\:��Ct,�F�!���C�à?��L��~�}�m�!��8F(p�@ h�5,>�ϭ�kq�0L>6Xs��}_�z6�Ou<`�c��`��e4l#	���Sl�5��׶�1-W��,�~ðL������U��]�n!����q��+��`����a�>��I��㥉�;��r]��Ԣ�hrj|���yn���8�k��D�7y�|=ȳ���8����0o��Թn��,���:����l�k�u�{Y��<�$;�`0$���<u,��4�p#�h�*��`�Qjkk�x7�ct1/��$F�Iq��Rn�P�6V����E���2���{/���k�ɢ�(�JGoo����&'ݶ���ޟ����GG'���H��¸LyA[QO�˟�k�|Mޯ&N�^�j��5���3l�Bp���f�q�k荎�����w�i���oD����B�o�����o�O_G�W_����wZ-�Ҽ��;]��b���Y�^�:�>�Ͽ߻Q�#����\���x��__�7��)��=Gz���{�q$T�[��l�|������@8 u�"x��XV-�N�3�%���lvvz||�˽����l/�j+5�+��.kK��j�j�Ρ㊱h�j�H��r�Z�B�c��cӍ�*5{C�QR�VkЂTE�j��dY�exg�~�|�f���S/�^p���wM�r�Z��#�&�V�q=0o3��Fc��q
��$�-Z(Z3˦�[��b� }Zj�A�I�rq���_�>�M�|v��1��$Z!�ou}��@«y�&f3�Ʋ���q5C8�֫��i�Al�.��Þ�2<f�+,,%�Z��f�;����x̪��Ա<�ǐ�q�(��δ�ggg�t��'#��c|b�lV��%��v���;:}I��%����o�b�v�p4v�α+�	�J�@v.;{���\��?94�z�x^���4�J��VM&�/�Xh	,ߵ��'y��K3M�~���筂�ۃ`��7�X��kI�iZ������ٶ�r�,תT�1#���c������l���W[����Ӝs�\�CE�����Z�&c�k�ǭ�9�.3�-�ǟ~���T���4��������5��>����+D�1��M�������&��ݍr�*�����Qs>D�~���ӗ�$��C�p�n^+�]����B�ģ�
a$�IY2��]����l?9��x<�A����P0�XT-�V�JRM	 ���X/��P�B��B���JK���V��c��w=�yտCU��\tM �(�H�9f&.VF�hB~ӰI?o�y�Wi"�s���y�a��H~Z$)�������<�-f�ĥ kA��<.�������ӵꮂ(��¡�\Wω&P?LS�B�yԳ�5������95S��U��R�D�R���N��5LMM#�a|2�d:ðI����t�$�_|�y|I��h�i.�9�&$ְ;�U{�sX��bDԄ��t�|�m���;[(.��oظj�i+�.]��H��l�D���s$A�9�!�+Q�b4U�o2��V���K=uO�Hu�<��P6�Cf+߇G_WKX&}O�L&��l	��p#̗�M�gs$����zZzj��X���sX�c)���������u���<8���\3������5����g�c������fz�h�@���*�z{:q�]wbÆӱz�*���?���I{��z�����@�%H����h�Yv�7�=�B�LO�dx��p333����Y�o��O2>'^�z��6��Y"����$H��E��PM��[�r�Ak�<�� �"�	M�*�uL�zfs��/�[��x�^4&D}m^�Z-҄�u� �X��k�i����?6�h�m����3=&aL��w4�i���7�'&&ۂ-�i��|>�m_:�Ʈ��m��<��P��i;�mBD��rL����(�u��8���cn� P4���m/��ĉ����#�af:�u�6��Fv�f�֨'j5{�~ϳ��8�cd����$��u��ܽ{���m{�����w��?]�jkCgg'��
"AV�!�J�;:I���!����d{���e�fg�x�[\!�P��؊p�x;��Z�ʿY���LMl�W������Pڠ4%�|w�������� ;�!�5&���)f���Y��C��Aj��4JI_�cG��ָ|W���>NIJ5,�߼)�C��8y�k�d�Mk)ŠaW�PD<� ��#�jC�\��Wk�[�)��]%ٙ�z�5��J3�|G�|���ѯx�s�>f >��H�X�2�"r��9�b�E�i|�FNҳ�=V'o�x��.����K�F��MKv�M��b�S�g>���k������k������'_�_���?-�;Эz� �u��q�*�,إ����"�/`rr3"�&��u�@�I�s��1��S��I�J����C�����m|6K��`xD��E�Z���´P�t�A�B�D���H{�D���tN��n�X����f��}���gf���g���y�h�Kt/� "�~L�RQ����j�r����8~�6T���H�g����,i���Lcl�3�q����0CZ�O�Z;���^'��C������חǧ4U�j�	���x<J�WA4C�l�J��d"����ֳ6�<��o�b����G�b�R�6�}ct��x;_#��I[#>4t<�G�������믿~bpp�n�{����o��w�}%���D�Bx�E�f�rC��uwwav&'��vL��e2�Y��	����LZC�P�a8�c����}+|Nԃ@���i2�i<Gby*o�v��_���;���� Ē�%�	���pD3�05�����a�2#����HX	x��v�2C(��[X��ƞ#�f�oKܟ�x�3p�9��6z����0+�"�#e�/�����OZH�>-LX�ɜ0cx���m4Y����V�6���F1#E
�&�#��@0�ϠE0��Q%fh��K�-FtG&'����QSL���j�8��1�G�@��j4j1RI���i�OHj�`A�e���=g���L�/������5AFCaeȑ�+�K�H������Fc'��h��i��F ���v��P��5[��_k�̛��ބ�C*(�%U��iW��Wf�9���X�o��� {��+6�4�~|���JR���P�G�5.O3�~�C� �m[���=��r�9�.m��fP`���������7k3M�L4̸��<���}o?{������3���<HY-/��j|�P���a��"@�� o�Z���ڕO�V"�M�e�UEp2Cz���V�0N�n����U�N��z'2�?b�P8�Eo���MBCT���$��*";=g,ʋ0��Gǔ��1��pH
F��BDh�"�x�,eb�0jD(!�V��<6A�3^=�V�IU�1��{ h����~�TA�\���D�:M�1M�f���f m\�1�x�Ɉ��@�f�T�oM� �&IG4�����&�,��qkX�s�g���D��
R�渥�^M��S��ӛ��{����F���uRm����x�xc��qm{(�V�h�F&�A��q��1�LG���!��+�mDP��1o��h�%1�����B!�b)/���:�ce��TVvjR$G{{�TW�&���=��xBl�*��yƧ��Aꢾá�<`<�SI!5y�8Bh��d2���x���L�$�4	��-��C�y�K-���F��^��9?���c��ƚA/�b���s�O?���9?=B�U���,&�g��֨c����T }���q*�|C��7��4�j7�f*��B- cc�� -��{�K�3�Æ�?�6�h��)֜'�����g�C0��CU�C�u"��]]]��AC�pؾ3#�\N�>�?b�`Ш���ݝ���٫���a�������8��ޓ�Ɍ��{���C���(6n��իqrhT�S�� \k�>a���0��NM0D�:\b\����������cYc�n�%���?xq�A-Ʈ���2j�[����ox6��_e����C�М�G��I>�k�������H8^j���>?7�D�2.�*����B�4�Ӱ���$4F!&"	�A/O��F@��7��*�3<�.'4����u$���6�ک���-��|(�7ȟ�-R�a��R?�T��6�0�QUl�n�mČ���3$Ї�Y�*��T�}����Z	�x'1m��a�>/m�FYq��ař4��,�uarz�.q�N�1]�"�'+>�<���d�s�M�A1XS�O��p5�$Y��P��G	^�g\��M�5��֟����x���{'4�ϚZ�)����nIf ��r[ƣ
ұ���#!P��ݝ6G������ݟ�HL��F ;*֎����ۼ�+�1
�z��W�uf��F5Ķ�?��v��ӷ�����i���'%q�
�(� C�^�d�%��`
J̅ݐ�)���
������_�x��7����̘�Y��wH�s�[X��X<*ЖI ������Q����m�� ��=�I��>J���1�/���^s�5g�"�R)"BK M�+۰���0��R�&E��E���w�(�gہV\�f4@���B4�P�^���~n�[��:�G���6�m��C�%�o;軆�+��c�b����
+Bq\�QH2!�^�4��T2e���}{�R��T4K��G����(��z���0a2��E��͏PP�E�J-4?��Z��:c�_9B*Y�t[�p�Mp���r	���b�C,��i˧A��mbt:O�ff��@3����F���� ����O��XL�!x̜�H�-����h9kT� ѥbs��bV��(mDw�E[$,i1-xj�������3�\cE6�g2���'F���߿ehh�6����	d҄�"	���p�a˖-xꩧ�裏�-]�(�g�Ɓ�R������wq^��j���] �7���H���Y=�ju�`v[�����4m�;��Z9=,kndVѐ��]%���t1����=Z�c��I����h?�y�bZ�*IQ�!
(h��<�&-Gu\�����x�0*�9�='��������$q�Dᠫ�N�._ǐ�=4�MĨ��Y����g@>d���i�|��7
���	���;��_�ZI�*ө�`�5DS0�1��a(f��&td��y�%�t�o|=N�ґm�mrݨ�Y<�g���L�sp �aՐI��h�1��$V�J��e�@0`��$n�(Fص���/�+�-]A7(�Ò����T'��=�O~�Sؼ�L�^��S؜�dx��D*�42��<�N��%�0>>#��1�y�	˃4����"�,RE�f��^x��o�)fQx\�9R�좕�e"r�z;Z)���b��U�V2[L���13�^¹�~&͸B����u�M7�Z�PX�UZ��q����8F+�s��4�xD?ߛ��	�a��,�s��kHiC�^N����k�1����Dˈ	����n��`ۆ��iz�Խ��fгOC���lMª5
���șY��sn�Fv�*4� ~��l=�<���M���j����0B&�\���|�����O
����T�6$&.��2�����r���_K���'�@�--�ʊy8�<K�i��_�����4�.N��W�m4�%9��dh�n�V��Nؚ���'~��N��0ǋ�$7��]���I_W_s~bG��{����R3��K�c��/��������
[TD����kzLR��9���\��JJ�5[q	���ݭ��L�q�y��8�|ҡ�>z~x���n��I�R�����D���]�!�ʹ@vf>g`ft���6u�wHC>�Ł�H�H��p87��E3���'N��s�����sχM�-E��V*"Bk��ٝxr����e�1�߇e����C)�E*��]����F���E��i�w�~1�882���� �����$�GM�b+�Hzc��>n��=~B��V�n� ��F�j0k4�����DZ{n[ۓ�b�и��zQ7i%����?ٛ��O�����+�P��Wl}���q��q�����>N�"G�HAI�6Ļ#� ������⍓ySF4�s:L`�
Ni|&CF��Ő�]�|g�f5]֘c#�)U䣜�D͔���g���%8'F�_��u�Y�Zg	X�5K�*��::��q����c"�fu�x�2Tr����Z�/���
=��W&Ӂ����ghݺ�Ж��g���|�#�;�p��݋�G����W�{��A�TA �|� M����gf�k�H$Q��Q�k�)�|]��~�:O�
�(�Q���DU������$�@#�pV>L��"�����ؓ���61���ݷ�`��>m^p�=���؋�?�3��=ߏ	KQ��B�����JL�<���d�����L;��}�1!��㗔�������g���}��`�F�y?Eˮ��ul���y����=�&#h�Y�<F�A�'� z�*�C�=�1�X<����g3L�aɒ%81|v��e˖���AW��@m(u*I:=��avv�cccK6o܂�C#����'��a�_�ĈrH�k���dO�B6���cp�+�����S��s958����XB��
/h�Par�;�������r}��J�Gʥ��1D�j�O�$�J�������\@M�i
��dφ�#4>��\Wζ�
�5]>�ƌ���Ee8�s��:M�/�C�g,�b3Opp��n�'�1�R+4�wd���w'����GTsa��Hڄ��	��!lȧU�I�!��3~�x�]�5}��N�8��8����w�ms�w������B5Mmcy����L"�bQ�c�q�J{�mZ+��++rX00�Z�"i��t���z�r�/�fff�G���%�F9rL�𑃄���կ���������m�܌a��e�p֖3E��u�V��-o�w��=|�?����.	��I�D�0�45�Q�t2ĩ�pǚ�!�����J�c�2R.;�P^a���L�Z5�䳺�H�AЛ@�G0��܂ڝ�!N�3���jԚ��)��}�Y��7���h~f����ԜC%�C�ܶ����A+��ߕg�h��!���ǩ��|�t�]��b�x�U9�J��sz�?ݚ���s���y�	��<h�Z:w˜��<�;t�Fпk�d�ji{����N�ãY��B	�2A�A�ڮF�ua�J`�X�]]8y������$-r>��QF�V�s���z�[��i�tJP�o^/�BV�BFrA�;w������"��!�=����Utu�B�"	x���HT�~x�nYJ��1�v+WJH����%�;�s�5��:����uẖ�ĩ��y��ҒV�KM�M��W��i��&0]R��WD_��hEo�u9@ٍJ�T�Uތ>׏���~CٟL�\@�vd,��~v3��Cjl�8ʎ�OE���̉n��fW�N��Y�z>���L�p��7����u�hUй^��_��g�o�l�3Dk����*���c����qn}.���*5==}:|ScØ����݅�L�>��W����d's�T:�C��-#���{�=�)�K̀r|Cz]p�Eb+��m��n�5v�? ���5kp��1����u��z�:\y�k������ą$�{,Pހ@T�&WJ�J�D�u���\�D��pA>1Qq>��Ҳ[.QU�ɑ[��T� ���\��7�9�Oe-����(CrY�K��5��:7��	n�I��X����#B�@Ur�bM����M��{6�ϒU6<������G���!��������'���xSWnܠ���ꛃf3W�sɔ�Li_a[14�2��-$���gݑJ7�.��M2
vN�3��V쮭��qXwmK	۩��(M�1�T/	�Pp��ք�|	��$킑�?�1|��� hx�{q����g��7���=>��0��^�Q,�I���듭�E��"�v����bxǻ�-��^���}Hc��ߏ��i�"� }&ہ?Šr�hSІ7�C�q�&����b��b)_I�&U���3���{ß�_GR��b�iK��m2�����	_l�a�S����"|Hp�e�:S%�lK>>����x�\�60���^\,�ثRv��ݞ#���Ɯ��g��Y�s�Fs�s`�$��4�fL��j6���
��r{�Ze��Q�]#�u��L.ѭ�&*�9�~B��+Bvdm�v�a.��x��+�Ш+OS,�@�%�T�����`4�4M�~�`l��=w܊bvV�t<̉��L�,*��r3$d�$����v�E3B>;�'d��,� ��F��9�ozz���"�(I���nK.�#�ټH�%��I@M��l��"�1.���B�OB�/�2�;
���E�V�l_[Zx�e`<�33�b{�����^
�п��3�9���n������7J�����~<s�hٴ��q���K���q�X�����pp��D?�p�1R�Ѐ�Mb,/�
�����:��/���V��Bk�ϩ��(x���D(FЏ u��S�ǌ"-��L�
C#�t�ܺ��@���"��C���EѪ$D��8�U˖$����Y�w&�*"N�W�Ob��q���sLJ��3&|�]���������Uv{{���ѣ$��]�L�!�HFd�(6��=C$��o4;3#����KF��e���Nhk㜥�MJ
(o���sB�B�lXs[�`X�:��t��gcV:*Jͱ�Te�*��D���a�ƨ�3&d1f�槮SD��l~@����]+�\�8��K�g�tW<]�0�6!����d=m<k��^%�6��/�7S�Y���H8�@�Ag7��g/���+��:��I�jC��]E$A� NUJ�:A�^2h�hZr�0"n�V�6�`LRl*����/$�����������=��3����fI@�X�2�	��!N�T������=t�333��	�������&���)h���+���p�lFl��B>�܍�+.{Y���q���:͑*�!�����Uz��(�D�*�WI	GJ6�s�/�HR�UT�@��������
*AJA=��Zy!xf��ݳ��mF�%��l�kѭS�n! �Ū��F���[ƧOr�k L��(�̂E�0�kpI��4��;!��U=�:;��E�X�;�5�</��-zbg�pakD8���hn���t�|�.^��L�%,���t&U�����K�b畫�
�g�M)5���l'7�E�i��v]�TxF'}Ka�4���R��:�}����Ę	H�8aî������6CR�abb
Ufb�EP����}�c45��)k��ىR�Jq*�DOw����#�[`I�jQ�yp�� )��_c|�8+�5��u�U١�jL���^w����_�ݕ�8ǥ��Y��t��?u���wp<���z�u�"ټ��������K�Z�%)=��wf8�7����m)�ӕdry����RϟO#�G�=6�z3D�ᵒd�-�@�k$0E\��ż�1[L���$�M��ɀM�t
�]�O�#�ީ<���CD�1b `&7�R!(~~�-K��IFo,VU1n�`*[�Zq��ա{p��*3`"��)%���'/#���������kňΒ>q����t��2������|��z����y��4�<6n�(j��'�	���5��m�S���	�n�r����y;r;��&�Ժ�J:��y���/�㨌Mv�2��y:^�!�&T-�Il Լ���~���*"��g�R�Ѵ7I�g��Y*� ^�qԩ�"�`���f��[�2G���)q���ۘ�J5Tn0�C�������6��e��9-�Oxsr��VT�4$�D�'W*-�vnL��������@o���e�b�3nO�����EjrRփ#$�H�ۗ�L���i��d�q�vlK�%e�=�:n���`��	�H3\�����{��e$�!&؉b5ӝ4��4����ZwOO�N���[��d�%������b��T��-Q�lToL!8K%Iq�yg�B,Z<�P��מ��gw�Ӭhy:�ĩ%��V����_��w�b��jh��|���m���A�Y�KX�<�������շȝp�0����Noܥ�m ��3Zu�Z�h&��P�~-�t�?�)�B�9�tvc���6�^/#`���3i
-ԥk��N�KR���Ud��b&;����	z��%��KtnI��b��.١d�W�"���W+%�?�]̀�Uox�c�<쁫��+i ����q�e�4K���a��d�S3{p�	��t��ӡ�9�p���굫�8�=�M��z�Dj���$��X*�_"��9�*�Br*P�\��34%�,�����Ҩ�me�j/�^l}�?1k�������R�)�і7�:�Zo���y�G:I���y�Kh�&^��BLe��i�V��;�Y�A����-;��D�R]3�4_��;���cޤ5}8�j�]����b�T�;��ػ�k�ז6�A�S�D	�03S���)2�j(�|�]�b$����<K�ʢ��R�P��p�Y4�}�j��]G9K���tV��I΂�-�3�����#�N�����/ˠX��^���zUx=���.:7E�ab���G�m�)ds��$����aq}j��Z=)ŵ�eqLX��4SRX�kہ��zӝ�k���T�h0*u�\Y�����q����wq6}��1G���-�s�v�i2�_���4�K�O�6<�a;E���.�F��r��c�,.U��P� �<�Qu���W�ɐ��n�2�jS;H�'�u ��[A�5����1�{ԑ[�=0MFbc����]�[RCB�R�D,T�6�	����{�h'��� v������4�d��6-A�+�j�M�=��	��dN�<�QD�i�f�VT~[ݩ�{`)�|��%&^y�%����ĶǱ��1\r� �^��z=R��?���s�=��i"��DrU��<�֋WdB�m�&.���ԙV+�P?�TI���H|m&M0*b�Iq�Ǐ�^p�E��,�$�w�0��4_�"�?�r����̇%M�sU��|���+i
^Vf3�Xܥs;Yh2u0�K�����J��443t�1�v�[��>n+G����8ݴXK����>?��D'�'��*˫�0$M������=$���p�����q��P����%F-�%���b(d����`�H�s������e�p�La���+7151%�6�a�+�Du�t��~C�������{��w^��z#���tQ/}t���R\��{ѻ,���ؿg��#���9zP��Ϸ��sh�>�����S2T�hG8YM�o����O��|�F��ѐ��Kr.杯!�-��� �����3��8ßj<�f�c��(��js�A?o��́Ӕ���2��]�����iI�B�r�R��k��[$*���Z�-Ϟf��V�ڴ5d�׿���9@��Qsn�VO!i���)f$�p=	N�;�F\�ό�@����$
�CH�9�`���AvX(Us*`�7{!_"�@����KY�X,8�Ub�A+!���]?؃��^���1N߸�������|�#�чO||+��!Jx4^�F�DH�YuK���ͨ�ʏh�J3XWIqCuЄ,�ù�<�^M������kM��)�*e�nJ$!^CE@͠� s�
'�=_��5 s<�4��%����&���l�	u��7n~���V��2+^,�x��Ubˎ���+T��:�m����h��Y�j�at]=���6w�6=���[²_'�<�ő�b�f%�W�Ӱ��
v��3�*<��bL[u䓈��	ģ9��5���*�F�����:w��)���r��"��J�'�=��b+�g��Q`�PK�j��jt��X�2N?x�}�|F��q2�6o��M7ޏ��z>��m��ߥ������{���m��e���6�	���J��C�zQ��[������*�R���4U��61O
���@�Q/��[���VDz%�}4�@�����3K -ȣ�?4����ܗ`��?��%�Z��{s�El��E3��j�_WݬM���z��oC��γ	�{д���wh��s+k"v�ռ�D��q���s�ߓ��*Ub�R�G�=�n���`ܑ&^�. c7ًh�l�FCJn�B{� ���� [��1t�=�T�Bx��dRٕ�ؗH,P�c����\|9�_��u�A����3��#���u��O|�çcld7&�|��� z�:����s�P(���v�i��<̫&XIO�8���`z������t��ا([��!��J���Ҟ����JyA*^�0�g�>څh���;�)�D�M���< ����k*�d#Q������Um2\S�9��⹚Ik��Ʋ}mW�]��r0(���Q{ͮ�d=�2DHt�i޸�6$9��M���y^�:���v�3x#D8*j��}�n�f�ʁ����2a��Ot��1ۖ`w.3Ue�Gm�8�������V踲�v�pT�==?��]���5��%''�2dR�d`���ޡ�����eG*�BV�ޒ!F
s���ׁ��2:�ۑ�O��_��o���}dgǱp�b8�6z�A�;W�)�y^F�[2!�����E�z}rOR�v���|QM�8ҹ���$r��<��%�I�O��#�y�8-�7�z콏����.�A�������n�e�I��~{�����q/�H��g��S��T���8����D@zc�&ª@ͅ+���W�c:��̙�R��ƭ��>F��X\Өq
DAz#���[��ʷzC����jE'q��s�j�";G�t���F.�ڍ�ښ�roZ�cf$N��<�t�H
S3�R,�#B�l���0(k��_f� �=�{��+�Y�u�m��0�5�X�Ă)"�(ݣC}�IWg$��u	z�`�s�Fh�)l|���X�&1뱝����x�e"H��؁8>��귝���4ƎM�oz-�c7�Ǎ�Bg���T�����L:�f(/�!*�0[eu�Ú�)bYʝ89�檔�P4"	v��I��|TarB\8$F/C	���"��Q�O(*����D$\i��@"(O:��s9Ia0n���N�b�G��Z�(��)T�e)�f���H3������	c��x'��L���y9�����'>�$i���XuU^JvL��t_�g���4N�/��ӑ�h|���m+���{r�#�*٪K��k�MKJ&B�0���a$�]�.b�)���M�D���)�I�Di��G�!	�M��Ć	"ȵ��r�bE֕��������"ɛ��F%�õ�i"Ȝ����H|�[8�Č����|��G[�֒�w��"f�C7m�ǂ%.��O�w��])"ܧ�0�hD1�'��Pd49�;Js��u��gі�g	�qh�A,�A�<�'x�]��s��_���ތ�}�l>������89F�a|�vo��I�����h��^P#8S�C��j�F^TgD�]cd�8pe�J�/;�EհO��&)�砚�h��Mʎ2y�<'�Yd@u�~��\�%5�ڨ�$I!nE�HcZV�\���yt�L2! �������es�b�=:��&u�.I~����o���׽� B&�����B"�03�4�F�k8��#�%�U+���25����<yR��S�����6��w�mQy�`:B�$Y~�	��4�W�9��&� �`��b%�RA"�	"�NqO������a�J5'E5�T��{F��@:C��Τ�4SW1��ў��r#��%���Q�r�:ҹbrxRn�8;W�%�O���=�,4w�,_�R�ut����ⴵ�K����}]I��p&k��9��F�&'N���Rޓ��zi�*�t���.+4a�h���z3Bo��48y�D4Ɲ��Kp��W�mߦ��S�z~ǭ�;A�!N0*�����Ĕ����������4������,�c��S]�o���uf����'�s��3��t���$.�ŀ�D�5�]��� �	����z����TWB���4$�o���wr)(w�����m$���ZUސd*2�d�&8�D�L��0;3+���w�ٶL.��JRzH"&��f�9UA��l�X4���i�vwblhH��N�%>��Evz�}]򂏨���#����8��g&Ӊ��O�܎={��:Np.��KN����1�l�*���m����&%�)�ظy��>�����������7�go==�4$D�Y�c�����������Ё}� &����?�L�u�4�q�l�d15:�:i��Nn�[�v<����<��la��q����=�y֜�eb�8�� L�W��m���$�{�r$����pqp�Q|��Hu_���g�|�����x�;� D4��/2��ÊU����'n���?�Ǫ��0<9���u�!���C:�$�嚡qVh�{ӵ9k�*�����uc�������}|��:�@Dowww�X�2��t�6�b�rn��O�pjj��'��c��b�A�\�B���4B�8�͢7�M���$	"�όbf�0Nߋ����/_��V�����DEJ�j�H�2$U�(JD8J����.�d��L�������&��s��0���B�-�P�E��5�]�߆{�ǎ�@߲�������c�NH��Jsd=EZnfjZ4E�{��G�����A&Ek0[����寓��R�M���I�ep��7aۣ����5i	L���va˹���/M�/�2=;%�ϲ���[�Ç���gb˦��ȣHG������Ż��Nb�Ř�����6�g�#����}G�Ƣ��|i��:i���lî������ J�^3�Y.X$4�%(!��G��{��.��|.�H�M;i�^b�o�-FI�\��kq����Qq��k5�%���ўg��Fp8~�8V��õ�ہ�|t3��)�s�^�|�^|�C��uߺ[/ƽ?څ����x��g�@�篿Q����F�7@�[vpū�H��q<��c��/�Y\�����5+I �	�Gv��*��\B4�����,wwwW.)-Y��T�:�*��d+�|�$7���E)7��/�L�av��-#��Qz��8
�Y���R���Jvhv>��a~�#�{;r=��]:�c��₋�$��;��E�My�����|����a�wP%]�,y��/߿��q3�u���9��t�x�V.�+�fq�g?��G�����ƞ��?�\��7�S��V:vL�O`��%�8lq����<r���Adb����w�6��8�w���t�>L��z'��g�c���|�q�@J<)3�'�!�x������s'���XAa@v_ON̊�X�ظ����ı#��p�;�w����M���b�U���n��b%}�ط�W2����~T���t�:���o���ZҎ1t|^wg���/~�+8s�I����L�pز�tt�2���;q�%`݆���Γ��!P��;��>�5+������ũҝ|��{���=�UKC\��3���Ż�}�wᕗ�f�0�Fʳ�~����oD���m��[�#-�W�_Vc٪��͍���X�c��p��I�H8l�4�����\����l+���_�u���L�ܶq�ʕ��ق����~����ع��H'pښU�Jn�Ԯ�I2H�T�r	R����!��}����]���~�r=N&�"���ڷ�I��b��W"�#˂C�N�0(`wx�X3������&��B�Q�qrx��������ɑ	1��{��������D���f�6�Q��1�rf���o�.�k֭'�5�͒6��L���݂E��dc����ޜZq�V.�}�>�_������W{�K^�{��~�x�A;A���4��t���tG�*~M�u�i�. Gp��xf�i�p��nOπ��>t��r��� �S(��}a���V��$�-�lv�ر�� NdcOO��:������5�b�}#'����>�g���;�y	jr8v�֖�N�� �D�2&�]���܁͛7�"F�=�+S@Ħ{o���ا:{s0��"�Ր��7��x�{���_F����暤SW�	`ɲ~��>���������j�;��~|�_'"?�ի��s�M4�+���x�;_�];�Şg4-��w!���W"l���w'[��Ŏg�����4�����ů�����|3>�_cɢE�院�=r� :2mR]��Cø��-X�GF�[�Yo���@�9���%�X*�ŭƒ���d:��#��˕������d��s��X�t�vY�d:N�?���r#J�6�qIK�$�ȵr�r��m�?���(�.]�|)�g\��#a��a8禡^tR���|��u"G��O~�|�k�(��#pqҢE���7�A�[[������j,F�j�c��12v��83 Z!@v�f6�h��R������՝������0Wwq���8�e��cjf��~1��^%bm8z��K�!�dW?z�Z��Ix��5�,
�`-�<1�����3�16r�l���Y���fМ������3$��#�F�ܐ8�8=�U/���Ȇ(��捝	���	:�[�X�#�r�舥�(q�������/�=��a�P��eA�I"�M�ˏ�J�� !����� ?���c�N���ItwP����X�d>�q���A  �Lq���������?���>|!��͛��kށ37���W\��{�A���$�l�>�wA�*��n؄D�w������o�>"��b\��ޱ�)�1f㙥�b2���~��$I=�+��kR��w���2$)JY"���h� =;1�:q.gD;�1��B�8��g�'�~+Vwz/ڀdJ;vLp*K��I�(a�6�A��N FҶ�p���<��}�<~�	1�,A�6�;I����e�4���*�hT5'`������c�Q(�Po��wB���`箧q���0L�n'�
�yu��ɶ8N�Ģ��������8眥H`�㽶��4+dw�6����IafF&;Mp�:]#�UͶ�8��93�SO�D�P ?�;o�������°o�,\���c�,�<~W �ɉ#��cI���a�1JzΘ�v��h� � !fm#Z@���\���&!�˖���&#��X���A�4^ij2�gB���/Q�0���n�	��W�nD;Ǐ[Ĕ��=��+I��i�s��6ه���sH�O��K2�_6����_A���ec��/���O���.{+�Aҥ�%�&�,�U�V�R|�]	�������YӍj�	$���FO�a�8�N5����G^4r~�ß,$��23�h��~uC<���	�nb�v��/:$(�_�crlA��I��ս�K0IZ��C©0]ʥ�� UI�H�v���Y�t�:9#nX�v�$���[6l}���IN|��CPL:ʓv��}��8��#���=���%H8I�-ʳE��:ڻ�ZY����(�I����Y���x��M�WL��>��K~�yZ�H��БX�y��t����!�O6���a,��W/� "�@�.��+�"4f�UǦ�[į�0�a�!�]����w�H��3�[3�ޮ��ys7�L<YL��k��0+��:踳���'��-�2$�m	�E����4	��I�V����.�G�U;b�ի��G�$x8-�ͳ�IqQ3��t���&�Q'{�
!�b�,��_\���C¢�j@�ȜطdQ���8�!�7�e)�R	���%�XDh=I�^��p|#��V��m��9�D<��d�['�"�
)ձzI;~��Yt��B��~��]we�����q��::3�HPuuG@�o������������~�A�_�� 9'�xo�� ��?�h�U��h-�J�l0�����,��4�&�X!#�ZR����Y���w"���-Ӎc$�a���ea!n~�xo������'R�8�W��u��w�Ej|-F�M��D31���t}�}H���be/�	��ۿ@|��)9��T7-�������I���˪|d�D
��d|-��Z�]�8�F�W^BZ� �NT�~�D�}=��d�FL0CC�p�����05=BĴ��������p{�xHu�sLҢ�YLO5p>���xN��2'M��m���02|]��p}�(ݛl�ݎ�vc���x�y�w͑Z�
�5��^�񩝨��H���:� i�|I�^�T;���!��`t��}��W8�ɚ���$~�������?N�61�Ъ&Bg���dO�IB!,���8H�AԷ��É� �F>v����d>�$�L���U�6��J�苘�_Gϐ�cblm�(����ҽ�]iA�uX�Lc�E�"��4	�C��ׯ�[)�+_=MR�m��M����qt�� 1�/|y#���ڭ���E1��˟���t#Al�e����$)� ��������CpdT��zPFQr��n�PzҋH�,A^�b4- <;H�����~"�Ũ��f[aQ� ff9�H�=k�yd����(��1Ż���8�o?n��X�`1��<�{��78(Vn��N�hŊ��G#��.Ho�tG���_�/?�$�Rdde�qO�P̕��R-�?��w��I�	��Y���z�ۥH��.�� 3M"�
I���
λ蕒6�����1b�$6n�;w<�x?�Ug�Og�]z�iο����%���6CڭJZ���K��կ~��o��"�!C�$d���:�n2����?Ê5���UI�e��l 3F�B�����w�C_���8�!'Z'K�����$�q0G�m!6S���&�Ա"�O��%C>w\����!�^�o~ۻ��I�VM�1S��E�77�Z�amQ�`e�VK�.,";�̛���v�������8:4Ms���8F	22��8jm�mw��&mA���� O��ٳ���^b�*�O��#v�+N����H�Ƙ"�O����ĥ���^��se�X��b!����<��ɸ{V"��X����PeL�)�$�����2�1�A�)�
."�$zp��F'�D�CR��o$I��t�
"���Q'�H�H;u���CG��/ǯ��V&c�sO�zz��،��,Z���虂gـ�9a�����w�I)W=:A#-�����ob`�"UL��9�P-�t�cx�{އ�~�:�T��0M��6�W�����ʕg`2;E��&���ҙ^,[��4�,��G�JL==��ŗ^�K.�B���W�U�%�2E_2�"���챇$� ���W�W��h'M�o
�#h�!&�7�8{��Qs��W�Y�Gz�Bc�y�ϧ��_����B�-��@;��QbDv�v
�2�a��}�=�v>-�	֖_|1�>�\�6a�����`��pr��>���/@�T%�4�0�(��\�)�_�f~���$I��5i\�*�6��N�m�:~���%!y˪�NK��0i�d�.N�R�1K���$�^�xD�(q��ln�x睿��Y���\$�"�9���ޘ��3;:�,]���L�%�7�-������������}=x7,h�c;p�do~���������cC��UQ�A7OR(���ه���md�F��%_!����pp).��UD�dX�g�h�K^N��
�͒����7�����v<��c�1�I^�����sϕ���fs
��x�l�JUJ)������n��a۶mx��w���O��U�@n��hy���[6oŇ?r���6���$fݦ����$�f�h�Ę�!�T�N�<���Ex�;�-};9�6trg�ǜCdH{� 	g�]"�0Q(� f��K���[��'����~�x$��قdy�":�w9�]�Ԗ����:�2���21�9򮊩@�h�����Գ��LPbXr���K��Ȗ[�.��_�&�n��+i�86t��� i�	�Y,]���o#���(z�"�1�����{���Ύ���[r�,��`�"[j�`�'�D/�YzƔ�\p.V8��B��;v@l�
1;5�=D�k�\��=��]:���liX�j'	�nR���w� #�����W^)Ҕ7�@^P��rE�
oxÛp�W��� �8,�FF]�Ƌh ��c��&��
d3�!��Ax5O*0O�¹���א"B��=g��h�{�q�؈��-�#�Y���E3�?}�DZ��.!����Y��Pǁ����$��-�������k^�z����~@ܣ|m>�%?#?w�4�:@�>�(�U�!V�Z+�/>'��!)n��}��M8q�(A�^��#ҷh����1 ���mq��W`�GH��䚖�6��@ۡ�Dҥ	�,�1�)m�> ȅ�	Ҽ� "�f�i�����8]�Y�Ǭ��g�ǅ5N=�l3��G�@��;:�zd[��#�}�wc||��i�6m��e��i1|rBz�rw:N>�U���^:�Y�[����"v��<��'O��+.êe��Mu������Q�;p�d���=P+";=I�b�m���1>qB{q#�p�ƿ�t�H����>ch�jW��qm�L�$��؊Ik399���R����ݍǶ?�K^q��������a���?��g��Ĵ��|��8�/n�O��꣏>�����
/�U����"yA��u�cUo�L::3KD<HR��e�%�t��ja7k�$D�0h���)LΖ�12�4!�?r����1OvEZ�����C%�����dU0t�������[^�m*�iltX��I���+�T���XT^�Ό�F1�^�%HTޟ�a�%� BY�p����%(cccزq��{�� ��p��Č$���h�D����C{��N�٣�+p����$���g	��7�C�GI/�c�咮qͧ?�_��w���X�d!.��g��W^qff��UL
�V9��H퇉!7K�G?������7ѳ�fW��_�ܭ�<-";�tf���ƹ眉�=�����{�^�X�@��W7�� ��]��W�7p�Ȑ@�81t�6��^�x��q�=��k	>���~�I���p�?E�ف�ĉ�#���ߕA.;FҼ��q7n��}�w�伿���>����|����FYb�t�Ɯf�{i�#)���/�E!��l��¤�*��j.:��X�.���W� �Ds�=��d"
�׿����b���R��<�|j'���b�(WG�L��/���M� ��ߕ���3��ɇ	^��Q8Nֿx)6�}1�.�L��uB0H}u�zP���w��^��4\�����[o��^������_�^q�$��ķ��q��d%��&q'�bI����H���,9������T�4�bVr��㊤���;�/��6�ecp]����q�%��md|B4	�LÓ�N��H ���/}F�Fcd�������ٵx��*΂]�������Τ�$�Gq�U�&aS'�މ���)c��a�5=�];���?��O� �t��+��@�����5������Y��}ca�}ؽ{/�����O~�A��JI�%j�U4�����ށk>�!i�{�%	�u���4�=�<�G�ќ�� {�{�����'�N���7��w�E[�":��7"-��]����j����܏���=X�8��#]��8���<�xh9V.�����ҕ�$H�H��;��-FF�x��߀2i).Q�ˍ�A�f�~;��s�#����D�[�v��[���{+n��&LLqS1��N��m:�5;�z���6�J�X#x3N����߻�x��_�s�8[�>���\�Ti��-��0����؃�E���A�RX)SG����G�y�˱z��b�E������\�"�����ؿg7��p@���.������$�^!m"�0�g]G2GZ1Q3�IM8�Fsl���o�I��y�/� ��b0�$&��a-��o_�-��'?@"����@j��t�F���_����b�\n-DqfF�_ȍ����zЖ���܇��A҈'�ֹ��G��_��X��&ö���������I�����J���J����~#�x�����cc�`X�1�3�;;n��>��	Ff	V�2��$$�ڗ"@8���Ez�e��%8@���ӤEC�p�Y��ݞ@1[Bn�B/��,��	��'�/?�:>�����FG�K�,�5�����̞��_s*E��د�x���k��?�CG������ұ{3DCX�݇'nن(	-�����CX�h1���W�#{I(,$�\���Ȧ��]���^5!i���nU�2+�/	p�aN�����	�=Ӌ���H�-�h��O~d��Ё����;�p�����n���3���~O�x���8J8ҵ�6���
�>vz��K�4#Ud=$��� =����L���A��,��B=�II����,_v6l:���F)��w`��b�D�9)F!��3C���=^�ض��ؽ{�Hof��^eF�<���І�N�{������#ْ�i���+���� ��@��ޣ���A[Z�[�K߶���]�R�вI���c;��mI����s�씾�Sē��C�������\��&#��+W,� aXii)���h�������76��)d��lL��W���NC��z�ï9�L����ɾ��O���}_g+��%��7��%�$���rz?����tX�
�`��.S5n�a ,z�����(卶8:�ɭ�U��L�q�����y�RB��f2Ɵ$�?�z�vf�ʼ����-�#�aq��?���ށ��Ff^��6��x.�{�	,]0�h��eP� �D:aTy�ʊ|t�����p퍷c��Y8&�m<�	�޹M�����9h���'y�j*|{:{	q�PJx���T�T�Ƥ4�s	���J�9Ɏ���k�m�)�&�De*����c�h�z���c"�8�ȱ���t\PIp�Z��٨c�M�GZw��H!��$/���#$\C����Cp9K�B1:���@iqF�Z���QQϛ�<=��G��
űe�V��	��%��21���Ok��$��f��P?��l(��q)�m?�dW_��ʅ�_I�,)�0���P��C���s���.�hj~���H��ԉ*3��s�?�ˮ��gS"^P����۷��ƫUJ�y�I��?"�Y'5���0�|�6����ǟ�k���.E���B�bI]�$��F^RUcö�;�t�ͮ�1Z[c���$����q!�����%��GGQĬ�j�|���S�Qes�4�a^v1dhb��H�/�MQX-R�K�e�w�!M�8Մ����>�8�����&�B��g��"�9����~��n��Vb��_���}�q�lr��TC�5�-��!�\!�/��S^9��ؤ{$��	��H��l��^N��L=L�w���Qc9\���.��N�z!��ĬY�(+�E��S^Qh�1b�Tzh(ADC>�	�gT3�M,Z(ݪ��ȓo:+�rz0����y��<�����-��#a�߷�8���2�_VY��$̋vם�ĢE�c��S��Bf�X>�|�-[����o����TD����'oT�^�Ru���^x��E]�W�E(��^��� *U;k�g�d�����i�.O�洶�1���:<:HǶi����Z��طs7o�U�|��a�4��c�ɇ=��D.�ؔ؁��DbR��l! 3��X�ڻ�l�/ʙ�b��V�.-+ 	M"8ү�������yE(/�b�906��9Ss�2~:0ԯ��sEL�F��gK���8���z�z4�.]R���Q��N͘�n�y��p�Lڒ�������dPKε��k���w��k���e6��=:]�Y)&�|����'�-�RN��c��jJ��HS�:o�`t���JY����l���ǴB��C鎘�wVT�<��!���NF�0J��.�����A�_�V�-�m"���h����0���]�6�S��y9'��H''��`aQ?�b����}����dd/�������������]�]�o�;w���}��*r��҆%��yV�fI���y$s̟?_aЮ;�z#�ER.g� �5�Q.W>3PD+%��-�U�bxpXO-y�)��͛7��H���,~啍�U�K����+?�L�=9�('�����0@�#�k�(l��:��HΜ=s��a��&��-�&&�:� Mϩ�‟X]�\8���u+�l�����?���́��<0�dGƻP��_F�{� F,9i%B�2�A�wfG��Ձ�с��|��T eD�	�ڂ!��V�3�f`ߡ��'_*�( '�U�_�G��E&�����qrt#�1T���1�"j0��O��	ԖTj3����/6�?[�~5U�\2����Չ2	�94�B�r��4��eU����\HK�2�=%&�3%4}�:��"�+��<��d c����L���5�U�۷� #�(L9-�m~�]�4�3%&���N��aD���A��wx�b�ٌ:��=؅�]�ϲ����� �x��q;ⱌ�0�Ӎ��:��{��C�`.[����'zV!�_�eAB�����AA<^`���=����K��H&pH�H�DO�L��\ ��C#c�.��|�
a~^oa1�wt���R��� 0$DJa��uhy!���8���`%�{�ԖW�Ir7H��ꔙ�4�����	��ڽi�1��r��/�O}��c�.V���T���	O�|���>�]��qf@��dTʟ�}��Q�m�5$���c�g �5�A�A,]���:�S�A
	U�`�E��(FG�D�,��B��B�b-w���������@yu1��{ըƥ���]v������3�yF+�K�If�5�f4ј�-h72�g@w[]p �]u�.�����t�d��U��zݸ��K0g.�ڄ��3j�L&�r��J4xݥm��&U��r�)�9OT�]_���ɜ��/�ʃ�,���S��<�=�7$��E��#A�􍪶e,a��s�'|QI�IT���8Nb�3��-�W��0�o"�����J�af��8��(b��㩧��A1�2�իW��0�����h�̱~�:�b��e&���"twwb�w�2$@��xc���r�:�<�\(9@+�k�DQ[W��臸��ϡ �C���@H�rfPRQ�X<L���S׬S�3���T����]�={#|C#4�!:��3�h
ϐ�g��s/����p���{����\o��u��?��f9;_{|��~�Yр���8�<��nr,���Ui�B�H����HfzɅj*K`��u2��q��8y�y�"���|FzB�>�X�ׁ�b�����;o�o�í}��3q�g�V#���y�ȩ���<�,��b� Jj�1�|��:��*p#�$�J��k���է���׃N/�Q�h���JWae�h����c��f���!/����ť�(K��BO�-y�)h�UO0{&3Y'�T�D�RA�bf�i����4���@M�X�*�7�K�ı2L�m�nUm����G1J��k���/� F%̍y���):F�,%K'��ы�%�9�9g5l�H;��i`�9=�� �����n�%/ųϿ�;��L84�f�,Fue�	�	�E�肿U�d
#��ޑ,�a���hjjV\)?S[[�^BI���PQQA'��ݻ�uc�P(-�cc!̛ۄ�W�E}C3ľe�Ō�DQ�f�����=��z-��>�/��W_��������a��?�#�C${.\u�U��+Ǒc����B�R��W]���z��V̤�NԟekL����,�%�W"��ַ7
�38,\\���ۈB^����}�"8 ����e#�2Ҹ���b�9c��0y�.��"f��ȍ�&\�kf6�i6���"f���O{�n,����{z�\A���>��H�d���R�Շ�G��K���D8��u��P����c:�-�`��EZ���=�E�&[V9���֩�n*�{�Ԫ��5[ӺW\�l�2E6�i7��ܘH��WG󙒓پ��D�=�H���X��O+Y��W~���Ai��W�=��C4�<���@�֏�-�	�*7��S����N̚���8�6�"d��'L���_z�h�;O���q���D�V�%/�D�칁[#�NQf�u��ie�ȑ#zQ�����/�2�8���	�	3!�rj,����!l{o^{�-�ϐ��^�����L*��]��	�F�,F�^a�s�و%KV���<�����桪���1�$M�t�a�'Ɖ�s	c�P�-��3����n�g�!e@&����*����]\���K�=z�C��6"&4t�����N�VΓ"� �7���j�fi�f$��?b(�	q��qFf�k���eI�������,:� �l��9��"F��ѯ�m��2o�"d]�h����>>6��J����葉�HW�IO�6o��lj+V�����O/�>�hTJqƘ��X��Y�\Ô�yJyBv�CV nZ(Y� �L���,YgG��$�9M���E��QVZ��<ڥ�u�(�*e:?�+b����X>C?�ՙ�xx���¨b�4�xM0����%'��δdѭ��Ih������Њ�f�cb�'SQt�pZ'�V�:�F�����F����Cb*�P���fbrB��D2ݷE��d��o�.!5dy�2d$�B�F�����]$���vq��8g��I�א���
1��Cnb�Ȑ_!XYm%_w����� ]}z�t���:��
\x�e*E��!�i���e_u ���c4��HH�t�8��	ǎ���t�͘?UN3bZ�\]|��R�,.Ŝ���:1����5��K:fE�2���=V��{U����wqh�Am9��i��,f��!Ta��k���$鄢0(�K>Ӝ��x������� ����]��/��F�}�R����	�E�D�)��VWV!
��-o�HK�^{ ��ȥK�ˮ`=�r����V��Pd��3ߦ����0U5��aJ�_{���M�鞱魠�2�Ӛ�fY�hPB�ѺO�zzSC$2�ZË>�i�hg�����r�����售��2� ��\YQ��en��!�AF� �P����E�2~�K&��~U�����aG���h'��Eżİ;ۻ��y�
�����jSc�L�����
��۲�]�R�%��0���BA����C�Fj���d1۔w�;]V( Ѯ*�R��=��Ö�^EMM�ěz�r�Lθ�	?_+9��ʚ&����>�C��Hsp`����s���}�����f	!Sn��T�����?<��>�8�N;rMi]8(;�O9}.��F����(����hp\�Y�M8����~�!�x/e�籧�"�.ĝ��,.��Zfb���띒�1���͖��]�����Xx���`�ض�E<��C���~HnU_8�ڶRi���AV#�z��g��x�?V����"�M��c׎M�����~��hWY�p4��"��?��Aw7�BuôH����1�-UE���ͦ��Yqh�6ʟ�.��"�1����#A���W>��ͭ>L��hS��T:"ENĘȥ�����%B�.�^3��_ /�p4H�]:��䍑%�iQƶ�g�*he9�3���
J%ӹ:p��o�~��v�#��#�+���L���^o�zEE9#�1M{�%����4M���rQV�\yb�FH�{�`���fwK�;#�t�ʠ����QL���E[�^x�yؾ�-H6��6��8�K��G����y_o7r�����ձ�\�IGa�����F��/ۈ���(,[�aF��7"t�ǉ?��a<����	6���9�V�L�y�P>��1�;�<K�6�	�#aܧn��<O���2��(`v$w��4�u�\���^ӢB���7�K_�"�m}G��(�BY9|Q�	�q���/�=Orֆ@����3�\����5T��T�/41��Kj��� ��|�gDˑ�l�x<�*'���N�0�O8AV��8��¨�k��Z�%����T�nRϗ.�Ⲭ�����>RF`j>"C�˗.CYI)�U�T6BfH|E���w����b�~�s���M��N�;��e��t~:y�G���7	t�.��|>/ɐ4���|�+_ƽ_���K���z����s�p��uh�]gw��~�8�x�\̣GZ5*� ��K?(_/P`Ҝ9s��d:�0����>�E��*��2S�'8�aH�T����
���I2�V��Y�'���z�9�3�]qխZ�m=܆e����5z;��v���`��q�^c�6#��O�>�f*):Y�9�	G���߈��N��1v�Y�r̄#�C�u��2l��6��T��F�,�·���4>�� ������
#z���+b��~���v=
\Ez�"Y��t�X���u#���������M�Ä/� ��ߟ|��|;�2c��i�(�������IN�]��^��DlR�@��K��~�v������*��
)�M��F��]�P!�)�����ig�ڐ)�|��B8���L/>'O�1~o�9�͒���%V_���rz�i�=��.��;,�W�7.:���eF/�KԪ��z��"C2\7gR����X<����m��tQ���S�j�8��x��v����2BLj@�"e�U;�q��jQI�����!ƒ��b��]�tA�S	��իO@)�EL�>��{�+�ذ�Lť���3CĽ�8~l�:������	�R$pc��&�8���ct���5�*+f���/+l��b���6�Y	����P@e��w���#Z"��*#�!����������
\K�H��dGa�Ɋ��.�z�t�0���W^	%�V��]����f��_;Y�4��7q��W��� ۧ�̳�����햍��h�5S���|�L4x���$�J�J����dۇ1�	�ZZZ4xv3+֔�5���R
�M+\Ϊ�3n8w�@�ɮ�Jħ��Io�L ��8�/cP�}�1+���8�dAb�r~ 6!�@�9b	�鏶p<'�IJ�XoW'��H_���{�^L�}�i��P妡�th>D萤qL�&PU�q�$��t�V9W�Ф���x�6�$.Ri���&TeY��<��������{8�³���P��ё1T��a��m��\�J�����$)'���uTՐm����#��(��O3���I��!���E�@��������j��m�*J	�B��I�ЀIyQ�#i?�1�O�t�uw�����j�̷�"29���0P �d�D��ǣ!;چ�KW���H9�����1�~�����%�p�-���F	)6�Rx��a�<e��>r���v��&��*L)��J~�y�|����"Y����^-:�xfP�9��{�#'�h\�q�cCJ���`5��v�h���sY�.�2"g"2��kBg�I�s�4�̬�AH�&E94t���B&��#����--�d"��ܬtD�;���h�	]?��]�%ۆ��6+������{��	�TA�P*C��m�C�����F}C5lV�*MX�n��{�r�ujqG���n�p_�F�C^*��4������q-[�['hh�PI�3�t�J"�M�A�V�u�-�hn��}����K.$^ղe��d�7@�����Gu*���P�1[Zi*�6d���V�i�qo���5�k��qG���8�¿PZV��"wI˖�1o�"m�+�͈�H���z�f)�Kj㒱�}�$�I`�fF�}$��

<҈�pXMr�iǘN��u&Z��G"�LV9��!.�`�A#��[HZ��*u.�L�����q��c(N�91(s���[;t~YtL�dfCJ��ܴ*Q�ⵐ�>��**%,��V�DAC"���l��
֨�b�f'y���XE�A�����H����h�l�	��3#���PyZ�w����A�g���v�Ђ��,��Ѝ��n��Z��7c�.e֟p�sL;����/�8��I��˙�aP�~$G���I)l�޽h���$r'6^z��F�F�ڔV_�$�2��T̺`�Lެ�<$�!��͋%Q�M��^���Ct��8�$��GO[qaB���8���ٓa?V~���.��\��*:j-&Q:��ރ�i �8&
p�����LQ]]�'ֻv3���~�:m�k���IF���n������� O�-�˒g�!�w`ɒ5ho۫c�["�c���-*��&�ԇ�?���:Xɝ֟����OĤ��AÌ�jI"+伆(�ѭ�����L�}�L+�qoo~Q���"��{ND��k��'����suYJ�Y���E�U�*ǕW~|��t��x��UVT{��eH������A�#O;q��,_�7\s%vn{��_��h)������?&y���˼��hH�myf�F\}��x��H��2E���àfa��Eqe5f�^D�b��h�E|�*'�� ��,%�鍫�N ���OF8���$Y���9!s��z֢�k��*%{��i���PG�Y�pX��omڤX����a���2M3k�؀g��g��2�w�¼��?#>�eq��QP�Q�������),B��<z1�L��� ���x:���ATՔ�@�a�v�i�g�g��܁5u���� wf:q�p+�F:�����'�ӏ7^߬p��P��w,�[Wf5�Ж�'���[,.:�֜z��<�_O<+J�udSd�%�O�ɁX�ۅ��V=//�W��2©(�e9�1�'�kO]��?�k�튫�G��0�ݲFsT��<��Äy���0;q��7+���`���~șCMm->s������QX�yu��&%���
�pƆ�t�C:L���E&55hj��cm�ؾ�x��E^��*K����f�o�s�>K�K��$�{4����v���Am;�1Vi���ug�řl�0zr2��mt� �oժ՘�����֊Wec3�QB���(Uk֡y�VB��f�у��K�����.z��l�4��M��S�A: d�I ��bt��(�8p@�A�:�CC��ߏ�g��������������A�81�l�E�T;:��ۆ�:7�/��IB�t��j�o+f���3�b,<N:�	��A�8c)"�5�4�\��	�l����`���׌O/]��+V��o���Gn>��q=Xͯ?��'��֯2.�|;f͙�F�o��h����o��m2�j��Ԛeָ���v�Ǐ~�S45�GeUٌo~�� *@}�L|�_"�L�k��$V�U����q������@H��EB���2�w^�q]�1��v�T������Va����&��qU��(��~�h��H�Jm�,�1�y	E}�>���7/������mM.#�h�¥�䧾���2���CA%�"e/
���_��{Z00�gf��I���X�l>w�=Z���
Y�HWHw����A��g���^y{�Emu�`�Ã姜��g�ǌU�	��P��%��*a��e̦�O��rlPϑ��}��`)6n���ب�E�S2k���y�<.'|�^�Tv��ԖS]̮#�^���t�g���PB��q�s�ka@�s�
S���鎸�����A"Ų� c�0�;1�Bv���\��$�5e�hLMn�J=�'D*����T�+mJ���uu��HG��]�n��x��7�_dV�@1\t�X}�z4�Ƌ��,��n�Lh	�M�������X�v���<�s�Uʪ�k*�_�r�����rl_MH�ֺ	O?���~:�ѦNsֆs���~��á�92�����tW�ܘ\fY����䉦Nv�zKp�g� �/V�R'�oL@��8�=$��~���M�����
cْ�XN���ֿ�핑QJ�%n�� ?��|��;�N���	��1�f����ZL�IO�.\6���袒L����Cm�E�II}}5���=�G��G�M�X��Ю3���Ϙp�����s���&:���D\x�-� c��fz���,��L2���Ӏn��N!bG����"��u��,��3��Y�����IU�N2�	_�a�d*��}z��n��1���9�ä[��:�h�a��='�d˓�j�����I���BѦ�+NFc]#���X��.�He֋-Ds�ɧ3"��{�NcӒ_Cc������2�H�����X�X�ȍ�T�č�}'�9���^��5�*&N.Ifq莳�֪�jV9�(����뮻����F�|�t�M����ψU��z��55E�M"���Wj�">�s����봘h�JD.���OVX�2�%�2�g����=��c���o���H'f�3��
�Y�T0l��+%Du���^|�PE���=�"U����
=�!He3�n�d����.�̐��S� ���Jn�8�|_2C@��n��̦*�lf vW�����y���אʡ�Vk��-��5�5��Ņ^8����l�zڞ{¦�A�m`u��
1���׽�B�����B�)�BO	��u�J0��3�s-;�T=Ñ���/��]�!���Ǧ���s��a�4��,}��ӌ1��E+:�:UN��d�VD�C���^M,��8
	�$�������H!N��d�����H�p���h).0̛�5����9/zQ)�%�z#�����E,,mu���OӘ��0�%��ȃ�4DQHdd�A�(��I�U���P��Q�+���:�U��K�김��D3f4h$����~�h�H_<�;Ǵ��W�(�UR�%<�׋$(�(�4�����イ޴ a�l}��uFF��*�*9)N$��C�Yi����M��!I�r����߫��wﾩ�4F��ݰ#�Iz�e�����ݻW��d�s�9�Qѥ��rS�y��P���)Q�~����;�?4�x�5�a��T�x{����5y�"�Α���f��~�.�i�*آE���[���x��!mt��VL�%y����f��Ν[p`�6���'Ƹf��X�hf6��Ѯ>D��E6פ�A�c��MZh=�o���9D����`��'㺛nc���fO�ӗ�\�U�Y'�|`��d��������i�d�4���C������#:�3�5�W^}��z:/b��oI7�W�%9K���<^����s�G�VS+�jQ~��������7�\fm5f6. ?�bl<��HF�T�P�(���&�سm��A:�+W�������EK��4���Y�*C�̗et!:@��,�b�ۛ��2�,ItFinX�j!�r���!�
�{ڏc�ܙ�����B��ב���<��2r�U8��#���U�}Pr�������n�\�'?y^z�_|��-����q2o�i��%�0B1�Q�h,X���^�~p��;����#����q�=w㢋/�e�GdC��,�����Ƿ���G�n�q�-Z�y�7�ag�[���*OHV�$;-Vi[/P�������*\��T�Y�G�����i\w��򗾉ޞAԊD��m���r�e�֏~�Q�%z��	:�9�7^}���)�74����CZ��F�Y:��_�=�w�x%ńIQ?av����?������<���Q���T〈E�r��-G9�YQ(I�"��z��൑�]���J�uA����Gk�KF�����&��&�������7���m7߄Y��˗,g�GBW����0��BW�����߇'��("$A�E�����ݽ{���Wp�uw2K� ~;F���� �xH���
,h;���[�x�T��hy����ᚫo�g>�9��8�������5��Y��7��Sh�صk�}lݺ��:�����[u���L"���C:և��vo�+��7b����oJ�c�Nmo�Ѹ�o��äs�\o������o��>�����([�:�;����9?����ddTj�"_�}�n��_�yh䓌���y�4���s,8��s��-�qG��V����w��������(���W�g}])����w���~�z��L-k�Ԯ���z�)��ODeY��l���Lve��Yn<�K����s/��!�R,1�v�n��f~N���A3l��S�-��/��yP�Rm����R���3O��w^Cy�[O�k�*tN���4�^O���_⊫o`��?)L�M?x�,�S�u�9D�G�qI�\���Jv�L!��r�ş�'����&����l���3���M)+c�c��ϓx�ه���_�=[�KҨfDn&�={_��@s�'-_�l`DA~ZIn8�Ǧ�~���.��YT%�I|hw���:��G��(t'�k11مy�e�0VF� �ÏH�����08*C5�Y���t�����啛��ݥ���ݽJ�e�^~NNBO[{zV�El���6?�$�z���;�5$"2֙Aue���`�w��~�x�g�)�A8�9���v;��s�b۶��o �fT4O�NQQV���~������oR�y�H�?!�S�삦I-^nd%����(��/��"N=s=R�����r�݂7�}�]��<W���$��ω�y:��a�޹�VgU,��_vɕ�U�i�&�Ty��p2�,jP���x�y�W8��t���x�M���Ζ����tn5�|>�Y�C�͡p�� B�\��i֬?��΢�[v�^bv��sG�%�m6|jtv������2�a�(j�+����3�&+a�Mi0��� ��p9�U]Z�1�\�{��Z�&@���Ԛ�%~�4e���>�,C��Н����&���/��_�#�_�Ab;�ӊ�:��pKW�� ���}�0wV9�}�Ta���삐�L"�j�A�����{PH��u��.��S[�2��{�6]r�ZI޼�49A?^c����΃Ő�I�g'Tq���s���W^'hЋ1w�f���o�@k[�����ghz�ZuGW+�鈁�n�b]�!�K�q�"ě2���Qr$�x��+�c �{�3���h�B�#l��F !BL���)��
*7�|�q\u�ZM/�u��Zu8H���9U��D^g�1�s'�Gq�����B}}�rq�q�ڷ�zS���� ?_�{U���"�#�t��?����H�x�^_HC7���?��<̣�x���*�I�S{{?��&B�#m]�`#vI�(|��A�qh�n,\Ѐ����Ԉ��������rOj�F�hm9�5k70"5j[�&U�����j=��|f��= 3��k�/��+Tl;܂�O�@�ͤ�-an�r��]q��߆��\A��dY93pzJ�E�r:��0��?z�l�8�B������"�HI�i\��ecJ�X����ũ&!Mb�o1^y�Q��)I��]i:��#J�%���&�!���/ҥ���R?�;+#���eD2��E;��¹%X���x�OO��ͯ�K�F��.U��U��N�p�|,��i\�H9�b[�n��DO>�\x�������j�cv0�Tp6��C�%F�xZ�q>q�?��$6�{�
�����_��0�x�5�!Ҿm�ꠔ�͎�NM�$���0�|�1f�[�~'��Ɲ��K�#�
3�x�h��F^��$3J��.h�]��ɨ���Z?�^�I��2�j8u�V��;s���	�3���Z��BI��;��LU�QZ&������'!�Ǫ`�Q#r�m������'iF�3��>��zD���N?�s
�$!�R�j�؃?0�25� 2�#�~�Q-'9-(,���m���0�&ym��<(�exhH��������"�~-ۖ�̤�#@ W��lI�S<�<�y�V��?o���}�u�h�vttثjj�b�G		���{i,����aM�2�a�w8p�u���&�����M�N�#,�%v�%j��蠌�=�"SD�
����Q�2e5���$+#�B[��$��r���"���P�Vit '�i�Hxݝq�a�;�QH�<�+�9��hK���}�������v=��KU��ȏ��v+����!|��L�a���U�xR6ӧu��@�Szq�G���M08)���	FHh�tR��P� ���qm���ޔ�a���ӤSܠ����#Y�a�|�nv0�1.�e�1B��"�TZY���'E��3�7
i,cpe�q��zj޼yZZ�6�pX�q���4։�nq�3{�-v=yA0Q�;��:bp"����@�4I���
�l���fr\
i^���Q���B��a:FIU�v�� ������tH{Qje�ij_��rey$�F/�-�[����Л<�t_�j�zG�ۖ���#9_4�Ngb�H�Į۶�];iH�d"*��4c�.���K�B��<��碄���c����$f���V��N�%���	��B^<9��JGc�b�|NzzN.q�)Т7C��1F:F`q��@,&��y�s2#��pQ~"���,���Mc��猡�ح�lv2Z�O&�fJvx��f�p�J�~*G�Fi�v�^����'c�I�.)�j����:�����|J5Iz�t!:�pȇ��B�3���|τFr8y�'���/?#��4�X��(�,��Oh�``����a�\��9V�.:g#J;z�[�t9u�:�&m/f���穱�{��$��Y�TF���Ǉz��t��(�2GDf��I���ty�����e��|�
�c�*�|�ںF�s�
�zh��|�v$yu#48��H#�k��%��҅�m*�3��Ѐe���������Fy��P[/���qHԇ�t��s�Ĝy���U�Ř=Q���	a����zЖm:�<��t�B%�:.s�X�p�����=���I��{�e�d
��&� ��q��l9����G�����2WAjs��瓿�S���;����_�^s5R�v��&i�f;�ب{�Qoт��ػ�Ma�$�r��ԁ�-��� S��@mĪS�����ʊ�p��g��?��v����n�b�<U��%�zJ,;*�h�b�i��c�������98��]m�5��0�Ȗ����b�!��.'o�[U�Z��,������$����8�c�ò8X�r��'i���� �L*L8�u8z���uA�D�8	��>��"w1���_p���0�XO�eH��P+�	�c�_����;��a�\*9N��ߓ�����nĜ9�e�I�I�<�,_�p>V�X�-ｫ�
�u�B��,8<4�U+W�?�	"��v	����Á����}��p�?��m�"��NB�����u���7�!?�3��8!O�`j�����㷿���L9��7��^�NET�c�^��$墄g�E�2{�'Cb9�lg2f��r�$;��=}�r�L��džDB<'��U1�?�d,RRZ����a���F����ĀZF��GZ�n."R]t9��h�0�N��u���=>zsiR"�a�`!_��r4��דډ�J��Ã���fd�q�2f��)9���8F!CiJ��p�ɀ+��!�>i���LJ]U8yi���kw��i���19N��*��uX�t�.B��牌ic
���v+g��"2�'�-���>4̞�sϿ����~uu�n�Iq�M������������$���k֬�}��������"�p�F#1`����k�BoO�E.=��#��>�3y��zG��<��S���1�
���³�2j�Ta����h�9�_{֟}>�%!��bXhf�h�a��A��݋���b��AU�Xr����>�9>=0t�=
/�HJ+k��`���+n��ｅ�-�>)����Y8�|�!h2c�sf�(^�i}�l���8��eF	�P�!�����̊�s�Ÿ�3�UH�͠!]EZ���Nx&�_2�HK�W�!Д�Tw�^�Eތ��&Ԇ�V�����?\~l�>6�ϗ������������8�a�����M�ߊא��UXVv����Qמyz����^^�F�<Ѓ#�:@]�b�:�������F��^����V{1����d�o	&��+��+��j��h�3��ҧ��EZ���3�Ì<�8���p����Z��-hDU�2仪��˴4�$ͷ�u�)�ErgGyuz�0!P��&1�E�Ǚ.ìً���t|Q�$Iר@
��l��1m���_��
�qg�~��M����/<�����Q��7^t5�Z{_�GZ�j{H]c��ˑ��۴�t2k�U���ilr ���T鮣c�@ӬE:s�HWc�̙�L}��(	hvyHEy�������o��t���"�ᔈ�	�ommSX'�b`R�ҁ�~��aw⪫o��W\�`5?�s�-����K���Ȼ$���3�uuu���M?���w�����W�[�K	4K���#�mk L���Y9��eN�E{��^�wJ��yA6#�r��r��������UQiX0�vP:]6Xm&l߾F�ٳ��w܁��)M�a�E��/ة/��-;�L�
���s�N:�"���G��'¤0�!~͊�D��R��b�(,m a�8��:/N;�Q,Ǣm̢�c6@O����	K~��R�s/?�xz���~�����.LD@ȓ tqj�ns��`n:�ik/����c���:iVRT�Rw����3$��|�4/~�i[�#~?�
�_w���j%��u9������e���HYlR���F<$N�S�s�ԛ���"-G
.��bY�d��K&��,����]]�	�	�n݃�0�s�����L[6��J�k�J>e��x�ꌖ0��0��DH�h�̞�Q����\u�ā�ʳS�R�`#pV�9[���@H��?�:�@ʙ��d"�Е`%n�����*'��D(,]��r$"2�&�.�2�)=Z��i�x�ƛ4����TKv��7�:,WGpuf]�1+�f��Rf���Z�`h����ɋn�%�\���Pޔ�ٻ�)��������� ���7�u��$jfӠ���FȜ���r���S.��X.)�����O�&ٕ�� ���E��U��v��b&��^����� �f��i�t��V͢�Ԙ��!f<&;rI�mv#��#}#�$�.�f{I��p��:j���@1��^)\�ح9:X�s'�	����Ց��RE�E�a]2.*d�j�<��7oR��պ��ˮ�i�qh$��yj9�z��D���@?~z��u�{>��6/��"W������LN��[�����R����Cޏ�K�>k�z]כJ��}��+*�٤2'�6!��/��gx�՗QL�(ZOs��&t���,���b��Q���P��D���߰m�l{�nD�չMsএߦjv�x]��t�E�uE@iI9�NY5�X�J��Z�9z6e�:e��3C�D&�>L�������L�����T)��Lؿ�Ya�^d�
,� Өֺ�l�g�{x���x��X��I/�u$+W��Hl�*;�RJj��\@'1�cK��h;��o��狨J\(@ss3.��:��\�FiE^�\�>��)�7ӱX=��c��8��V9��f�[��Fr2�D��~:���١0&�"�AR�
b��]h��6�>�i����^u3����6���\L��PB��1��QQ[�w��{�=�;�����D�s�=�:!�Dr�8T[�Q^�����ڬ��{r}�~�<����=��2�7��*�2�,q���	�$�a���F��?�$��N|�_�e(�$�#%7\:eX�?�1}�Q��r��O��?�)~��س;+�,�5r�,�"�UU!j�����˵A���Q��2*:܏o|��8e���7�Cl��)ϬM���Z�{r�	<�ģx���Q�u���H˝�����WH���ڷQ?��}����[2�$x�E�)�Sj�G���%��?H�AG�&�z��U4���������u��l�2g[|á S��D������n�<�A��Aw�#���ԓ���ʗ�o;/�o���ߍ����O\�M`ɴ�W�Fg�Q�����_=�ǟ�;��+�bP\��z�R2�!<��s605���ՋH.͌fG�z| ����q�����E���՗q�^�|�L�xq��p�ބ<�8�yV�_�3ϿR7��u�]OO�BUE3J��+7�={���t�*_S���#;v��-��¨�I�z��j�r$[����?�c�m�L�x�l��x\8t�_��K��7��M��ߐ���|E~w�`fc�J�H�V�&�|�y3k��RZV�4�=�$�EP&��q5|�Mڒn�f1���!\IC����uA���hKF��ٟ��#b�	=9�z��ʬ�&�ж�?��	,Y�����,I8"�(�����x�0�B�/*v�^/��IT���~�k|�;?�}da�H��S�)=d̢���lD��۸M9ٲ�l�@��0���ߗ��bѴ,��H� �����\��T嫂��ϤQ�����.�p��?Vh��t�Z���7�W�����&����9��O��Ǟ�Ƭ����z��ϳ5��N���]x���o�2fw�q5 �æ�����ڲ+:;r�R�1�(j{�v�w�Nw��y�^㌬aUKK��$��x����M$��`��5��.2����t�<�C626�7u<bF�M��x�O����/��U���1��M ��>��Y�xYVQmj������\�5�
��3�sR����mێ��G�br�h�jUU��A���jk����5�}΂�[Z�ꮱ'{g�ߠ�1Ȍ$e҆�ܳϫCI&s��W�Lj_��r{
�ض}�Y7a���ҳ�r�9�xc3�v�6�O4PJ#N��D��x��gp�E�{=jlA�����=+�F�i&�xV�_���U�8�v���ìyU�U� ;!���)���א-�f�ӆ?%���l���S�_ӎ1�k�Jgr�w#�����r�L�@?�`3������?��9��SQ6����%�����o�M�
��MC�DOᤓNGEM�F���UQ]���z��:��w���2�}�E�e�z�z��֒��ʲ�u��^�䓏�ws��tyv���������x]�x�鿩���7^GMm	V.�ˎ�6?��Gmu��
�CϷq�7~��J�6��YaM}}���VT3�b<2��"F�!K�"̌BX����Mn?ގ�_~Yኴ#�a�<��9su�v�g��H��ug��C#|��T�C��́��֣�t`�n����!G�d��J��� >���u[��{�-�F$p����Ps��d\L��z���~���&\��cڡ)U"1!ƒŴuyr\��Duܱ[Mhll������N'>B�ə�[�B8�AQ3����	:	3�!c&!���4k���ڙͺ�g:r'%p��#����I���"�Y4� �{>�3�I����e��'n�#C{�fg��O�Ta���{�q�?c-2�v��S�E�ͥz�Q60�$1����p��e��c�r'�h��Dyy��B�P�n;�wc��9���!�a�&��۷��֪!�WK	o�7��_�0V:�(�x�Ǧ7Aڌ��QP^�'Żv�EQq6��H.���Q^�U�3I�e+�~[/�"�3��������q;�x����|��"���p�W �RR
��y�0���*q����n��§�V�w�yK�>�J��ɢA�vGv4Qn���<d���J�U�&=���x_*L2�,��dV* �n����	���~�|�:���;���T�H��dǒ��)gӈ+��r� PJ����H�' �����$���&�e�Ӑ�"̬\ZR�+��^��S?(��3�%�	�QMt9�����ڽ:�$-�-�Fcvِ�֪R2��-M�1zp��-��;�830��pM����q�GryT�W�z�-}"i�m�9C���@��cGT[_$XD�jtx 3ʲjČ��v}~�^{��J��?9�(V��㝽8�rT'��BBM68\&f� o�}*�0��,7-g*��1Ih��=oQ!�	+�I�W���AR��n����qȒ�*:(o`�Bܧ"a�}+bc��Y�� y�U5��iږ�ko��I��=�����{���A�R�j��bR�F?��%O�]��E����Vo�!����?/?�r�j�9��T/.d�X�D�[8���L��HD��"	b��.��+V��3�x�DO�Dw9�l���a��'�D��C?!��jh�� �Q�-Q�K��"��g6�"�kB�3���Y�Q�~�M���̘5{wo!��sB/o�����1#7�ys���s��ժa8�qjׁ8@:����F��).��3�8r�ȧN��݁j���OC���_�u�P�������[{��,�R�0�S`�ڵğO����ܮ=ⓡQ]"�1;!�a�BCc��Ki-F�,�=��%�>���V�D8*��eF{� on���H�{���CJ���ܢ4�93g5���L **$��Ew�}��b"��ܤ#���l^�.����������aIf�� ��4�:q��m��'���ጵ'���8B�l_M(Ǣ�k���714:��"O#]�2^8��`֔f6�B��!'�rͤ�A���D{q� �p'?���@l�V���W1�\s�UZ�9D"�o2W�)�J�wuw��|�ޯ�3���d��ܧC�;�<��j�Җ  }FRM��I���={�:�\kY����CX<_����/~����Y~��Bk�A��hЙ��9��ݤ�T��FG�-.��/��?�����
�D�� ��P
��Y�`���h��R)ɾ���M�(6Jg��/�R!v�'����?���S6����B������p�ͷ<�m۶n��,PEQ���x饗�RN������$�}���%�Ξ�e˗dS�x�)~��'����?��������4ZXT�}E��HΧ1o�|UE`ԑGE1x�Q���t�� 
LL�l�A��rLy�麛U� 7'��oJ�kPY��с���i��%$�MZ�FM��]�3�ȦM���8�z4�-\����n��'?P5�P4�¾Rm�,�%K7nܨeS�Tt�Vi�޾sǉ�r�)�l�n��̘1C����~`1H٥�~�z=x��n��,ߗ�p$ϲ�_��V��5%��sNGAY��a����?��aͮY��b<g�}6��V�"V�"�	����yș$࿭��;�H�3�D���D��"�\{.���)�S2r;���n�h��I'��ǟ|T�t��ƞGB����4�7c��s�X0��6�Y��:�{'
#���Fu �kV>����-��"`��X|`����S��ó����͛7�+�#����\���jo�������1�� #;�bPŷ�3f�������Bڝ6F�*��H{��3��O����Q#F�j��x{��F���p�ɫ�����8��b�\,X��y�_��+��31<�Ǜ�A��>��4���/� ��XM�#��G���+��"��p6����o�ͫ��b�6��2��D�)TW�����������eE���l4���y7�4X�O���{��耍���.m�W]q�
�n}�߁E��\s�Z��|4\��2�A[��1#.��F��oڴI��d%.��VkdZd%�O��EAQ��Z_r�%Ȟ|�)%���3p�g�Sw}��6}6
�#�/�g�:!���^z-�`۶wa���9g��@��ٽ�FO^��)mV[��)�SO?1bz�R��4��v;E��*l�p�jI�g5�s �f��Rz�HA@`���u�y���@�/�>3����1=��AG��!��9��Y��6QM�H,�u�Zn��I�U�^}:��z�$,���X��u�b�p��P�,�h&zDzKyE�z�}��1��ؓ��� �@���n�g�;��L#��uS}�0Ad@��D��]w}�g�#��ȐGC�� �1w�r\p����}��#�~�{SUY�� �=w%��"l{�u�6B��n��uX�&~��W�X�\NIf:�u�ܼ~������7������$o���n�L �M����6������O}J���۟��wgo�h��C&Ru��-�UʘaD��ݎO��)5N�~���z5!�ݔ�
�z�"��9|n�r_$+l`��L!� �.�]p��i����e%�3mQ(*�v&q���s�?�c�2m'ﻫ��o�+�K���P	��!�<����睿�����H��i��'Բ��vѮ��w��$�D�������-��Sd�`�Ȩ�<=�&��͚әq��ZUʶc4h����_��`L��Z���z�� e���VfGC�X��T�~���I�)ӓ`9�������%2�!��I��$�v*���o��P@��=$��s�!^���T��:PY#�]R�-ߦ3Q=��c���7ߊ��.M�Uu3Ո��<������C(.t�����׭���G�w�IVVۮ
]]]��:�4ݓs �(ATD��"�>*z�WT��^�  %���LN�s�����뭽O��^�I��Ǆ�:�����^;��V�J44/�g�=�D��4����̦��ʍa��Q��3�J�8���/���+����\۶y�t`^����K�c�h'_"9����m�\M���������#�js!��6^|a,N�����=τ�}1b��B@G�����_�~�c��\XG4e{���n�PDa��8d���i��09���:���2t�g�z�5�������Mx�H��޳{;�{J[��*�BN��J�`�w����r����"��i�z�?�c��z�)�N
˖���3�YT�mƑZ�0U��5K`�aR,_�v��v�����Og5��#���h�V�}��g��M:�W��}R���M�ޑ�\ӳI����n�ŷ����t��7�Q��3z��h�Yd�9�LL"����w��K"@26���V�W����1���XԥJ�c�J$q�5No�\t�>%Y��{��г��s;���V�=m_ԍr:��܃���,jH:��8ǣ�T�!˜�����ġ}�	4�_�1o�ǫe�v�!	iw2!�թB�@��\u�N8���R����/3='�Y7 K�jJˠ�t�>�\~�庢J�F���{��4�u3���s.y�ź���L#���{�B�	O��I�IW(��Ɣ	|KC3��<����կ�<G*F��.<�|\z�e��	�u{=ᲨhK���?��`(r?e���dnŋO_u-N;�|UIϕ�T�RJ��5H�6T_^z�Y�{��x�-z��C�v�Y5��׾qz���f�T�%u)oc~c�r}M�@���a\��w��h4��oC������(�UUi5aǮ=�3#�z��U�q�d
����P�\�[�NZ6NF�����=���v5�L!�#�XJ�o�%]��K�C��(aK��/+es:��\���蠶[���e��Շ�ԒyV2�|�?>��=K	o<���1�t.Z��Y[���0�|}~�Ûb����uM�X�|9֮?
'�p.	Z�z�O[P�c�ӰM��p/F_Epl��8��C8V�Ѡ��hn�BcS��!��&E�A絴h)��[��^�^���[~IXi!��_���qp�A�H��L���av��K�Qn`}Y#����n�}�߫r/:C��j�I���ˉ_��k|��o��:�vu���m ��#���\�/�ˆp��Fz�{�1�����ǖ����J__�1�%n��v<��꠲'M�[dd>�����ŏp�o���FB�r-��~������?î�{��/}�3q�.;�&8�AN�����15xK��	�͘&�n�c���՟�7}�'h%�6k��F��[�A�iK�P$x;i^��b޶K&���?GH��E�G��M���-[�
I�T�r�u�����
�B�56>��<���7?�7,�h�����ꈞp�ػo7���~/�f�~��	��Z�A�U�'�-ajl����?a����X�N(�Ui�#	�w��?Xܵ���������n���[_}_���E+Ioc��XZ6��x�al~�>db	�{�u�"����.WR&sԓ��*�3�(�C�O��!%��c[����އ�wvv�@��P�8q��7��_���lA"�@-�V:~�ӟ3�e�ɏ�h*O'�+����
�l�0錎wJ�N�D��Q�������M�}� JD��
�t}υҶ��A��2�"�T�ٓO>Yy���l�����q�t�XSS�� ����V�j��_�*��n=Qn U	GG����.�GBN��<��b�uͨtW��m[��c�`��'�RyM�"FL�������@/���r+h@`�,g��ud�W��)n���tH~~�F�g�]kf���R�W[�	7���C#��g�%/?أ�̢����t���'I�͒��7_�-8'�t*����ox/�ڪ���v��&����ĥ2xn�#8�U�{v����n��A��#J*�����1>�,2$o%���x��%	���̧��_�{T��F���0>r�}�ϱby;Ȉ6x�����_����ah��"�_������I��fb��8Z#*}Uڣo�Órg��r/
3n��q���H�j*Y������cd}��Dr2�^=�ǅ��i��g�8��l��ͭ���t]R�é�@yȹ|RZ��s���h�Sj�3�Y�[3����a-yz<�{u���c��5�6J��!t���?����)�j�2K-��w�u��U�f�X.G^��B�(
&fw9�xa�sX�v�!�BÓ(�<�����v�r�0h/�uɼ�t�z�MD�����S��t(��zyf�t҂�|H��$��r$��4a�>�6��r4≱ADK��W��r�.>���r遪pb	N�Bf^J�t>ʬ���, 	�b��wAz��Gr%ā|���),�
�epNg�H��{��*���L`zb�V-%޶�׶c��ON�H� -�m�R����k�V�P�]o���R[��nG�XJ�O~�n&\����03�����I�}�ȥ�L�fu=��xG�l�"T�|(���,�4;��6?�74��a��)	�"�&gTdJ�Dc�!um�|�A%��*?ڃm$,꠸h��.��{uH\�H�%*�si�u˳��9l}�U�w�9*��E�(1mJ,+��\J�ɬ�2U����d�_��8Ú5k�����y&���~Z�		g���1�浍Z �~AY¾>'�2|��}��{��1��*]HX��Y�:$��n�:t� �9��$�
�V�׻�Ƚ����k=�@��)J�3�Q��R2���B�X�%K���3j�쒬W�� $P��f�Ɩv��r�"� p1�)�W~L�+s�U4��*Elo'���������̴�>!Z�w��
�|�r����yxf��7����L3<�nT:�01�G����9��O�`6)SY�VL���?�uG���W��LJ�g�f�����I;�03|��u����;�q�4�>�]w,�)���ͥ�C9ٯ���	Է��!lۘN,���b&���$�JR��B�U��n��g�"���,;�IȉA����&��Ҽ����L=�$���編`���C�!��N����et��7��v����"6�Axn���D�C�k�F�ee�<�ݼA��g��t�9���m�+Vuaˋ��iu�'U/�k#]:%J2X�L>9>��^�D)9a��L/�q\��תl�N��s\����@�\S?���C��)F0$|��!���*�E?���Ja�ӏ��V��m!g�x0���Ҟe#�*�(3**�ƛt.?9X��U8}�{$2�q�*n:ߟ%2?z2/�@��|��`T�*�������<�6/8�;���?��%y��rs%���8���J�����i~D�����"���� )�	��ٰJK�� -�)F]�Q�UE��X�zuy��� �,nf�~7^{s/Rѐ�^ĈI%���D	�����9�3m�0Fx��w`���:����_k9ȩ-��\^��L�)�������f�Y_�W���=��F�єFg���c��'U�t�:�2���}*�F4���!o�C��.2C�S�u�r��hyxe��&Aq���"����T����|&L�(���"����M����3������@���+��Jص��]�S24#��4��;��� I6)2O4f�P	aH'Ss"�#P��ԎU� �O2���c�B���E�B1��K������A,Y�VK�R�=UmC�A/�Y��7K�����9Ec)�.����eG�W��.j����́IE������e'�=H�R�a��?O��r�|Q*Mo�	^���K�@��6diT��rm�a�b<B��F��,�&��!��V��rW�����x~ۙ��}*�"�9�	�����3ڤ�b�-���""�v�t?X P�fF�t.�xZ�\�t����|�"�B�^[c��aD$.���zFё��nOBsqTU{�W0�ut.g�zA���sq��F�K.��O�gu7�fhi�E:�0 ��y\��q��$��bQO�+�
zB��Qf�E�������i�jh�Í_�:��� ���C���?��|���Я�@eҴW��8c2��IǞ�3�<#3�!��KYZ7���lB!W�B���w�ӄ\�r��	�͢�����W����v����S|�ir�F�g�lQ���#NЌ`�ѷ4�����n�����-����Ui�D/��@um=z{G�)���'>��SSr�Y�٦�{1�����~	l%�5F�����?;2F�Qf��g����>��hN�~�y��c9c�e�j�Z*�4����-�*���Sg��韎,��#��T��&T�X����r�|�QǠ���˖h�T:'Ńe�N�שk��~&&G�K��L�"[*�ڵG�[,��<�XH�gs�H��o�+ZNtJ�Yl%�^���t�E�^�D��e��h�Zں:��+>J��38�$�����'U�I�a���u�tVoZM|��G>�肓�/��B��e&�o:�쳱�#v�lop��rUtHɐ���=�9���Ç0��7�����E]����$�I/���M$�������h�B�(��Q�ུ�+d�c$���a-���hRN\e�ˬ�vlt�Po
N�U3t�U�As�V/	umg'V,وh0ol�t�#�fp�g�	�a۶�(�Q3�$���$5�Ё<X�d��oH+�`r9���
�YԹ+WnT��^�D4'��}h�\���D%#[4�@�pV�IdXK��W�Y�G�zK�vcd�#���Ho�Ϯ�x$!�f�ǧ[t�y��B�[E)\�P(�9X8S��Q�y����XB}GG(+��0Eֆ�ݻ�l�`�ZM
)�j�I�na%3��L{.&���O�q�AϒF�ɿr����U-hj�!��"B���!#k�fcsI����!89���0z�`�����Y
]1�4l%C�3�Mh�i����G<���6�Iډ�,�;�с�c��zZ-��r�#�"v���AF�jTF�̚��yQU�A��գ�z)��j�>�k�y�Ỷ�4#�9a!���ᇞ���q�ZY`��#�4b9j[jTN'�!:_�_�|`o�N�{`�q�9dsV�m���W��è<��@>�%�.��,V�|��uh���)�բ��5t��\�D��&~m"�މ���,b�dfݳ��صMK֖�#�J��	T6��S�#!�±���WU���	ttu�3W]��O=�������C�Ʋ�+�Yy���EmC�{g�͛��q�>r�e8��#���c��:u���`ͪը�o֒ym��X�[(��d}��yi��4�YM�����2ʧ�ڹj6�[���B�pA�Y�U@H�t#F�AmҘ&	޸n��M����ػk/�8�L��zF��go��А��C�0�|���v^�!eR�'��2"������FzY2;3�����o-Z��yk�vñ�O�@T����'$�d�R�ku������To'�N��UC#�{�`�G�F8T���	�e��AIz`Kenb��h�uܯr2�d9��pW�jb4읧�"�s&x��eFSc'>���}��W��j�j�bm�)s鮕�Q'�������JeX��x�\����н`Vk����(
gFE�Z���f��T(���5�T/A���%Ǒv���e
+���2�G� ��ʴSV�S�h���{�ٶ�]Gj�V���I�����<�kwvR$�S>��?H��W�4���Q�E�@�dǃ���WQ�#ԓ黁�^���L�\s�L��~�ʏk?���Z�ɪ�b9B��1/1�2��Rϖ�x��w���Ӆ.Tm�0�5��NE�wt�p8b������\t�E�b!M�X���ZI`��fnvz�4ԅI���Q�V�\�+�1��t�S��J*�H�����:�_D6�3�K�Ih&�s-m+�t�&{�z�'���5E�l�a����f4�ifH�n	[X�s�t�#�=9�L����d(��;'����%�VfT/m�äP0�r�\8��ƕ|�e�9�|��%��5P���s�<1:
	��A�ٞ���8�jF�M�֖r����JDu�M�C��H�8��@a��1�i<#g\�Ý:�P��Q����I։2�c2<�hJNS��3X	w�Ji�yd
P~�T��}���PF2OD�紋)�ɩ�ͭ$�M���B��9��c��)� |m�iȌ���f�x��Am�۾��|#�9��6۵���A'�mE2���ֽ��׮]��?��j+̉'�e˖����	D�/M
�,��]����:���?5�R�B��ؑ���w�z:N[���%dya6៝*�KG ��b��pD�$�^&J�BRd���ؘF����
+�H�2s��Ĵ�("�(Z���SQ�p>�,��E�@���oO��,�� ֓s�ٽ�:f�9��,���QX��IӘ�B��i��݃��R=ď�-�kDeM��4
�Hr�-�6��C���ߩ�c���߃Gy Ys
����T������rL�B�l�D��d:F�!�L���9�dz�$?I�17"�� �1�!"a��XА+U��D���[t =eP(�H�GQ[����,d�'N�1�I����Ǉap������hi���,����8�j�e�Y��	�j�
<�$���Sy>&�,�ncpzͭ"(A���Ώ*_	�"B�.Ͳ"�S"��HG�{$#ػ��%p���B=����g�u.8�C�v��K2�XU�����"�%��}�r�&�շB�}�1�G����G�|A��'P[͟M��x��cv6��7�.� �F*�P�$�¢��К��W�v������F�׮~��g6�+�T��tD`�ǡ)]<�ྜྷ8�w̌"-M~[
�q��ލ��g�гp{���9��D�	W�	��B�ݘ�!��i=�f�x�o�p��ꆍ'3�U�Qj�ŜH��#1|��1:D��4Ԉ}_|f��"��ע��0���s+)�D��s�׋C;^���ݍ��v�م�����j����=��λ�������;jwZUO)������/#z�)-Rf��V`d��e-܎VH�����g	�����������w֪�����P�وJB�R��*�L�v`��S��[��\��� ��2�}�Ń:!r��h��E*'�9�eb�I����ZT�4G�z|����볨�1Z���*ub0�,�1��|{���,��*�!W|
����£��??�'{���A]�m�V��ٶS"7�����t�C��j���T?�$y�gq���o��3�cvVR�B�,oa~��5�L�M�f1o���ny��-�
��¿0������z�B���u���1�ԍ� C��r�(%'~�S�I��w`'V.9��K���14��(��/���	C*��z��k̒ ���!�ұ쨩�D)�ȋ��N`_"G�lA��O����ʤG��uၭ[P��+�u9Q��Ѓ�b����6���5��Q��$��r��
3��6���Ew{36m�$��_���L#K��{~�K>�Y]b�;i����ov�AF�VIa�J�p�O���k�KX��M��g�=KS*�/�@���^�:Q�b
�;If���܀��$��Q��g��^:�YC#���1�kXx���,F�w���0���,*�DM��c�AT�f����'1��7o�c��-X�ҧK��G��^!WyB����	�3\IwG�cz���݄��I���[p��_ACC�,�%�:[_yu~�¤ӌ��!=��j4S�2�_�������K�_w-��'h�Nf��W�h8��X�r��3��^�6U}ַ�b�}F��H��f�p8���O*Ohmk���ob��ᦆjD��W�2�nVUO��4?a���c��#�Qq
E^(��=��~�8�Ĝf���%F�Q`Do�,�I��~c/�:�t�����d���k[_��t�H�I��R�%��W"ھ�o��/��[M�jl��R[4Cg�'���p�(��n�43��D�n����/�C��RQ^��ld�fB��L��([�2��.f��}�κ��[�2C�P�Jr��e��HP�����"A��Y2���SYi"�H���T*���j���壱��� ��dUN��lhv���7�כ�����:.�Q�B!;�2��^"+#�l�!Գ��"3��\l�0�;�������� �;��I����}:������_���i����L���n]|"j�`���N��� Qȯd���g��G>�!����G�v�?%�Az�4��"��.��
��ҽM�Θ_�B�0g�o�>U�T0��l�/a|d�[Ҋl[�~���Fm�*���U�ᅦ���@l،ddZ��d/��D/��1�[n9C��6-l�3����Ԕ�Q�QJ�@��.�8��f��ɉ��!q�i�Y�A�J��f����̈́$T�bt)���C:eU2&�$�C�hm߀U�M���Vw�~+Ih몗�hn$�Y��@ st�,aJ�� ����2]|mD��IJ�R-�!N'V�}�>B�"=4��F��J��h,�u�R㖽ϲy�L�y�\��N~��1�ɐ�No��M��Gve�Fp����	�G� ��RG/�E����.�5{�M#�HB���D�H<�3��S7H��h�A�������aA�D\� d�!Z��Uq.�����������F���f��h2ZJT��Y,[�3�c�ͅ016�k�ʓ������H�@%}R9f�htN�X�@6��j�՞�
�,=�3!To��,�D���f�����j��Ywhy��&.�H�?:�=;�RYtQ_�����k�]~ �s9l8��7b�(˛]��X	��3����;*�շm�H�|)$BA>H/��8fiF3+�[�@�e3a�n��@�R�0DĆ'��c1V�Z�$�2�"ID7�Ic4cǛ�g����T˔�����#�
720���&���ͤe�p0��� Bl�lBV"9�>���m�ѹ����r�8.�`8�'�n�I�
�Ba�MqZi!@��L�#��n�� ?����s��9r�*�z(�?�PXUn�������@������LT!�K)w��t�vaJ����L6���IxVC��0k�CTVi{Ce���0#�Ք ,��q��tY��FQ�6@�&��N�j3Ety��/� *s̵u5��-A�.��L�BF�]Dt�¼�����-7�l]�k�� �1[t�K~�8� ���o��a)��<%�م�|�߇F���[���Y!�u���(*���ۉ]ݺ��Xȡ�azdjy�u���e�L-e�b��J�2U��Ȗ�6-�ׯ%lF]m�JF��x���0�;�d�X(F$�I2�@~���V@�]{{q�l7��t�^��XM$��v�����8�����W`���d�6#N�*+�~|U�V��@�W�qV¢L)Ig�j밵����ڟ6�𽬺���:�w���f�y%u>B���(|�6�L�DV���B������C��Th�3� N+����DDwXK�N&�|e��/ٙ���B��/ɂ=)c�Q�+kI�3
�B���W��P����BRK�V��8�F�yj������1�*�%�G4I>��}3�"Kǁ&��u9���If���%Ku���aáC�� �NNo #|��8�sUC�-hG.rBi�*�W�P ��)���=�7ٽ�J�ftO��U2���}h���= ��EsrlTu4dc��R���5�7?k΍��	�>��t.�)Qd�t����"V-*I��}
1-[�C�v#I,�+R�)�z*��M��EhH-�ڐ�'�5ƈG;�0�{�~�	t�ib�$�zfIc1A'M�q�%�k���oAmS���P���zZ�l]��Z�UȈ�Z��#O3��y#����i��ñ1r���g��5�����J8���g���xwNF
	Q|�5�ѩ�1���ϱ��B&螡�3�:Q��"��$�M��j�V
�BIɲ�`�mr�P�\Y��o�l��BdK��y:���m�jBL?���i�x]��:�m��=J�(c�S![�k�T2�	������	��5��\�,'=>�(�A�Z֒�\vFaO!��1G����Qd�ݪ�r
}�	'�����?�O4���׬�wtp\�.��b�Z��0�%D��*�Ì'#4j����)4��� � ��D·{9�����3�A�g�A����s�uO��#L�G<s!Fֆz�����&���p��7�猨f���0v�ُEK�i�e�}!�l�&:K�� �S�@K��V��Ҋ��@,����Ť�9F�$�o����Of
�h�I��U�:�\��x�6�ԋ1b��A�hR��G�@�R�
mS3U�h*D��/�֗��� ye��"7�`� 2�
��t:���!�2�I$cX&���� 9����j⃢�H��D���0�����/�{Y��i`j��i}���@"�d%�������m��C3�\��4v"�4{����͕*0a�.SI�Ks��<�h�Y^����v�)X�E�9+^~��;�4v������ ��ȝ��k��L��l>�^"��ӡ98�6��9:-3G>L�ֹx�%��_g�h6'�RE,��W��[T�H�,D%�&�\u����㢋/VU�ҕs���5D�������R�).�Si��1�']�o?G(�j�;�s��d^�a��;;®={��<�c��CG`d��`J��xk_�������U�)P�Ŷ}����W|K��7Y�p�0�H"����q8p�ƣ�\<�}3�*���Ɖg���4�rw�$��O�D�r��Ha�_��8�� �L �(�?,�.^�q�{/A}C3I��녍�Z�!������L��`/��r:�Wa��Ո�O:�L�fb���8�	�N㘔5���9Tav:$[u����W���Xܵ���.�"��d	�� K0������9�7��h�V�GO[ʽ�;D�ĭ�|��E�jђ2j�N9�È�����H�py�����A�
��A*�{���^�d$�k�i[J�����f7���ӛ��(D�._t�̒��[7��9��ix*h򴢶���d>'��A���sq�U=h��Sռ9>_i��^���`�с;�o�ܩCI;v�@��EX�n�*�<��(í�<�J�;N���* KAʅ؛�K���1[��&-Ʋ���-�]��¿ϫ_�Uӝ?P�E;��yVuZv���N.��L�cX�v��(�Ā�4d�ڛ��QA&���TЊ��P�2�R>����n��I�>~�-�QD��TVk_�]���.��"�"*s������߈��LLM��A$Wk�.	F%��BKr��&e�*-Y�H�'>~5��&{wo���t�k�\�Ab�X�s�t�a��(m��'Lo��ǝCC���>d�ZΊZ-#5��.Z�r�e�7(ɞ�9>ga��~?��,V�i���z���G��7�t�5���Kf�LK����Yַ6��z����	Չ�V�Dt�(�� ��C�@�I��k=L�6�=+�CU ��b%�ҵ]N�T�"z.�=��"cCC�Z��:�^nn	�ޮ
:��W�RrѠU�u�վ��>�Y�5u���YO!	�z^y�h)�5�mm�>�2�!D��.Y*��9H:w��,�;)]�܎t-K� ��Y��Gm���0o`�ȿ���L:SR����c��j�H
ĈF"���Bg{��Z���rI,[},�I�V8�CEjrznBu/pI:������X�v�*Z��sH��Qm�����zms� z}$u��g�^�ll_�jB0����Y�*���JYUR�`���4�$oIZ�Ě�[p�q'�yG��L�$�qXk+Q�"��ϔ�9\�Dcg;�C1����-5X��4��1�'�f�xԨ��lrd�Ҟ�X<����\�;��Ӣ�Z�3����N~�M�C"7L�����d��ƿT�d�ܯ03���F#h"G>!'���If�Af�I�r|�f���i�k:&�7vZ�Rs>R~����1��	鐎���i�5��XL�m��ҩ���ͪn-����*�cSx�ɿ��W^�,��<o)U_q�'��o`6�@�dCh6��;M�m|^Mz�����,a��}��Y�s�QYѩ�6���J�1hSR���
�:�y�����B�s�K+I&˿�CM%��'�b�����1��/_܃��zC�.����|�1I]e���0���c��x쑿�?���}C� 	<��#q�I'k�l��W�	��Ѥd�DU����cýx��q�=w ����Dy�*|C}m#�I�����w�O�
1Z>��c���3��g��-�K{�┓���������Ųr�����nMR<������?�ǖ��^��30K�V�c��%��F�������@SYS��t�>Y^ߴ�Tu8�������@�x[�8��c�&��&ly��c�� Ο�Cj�����*�t9*H��ѱPY��p�00���^f�8�άb�9���p��3�4�r$CQf{�f#�5��\/��.f��Q�!�J��4�*����!B �A:9��vӺ5xc�����0CL�@�dv�}	��݉ǟx_��w�b���I0��c	����-�|�<p?z�~ {vm׳����w�7�����������Di<�3���}�C�ba���-M����[:�R��^�[�,��׎����b!����c�����{���d���N���сuG��*)T�ѹl��\x�H2BG��������b߾=x�'pݵ_b�܀��}�j��\���##�<�׻���~�������1z��ߎ����w���E��-Y�V^�M��=�k>�9���\эO�ț��^:���0��ߏ�^}j�pܐ��j���Ww��o��7wण�����q~͢,��U���=G�%���YB�r�-��E���a�k�s��W�ÚE"=���
� �]�H���7`tNZ�|�}8Ի�d� ��zPWf!sL3Nbtvqf��V:�l���B��u6�kp��~C�Q�Tҙ!a&M�f��YU�EwU�IB��nFphkH�T���-�����x�Z2m1�h.1��Z�IQ�3�u ��I������8���Zĸ	M�d�(��צ��~y�O��Oζ�cA嗲�W�6#����������=sX��UyA$8�j�[�nǷ��5|��_�
*,f�K6J�&�}�`l�\(��FFfX(�ʟ�����;g�eJzCv��/�b�ڕx�-:k\]�ǣ{@�K7ވSN?[�*=�U�������|Az}L�EOgzv����8�{��V�Z�����t�u���w��[����:q��ݜ/������/�]=����Ҙk��R��/n��*��޳03���4sY:�$��Y,]����9f��rr,���^}	w���8���1;��Lr2�2�bԯl�Sņ���p���`&Ql[Y��e� �AUmm�O���]8$Q�Èі����:�,���|�)	�ӄ���;Tv�H㰖�+�&a�-Δ�Ps��v��KBJǐ3��:=�3k��m%�·����+0��rr�Ɔ&U�hj"��9'�u���Xl��3�Cãhm��Y��	*�]��wv���9g�b�!�{(<#�V<QNH96�_�_��:#-�"���Ӊ�}�F~^w@�+���됓i;��C*�����W\����y��I�V��o�$b^o�������&�a�����8BCc��I>��>� 6l\�=��"S�ޑ�i��#�x����6�<��\���~%�������ߟ����̇P�ʀ�u<�䣺g�c��2ch&��fhb��H�m:�a��������aͲ�ط}/���� >�>�#����Ք!�l$�\��N�Ԝ�l�/����F{�����{p�I2�[-� |/�}�>��܄ #���x<2a�������YM{�Ӵ���)���8_7�7�|�����]�bjte�q~6��]V�;��`�I���Q���"�{c��=DZ)����xRU�#c-��L�[��ϻ�p�HÐ}Y���g��f�5�g�CXD���2=X��`3~��?�6iC�_U+�'r��'�NË��B:�&[�d}m�pLW��u�1~��X�����T!�3}��8�ԍ�7VC�v��9�����*��%=�����s���Nd��ȉ��=x������y�!��ɬzkS-�FK��m}��}�Ft�lU-XєjR�ذ#�/ꀪl1?�vx]����q����lVk�/����t.[v	�ۃ�E���xm�5����nƣ�<��n:Q�Yd\�~�:;�t��L���LjK���Z����El�PN;��ԐI��������TWT�����j052M�Q�)-ؼy3�{�����8V��N�T\�,�|y���ʍ��D"1)�Ms$��q42��W�Ӊ����=�>>G�j���kc��/��z
U$���:k����l$�H���7�߹O=��VQ�Vŭ"aBN��Y�$����p���(չ_��g�`M�������GÌ��Fըg��zF�H�>��g�����	��H����YU�3:/K�R���U���Xu���\�jNf�i>��Z>��Z"g�F(�����ڶ�q��'{ژ�]�r�&����T~bd�uMz�^�͚t�T"�{��	I%�H3��R�p��{t���E)���9dQ�p�3Zg���úe�LW��I�����/�h~8�T��.ԅC�����;:��%�J��H����,:�)o��"Y������Y*���mzZ���%�]��5������Q�'g�[��	ޖ�Ņ�&�?C�#���?0����>YRQ[U�C("]27��+]�ɤ,I�}&��t�>ɗ����LN����H?�D��w�0���o���#spT6Ȇ)���u�!F���Rط����EL�4���;LL�h���o|:2���4����J�p�tp�L���f��61 �׬*e�\&�a.g�J�˦�B�N���$�g���[�LXPْ�����`9��\�L�Vj�RZl�X�畦�8u�OJ�R�\�������VA�f�Y`+8�RF�o��a#�\J� 8�D2k���$|N/�6B���(�jk�\��g��Y*����Yk56*��u#4��F?��ȿ�^��S��S6�־#73�����,W�w1��p\�DX'�D�h�WvJ��-5��;�߽#dS)W6�׵�r\����L�Y]y�����Œ�k��H*e�����e��$!�js��^�><d������&B>l@�Ǯ��M-���6��32�H�S�v�t�*���4�g�%t�T��2�,�&/���f��jm'�EMU�~6�h������[[t�H�D�DT������h MN1=6�����w->���G-+u�Qmc3��8�NN=�Tr�)�Zݦ���I>����b*mV\)�C'O~"Z�7~���r?��!m"p�h)��"��G>$� $��y44��	��{���}�r���H��2��c���(_���htb��LH�ׅ�^s�g𝛮�4���ʊ�t��&m"���DoqW'R̠".&��Z�:q��p�A��qxe��R�hE��Txt���3W_�s�f��lxN�1�І�G6݇
B���$��t���M�wtc��0�,_�JO�ә��.�q����^��0b���>5��%G(w8%����k�W02<������=l%.#�`K�n����a*��#�����s��y��%$�E�_�U._���=��#�zFI�r�Fg�}�.*��7��gd0�XPZ�GHv��c3A|���4��ڵGG5e@\��n��{��7����1b}�Z�0B�u�4���'>s����3�I˨����U�1�Zp����6�gi������o�����g��M ]�=!�#��jԆ��h������S�(��G!K���`�����sAG�Xۢ'��/��_��^{-
4�F�z��b`�M���o��$���$�2a� �e���c��C�.�RPQ�xD[��x��p�����Y!Ѽ	Y5�X����'q����J�F�D*�+�F	�6n8��q&I���	+;a��d�j�oތ�>w�E����*������}Twgê{e��������p�����%�$O���Oᥭ۱r�:|���I��i=ܳ�L�C8F�,3A��k'�[#���x���wt{�'K�d[F����v56YHWȦ�t�J��b����]�����(qksF��u%Љ���?��o�f�푉1���`���z�j|��ִ���]r�b�`8����9�T�X���_�i��`8ECu̅2|�k_���C}��]*e?���Ez�w�n�������f�;��eJ���/�����/����i{dv:L�����Q�+[wa��otn�=�л�U����uW�ɛ]�LR��LCn����0J&

������8S�l_�?��Zf�g�� ie#_�s^z�L��dH~���Z�W_�ic�l\5�*�n�:)�~�ySg��3)��~�����eU�����|f�d���:j﹜��҄p�ի6����ؽ�u�P��I���)���c�;u�|?�wyJHu�DfF>�l$�I��|�a�VU�v�ֶ%�~s�E��=��HlNO�E�H�^��Z�'���>�({nnjřg^�MG��KV0�T�LG쌯��"��^8�����m'�_��A��p�/!�M����&F��������!�`����Ќ~��t���}���M��E�H�Pv.Z�N~v�xS[�[�\��c�ڕ���W1������W鎱ޱ!ř��L�ڷo�K/o����'������k����>�����es�:�%[\|����Gpه/��O��aF�A����T����P�D�I��ѳD����C�ON��܁���8�w;�a�^�����r6�YW)�����8��K���ERW�2����clݾ�����f�0�/_��9�B�E���Y�o��1Y�>::B���M߻Yw�f����O�"�KZ�Fg+��*i|��<�:6#x9��e�~��r�}i�W����\\%�zbwXT#��c�ɼ¥��e��7o!,T�'����z����t�`4�s��c��<p��G��$�+��?����/d ����3�d��-��#���`�t�󋸘,~��w2���-��)��U���T���H�i�&�}ݬ��F�m(��o��� ��9ļ�r�x4Rol�4��Þ�{�c��լʨ�\�X55�#ݥ{p�]O"Q�&f����.���y�F7��v��1"Jӕ�N�p�&���\L���.��t�����!�?M#8����TbͫP ���ժ��@)KJ����pک���QW�>-c��YOT��7:Ї��������(s���^x����t���0&Qp��cvh��ǉʪ:F����d��aQ:�ҥ���ܤ;�d��[��ո�����rȥ�tF��DW(�ѽoق�g*{�D��X�ي)m��9Hc���f��u1S���G��8�@%!�&�pb�e"&S\��/�v9�p{��y)_kA:g��_�X]�Z�ٽ�2S�R� j��#���눓�e��:��;w�Ѳ��\�*�ȭpV1�;�:XFh��֤��RȐq[�,�w�0F�<)�7�7NSSgU�}��VT��Z����k)yn��b�֑J��JʘI���N�.�#�m�����1j���Gnđ��kӛ�@�é��A^x9v������9@'�����+�`�7ѫk�D�fכ��kQ�;'��2d���=wh�OV�nX�^��?3Đ����ؤ�A/I��b�,��֗1E�.����W�ԝ�c� Һ��Ub����4u��iU�����v���W��aN���c�Q����x�sߛ��V���e��tq��1;���x��^���E�ty��Y��˗�T(����H�*,�>���3��% |������^�g���6m؈/~�Z4��u;L9�΄UF�4��$d�����nՔ�"���'w<���T��)�����ɠv������B�'�x���*�%��R�;��Sp�5�'9BF��D��{�H#���F��/�<���ƂC�_�Gq��G謓3��MfD
��!��\�MX����q߽w <3�������)|��H�����)DW�2r�!�Q36����%��X�,��J+��Ė_�:�f62��q��e�꺺C&�)�/d]"�;M��y��rr�)���`$����"��S��������%K����^�|��LF���篻{v�s�G����Y���t:��qh��јD3j���qtb�0�_���?�RW��C�Q���	?��&�/,�D��[�l+Z�ʥMX����ڹ�v[a����گ���RҪ�T{�A454������⿾�]��j�8s�~����%8��p���Ȓ�N}5t���A\��s�����ܠzώ}�/�-����g��1�"�qy�^��m�8��3t�K N��R�$�����/��S�駞R�'U"���&il]�{�?�7�x�*Z� ��4>��ؼ�9���_�ZY2.��2e6;;M�i't�����8֭Y�ٙ�A��E����a����ˮ���3#����!;�d���;���n�)�[j�YQ�짃F�o��H�E�Aޓ�zn w�\\vKK�N`��C�a������T�Q�r��Y�px&_r��}�% +^�6������a2�yL^Xҙ��ɬ��,����7���R������q�o�Ӈ��r+2�9] a�k����}���P(G�jV�'%B��}uc�����������M�8V�}�C�b�C�k�#tY�:16�O|���w���N9Y+T��iB|��:[��k�A��]��No�JY8H&ۏY�[��&�ۏ��;��-:�)��S�Bϼ�Q��%����`�Ms�P����^��} ]?삙� ������k����
��-�Bf93�F����g8�ēh���N���%L�֡��}�K��AFf�Q��1��cU�=��7��e����<��p��4�!>3n���
O��i�^9GH���_7��)��7|�������D��df���Ď��u=|kkk!�R�;�c����N���Ӫ�z�{/��L����`Yr2B��#�b�nf�jO�l�9|�N~�~��9�U�ב,[��Df!h�U���%ϼ��S�_�B�U������#��Ҏa��8�ZX)U,��]�H�ҩt��kĐ�rb+�$��������2�<����Ie�����'_��߁��{���v�2B���@���woA���ǔ/����KJ�C�\�n~����߬"]�����ࡇ�st�٢)Qj�r���\"�If��7��#�:�Xn�O��%�������l\FB>�����m�(֐����߰��3����tI�Jd�y�����!�E�L�T��}d�`�`w�T<��{�ť�X��!�������Ҭ�V���L�6j���Y�"¿����/~MN0�;���,f&G��c���1�ߧM�jm�Z�@wtu4b��jۋ����2;��4�?���JT5k#��Q�k�ז�T2�v>����\�яc8V�ho%�݁�}�|���5��"*N��+A/�2hi�����I���dW�<��AF._}��r�ܝ&���체�ˠ�d'mg�к��K���}6"~Q�?��-�Y0l�(���4��~مH/_j��=E����X�#��w��us�|I���a�X���e�J�����IF�aM[������Ri��]et�������O}F�.9]��i,���/�>9�H�S��#P��Pi����.�X% U�T�j��E�Y�9���=�QOR�j|�Ձ v��*$@H�o� ��au#� HD�gĪ 	�|�=8v�jjX+R`��
����0�����.�$�Vvw�����| I��λp�'>�I}m���ЏS�YE�5�3ж?I�d���N�  ��IDAT�E(��s�PUPe^f�'T2G�.I�g���Q�I(8	�ۥBY�H��ބ<�?��bú�&f����d�&��)'�]��G�ӹ�8����A{���[N���=;eT��p�ܹ�N<d�j��M��B��ك�k����)�HP�I8�Ղ�o�#�� �<��,_c��n��N��B!��^}K��թ����	QB&o�I܋.jA�
&�Q_�rޮ}�Ѐ��|��Xpa�᝾��#��KA��6Uڗ�I[����C��6��BJW�J�/CR,Q�UيC���fJ��dk��Q��]��H�i�I�[����@ʬ�(ODbIF�Q4�6�I%��PH.H������Z�U�%��H$�{�t��J~��pXU8d�]��:��1Ի�54�ꪅL��{� ���c����aTz|�=�ePY_����6�j�zE���%ዧT�H��ʺZ����_��ITh�V�C�̈́����Z���*����
�3�&1L~QS�#7�C%ў%g!���UYFn�RQ�+���f�ۗ�-eL�g�����I��.�I�iLm��d#N�NTc���|(�?�C1���m��!����'"��c��ڬ"�B/j���2���e���I�V����GN�����z�/�:�p/H@T�E�IJ�%�E3�[�a2-^��������3ƻ�F�!^kYy�hQV딙1�&{Ĥ	L0���=2�V#����	�Cz`#Xʤ2
(v��u���$�4\i ��|���B*"�#S��[Y�Ѡ�7��0z�.��7�#OV�m�FCV��%-o%�,�C�r)+D"��T3�i��I�%���m^%w���hk�T\��j1E��o]�#�5#:�+8�kHͶ4�.3ߗ��ZT�r�r��ߧ��D"�����a6)�G�f	K�t|3����aAMkF�֬Z3���]B4�QyM�46�Z�W^ކj�	�b	�v'���D��(�[�'�_����S�6l:���K�=6f�Q$x�.�VE-����(��O=E#�p�����V�hn����{P�̕+�k�r��IS�"şgPW�.9ߐ����d�ݳ��g+�C�p�=*̜���et���v'tu�H�(�m�Щ4�B��QKD�,X�oI9��#�ۗ��������^�7-V��b@2�')K��$u����<���.��r�S��:�m^��P&)�7K2��x
.�M�X�l9�<��v2�~d�oO$2�b!���c�jLr���Ä��֤��٬��KC��4���Z4v��EG4i/�\<����55��~�F��*%�^B2�z���(�FzH���##S8�F��3��+� [/_ڍ�����+ϣe�ZU� ��f�!I���uGi�rfl��ag�s!^?�ŏ�gJf�]�*����'�ܵk�~�/����"�B~!Q��S���Y���fdlH��~��������\x�{�N�:2�gu*��x�8���h�����FKK�:�4�y�~�73�d���O�L-�y6f1,Y�w���n��1}��"'�m�vO��gW�_�@Y�S{"�#�Œ6��3߃��a�a݀d��-./aR��e��+�@u֭ۨs沓:��D���� ����Ə��F�H��%Kr�w�16�f��%B d�@6�n��MY��!�B !� �����ݖ�޻f$�h4��ɰ�|�>��c��̼�{�9���l�fEz�#QD�J�ZQؑbƞOJ�_��-S¿�Ɉ��a�z��b��	��P0L�"m���!+	W\u��[i��)�&�Eh�A��K��f�|���UV�[�\�`�ړ-���wx�3l�����}~��^>���X#�����*�hG�Ԣ��ny��a�`���i��ǟ��Bye�)���h��Q��aK��W��7��<���\�\e�;[ }���=g�;��T	մW7�h����t�zt���v]pN� 3�2��X�to1���J�Ųh�	�`��`�ࡽ�C�p��x��N����E�Y��oN�ލ���^3",��_��+���܋��r�T���hJ�����5�Cc�l��I��w�6!o��w�{�y��;5�� �ij��Z·������C�;�F^��q���U�O�����?�Ey�<����3���5'��k��6��n5:�g��BNA!���z����Q����7�3vb�ٛ�NFaq�m�Q�HB�.�
�1^�L�&'�$O�P$�cN.T;��ӧVds:u���s�D����'�_�����;[T%nT3��e��y���/��o��F�8�y3<��7o!�`��F}��˱�ep�R�h�1ހ"��'U�����^���~��L�l��h�2�r�����E̸,Z����y<<�a�5v�~�0�w�����U��yE�O;m#���&z�"+CШ�u�ހo�v'|>F;�,Y���xrLj}����j6^y�ct���F��P+��0֬Z�}�;�c�;|� \�T��7�� ��� ��J"�)y�����Mp���X��"��WKJJ�K�M�o#��(��ŏ���}g�Y�A�����/<��-B��0_;f2�2^;P��w�z����w�û�k������p;֯_O���Ϣ�����ͦ�����m<�<�����{62�Y�\���=U��Mj�p�ZG�D�}��,Z��ЉO��=zB��\�r�>�b,Z���3������X�GaB	%t�'	��@H]��2�0&����N��u��<��~���@l����?�]LWר]�>@��D��,=�65C3̪�PV\ER[��]���.���E��!������1����X���J46�Y6J�^^�l�}!U�h�<��8nLm����u��s���C�M�Іo��pme�4#�z���%� =���^Sm׬�/�r�����i �H��ƒ5kQ���~��EH)`��1�0!�	^��ׯ;�]�������	g�B̘U��V3ʑ��v�2�U�\���w��a4Ŝ��P<s.�Htld�ȯ�ԕ}�кآ|h�i�H�:?q�N�|�L~���x��C��UCikoBG׀��;*$� �@ﭵY=}��e�97��[�ƗOw���ާo�\��N�J�W@�{���:D.�|���y���;��d�T��Oyh�H�JDy�z���X֝�����*�j��ͥ���z޺c�&� -\�\i.#���b���zh�$&4#&`��<��5�s��.Q3��I�i�2�h��<4�b��R�m��m��a(,.����M�Q�#Is��t��V�~�q>�,�Jb��~_�`��iҍ�C!,�T��F#G�kFuq|�H�3e�E%��V�K�g�u�~���$40�`08�eb�$��QF�І���J�[�G�R˖��V�(q�/�H h^h<B��Dɢ��D� ��H��=X<o1�����ߍ�Kgb��}��������eSWE����Tn^〩��kg�@74�1r��>0�)�,	9u���TUWۊ���D�,������GO��_@���2���f���{�o!'*Ʋ�kH��*����4��h"�,��zh8�䐭 �쀔U��G����=�O�d�;lh(�r9���݄��n��6�����ϟf�J�����y�,ϭ�n�#8zd�u�j���Y3��}�L�?����?2���>7~�y�4�~��Zi�D�o����hdO��ˇZ[[��ϖ�E�!�j�j�	�2A��[j�@��A���1��R�Wi�L_�ɫW!����}���nK�U��$IN7ɒQL��}��/��W^0}�Z�I]�,��P(b�J**+�C�6���!�9����O���$����A������V�[����6m�$�c4Z'L�:ep�G���_���?��L�;Ń�7^`=�*�|���:�\%8��M>Z�:��m� /?�
v��І�G����+p��� �(m-�<�QƤ��v=��������;$l��v�v�����N�=ej�P�j��p��0	���^}���R��Z���+&c����=r�,���D
�C~>�,����{��P����4������٤�2h����o�4�^��f[>_NE�T��];���/>���z^[&r��,+u�a�g��� ��J-ݭ�q8c��gx�ߺ�?�����3� �5.[�W]}=�=�|�ٽ�>�B�h�6 �`�_�8.�2�-G?S\�B<�k���:R�c
�"��Ħ���O<�ݸ��+��Yl>���&b�d��%�M���ކ��}�b]�noF]�ean��1�<<��CX�z�LR7���Ⱦ� =�ÿ�%^~�V�_�hox'_�NB&X�p�rSJ�N�c/V��a<8���w�}��m��<���h;���m���C��W�BkZ���,^kn���} �k���������;͛S�ѡ B|�I<���ŗ������-�����"�������Q<�����SO�8{0k�\tu�㞻��#��>�(j��-c���N�����yVv��sq&=8������%���-����7���Q+:3��m��?���yy�Q��(���Ռ���N|�������5��	�Ծ��Ӎ���8|�0V�w�u������0���݌���lܸ��FQm����8i^�OO>��{�Y8e���Q:??Ǐ7_������&S��㩞>�T�;��PZ�����طg�x����1����w�����gl�
|H�4"�)rl�)�Y��ԟMA����w%��!�rs��G��W��<�tt�ܼ�H�1��/���]gz�>��ɲhwXVf��ɇ���D~�!�"+�UUT�0��5W_�g���I�ŉ7�P�Ij"o8�oƵØ00?;��{��+�������5�R�K�2��P�c�6������z�N���53�N�5@����O�2���R�4�� ��G�����E��H�E5y�6�����m��c)��+w`�7��?`5�Bz�S������9f��:��fF9/2���C8e�J9t�FD������2<���h�Qe���`��$vQ$��m[���V�]ec�J�l:KCG�ly�	sr2x0�7��i��>�>������o���Ɍ���81�+/���?x�F����cv*K�h�4�B��?�鏱h�+����V�W�������1#����e Z���))5�����r�:̘������k-�5�j��������ڈ��D��̠��Yjz���u�M�E��� ��Z-��@,)b~�&��S�2�V=�t��FP�TR,����� SD�>���εF�ݻw��A,˛�p����f���>�-��0���\8R�h���8�^��uux���q�ٗ�j���
�)����'����?d�o�É��>5���l����n�����n���>��#�ک��c$���A�%i�>s.��=��ϱ��s�p�R� �C$����|�R]|z����>�9o��׶o{g�u
=�l��CYuz�A�w�fֺ��J��Ɓ�{QX��J���0̣�=�;n�:�7�J�_��+�=���V/���X0��I�L��f��8�\u�5��=�4���--M|�hik$�JGuu6
K�ɓP��P+	{>��X��$60��1n�u˖-�;{�}�H�4I=^�]����LoO>��V���?	Q4��ʫ��H?��CS�a���z??��R�ҳ���70k�B��|�<,#�c��7w�H���ح^c�)rJɱ�[������ʖ+����M���I�ǩ��T��o����k�j'�4���/�_K�x���,��H��b���ՂtO:>�_��>�u׿�@��=x�-c!�����QBl\������D��K�r��/��u�]Dx����mM8|`�C�F4Ӳ������j�e3R�8Z׀�W]m�>T��d�L�={QR��O�����z�zg��md�/�݉��yN^9	����i�.���g�������b/�t;��QHo��PA���q"7)�0C#$�i0��CG�����SbZ7C�����.��3�����[�t�e���6�(ΕX��fh�����4�#���v��n8�f�����;0<2̧�a�*�1Bvw��ܾ�{�z��tu��P���J�FCQ��w��4��Qk��QƸ��N�$1��=�6��U�mc��F�3U�ӻ ���IcUu;� ��3`Җ�O�����x���t�'B#�����6Ao���ǥ�M���MGQf%�Rǽ������7Ă�f�d�T�9"��_j��
�X��9�Rfa-c�A�F&�|ĵ�BY�AT��{�z~��e�����1��q���J��Fx1��e$K-|�q-wPPm2s����-E6��EIe)>��$��[IҪ��N��F3z�Q���t1���b(���oi�;3τ��˴`�td�Gx�K`�	����"ț�7U;�+�Į��<D�1b�qL�.�uK�"��������!�JvVY��#dtrY9^����VQo}�53���چLߔ�K=|m�9N�FR�;t��^����`��3���I���E��^)���o�-�d���k��˨D.33=��J���%z&R�6�|�FJq}�Ȫ�pOS�jˎ�T��/L���[�I�����X�'�ו$���P��v��:��ɶ�/�51��Rwpp�gT������ċ��7��`g����#�٧�J�֪�2���^��*�Tm!9�s��)'8��7M{����dU�>���ظ��Q*�PH7إ�J9�����Ǒ��_I����
�"-9Y�6#<�ؘcv!�Ӑ�zMy.[e� ��rެ�HM�3��RI?�� <���1�&�TVV�=��V�)�(�D��Y��L���[Q�kLb��.�<9�����h}!L!���֪�~������:?�I���U��Ԣ<�ˤ�x\&A��7U�'$�����)���G��#X1Ml�Ԋ*�Khٞ2BU5�6Ю�-A�;��:n��W0��"����t�҉���4Z[[�l�r��\Pѭ�v��[�;?2(�&t� �А�"������9{�M����ä�إ�^���}ʞodbКÌ��ZE�SVJ�G�Nr�j����B6��e�]�{��nӻ�P�Slپ1�ʨ��������ދ��	�c⹉�IL�����O��m2�x�R�m�$j�д��O���X�d��q���
MI�+"Dc�}}B��U�??�|\�"v�a��I����N1p��c|�(:��m�ZC�a^|��@7I�I�fق�C{�l�ɥ�`i�~Ls����;���'�)�2|Jү��+O��w�������<r*ᆋ7A���a��5<���$Z2f�1N/��/}	�>tj�+i�](�w�OO��s�I�-�+j0�ظ��'���z�t���ݯ�b��}4�ie�18H~���*��3֟m;����M�y����c���ы�r��6&��H�L:Q}Z��9��17ٓQ��y�����~��C�-�fB�s����}��k6o�l�9*4�_ł&�/��>�x��4ސE�'T��n^N����Ɏ�.�P�йI�`��K1<6���}�8��>	���@J�_u�fkk���&J��������w�1#��ed�b��L;��5GZ&����:���(��>!F�K.�̈=�	���1�ozy�62���ƚ���/���g��'�������ҭ2���QtR[�25�<5��X\?1CG�˟��r�iؾsJƅG�/�ìYs�L�cfa�%�,o^����څ�����݇��#<�ڝ���:�W>�'	�]��K�ACk�m�Ԑy�+�d֝u�n�x�=pe��+�#D���Z�3��"Z{U������i.z r���_��^}�9��������$���#���+����ѓʚ:e۵!'�W^s��Ã��¥i�y�
����r�|�X��d��I�l6z���p�����nśolA��v�,����9��ё .��R�:|���m5Hb|)�G;v�C�R��VT8��C�p8q����H��U��h:�`��53�������(�'�x��[J=O�B�ګ��o}�0skG��qbk-lt.��<W�Z��[+�x4���z+B�r�-������2:�@5����j�@k����Zl߾�E��1Sپ};|>n������a�0"���	6ۤ��=���LY���Ut^���!پ|�5�|�Ֆ���Ti�ƣf�2j�5�K�Ǧ�p��<��ӧ�s}�ݧ*�������CsƌYغc�ɡ��[�䗾�Ư�"s0(E�4t���&δ�\$���ʉ����n-����)�e�^��Yk0�Ћd�p8i%S��6����u`�ϐ|���~T?�w�p�����'�c�a)dҫN�;�zRM/���l��g���]�Ġ��L/�|Xt�\s�M��3�~E�(�s���ߩ|�sQʈ�H��������1Ђ�sO��|�xEɠ �x�f��
��]:0c�t|�o♿>e�þ~�	�*I*����Н�&r=�)v��y-�����7��}�6�n� Z�%ޠ.Z
i�y���:d�Wչ���Ν;q��!�R�㌙�f��R;���8�2.��yX�z��C������d��4k�k��;|ȌB��ľ�!��[G����oB�r�#��A^7�r;N=�t���!�(3#ˢ`���j':�'-_�;�[?|�G����g��o����S�M��.WbC�~"#6���/g�;��)�4�6��>�IJ�?w��o!�������-7Dӱ#�3{���a����kѶHr6q*�&�dR�kN݈�T.��^�]�&�Tzl�X6�F�7
x ���Nq�r�U�A��0N�pf�[�yQo��f�CrG�#�����&S�JV-"���|�����w����x`�qg��ꁷ����0♝E2拢�W�S#�TA�ן|cC�8�� #���g���*8l	W�Ĵ��34���Z2�t��\��^�<S�k%<�@��#5��ե�')�l��1�ԍ�t�2̙>� ��|BQ�رF8餓��A���/$fo2ܭ�OM�b�ZI/z��:zբ �R�J֙:n;�J�B�Cs�)����k�L{=Y�^q��A�����Y^�"��J�j�<�/9�3q�e��,�d�1�y�����Hk����x�ZD�,4;];c��L7#�u�_I�Q
��<����%��d���q�=̶{6f;������br��e��5k��<�-�'���߸i���p��g}�E��<�AzT�j���2&<>J�����$8<HV�F `Jqy�L��NR��N�����_�X��8>H��������Eh�i���#�$�*-/C��X����A����׾��vD(/1�sE����aP'k5�Ӻi���©�b�<�m�皨�����c2�rg����ԙ3i�5e�xx{�푧R�AGP�ݟ�2��[RRn2�J�ڵO>�m;l�b�
�u��v�iZWW���&��'F�Ki؇~�h����,-3Y��s�YVI�M�_?�>�gW�_r-o���A�Ox}��6:�ґR󡼭Z�u�D��~:�2������K-��6��/�����.�5���jI����m{�Ӵ_]|�R�PT+�uK ,v�Yy�j,���G�8ߴaS������kg�xݤ�iJb��`r���v&���9����!͕k��*��J�˴����hG��~F�ޏ��8�.���
�7�3g2
�P	�C�H;�<y���#��`��?��;_Ę��Pʉ[�_�+N��ų�GI��ťF@g�0<�yh�:�??�(����Ó��#��sp���a��087�5wF�e���|��R��z��o�e{�I�%z��W��6a�i���0��t	ځw���xEٙx�՗�����0z�@�Ǔ���e��&Q�kiW���;�a4�����M���}�M���+����12U/`����ҽj���p��O?�g����rtv���?"�r�����_n�~��j�ٖ�L|��%#�6
��ƃ�U�:�Ͽ�
�<�L�t����[��Iɘh_��3����?��7�z�Zi�f'y�Z/�T��N����L�JE��������V\S��F:�:s�i�p�y�x�̘

K��� �6���{����ű��B����%��g�7��v!�Y$�ҚSO��FN駼��_E��VZ��~8�m7HP�'š�����X8g9qx#J�>z���ҺhF1"H5l���$'�d�9��(�"5�M�����4����i��k��jQ�2'%%e8r��-���_�#ݍ�rV�+Acc+�^6��j�q��1c�)�b6��p8yH�Z���_��x3���M���<��㣿�Qb싯�����Ӯa� d&K�<�s4;�%�X3Y���1���|ؤh���oD=���5�ǃ�~���yCy`�9�]��6��z�W��(ŪbZx<dT��2��|�{�j�ض��8�<�Kءt��A���K7c���ܴ�U�A��?��E��y�D�S,�f$Ϸ����r477Q��'�F�}�����cs�v�H�K��5���ÿ�N��V�Dy��$][��J�Jp��Z:計�&=�>�-����v�n��n[�դ�#�l�4��b�R�s75�y\��s-�S���7ʦZ-9^e�?'.�200���a����[�7�o������_R�^�Ҏ�Nd;BX�|6��:z߀��57c0�/84g�e�>Z}���OQUG_O!z�� �C�����q��;H���BE�a�䗡��Sl�O8e=����Jxh�F�(;�~�m��'A	�/��#��	���S=�̚���ubC��t�q���SX�zr����NzX���<س�]4݅����4���)}�`n51�'�������oŞ�G�YK��~��K*m�d��Ox_9|�)Q���н��P��YۅDՑ+5J��i����HOs[jZ3�?�N;�B���uQcdܕn|b׮]ֱZG<�ޕ(^���DQQ��u�?ڜ�7�$����um9�y����4<��d-U�*+5�u�$�KͰ::�li�
]{��1m���\�礣���r���0���L���OɁ�QY3Ӷ�ʷODbV��K�ǎ/L4�!�wjY�D��[*qb���!E���5�%#��+���)�)�9sfم�k_AF��׿&2��� 48���<�V��y��f�\HҴ�Ш.G�yn�~�#�%�1�ׇ�Drܚ�$ ��#��~�]���$�=C���̰mC8�x�;�hPj�q�ީ�mb�x�,]~�U�����3ܖ�#�4i�;lݫoD��!	uR��O���{��� �w���)���HԈ`�j		�#�|'j*��޻[���s����Pc`�>;|m�8^�^�������C�6�`�v�dO�^Y#�%l��!=j&��*���MP2��V(��� ss
M�E�DQ[pKC|A2�k��W�#�����)ǖG������z���/��2<����g̚n�Dc���.���񉈣t�����W�:��9mֹ�y�(����.g	fͨ���k��T��Q��>:�F�M��3T3U ����Td��)�{����.���z%k�7Y�=��
k8DX�����3k��#2��>۾�r�Z�H�K
f��̵�s�c�h�ً��TK^��e����[�`�_������(J��`h|��!�J�-؂d�=U��Agz�y>�p���Ψ����]8��s08�O.�Gza:vm���cVq<���++������1�!EC>!F��L�!��b��J4�FIa��C���b�޾a����F�D��_5Y��;ڽTF��w��uk`�OCC=��?��d$�ԯ"��3��»�q����@o�M
jrOݻ��|�3thf@���caӆ	mQF��.8�"�A�E$��F���WO:T�-|�%K�`3�P�w�u�-{�q�3r+��[c��X���&X,�4I����2�C����R���u� �Ȗôv�a�BnJ�z�RRR�W�u�_�����D���T5@�$�6pd]���5��d��F�<r0
Mh���Y��{y�s�U_O���p�ϩ�7#���0�,�FZR�Z������,ۨ���G49��F{1Aҩ�Xg��l,6�3�7#C�
E�ɛX)���re!=Ǎ���j�����L�?I����g5�	�x�z���"������~F�d{SM�14�k�_�&6?�ԁ��2D����x�])�y��FJ4��xL�������=e˶6�22Jܬ�Ș�|F�xR*��#fO�	k.����<p��	+��YtM#�6U����A�Q=�ji�э���Y��(]K��Lޠ� r���Hi���R(Ԇ���B�EȻ���&�F�EFB�%4ܻg���9��8ő�	R�ț�����y���n��SE��RD7#�TM�iӼ���%Ȩ�29H�V�碹�.�	�|C��ɰȡA!s�D,2t%���-5��<����(��a�4��jS�`jٸ����g���6����C�
�J�/0��8o�̙�q�)k�9[�AϞ��MS�QQ̐炷0^`��Pc�R������â>�����,d��at� ���^�46��Hf�,B]s
��}v����/�COUX<i�.�u��,Oz��L`ޢ4d���������/B;=��Y��o�Af���U3���Q�X4�0d?�K[O�IFV�@r
�jg[�<��IE8�'��a���M�������#&Hl��,dpF�i�D:��Z�|1����a/�l	��{ɊR���;w�E�ʲJ�E���2�V��T,T$ҿ�sТm!�3�[��oR�v���6�+�����'�p�B����-�'!W�� H~a�e��[-���m�MC5��VR�v�؁�l�-w���v�?�`)j����̝?G�lъ���~��d�j&J��"v�����5W���V�p9���qF4w�E9���d�g�BqK�Z(1 ^����罿�`j���3a�'����j��'��M�����gR���ZܷG���?	�2�eá0Cp�zdGF�L���ц�H(%��m��EuI&:Z�M�H_2���ȄiYe(.����
��0�C�9�����N-B8��!�%L�"���IH��X�'��Ƈݎ��
ݸ�.��?�_��<�HfH�%Lz��Q6}�ym��M���.�E���4��˷?��h�DphU�4�.8c�7I��`�SPYU����jj��4�֭[ͫ����f�%7���٨�x�_DM�P�����*�m�N�VuhuXB� C�4TZ�{��v�i�7ir���Ɉ�����G�"�W�PA3�J|� �}Zw�:��H�䥹�ֱ�����W]�ė�|�5>��M ����.F�k=WǬj-:���ڼ�r<��/mf=F���sZ���k�;'�\�������c6o������6���oL	v!���$�/.��P�KH�$�3-u��O�$��=Yd;qC�o����X����lz�t��q���ӗ��7;v¦ӧf$ӣ�A�tN�tb�|z�n��JNE�| )������ɕx+� 6d��7
o�,�/[�do::{l�ީ��\x�+q��'�_�u��n��g��Ϝ�k���� ;����4��^]�az���*�>����_�������*g`�?B�X�Ј��-C�G��C��H�H�q�X;��_��n�Gxx�:�=Ry��b$T[���'��\��Q�]���0!^6�{^�u�����V0�K�X�
�-2Վ(�";�s<�������#>?�rM@AY�4z�U�O�-_�͊�jԏ���2��=���o8���w�܅�������bղ��ƐE�v9,�@ap�<B��������>8z�H���n�^$k#�tY��4�<vp4�LF�V�Ak{+^��o�u�Z��[���眇^���F;�B���$<8�o�.��ɳ+K�*)�DL�"6�~�*���:g5d�/�#��!���2Cd������W�W$T$���m�u�ҕp��=��Q�������KO��Y+�H��IG��ic���!��9��Q�|=��;�����~de�(�yJk�ѫ��E�u�Z?ш Ġ9�娝���ek�Ar�.�Mq�a�9p���H�+q�H3�5o�Dؚ�D��),~�_DE�,l۱w�u7֭?�P-y�<̞=״�vr0���Jd����Y^�&Ժ�g��ѣ��{;�B�b�
̜>Q��c-�ġ �(�d�b̟;��A{{�VIό�E�J�E�0�HM[$�� �2;?����8���s�5|�F6��<�`I�Yڧ����b�%���}{M"EY���}ՕU�n�bTȱ��>���=�JX�0&���Kqq�|ӟBPUZ�lj��a̰���h��22���Ʀ/��g�I��j�����a񢓈6|�;��s�dƧ�ri�J{�}��p����NL�NaEm.9��L�"Y,1���L�"���qVR��bXm��	B�˕qM�8�����d,=�5U֑�`�X�l�d�I�oڊI�Q'���C�8��JE�E;�R�)�ҩ���P�n�'"����0q�OAyI���ҳ)E10B_�Y�"5��q�雭�DDP[42Ȑ$�LP�W;�SH���WMj�0�>3�{=�)�^���*����/q��'�B(�($�>���>,[�uG�ȴ�X�p*�J��=a8^�+N��Z��4����*�,-GIY.m�Q�CoW�hK����p��*��N,N�0O���ô�%�� +�-ݦ���8!b�=͞��ɦU�ơ�����Z�c�Avn��|+eK�E;F�G�t'�:�����-��8s�]���E��\"�qF3�<�ԍF�ĕFx?=�r�h\��T;�R���G�H%�(�|�h��ee7��ktRqp|b�P�й�MUF)>%�8'�AHlδy!$M �s�\�/�k��!/GHT�� �FU�e�!���R�!>�����*��M��Qk�tp�x��>t�C�Z-$'����f�?��xV/����͑��ۑ�LF�H��ɏ��~zM5�EPX���a�vӓxx�L�D
_+m�b�l����6X�̧��6���砨X��
}�|_�뜜,b��xj�.���s�z[i����N��\s�&�Fh˨X0:JL��C����=sXu���D����b�G���H������������]gj��R�[�~h�_�*:0��S���a�(��5_�c�[ob۶m&�(���gBQ�?�B��&�O��=j�;f�b��D҄�c�F��dۻ���`���fp1KM¦���Z,�9�S[�mVY��l�;�$fUJK�MqPݥ�����E(ܗ�2��i}TJ���a��X���X�2yMW\qf�]��c�ƥ�yt��:���[9�$�5�W�'�FxbbrcN�G��ܑ��#w���x䑇g/Y���̛�<��@4� ÿpz�'� \�����������Q���<���$de�b�_1J��0Ҵ�M������k��D#��n�����j�d����4��x		x`5O�����ڀ�%D�P^U���l�9�.'�L�r~<%�^�^�{���P^y�|��!�vgf���~��k��M_�ͭ]����y�mԼ�fzc�t|���������_eL	�v�z��n�n	��{��E&��>����^K��h>|� ~���h�}����;6�?�j9�!a+����b~G͌�oF��-�Ev�57~p�>�\z�fS��g)T�h���m������q�:keѲ�ΞNC *���؜0����F����!P��^��*�)r��;ɵ`߾�i��M��^��15ۏ�������������6�j�`�?�ѿ`)��%�^i+�Ba�j�]�^r t6F�c�I6t� �e5���R	K����ѱ�,ӂ;��m����Á{	�+�m����۰|�2l��9�e�Hu$�l�]���&�%�4��B�y y���&���V0����ni���}��>̃Rw�!���9�`��q8�z紤B���,~	�N���� J����� yn̞Y2�� �F'�k�扖.[���P@j� ���Q��?���(�/CQN-�\���B��N��/��u:��'E�5�v�9�'�E��}�*K����W�x;v|����mipd�"��Ou���w�6���C��?>i��~mSb��V��pќ��-����G3J{���Iǵp�t[�����Xu��K.�D�����R�ݽ���[�`�R�42q��3-*H���'��5���/~>�:�֮ HU[[���C���<������
�T�"�s�<M�4��h:{9yr7y^6>޹���1�乐�N��%��m$���wY�x�g�;̣�p��$
�� %z��>��~=��a��D�����)>��ZZ���iތd��H^bΏ>݁+#)݃��X�h]���J����PV���ɱz��g��������JF��<�uğ���	�n~�q2ze�=V�w�1'����S���(��s����3�e5)>B�B���g7@�4��!bŷ^|9eį�Ҥk_x�P����cx�ݦǩ<��d+�ky���믽��.���	�7w��ւ��~���t��a}�Qk����
��ꫯbÙ��{�lz��?���ڼ�I�F��'�DD5l��]����,*�6*=���^������0�˄�+Gh^�����ƽg��a9kn�-B�aZ���K/c����$������j�[J2n�����K�5��\ځ������[�f�r������OIV�-��B�s�����o�V�M���Y��9�7�f�מ�ý������d�gϨFg���˟�x�*�{
�Tcp���S�xUR�^LBJ�J"�VN�����v'$R��Mw��$=M^������74����XJO��[�~�����!��*\�Ԕ 2\��u��z�H��B�ԟ�`p� <���I��5.Fp>�p����Y�ę�B:��?�e�T��t'"������Ƶta���h"��6�=�0<a����1�A�\�3xC'x홅���C�1�հw�!\/��E*�{= �M*qm08�W_~�&�2�ҭ1OU޼���d�L#�%�:����q�.�p��z�_z�%�v�?���1Lm#R�WdN��Ё�;e4�*6c����+�`ӦM�UQ�PB��g�+*�EP����99^>|���f�6���oiUɡ�Ϧ���(%��Ov}����0Ւ�476!Y����]s�β���Do}m+jg�$�)YAG�K��NO�g���Kʅ*ک�"���aSI����{����f{"F���R��Z����F�U�z��לe��	O?�[d%����?#��% 1=��/�����Ie;�Y0�<�.B���I�&���ʫ$e��&R�1�UO�B~vR��ۚ�� m_��O!��dOH�� ���m��o"�g�����u�C���JRJN��dB�8�v<%�F B����J��F�f�碳� J�$ٚ���&���{lB��jDŴy�.iE��<4".DSq�p�	պ�J�U��wiI*Љ��R�5VP�liН;��@Y$�ϰiE?=�����pzcS�qߨ���i^R��^��V���D_m���`zB����ڶ�r���j�&�$���NeZ��G^Yj�1�d2���+:�¬� �����Ri�����'#1,�(N�X�2�~�<I���bX��D�ڵ=4�g�8����h��(���@O�#�Qia��%YYƈ��aKWix�g�2<a��:`��t
�~b�Z���D�M
���(Yd�E�9�'����OU�52���;�y��p8K�^�}��iU%���f�a�T�Q���2#­|@�1� �Ӻ�m�Y%���r����9�&1$J
=fY�IrZj���uy���n��aN*Ն��#�]�֎�-�˟^��?	���LCw�����W�_[���ܗ�y������E����64��1����;x�ڍ�hC:�V�qYPGg���Ղ��)O�,1PTRe^��3!^�q�䤈�,��f�أ�ʔ��{����USڔ��y�����WPqK� �=Tн���H<4�� <��E|]�Z�u0<YnK���i�ڋ��x�zd@���܌s�q���k�����4NE�N����R��L�F�KL�1��	��4�,��Fg�}��y�m%�Z3�mi���(,������J��MJ2)>f$:B�҄^����!�����N��sؖ��dw)��I?�E������S��Պn�oa��&&2����)�l	��������<��3����x��*fX=��فOv<��l�nGyp�,��P{`6���̞�9ӗ���гx��?�����}d?=��
7V������^�<�����Ə���"D/{�g����j���CIG4��\B:r���f���H�*�y�2L��N�9A��t�x�W$�>	�����6�C�1����k��O9�C>�����h��x��4�T�T��Xn������-�Zܷj��2� I�s������yIq	zyM*0��mje��Y�{ZYQAs"e�<��߸?�������0"#:&�Ȇ�����7�|����Β����:{��5!�I$M�����|"�S�]F�1]�6�ϒ|����K.��7_�[�.`F�(��ek{֜���[�9蝥}��r��W���������}rl���$>��F�'��.Kx{�{�L�^�2@!�]NN��%��Y"�[�dS��2�D�K �A�zt䩺�����(��HJ������/�
�cO��u�(cƢs��78�BO����!ۄ��ӋO��`��K�~�:A�D��k3�!%-sg������?} 3j���X�0:�i�7�z!1z��D�[�<��_�b9�?����y�rH��Y�ԧt�全�����NaYȓ��`O���f<���G��T��-EM;q������OFSS�y=AuI
����{���܋���(�/�p���RnFE7�`�����)���./�6�=�|��>"DH��!�BeQ֝v����㝕����W�EUO�5	�ǟxºF����#����r�Whl��9:&�_�l^��^n��6'������Gݫ7�|��0�*z�Y����sχ���ǎ �塳J6M"�6�q���M8��-M��4�i k(A�5�x��7��O<B�ic�#��\`<���l�^������dJ�	��AR�r��(v�35�xT��E�ڮ���M�c���!ģ�T��civ��.;=��KR�D�����r;f�_���#=������+�i�O�3O��k�y3���������x�fb�\b�vx���P�(ʲ����v�����PIR눢�)�M�\�ko���{�^y�2IR�v�S�M= ᮨ�������(IX.�6q^�t%ν�2r��k�],wJ�&���m��ΥW�ì����O��at�^.���PQQ���`ͪ��$�%�v�yѮ�l��0��WY����"	���;h��gL/�g<�Ľ�N���r�6��Y���[�b� [��i�^�:TO���8k�R�H��#�|�W���g?�!��ѣ���bن�X��\��)������y�b�ר*��|ʔ��{�=k��t�E�η�\�lmo3���-E���OF��g]�W�E4[�H���5-Ʋ���ۧ�R�I�d��6L� %(�jg�С}�eG�w,0��+�ш�EiY�ـE!����fFTDY���#�d�&��:ty��G�'9���~MJJ�!��g���3��&��55ڃ���˰�;g�JSPC�T+<B�1f2�m<Ϧ���
e 2�s1}�\���Z���c"����.e<�j��a|�?E'����~���x	����{!�Ph�އ��C��Ko6�Nĝ�閻b;��ӏ���EqI�io:��㪶o5әHč��6S���[q�闢������x���8��z���R-ߎn;t�nt#w�`媓�f��&��NR\�_b�+V�2�������3�0. G�tѦ�ɻ�,�)C'R����<��s_�0֝~��B*�d;x�Z[�ͰD��{�2�!Q���ݖ-�X�럿�m�y�!��NF(���ȴ<���4��;�X$?�g��-�W��n�kX�},`�G!�S�T�4�M��4��4�@V��~Dg؀��x"}�L��
��v$������0?#�f&	���8ܱ��폋M�M���7	��E�S��{����Su����j�q�4�f뷷�h�u�:Ɂ��L)�n�����8�����N�����a
2r�Kx�?>��"13��h
�z0g�b|��cT��IH�f���p�TW"22J�Յ�8�?���7*N��é���6,^��9�&7�6��$t�v��-%�i Icd����4y�d�eų,�?��$�^�����r����2ܻ3�`iI�9]B<L��0w�b��1�'㫥����6��C�$��Y�1�V�X&Ԋb���v(U�UE:M�?��H�U+C~^B���X����ԡ��d<��5���g��{VQU�9�fc��Eh�1+âyf5��(&��e�����ub���A��Qb�����E�O�י���h��m"h==��I�N���Ǜm���"TUV�ȡ#&�����6�hT�[{�z�fL4����gJB�8jSz��2�Q��m�3�!JS����r&"�4��6����vUlu3���'���	#�E�K�H����2�bf�gl8��V� �k�XR }$Z��$�S�x2���W_Bݱ�<�Gy0�p��Xw��<�v�㑄�YVV�y>�̌�ք�ч��Ȧv�%^]t�զ�Zɰ������5`��إN��T�v4��Q�X��wԙ��(���ճ'������>M2yF�T�)�	��o /��t��z�<�w����a��P2�⃼�T��/� ]{ݕ4�!o��G�t�b[����'����b�L9�'�����3���	�����ߒ�.µ��@5�Fhuo"������I6�&���/ei[��F�����hk��CYF(���Q��O*#A��	�Lv��V��/��\\y��6�0����W>�V�q��n�G���
^�3�Z\}-�)at���/Y�o�c�G��x`�F9�c-�e�ؒ�������f	.��>I�]�z2� g ���+��j~[KvN�
��۹u��«�2����N"�=xt�G��_����l�dN�8��Ӂ�|[^߆K����"����?+�7��Y�/~x�z�z�����ol�Eմ���?�ͷ^����{�MĲ=�FxS��6ޘ�o������=ĸ����ZA_w���g��o���=�4t�t��@�k�c��W9'^|�14=@�ы��5Vm>�>��D���_|b�1���M��E��ô�b<��_��[�9�����H��ۯ����}�s*�q�7�C��[�k:P�����w��W�I(���d�[����k�>���{�_=��r:�6#��#>�ނ<|�����;�HR��Usx�q`�^�{�=���_��g�@���� U��J��3��Z'��jp�X�
�̘z�Q� ��n�����(��P��?}���R����0z0ov�x?؈+���ϩ�)i��,��(ǚ���+x�O�b��i()t5!�{���=س�^|������g��j�KJ��V�]u��ԙjT�����/H
'�W�:���{�2��X&�����N�2�3�H}M?��=ن+�U�UW��7�0���sk��N�4J�NbXUV�������f/[�(�*�jXo��/=�׹����cZe1�`�S�#������oY/�B�
,jK�Jw�'?��x���?l䭄���hj�?��Ω!QNE�1q!�67;/=�$���G�7�d�-|r�t4�a����� �j&����h"��e�����x����[:�`(���m>�-:ۛ�Ir1�W]��3�� �*J��/Hl����\s:���>�L2�����~���S���ɳR�
�����o�k�4ّj߭�
�CeQf�(����￉����g<�G�M�_Ww/>�.�c����M4�5�2�2��9_8�3���;�0o���F���\HN�F�g���L&�q�W�ž=;p�iy�1B���[L(XGn���/ҨSm�ԑ���x���!4*Dc� ��'?Ư~�#F�<��*�ظe�<��v�e�vЕa��5"�vN�B��ɡ��SŶ�MΙ���b�r:���:aC ��W�Om��j�1Qχ
>�J
����`e�&o�7�^X���o��15�ɑ$d�sN���ن�"/&�L����ư�#Ņ�����v;| �j���S1�?l�L����lz��0֮\E���n��i�;ﾁ�.��!?hZ�%�n#�Y���K�ܣ�0f��ۈ}_oz������2����\��۷~h]����k���v
F'T�B��(v���/��͗\`0ғ�� �k���̬\���m(-��@�y���y��|�/]{��0�HpxKJK��/V�p�)�Z,)�e%!I��!h��Ҍ�#G1�I�� nt���[ǥE�Jժ����!D��6��������'�vX;�'���˯��¼�.f׽9n��I��<(%�w��;�\B�Q��#yzA#��z�֔�NM ��&����Ä��;:�֖7q�Wn1���t&D�4�,��<u�Ö��ۘ=vL*XL�cq�)񃩢����x֖��T~��555�;w&� ֬YeJp: o��VbI5�l0�G6ayI����&4����b��Zh��zV�_D^�
F�I���H����R''�A�LF�ښr�ۮ=�<k��d�Xh�����0=g�v'��:�Ju(\�+M�f������a�����J�Xf��̨%e>*MB�
�ʓ]i���M�ڑ���Ho_?V,�M����� ('-�^mxCqy:w��ܲt,�|���ۈ��^z�v��WTR֨��������m���H``���FFR���.�=��Y�b^��,/) ��@J%)K#���=��G���ٳgы�ޏB�`-���6���U2����=q y���Y���$-��'޻��e��ٜpQa��8�	��H�σ¢L���;F�G�~~f�� \4�@0Q؂C)]'�����=�����1)r��HVR<����M�E���R&G5��9��l���H��6X6>nI�ى�Oi��|�$��NuD�ZEb�)�-?�!��#��. �� =�ǶTj!x�7/$jM�aKA���σOIH�K*��hh�|����ɋ��T��U<�p"�Xd�H�gM���{0���\�۽Ϟޥ�Q��,ے-�mܰ�Ml8�NN �ܛ�Óܜ�=i$�%��Bq�E6.�-�꽎F�{������_kK&�	���<��Z������SgX����i��S�*���N���LSKu&�,$�ABR�"�PB��Ī�l68�ϐbD�p&k
�*ӱ��X������e����q�#���Fqy���^�k�B��Tc}�$z4RUU��]##L��R;Zdi�Rj �ʂ)�<@�� �|��j�"z�z$�#J�!X�h�JI"m���U����(!�Χ�c�$��j
š$�s2���[T�67�6���,���n��˓� n�&�U�Y33��G��h~լ�MF� ��va='��"U�+*����#�kW��Tք���N$�tG�g6�th�zs�.�`��5��'ׅd��o[3��){���7�h�4�.��B�t1a� M�#����9b����6�F����[W���	�cƦR驐X�Q���<2=H6T"Q44�)˖.� t�x&Tʧ3*C�$.�I�&Yǩ2n_D/I�E�x]��*�������Q%9:>D�W����K��U�z��?�8������PD�����f��J2�j�9�ͽ�%J�06ɢ���3�0>>�~P���R)�ɼ̹�RT'��Pҍ�Mʲ�wѩ�V�[�`1;��v���̛������JR�\��454HT	���EF�L�O��=�����3�Ѡ�G�7e�1�9xP��mmk㡻T���U�!{���-�m��əs�Jݦ�`l:�!.[���:<ud[��,�푖�z%�Z�7@{(�J������R��Q"���ֽS�795M��f�%���X�ae*��pTl)���h&C@������m}��YЏ���/Y�&�캈9z�	�� ���C�$�x��ߤ��tC�fH�isC!���ѽ�裏*��I(���2G)��RV�&HHZ����5W��5A�s,؛�����)o�xE	�)-�+t,\ ��ƃ'�,GX�d�:}!��U���pLU\���E258���D
�DÌ!'�%ɌLI@?3�u��I��drT
�Mj�l��z٥�P�P&<2<IF��|202���#�^�!=�0J	u9��П�,������bjeLͬ��(�Q����U�4�e��E;{���w�u����}K�k*��͛eh��,���Q�}�n�I�<$��pB���<�B�E�>HG1�>LA��Wm])�u�4q�l�w���5J%���/<�Y�պ�ɹ�jo3+ �RI�G�/jv��|W�]1����A~�A�1F�}��)�6� ��j h���6� W�Y~􄃠A+�x��f����w�W�h���T*��U��|�3*��OO��HP[���{��I2�42?�rVy�U�]*��S��h�N:+���;;;��Ӈ9TYU�7+�T��>��r���R�,\�I�Jy���*y:�Mת�ꐡ�	¶�y|L���e+V�m�9�BZz�3{���+�(��GZU�C*�KA�Q�N�ǧ>���/[�\#��엧����P� ,�޺�rY��2Y�v5zc� p�cJl�_]}�:"�TI��{����,�4X� ���ʵk�$�\�ֶ���Ò�K��w= ?����^3�s$��J��/]��K��%���EZ���O-R���+(Y�A�ܼI�~�Ie�n�2����u��U�M�ġEbD�F͘>��;n��?�N&I�E���GN�����Mf!t���ibOy<��=,�5�D�	���Vٳ�+Eׯ�(�����oPϳ^�~{����*�7��G�Q����-��aZO6?%{R��"{�r�w���8�%'�
|^�*t�*0��ӽ�z�����_P�ʨ���9�����I�H��E%�=CJ4�D_����덊���u�^!�9 \(�0|��$ܥ�,+g0��[na��MJj���4���.���ݧdnzN�,�"{�����	�(�������m����v�N��)��T.���H�o�*�P3bq5	�V[g������%�:dy�*��q�d��e��ﾇ�״�Z�Jl`���heD�SM�+��Ns99t`�:�SRS��_m��^�N6nڪڠRטP��"�
jz0j&����7��`��W$��Sͭ�2ܽw~H~�OȂ�&Ր=�Db6�Ax���k䲕��w��ġ��B��M��ֆz���6���|n:��7#G�f�(�V�Y%�7nb}~T 9���g���0+�}���m�߭f�<!0�e��-��ʙe��C��e��[ rIp���'�����{�[ϵJ�v�vۍ�/j֌�\Q�W�3���ɧ�R5F����-����ɣ�q�e,C_�f����[Ș�ش�_��Y��7�Mi� �4���0��2�oALӍ�"m`�M'&��� ��g�/W���e�b1���jJ  `�����S��p�ͦ+�06=6:I`�\V���}DJ��ՙ�MRIX��9�:$7�_֮٬Ri�ݔ�]'U-m�2�����a�E5�\R�r�����KK�����(�Չ��K�ՊY]C�J�>����ʉ�g ҕ����;／&���Pƙ�`4�0"d�ơ�u@(A]c(�w�M�ɕW�S�E��QILԊ ��S�֎V�=?�&�W}��8�=h��^�\V.],���t A�dVd{U���8�Jh�G3=�#~��mٲ��2JB�0�i��fi��&V,
� U!8�T��d���r�>�:�����yZ��IKcC���ˬ�;Y5_���.gt.��L�z�<��22����ʈ����������ɢ���{8x<�-� ����g)�э#�C�}�xP��ti�0J�e�@;��7�a&_�XC2i��,���%3�ިf������� hL�lHZlN%�=���cL���R7@L	��=��jF�,�f���26�g�U����w$y*����"{:3�-.�������A�c���%��i5_<2	�͆9z줙L8e����E�a�����bT��'䡣��&O�T���B�����0JWM1��8�PҌ���I%���F>Si1�/S�V;t��E�&�qG_w1������s a�����545�	a�0[�𡣲��W��cK�Gԉ�&�0wQCЁ�^3҉MDL�Ç��fޭL�+A���v��Y'��Jo����9��C �%r��7-mif �<#G7�t=+e]�Z�|>|�>W(X!����\��x=�׍�IW�aj�5��S[đ�%�P��~��:�f3�:*qf����� 4`eD�����/2��a��˚��b�K��w� -`�f��&ª]1sT�T^2#�b�6]KI��R�������M���+#��8%��Si���^y��%�:�������{jU�b` AN�AU("N`��<��S�'�H*��z9r +�yr��[a��+�DL�P�ׇZ��]^{�Yy{��J�%ּ ��aӕ��oP��w(�:s�(�˩�Gާ��ɋϿ(�g�2���l��Fٰ�j59<D�ce��Z�74���ex�G����G�S����JOhM �]�e3˨Q<��O���~����'�`d��`3C*��_�O�@���͋�%���ꄶ��|���O}�TV�D������r����=w? 纆Xڍ�xu�@�C����=�3�9	!P؉�{�k�QG�.ֳ���e�V%��#Q]gL��N���_�z���FD=�ʮwv*sn0���'Acz��bN�?�D_�<�[z�w2`�d<�q��%ұl�:��!�=�b�Z�鶣��)�ij�6llh��e:q�K.�4қU���.��lܴAFa��F��_��|����^�<k�Ϟ?%�,ӳ����wd��eAs������0X�/5�z;�)�/�P�b�u��֩�ܧ�3+u��t�; �=G���!�*��=�TQ��uJ~�O'�,�C�M�*u��g*�u#J�66���ʏ����ׄɌbgVU4ɨj�o<��rǝ�˒��T�^���{���T:qP��ͯKk�<5���QuB'�;��gGdR%�ͷ��BD8���Ѣ�qd�O������Vb�I���;XK��'�����������c�u=* � G��/Y���&�K1��!У��z�A��_~E�,_$'O�UӢ��@~�G^z�yy��g��	s�fuo��NN	W���9�'�E5W�|���1�<77�kp�Uwg'q�jnݼ���U�gCC#�³O���=�}D����TWp2���Ӳdi����vy��(-Q�*VF�U�業`ƣ��sOȽ����kX5�A����
EQ^��M�O)�bAZ��A���5��L#�]�Ϙ��Ob�)��������-�S��s錠RkNl-p2�@[�h�|�O��*�k_�m��CT-��.�������\�RRb񩭯�-n�^�;{�]uN#25�pe�L�M�[�=�nd|rD���+�I���)%�0ofh�L����wr�=�H�ج44/"���؀�(1y{ǋ�PdRqm4��Qj%]9x`�Wę�H��J;@����e	z�W�L0�U��5�!�����/��ˤ��͔�)����SO��ħGU�;)���쏩�<�5(�ʇ�j:�z�Ⲁk�o��[o�cR ˜"rh6*j��ᐼ���j�4� �Ӫ:�,����Nd�+y�E�J����P󵶒�(�_�$�l-E4}
����}!���j�'�2��&�V˾=��_QW�� rH����8佽;�\��S)�V�n����VQ5�����*�p�6�M>�۳K����$�Sl��,fQ %����zkW1�K8�J'�,bo��0��&�i���L���a"It�]?p��?@���E�j# �m:<0.}=���m^�mNUܤ���+��\)I=H����~A���R\�"?)����-�R�JB������RɂA���z���V�,Ɇ��Ɏ�vɶ�*�[/�)�d�5���/=-M�a�8��(���%��P��HMeP��#7o��KWI\���PN="ݧ�l�\p��*-=e���9����ޕ?4O�p�Q�4hp�����U��	J��tR!��e�V�_y�M���[e6��D;t��I�!�N[�i�[����gN��"
�o��o�g���c#��7_U�>LL�&����R��_�/=�g�{(����Ԡf�w��8��31�nql��A�,�������Ï|BM�!�f�#G�ʹ3�Uۇ�����5� ��2�CVF}r��Qi[�X�x��yq�7bP�7������V���B�ݐ�����s����s�Y����BT�,��]n��j�������� &��
B{����ۂ�A�6�/����@o~��vݧ�<�C7?*�z(�u-���d��wd�:Ic#3�TWI��p\�~j�����f�!�^�@N�t�{��!gϝ����&���3AgaZ \��x�U��j��$70L�3j&,,�٩��㌫@ K@
t��Orj:�1����'��$�����)��0;�'�E!_D)"��]��%TQ!�Ϟ��a>��P���M/0)��!��~O8 ��jUf>%�Y����`w/�M5ڱw���f |�~�i�5Rp|z�ɯs��ōp�:�+Fe�L���5��G^?}������2p�p�`O���
cmQf�gl.���O��X�-V�%���x����Jk�g�f8[�=��&Tc�6��D�r� /�&�̌�kxF�&&�:Z���-Wo�HF���B��� �;"o0�1"�K���$9�ΰV�@�
���ϰ�À�yO�B �d�|>pɌ����Tjvx�?�~����HH�ޮ�9;4J�fP�nZ�� �t�H���[m̚���%�R���@��ͧS20��J*��:b�E�j�D�JLJ��c�J0��v�����C�uFeb�>-�s%�g�k�#>�O�A9t|P�%�
�L&��?1�z�bM3Nu�fd��i�Y �*A�[Q�� .uP���X�!n��;��l&�v�S��u�|��A�K&�dEn\ttdB��ODp������&����M����`?�s i./0ΏqO��������0��C��U�P�@�i�������YSF�(���(�d$Kr0	� 3�@����6lk��Z�2�
�cu��Դ��Iʯ�������Va0VQnг��0�d��b0E�ʌ�/�cy��o���9o#���U35 ;w���M�l3��e0J0�h��1C�0��of%�ds�����`��t��D�е�.NGTq�\:�r�K��҉H$����8p���sg��5�l�kL�DS����v��*��\%7�x�����r��W�94,]tD�����,��._�x�J��G��)�1�YU��9H�<��
@�v�E26�Z�XM�Rt{զ�Q:!�;�2y��?RS`L�'��7�%5G���70'd!��|�JW��5�͓��	�)!E	A}����2?"~%֣'O�#�e���F\l�Qb(G,1���V�w��N�PJ��wzbJ�����$ e!����>(���g�)Q2�b0�p������z h2����r�-�~H�����D�6G5��X��	���j�^���l�F���M�qD�j��]�l�l�YՀbA���	�1�{Эu֫=��sAV�{8>6���[�T����:�L*z���M��߶@ͻ�f\��J�>˱�d��:�Gl�K3D�
WhN6�c2��!���NR}��<QE،cU��e,9���I���tS�yMMN��dI0�'��Qd*;d�ڵ�Z�R�������J��/ɪ�R]k��H�LM�u�*��n'��e�����R�#<D574�H�[��I�H$�*%*i^���OJL�����#ʖ��[���q�����ڲ��tƽF�Ɗ*�J�9���d�שI���>u�����m�|�s�+����R�DՊ\�2�f�_����t��;>�l���� a�"��~���/�>K"7{l1�&�*��*$�}��_?�(M�7((_���,_���#�<"��z�{�����6��|��e���j
M��1r��(a=��9����k�(s�\E�1����� �&�ԩG|��n��M��>����K"PFs�x���s�**�ifU��SK��5���o_���ٟ��t��Y]� �T����浩�S�Sg���џ��;�0wTCg�Y'o�f�j�)5������G�U�t�d/:��޾@�	 	4��G�,@dش�>d_4j!� |%0L=JV��~�VM}Pekk�o����[�|�)��U%��,������c�=Fb@���(�Us�[>���)n$�?�<��n��n�U���V۳�2J)Ƃ��F_w�M��K�ʱc�U�֑�**�UDu7Ȃ�K���!L���cSҺ��~��nd?��3�T:����0l$��}�A���;�O5�#)р0u�5��l�<��y���	U[��8���n����HT��j�V�j�C��B4��}���~I��տ �v,]̈$1�0�qyt����v�����qj|L�������f)|��1�DʠH�XA6_�En����g�=����G��~��!!LLN��J @u�TM�G?!���w���H�2ΐ�C��d��7]�(VZM#�24� v`Z2���������Y]��E*YԽR�k�<��do��L�� �cFDP�WI��k�ɫ��̞��I���1>1#m��>	~����;��V�����Tfh�窩��犬q��' ��,�zn
�~VF�'�B�4�9p`���]^�����~���;�"�"��]NG�@:O�.]v���W�����=�tV���eA�fRc�"�)'C�)uX�%�~U��]3�0+��[�f�t,Yav�Mq���wI7�3��1��^YۻVN�>�C\�j����.�VI1�0m�aw��N.�X(��r�6�-��������ÌouM-mz0�8ly$}Pǃa#K�������d���W�������a�@�9G}��p�y6o���BP�j���5@������Q!����(�����|��Y�%�0W�p�6��I�ɘLA�9iz���_�[>�a�u��o��m������q��jeD�R�JG( <�
�]���cB0�`v-X����`��>�N��(���o��D��p�G~�>�I@�(�Y���)�N5={{�3�"��dMQ&�h¹�Jc���$8�3��B��FeK�Y�5?�F��O7͋��-7�&��{�`oy��La%>,��(�&�m�jv.�I�����%@�/H�7 [LN'uC��HUs�C
�>75��%ϥ�)���A6^q�;��(�k�	�s��6�~���!�R�%��%˥}�B,"�3<6.��@]t����Q��8����y�a�fY�t�� �i�v�
��	*�j(��{|��:��V�\#+V��-X������`,z3p0(�CB,ɥڂ-�J�����@�VOҘ����3�{|�?s_��GG[cC3�����W�
��${�yO"��g��2�<5�,�y�G��[[�h��2��+��p����n��֊g��� �_D$.�#x��PtI�D����<<�;��_(�u�0qhvր ��FÄO34dN%FG��f����;�Y��J2��0h����nw�I!���M��Y��]	�{�yx5~]hҨԝ��kU	<@�l.W�`HmC=��\�R�����H\�8
�����Q�sv����H�|fv� ��0#�2�XH�AJ�3�,����x����$Q��UՈ>�Ԭ�� >w&����G�%G� �B@(ky`B$Ri��q���[FGk�� &�`M]�Aϗ�u�'N��}���Fh�4Q�3�-�RD�@��5 �~M��x�s��f2���c6��� �Y]?�
�� $�������aqN��bE/���9j��"B��aL���!(�#�n��p��4�yP皰+%>�{�07�]1%	Ql�������`Ϻ{��oU�5|��̽t��Ē!��.BàtJ&���w����e�x�Q#�%1BN����&��jd���@��2�U�A���aJ�z�kP������ǒ씩S���e<�Jqp@m��$'��؞?6"8�FU�����	 ��N����q�0��qe<Ē����"T��Q{�v���֚�`�BPm�@� ;��z ��,5Nq���#0�]#��0�� ���IxE�h�8AX�
�^��81>N�ճI+�@�E����w���'�P�T����I&`a��>�a7�÷������Y�Y��T�lG��(�Ĺ��4���v�z����\��
*����(s�b�:�,�@�D},"N�,��S��`��Du3�����&�(Z�+OU��Ŕ^�8>Eg���)$�2��7V�f3�R]�a(\z�&�RM�w�D���j���ly,���pF��!��z�w�� �A��nR�i���� ���u5�ah9D`6 ��`�*�VC���1�gP�%:UsCA:[��#���@���K�Z2g͞��đHb?��^`^������G�'����٭����}=�I��~H|j-���b8L0Ըj&�m=j�є�AtX�'����IJ���r�/	�"�sb��4!�1��E�'?�vú�c!=��Q����U� �kT�>_�S�'2�^]����ա��?�*���dg2��ܥd�
���G�Q,h=��bt,�EȜ1��E�	��`�4���.���$Ϡݝ���|�R�L��p6ikTB�h4�[@q�@�)���}`����$�n�gU�aca�D����0KZ�Ŭ2��C/Y!.���*����p��Y�2\�`w�qO���u��T�T�bVh�e*1���Ą�K&��qgɪI/��>oI"Օd.�}�
�LRL�d�e���=�cw���B��LZ,Kg�<�)�L:�wD#⽠�P���rjd,��67y��*��m�k#��L��6{p�6[�bUfڵ�0�\Vd�6p^"�C�3R��ϲE�5�>bVD�i�tY�� f���4
~g��Zё��Q�a`	2��9�y��nC�Ng�8�%�ȟ����/Xg���s��>{,���g3��}�)��Q&�3-t�vD"VU��ً��
H�$R칸9�]AL��u[^R�ͦ
e´7�\?b��a�SB��فg�6��\d��񫜟��e�Y�fڟ�8L��j"�����8h�������@��ɂ���h�����ʇ�h0G`������#@c�0����s���(��S��5�a��X~w�ALr�EԊr;c�&$���0>�*j�|�AM����#h�y�g�c�߸��C��4�_@�� ���ɸ)�3�NT��,��_iaG1y\0����"�k1�.EC8W��M�����pr�#pߩa�l+JKk5#�B<�t�K��}�����5�Q�Sp؄b�nہBi@I��0��B�q�^�ep���a5^C��*�d6��>D ^e7l�m,�@N2`s @3(��GD��Ļ[�æ:X�nKA�l�)Z�\ �y\���5C'���S�b���벉�F����I��2��3�?d�/�x�p{�Ņe����S�~c�����]��4���/��6c�1`��߂�Ρ�!�{�)�J�w+c�k���6ҸdȤ\*��ۃ�Y�K�i�(DV�q��O�~k4{\dO�P�0`h4F�j�N���&����X���iZ��jN%�b$q��A()5�� { f�Q�8xζ��Qi���q=yH�,����k[b	���0v]t` ���D�CL��{@��3�A�b�[B��删"�j�NKes�"ui��)8O�:p�A�������:4 ��RF%Kڬ���|҄)�6J<�@��sZ��%�ctcT0M&o���A@��ܮ������[�""�؆&�Y�YY˴��`k��iz�Mm�A|�}����>³��� ��`��9�2����<�#Hw>�4N�0�b�G�8�bm�y�*����n�c��s��0��h1����}���3-�{��O'-	��?v	x�v��5IeeÒN?##�C�9]�n���Z�i��:���.��fX\ɘk�e��%6��Q���
�J$�~�uH���$�e��LSr�	�����h�2����"���{��=:�a5gɲ�/lb*�����bN�%��ږ"��^
�f z��.Ʌ���Y�\�����$N��F��m�_Wbc������x��0�ՠ��nXO!W�L4G�0����i��b�B�^K���D��辶�q�/Xʚ�໸��I��{�$/��Ͱ�ri���[Ʉ���D�L�t���l�x���s�fg4Hڅ����(Cǽ;;���r�J�	\Y��8d��O]�.#�}�v:<�A�4���I�:��/5S7���a��a�Z8,��n8$��Q�¢N`�9���|�Q0�M��a�rem�ʤs��&�>�4��gҍ�FR3�b�N8L���Lq�-y, �������bC��o=b�5@ =�[	s�6y�����ht.IQo���oi��r�3s�;c���!�Q0���d� hPZ�N�˄cK�d��o3eQ��zʄg4��{C��/�aU���00>�=��4��qm���tY��<]ֽ��r]t`�|���:�a2��/�H��B�A�h��Sr 8�����
�G0��`@��^b�H	,�+�*]�v� ;����Gl�x2�Y�����h֨M4�;MU��Z+Y��F.Ƽw�9�I;�S@���3@��av9-�c�n��d��&����G�� ��h1��G@�����刌�F�>´���vN�����߼!^��Ȯ�h
f]���Qފ6��.���~��8�a�21!�kEz�Y3�
���&��%���8���#�Rն�m;��\.���mk6?c�%���-�7�d�Z�:]8��y��h$��P��Hۣ��H��lʙg[M��[�IjaV�r�KW�g ���)q�r:���n �h������P[[�UG��X-�F~�#�)Ý��7Gυ�eԶ�bq��'^oy>���Y���� ��D��J�yT}E�p�~S���r�T�s���Q�!�p���HN*�b�L�{��~��yӷ�&�[�	��<��WF^�!��8����L�}�vӌhl�,�Z�s����!!��P)i���D�\��h���:;�&KN��Ŋp���g9�H���"���I�*GFl=���l9|� ?�t"��4��Ĝ���U{"����	0X���f,Jqs�!2��ꔤ>�����$�B�SC��$ijED�ް����{pc���M;����Ԅ��F8�=@�I d��I֥�.���gߞ�޻w��	���Bʲ)�������p�O� SL��I|�`���o���fc3�W&��b����h��S&!Z���4qt�dvz��;�
�E��W�\Vy��,;	!0Y�J�����!����*I���w�ҁm��u��c�DcC\�o��2k��r6�&���$�<d��E(F"�9]��/DD�U��41Q8f��ơ-4OM�#`�{�^�;�2Y>�MĎ�s���$1`0��0fM��̸�2"���� 2h �L��D�`]�M�h�>
8��mɘ�^"oX����nO#��y�`���~$�^��������*�f �j�_uEm�;��qp��2%���3{U���n��=|�k����̳�|*O���PM9�����%��03�@@���%�jUU��i]$^ ���K�ԧ��"\<\�ryс��ì�J�V	��.J�,	،�-Z!Nض��(K<X,V@�"D�7��<���5��,���(W6�T���E��M�p��s��΄�p1D�-G�p�=.k����~���<m|��|~� ��3���ޘ<����U"�A���B�pҤj��.+�b�A�`���4!qH�T2U�@�0Z�*�@�KK�Bh� �R[Žu!jXppx	��LL��v�a�PzC#)�@�A���|~	� �,�ߦ`i�$�(���k��Z3*#ސ(5JF��RY�,�`C�ң�5�!�*dP��|�����PwP˗��V�X��;v<�H$�a�����)yr���V+�AJrHH�,[��p�+��&T%f�	�R�vX�u����&�__nas3u.��,��)��9���`�$	��}��
F��IF�=@�F'pWY��LQZU����2Q��e��M��0Ȣ�P����(.;z���(���XOP*C @&a��ɆJR����P��v�!��)Y���@{U�V��`��N~-��h0��\̊��Lx��D��@B/��dh��`ޠw�ծ(�@"ѰuQR�J5*�Y\���
h�l���Jscn3�����Ř�VH��}q�\:�jX�'�` ����H(����$M�R�O{|j��|���̙N�AmS#��)��	y��=�.Q}�h�+C8���I�#���h�韦�:::�:t�x,��鉉(�Aq���\���<�a � �㝝��[��ZZI��;P�f��ܹJmi[��B�)640��c��S��7�si+��a���#G���(i@X/OX�
%	lY���@��!� �2�N0��MiA�3���Aj�9�
HU@�� ��
'��17�=X�)y0v4P,v!�R�����x�ɚ!�|�jjb� ��F�+�A�V���Y�fd��&�`�r
�ה]8�2EtxUA��Ω=�``��F Q���8x� ~x�W��a�"�c��AVς����r�F"�'�s
LBy�2���*�9f�"�Q�g����655F�Č�8�W�W����(9�Gs��*�U���F����sD	���90����Kf\�֭{�董ߞ����]�Ci_�@֬_#Y5���8��g$�t�Y��$��W�����t��%�䵗ˑ#�T�(A�j�V�~�� h����Y� (��j���"R[&�"�F� ��ۧY%�Ϟ�����\�t�[�;�\�i���Ijbz�*DII��č���A(��f�+ޛ	E5�9�ݍ"���Y�	��?O�5&������3$���&b�ɖ�H������|�4��B�$|/0$�dHW����ѹ��mbB���.�8"S4�l�{`� ���<q[[��ņ���	���t�"�n�{�]oI}C	���@��ei�p@�f�2L�����m���%f�����kxU�n�b9�M��	�_�XEs���yik_�^X�eù� y�p B����.�쮭�U��O=n6o�<*J��_?�F(��>���GX�a�`L�<�\�L#5�uR1:B,|l���/ɧ?�iv��r�n�<9|�4�կ��ɏ�ú�Ͳd�R?|�uŬ_��A�b��]n��&�ĂF!�OŔ��0q8�p`�o ���je�	�y�w������lK��f��r) ˸�	N�q2DU2gi�$sh�5���r<I�L� ����V_�<�'�,/i��Al�ʥ��$�c���Z�t�3Q��ć��	p�7`6��C/�a}(�%���#f�4����K �W�>?
x���K ? -�/د���E�����Q?;�BD�� �;�	@^F�� m�<�����>��5<D!oY�^���6�/�_ AeldH��G�
D�+(u��ֳR�/��l���&l)]���1B�Q
@ Z�z.©�O��'�廬c_ޱTv��MG��ϣ�oϞ}��s��C}@|ʡ Lr���ԜA;C#�+Uh�>�Ŧ�����PPc4H������^#�o����9³$p�B4R��(1�j8G�C%�9���(qO;�I'�T��q�#S��a�ä@�����λCR3�f���Xd��kl13�����g��!�ѫ�`�'7�	8)vk!��"��$�&@�Cw LS�(uV3��`0���u�<�F܍�z������G����6��I��lij�gN�>�}�{�u�q���^�%tZ�o�ۄ>��Jet��ggdtx\�5d�0�"��k�J��,�.�c]����{�I8��E%�f�/\-<�	Y�d{�zfx� ��|��x*(9{U8DU��ͨ@)��Bͫg�s�M���e���9R��j�ɰ�_�M���V�tN��|3�n�ܮ�{}��X�r9�%dS���jc��H��>���I�������Ɵ�<�J�e�tT�!�j��I�S��o��SM�#������%��)���׬]-�l���WX۱c�h�G��5^q�4�`������H[M�� �3s�+�k�o��U�s���
B|#�@�/�X&G�e2��,����$"�5j�2�A5,�gߞ�,�^�~=�`F1M,�A`J@kA�y�TA�&��k��4X�P(4+*�9ZI͋���L�^�N���ֆMB��D�~ۼV�3��-Xܘ��!E�9�k�V��ٹ��\�XjTc,X�P��v��z&��3c�n��N"�|'ɹ���j4OQ�| *��u_#z�,��I5�Q�hU)���2��׬S!������0AR3��K�4K� �>n���?�~fF@�����Ib�'M�@WW��_V"��XL���=����P�>�,SS齽{�����Y��N��xρ��'���L/�Jȝwޥ���8D���8N���Ɯ ��0�\�~B6_�E6n�H\Q8z�̧���ke��MR�(Ϙn�c�y��wI|���s��:�Z���Mc<ʯ�~D�<�,F�����w��a�a�@�n�z'�W_	�_���(���#��~���v�Ю��Q�`t�CP� f�]�u+��3���e�d9��
��<�L�ƍ���U�Y�{�I�m1�B��硁a��o��nذQ^Q�	9 �]�T�~Z	}VR9�S���]���+����E�4�k�g�>��1Yu�R���JP�d	n�x��P�(0���8C��<�Y8�!#*LjZ$���� �=������\�r�7�)��Z������<
��0�V._![�\i�R�dH�7�x���:TR�o�G� �@���MG���Z9����{1��A�@tسg��|�e�	��L҉�QaBY�CK���?K��	L���P�8`͜޼��{���ٱ�D���H�:���0����iU��vw�=��O���w�T��.0�0�����/���@X�Bs�&�4�#fО��s�l�|�;���Z���Q	������U�_��|3�֡��կ�A�|�?���yFͼ%RS]G_=!/��25N�h�?0_<��[W_�&Z�,h��	; �����^jȅ3ҳt�j�5S�1�p�J�^R�o�=�g�T�A{��~�5�r�-S��'/�FG��-I,��:���$��s�].���o����7e�[o���po��G{#��6�&Y,��X�wȡ�����3'�mP�p��w�ɽ��8�u��!���ۃ������7��2��zp��C�����]�vɻ�w������5K +o١��٢&ǜ��l���Z)��5=����l��������>��0��6mb�s��l�Y9y�#��6l"�<u�<�ρV 3B�A����$Г'O�`�<��7~oW~���O�-��N��ň��\��Ѭ �B�P�>?��S��]4�p��2����!����r���*]1���A� &vù�Ȏ�%t���{d�޽ A��;Ьb�?��z��v��ۮ�^�\��	p2`Z�Ͱ �߫Z���O ]C��߿W���3Ǐ�y��۷o'b��`~�&� ��U�Mf%�F���(��w_���埾�-��3� ��x�|`������O��u��I�ɳ`b({�P~������{�e��,`���d�]��Q��Q��"ygכ�z�Je�&��C�����8cj{4 ?�i�K	�v}M�n���DC� ���>��m����)�}�~9q�$���p�����քJ"�T�@�0&\եz��t����ٳJhQ���d|d��F���ˊ�Ketd������k�:�D�� TP�
�����<LdF�����㍷����˗ɧ�q��;���LR̫	�������˖�qzb�N3��P�Tg/����x�@�7�x#qQ���E�+� S��2���+/�Ë����:��De�WH�n�x�~`0h$�@���#��t�"�� ����hb�V�ZM�	{G�4s�U�7_��*�{��ɷ��M2¤�u�|�Y=7���`$.����8��ڽH6�ō�΢A�����0�:T�]��C\���ƨ�������*3�*����x\�b��%?�R"�3P4�,q�~��E�p�~]@�8�=*ж��T�N�ا�]��(M<��� Ã��L�Cў�����i%�Ԥ�d�zp�v,����c���0v���z�
�|�F6�#���#_%;T:���<$�pį�bL��nrX�!K鉃��ȜUO
�TL�L(s��C=$_��_���GeJ&w��� Ni[�R�Q� �Z�j�|�Pg�5&��m`ZAZa~ ��]w��P��>+�}�$z$瀅��|�E}X�}�H����s�<��(Q����A�,^��C����W��o��'y@�'0܏R7n��0�����$x${�32�?���[�r)%?��˕`���%8�Q� ��Z�'z�AQ%�~�"(�y���W��[Y���`�Wo-q�N��$�RB;�������0�$����o��
���n��N�Ǐ�	ݛf5i�*�'�{d�l��nY�Rf�)Y�q����
�R��t��"#s>_D^u��8z� q��R�|�T�@w��{:9�n��g����k�[����h��!Zݩ7����)7��g��_��&�Tw�����6o��%|�R1�Ü~a; W ��][[���Jr��?�j�=�&��-|�y�8�o��LT��={XJ��������L���� i�>w�<�����a�����'��	Y��U֨m���x�BS��5 �:ϝa���]]ݬÇ��4�^`���!�BF��Y��׾�U���+�F��e"(#�H6�3���uݺ��7�4A�(����"� s��d`����h��p��ٟ��Ҧq����X�K�Z�x�w�/x�sʸ�-�~��B0=#���C{��A6�]'��Z�����V	�����d��v%�S�� ��xl�K���.4��JM�ljFz��3�ߓ�5!�:$�JK:1Ǯ�Z=��T��x�;�R-���2I��!._-�%��m�L�fU�2�����T�L�����p�ѡW_Y/�_������*�L�U�iR�ת��
�&m_#�}���wߛQӨ������#��a�}��r����|aͳI�4cϐ�M�4�*J�1i�9�Ub*}W�X�6�:��|�A|��a6��ɡ#�eD��i����_�n��;��ww�~L�UV3�ٔ'$9�ddt����F��7����A�x�G���Ѷ��@�
�� ;���Laf��qk�\FBZ�z��ۿ�lCB��'��8>�O�ɨ�[:�Rmr�},�FT���<�d�}{ޓ���4�~�]mu$��z�M���w�D�y8<2F?����1�P-R$�ü��K/��>�"�P�bt�A��WS��]��B���|���舃i8>1�*V�C�`��ĕh�U�ի�Գ�c��*���M21��;'�j߇���U�{��ȫ��>!��O}�q���X����]H�����rG�4o!� @FGGh�Q?��nf���_�T�����F&��+١��1�ׯ�c=	 ��/�ڤ^�Yƽ{�����e s�덑L(��� Ke��J6���*��W�#)΢K�:F.�����|�����!�V���/��A�6�7�*d��Ң>�;ＣN�jT;��!����9B1�ؘ~T;7H��s��]g��>P$m�-�Q3����y�,��=���:r�0c���*�!�Y��Ε� �Y�&õ�^���η�R�e�?|�L
��)�����@��z���9Y���d�QJM`�hP�O�1��t��1"�+�B��X�̹NN�?����KF��R��c�	��[x}N�n�U�^����lN�BQ�N����h�i���bN}�ʒD*��s�y)�U74I��f!���g3R�Gw���3$�y�T���� =��j���y3��/�e`{KqP쉵��>G��Ynw���kbο�����=����b@X������au#���x��EB f�~f�"��(�*��&�H��f{��E�ٲ֥�Z��G����
�ϐ2ޠJ��J�Q���aUI���mAU�M(F�6��@;!˜PIsl߁�dd|�0,�0ӯ�&Î?e����I�t2Ni�IH�믿��&�� P�#�L���$Fh���7��!��i�)ͦ��l Q���'%d��DyY%7�FϢ�e�J2�j�_ �����\ ۹쵁�qR#�<E�54Jlf�IK���<�ك����)gՉF��YM104���"�}
�7��̪���D�º3���Qm�)��W�\	8�8�*��jħ������52���ϟ���C�9���tL�����,kB�j
�~QF2k��M�N�Ȑ���������0;QVtxC�FXض���/O{R�s�P.׍`�{��ZLh���U��&jQm�dT���H�T
e�G'�ȡ��4|��]4��h4-�*�0ѓ�Q�W.�`4䊫������Ij�-�g������~k���1�0�C�i�,�D�~�m�����q �[n��U�ӂ�� 0��Ĕ:f^�'PW��$��C Q���2��T��!SG}�ˤ��:j�'IX�i)���]~�ꫯH,�d��	+�'۶m#�!6��'��%=��U��y�X�`�N=���,�j�V �l5X��z�*� L侘j,�0��r���w��#N�n��A��FrqI*S8|N�~N���j�n��J��G�&��ő���\n.;�ɧS�P(77;�KgJ�@�V]S�Y�~��ٌ�X(8��K5*`ԟCPX����3���A9��a���kٚ�?�������6��&���LZ2�9&I��U&;���yD����dE^�
W��=�I'p���o�#=�'��Hbv�v""4(h�gb\����O%��J�0����Q*؃ J��N�,�Y�p�"������C���ݻg?5�+@�@�\�*�3k�DQ�j��E"L B��VU�{I���P�F�馛�x����b���y�Z(�X����f��MK�,���&o�x��e�{D�uv�43i�� �60�
�ȮN���~a3h�HHF�"��D��.�׽��v�4����Z�a�.��N.�hY�2�8}5�S����R�ڳ�",ѺΝ�ܴjB��U�)FR���[��������������YhR���֭[c������IL'���������y�-��L��5��]ۮ��;ǎ����ٙ�}}�~�ף���&��U	g@u�8���h�v�RE��r0�*�����IO&��o�B��yN�uGA´lݪΜ6��=r��0��@����{��'�$�|b�w�I![��0�׭g湧��q}�p��M��ݻ�����n����ij�Gm�%ł�[�=0��#˩�� ��y�����e.A	�]ڨ�u��1J���-��C&ӑcG媭WRӢ�&
����y�>�駟�M�6��U�Y��߃����s&O8D-U]e�wb���Γ�^�N���2_jk�� zD��@�0�H��ɞ@�:(&��N��s�Q/��pQ��U`.��rπ�a@�5o|aI��klRB�s�/4J$Z��:�1�=?+��o5G�����O~��{zz��}�)��LY�/��]~���׻'N��v�r��t:�u8�c���B�:�HV�b�L.*fKn咂�盫{ᡀ�鬯������w�+����w���,: �>'�M�Jd�x�l�$��J9�c.�L]�0�gϽ�cF�n��C4�Po�I��m���uN���N�A��{ͪ�Xk� M�1��*	q<}�u*��'�ƍT�#�u�0�@��-���W�����I8$�<��SҬ�5mLSH�N�GvYƂ�6�Qm����#�����[(_�7%%Jl0ˮT3qP}\�#h2���'b�����\�m����!!1��h����O}�SԊ �-����)�9�5�6��m�1��]�T�q\N���V���̥ٸO��C*`�~(.�$s��}��j�:�-mGd_��"���t�	!�����9��ѥN۔���'~8S[�Ⱦ^\P��j%�wX�|�,loU����`ä�ͥHd�}��g�ii�ǑO ַwA3\��;ir�\?�±1Ge�~�&����������M7ʙ3g�0�6�;�DJ ����+V�`�*{@D���)�Hl!����zo7�S��G����&��%d�1�ɷ��6m�@߁&U�Ù�	�w�z��Q���}��ש)����'�R_j��8s@������}��O<-��}�}���gR�d�_|��U=f�A��Ƙm��D��E�O�p���ep޼�Ͼ���2�{lq�ҳ�B�������u �(�����\�l�8�K�T�e�5���-��wp�L<Q;���m��E�j��U�Uݥto������3�/㚝K6`�NZ%-:��j9�Y����QU簐�^|E-n3Hj�:r�U��M��b�r2ώ�ޖ7w�m�p����m��Ч&	����L�v �
��Q�M�
I�Z�38̈��K�s�� �D�+;w��߃Хe_0S���-��ǽ1����U�0%���4u����(ߞf6� Ͽ�,����7�l��� ?0����	���>K)�Yl̝��i�Y��7	~��	��^{�uٶu�`<"hp����Z]�	v�А0ˠ�.XLm��J>������}�����3޷�L����?hv	�pJ]�Y\U�D����ߕtV��q��/LW5�Ճ��j}6N���d\��c�2������b?�J �p˭�J,�2ǆ%�*��j�d�D�!S"�޵[�z��>W*��V@�L�)���p����P�
����} a�=|�w�y���a����ah���"����hU�/�LbCb��[;wH�:� BHlV�",�|9k����s�ބ^���wr
hC]�C2���<y��
��!l��7��E^ 6<4��v��I��eòc�p��Ԫy��s8�7�|�<��3���oP�$3�r���;d��5��D���o��ZȆ����zX~��%˖un��x(�qX&4�7��m�O���/�reX���TLN�:�:��Y@�����J�
(���Ff�a.q���,{м^�n""�ڿ�(/ ���c�
h�v�=� �-�!lrSF��id�R��*爑��������JX~����{Ӭ������:-�g89T� �h�A��#�L
GĊx9H\�S_��f���7#�T+bM�[8�x? h��/Qm�	������C�OX4(�-=~�����kL�K����3�+t�Z{�ܓ6����a��+��Og���@�n(�y��[���w��aƭ1D9",�@�7�c` �	!`���-���	7%2�F����["k"u�kX����'��D��n��ǝ�&sM��`���]	
�y�Ȧ$�`2@Z�-��#�2��T�446S�y���
����H�( s3��8��!�|W4�@jcmP5Pu]��$��x¬̬��߁�m;�D�S��c0��&j�h���$�p1���k?�`Zp0��C�GG�j�ʯеz���_{��I��O�p|�_�#~����!����h���jl<��$k��Uvي�u�e�6Us	�����, �v�c�@��p�H(l��Z��ք����D��A���a��UBMG�ib�v�q�lJ�����U�h$�lTd���t���86�z>̗�5�
� fD�8��2@��4Ӳh��/{�oJ1����&��cna�6|����Q�v>�n�KC0S-%j0��
��7G��Ϧ.^@�&>Q.*C�#���p(�7ɯ����ܓH&��]�Vy�[}�K�>��㪮�΢�5A7_NB�W���HO�9o������	y�ٗ�O����Ɩff"�U���i�T@xh�'Pm._Fy�Q�p�!�&��Bv #T�d�&w0~g�c�|V�Β�B��GM��� 62L��?\�:4 ���;?�S>�`�fs�=�R��>xC��_�.kf;Z�f@�vk+����/�cW��ݦ�,�	��t��q�L!3T� ����ژ��I}~E�~Ů��.u�av�e?EN&�5P�?�n�����}PU���G��#l�l2�a���i���'3���S��=��b_�ς>4�4\V6Ղ?���8l�u���`���u����A`�������e#`�'ؖ���x�x�2=��h9k8"|83^�]�4B�3�Tf� �����?"� ���e���(�ڎ"�b2��Y�)S�7~{�;6,����F�����O���9��;�W�jln>u�왼��m�`�>¿�@�Og�G{���:��٫Ծ�*^d���8G1��ћ`�8�U�*�9"�a���jxGQ""E�Dɐl�A���(3�]�?�C�9bUM Dq�J�u<(����mj�����QF��������#�e�[,��?o�6���*�E�f�E�H��3d�:��m���FD���2`d	3>�� $�UJb���yHb�B�>H��>6��p�!��=���(��NMN��}�)aWH��I�U��Z���{L�����������:#�R��Ў{�髾����q:�lI$g�ZS]W�{C�T�������T���1F�JH$��L(D�%��|=L�ڵ6�4�_	��eM����ٓ��/�Ϣ������)q�����/X&�2ٜ�"������e��e3���_���3��6���أZ��n��2C��'RI�����+��������b���H��xZ��A��#`h����X�v6�52�kpa�m@Ò����z�;��W�R�Щ�0�묷!=�9U������J0�m�6ca�/���[��ZXХ�^F_�W,:�z�(ttg��`��?p�B�����˥����A��[
�;_>�J�\1_T�_t!��0/����τr�bD��W�WfPZ�{�9%6�~'�1�LΩ�q��Ig.�se�i��`�����Q��T��J�N�[פ�,8�(qb>��W����50��qu�A�o@�{�oP�!��_��J��H{%67+�x�jc��N�8�����ئ!��%!������{C���t���;�ݴ� �����i�P���@ą���o��,�z�	z�{�^�z��Z�V$�
)-��ڝ1v&=Fq���HV����.�3�A��b	�fN&���Wq��9�c�����H�@d�7���x�#��o a��!��h���(��m��]��m�Z�*0�R�n	�F���D����{��<GY�)ڢ�����:	Q n�2
��vJ���R`_��D=�cȈ�|��H��3tV,�����6�~�`�`c��KAw��+�p��X�ڲ�-x=G����rŲ9!�h%\�(�Zk)MK,AИ�|;jZ*�i��w�m�;��.��ֺ�SL��"Q�����<?;K"�a�1�(d�k�a��	�1��MϵI���S��[��0z��V.��n���d2��[����b��,�Ӎ*��)<��H�-�cs����ǆ���x4Ƣ��z��Žz|�V�E�J�P���a����Y�N!f� �N�W*��^ r?���~�J��WW�f0]ܶ�uDD���A���'M�
鰝� ֘��1�N��Hy��H��>�Z�������Dw-�#�t'<4�l��^�jB�a!A����� �WAwTX,/�6B�ؓ�g?�~�R�u�ܳ{&� �=�=����N���=��GQXg:�^�r9}{���Ų��`,��� ���ppxBA{���m��᫪��p��8(�!� 8
���;�0^b�SY&9�\Zn5E:a~    IEND�B`�PK
     ��Z�9M/�  /�  /   images/0a03a94b-1490-4d51-a356-eaee23e4f5f0.png�PNG

   IHDR   d   �   ��<   	pHYs  �  ��+  ��IDATx��}�{�ו�{���,KF�Ifv��B�i�t�N�v:m����t
3�R�)e�&i��q��$[��������}G��p���'��{/|ߵ��2���?��������PȾ}a0 �@v�yy9��hh��W^~�W$`wؑ��	���k��1c�� l6+��L&���F#����W���x�����kL��"�;u��J$L�h�Ǥ�_>QO���yN���WB�Db�.��3���a	�u��?Q�������?qmN���M�uq�.���d�<��<>aĵh��a�a��f��j��k�������aq7n\��מ�r��m;n��)u������?!##n���0Gb�	*�����јܧ�g0�D�EJi*-���8y�&�d,	��A��|L)��R�k�7]S���~���E$]R�}4��BI����+���x��bA8BC�%`�Y(섌��1Y�M2'趢Ơ�6o�#5iRc3&d�fJ.++Y���N���`xx��Y��B<�	5������?ٽ?u����P�����_���ͯ��_�����6���{>k�X/�����.WjGi��b4�jL��Q����Ѡ�D!�M&���W��&Tc\���&6o�� kD����/�'��8��F�d��DҜ�Je ���D�*4j�W���=#���G��k5��T���U����$��x�Ƹ���AiN��r�^����C�w6+#��5N��P�
�\���_�kr��W9�a�Y$����P(4�31��U��#%�&�?���eQF�Yƕ3�ei"��hn�>UTrW�F��S�G�q]H2�7��G��=h��A�&�_��͚I/G2�)/���I+���,FW�ѼQ�:\w�v}rd}ݻ��*�4�"��:�4|~�钢��g�����=��LQ�O�'C�`(���+����hok�c!�é^���U0���é����kԅ��Q���1ݭ���LZhRyFM�b�@�ԵД4��Jr�bIf�5�h�LL�0�3�1lJq�Y�O�A~�2�+�����4�C*��1�ͦL�m�;bq]�q1�^�2DQ,CD,*��l2�<)Iy��a����p�fN�GC^	G���J����;h�͹�`�47/�����<���{v�v����i{OW׿�c	k������b(��ADU��j�a4��a=@��Q-	����Y��T��z���p#N*F����(*7�`���{S^$�ǵ����+!��I��x�R�2���4���n&��(@.jNZN�٭ؿ�?����?<�`8<��o����]!
]1dى�f����^��?:]��VW׾t钛�:;�T��e�紺\��h�z��qB�UC\�$}P=<�a!)�$K�%#4�)+TsU�P�(C0Q)��!D))���E|_R�IOS���c�"����QB��6�M���C������<5&���8,L�I�S
��G#2W���k^��X� ���d��(+p��wM���ϱ������B�%$��|����Vc(��j5������ʽ��2�jPa*#�,��&i�!����`��D]%^S��9��&�\}��ܓ�B�����8z�JBGKɰ���We2i�4�y��_ݧA�ؔb�|��^=/D��H85����>'P��M�	������│�ؔR#��r�;(7ih`� &}�p�R=���X$:�?��K/�!j�����<��������X�ਖ਼�#�鉰`!$�����LFw�%���u(�ǌ���Z,���PN�d0^V4(*�1�4�s�I�����/-$�X5���J1�@���3���_T�k�%�P�b0|�)��L�W'���W�sC�^�y����R�ۨ8��k��Lz����N���Y��݉���7��W��U拌���.G(�G����J+�plN;����)�	{��R���Z��x�!9�"����ĪO�hK����H$� Hrq}�r��s�K����@4�Jh������d_=�j���k�3��T.��dV�r=�2�ə'Fc��L(#��TH�TJ��@]���F��T���	��x'`,4dx��iK�Õ�_��?�	~��c�����j��!>2�U�ף��[���0���t�t��gZ�0Z5 1�2SlM8���$G�P
��V����iV�}�u�A�s�d]B��܄�xM��JH�9׼ͨ�x���5�j$�zƬ�M��j��(�e
J''�=�(S�ِdG�BԠ�Aa��bCh|��`0�"�q",T�+'?�B���y_z���/��ņ��+* #-=y�d��
/�����}�V�@?�Ucd��x����5mV�Xq�)�ay��Q4f�� �N���+7u��td��T�����B�I��ߛd�k�8Hz�ɤ�%m|����&�3��5Mq�xB�.�dhK�_%���Е�(o$i� rD�2������3��b&a��`P����#���vσ��_VRRV����\��vwubl��9y�,.@�ӊ��a�e!�
�x�p]�/��j!Ȣ!%�]��4�	o��j��6�$Η�ğU�M�)D]h�����Q��+qGєm���E4�jaҬ���6?����N),�<\�;����@���`L�!���X�dg���ʛ��FG'A΁3r��<khjjFWg;2R��k�x�8���xI^~!���p0���B��M�R��z�(���a�N���1]9�����)�/V
3%$�)G�qݳ�E��T	�4�&��L����=�pT��~��w��¢�5���1!����c"n/5�M����[*���W`G�����<a����Q "�YzzjN4��$
��r���N|�Fb��!
Q�|������ d�Ϝ%aKA[�نܼ>,Y92Q�^�3���+�W��tT$�ArIb�S$)&b�+�h4��B/2��D�Lh�)OL�y"��ŌU�G����eH�k����a������<Y�&�sL�eѪ%{7�x��P<��.�!q8�尘B������6�83{v����Ob���F}�@�MZ�)DU.�}��\��~�g¦be}]���x<�{���&��	�́��2q�Դt��NZO�PPH��h\�])l
�J��L�@u%����hR3k�Ob��F�aM�4?W�R%�x"*�'Y�����5��y��aɐ$�n�g�*��������¨�א�"D��&8�|�NL�3f
�֨D	@��P "��b��&>��O
Qf��mF��!���u{	��s�ph�!�_�����s{(�˕�a�HP��3����N�������'<0r�^NjbbB$�!����I=K�iu�A_��^0�Xj�'�{b��Г}��dΉ�ϾVԒ}2�$c�Z��I8ѐOL��RC3H�T����i��ٹ�Izy�JsF��!4��46�!���3B6�s
�T��gb87�4h>�å���q�jI�w�0(d��O�	�����g�t87fg��"��>!���&!%Q�nJ��^Ґ���_�:�D��u����/�/��F�I�҉TV5Щ�Ӊ]2<����	�TNJ򔘮�����
���Z�|#���� e�4 �N:��	O��[1�e�
�G9Sh�!��X"�VJ3�'fW�;�g$d�ȮJ/��i�p�m�jE� r3�#�2�N���4�}�A��9�@�U�SE<���&��Zu\+(�R�!�,G���Jh�E���8%<f$,<��Р'����UL=+Y�P!M=_}��h�֠������$��+W0:Y�L�P[��J��g�٦�¨/�)�$HMGpF����/V��%9~@��5�a�`��	:��(d��T<�^�J��2�����Q'��|j
���C������Q[^L��b\JJ����E_�0Ȥ�%JbJ�+��	�t�STm�U˺&�i��*�Qgʚ�'�
�dW��X�Z�UbzD}r�!6Ǔ��a뫅j�Pe[��J��w���8�)���J�I_ZԔ�Mlj]�  @y�Q���C�&�Sj����C�{�!�	�i4��f�6F�{�1üSG}�b��47yH}���:��|\�4�\����t����^�*"�V�'O��S?=16�R�EwK�x���k��y�T�Y�
#I�$��E��Z�|&��ص2� ��p�����|e �'���paQ�V�,@y��P��%#A"��Z_W$R:o�J���*�âx�ũ�u�`��L�e��Nz]ħ� "q�\�jKjj����c(/MG^nP����^�fb���28f��j�� �\s�z���������e1�I����(��\�-��pZ�z�H�AS�ɠ5$�ܡ�z�F�����}�Ѡ��ԓ"^�.A�`4	�<!!����~���-��}��c�b��(�8���HL�P
q��gr�&���C6Z�8|�򛄏�Y�<�+j�&�0a��bHwXq��~�]z�.�G�����B�Ӏ���x�,�2�����2����2Ջ��J���h�B��ĵɩ�HT��p.�dX��P�#�Ԡ,\ج��+�1��"5�D$&��-ZyjD-F��$jkJP"CL���E��Vς1D%h���⠁�Х��y���`�f����D�ʒ����hAr�<=%�@@�Ȭ*k��q����H̜�ݘ���[pYRd�T�E����=����Q&�+f�o���|����k6Wj�o�~%�W�!THB	*��E�yU}�ts�.c��T�0 ���,"�p����K-Q
$�Ŧ8lD���@HdL-��v�Ec�VF�|OH ����1�Fie6+Q����O��x,���NZ��D���E����1�?uii����Ay0o�jV>74���-�\�˧1$�%?I���w���J��V�/�=�;�2I���fʦ�Ǝ��ҳ���ee��
)F;��*���?�MKɄ�m�g,GZ�	�_%%Y��Be$v��"�Z8]���O�J+���4]����c��T�΄�>z�Z4��z/���#��fΚ���x�&�L�Ӏ��?ľO�����x�(���8��ۯ���������;1�a����	-�8�w7گ^��pp���ͫ�<c#r���j��ᱨb6�l��D-!�P�M�����Gg�El�҈u�7S��b�����? �'���:3��b��p82��8��{��s���`�
؋���7��͢�S�LȪPh��g%p�)����RR���C�a@iAN��@eE&�e&�,�ϋ���:�����Bzf��c�^f!g)̙��(++S����WZ�����@oO~��_�i�$�
]�>V�f�K�t^�ţo#�/���KX����ꥴ�N����i�D���<ݍG�
�5N
����K/<Gk�J(������OPZZ�gƱ��wq��G�t�Z�烗�v�(*�ǩ�0�����j"�CG� j����7 �s3���"���TN�g�`���Bd�9�ɉ~d1$�A�^�@ސ��o��a2��{��?>��lc}�C��ݷq�C��r��cX� ARǜ�F���˩�a�0rL����� RR�G~)Ce�I%����A[�f�ˣG���ӼEO�+p���҉��EFf��jK+'a�E8w�$<�p�gq@q���66�<���i��V�$nq�1As��Q��/��p��1qA��l�.�O��w��o=&��:s���$ɘ>�0-ﾽ���
�;G��ˬxB\/�|YGW
���r�:Ê��q���g�váǎ�ƹӧp��$-5�B�+��Wq<��G'$�hH&&�Bv�LѰT��f�g#5�A�l0�7��qX� #����Rk6F�p����"!�H��CZ&�Te�n;B�T&�z��4 81�:�5Q�����aT�ɉm� �	���;�>��O0TM(+;W��b�~��q�9��2a������nу�9C���I+𥳐��J�;q���t�r"�� ��%��������艃�?y�
��T&u�J���]-��2�%���ԥf�� �-\������ �z^~6���pBẲ���C�֎��4D�A�͆EK���7��6�^�7^=	�W	�spfcå��ߌX�f^{��C]³���t�F&���������Z﹣��D%DR[�(�cEI�C	�xeM�71���Q؝F�1<�B~I�tUST��B.�"Q���DUM��J·r�Z%�A_���L���7g#C�����n1��=���>df��v�̝�A��B<��o��}'��֋�|'s�,]�B����n���������ػu�fl���z��rÍ����d��Ø�d=�͢{QZ^�96��a�B�r�Z�Ϛ-$Q����3o�ŋ�-[�s�/e�"�p��V��ʵw���*T��%kQR� esB"8RS�bÝ8}����07���F}O�4���ʷ�رq4_R�HZ
=�b/3Y��#���8��[VL�"��qNY�.�ĸ~�"Wo!�֥)���*��`�<��pPeeσ�z��H�P�W���
����Hۑ�=N�t��0�򋑙�GHL.C4����:ڻi��()*8��<r���~CÃ�x\YQɤ�"�[眶2����0<4Ȑ`F���J��C�5+7o���HMe�L4��Dn%%�X�z��%Զ��hz��x���3�b�mX�$��zl�B��S�Q̙=Ki ���V+)�qw/�?A�eź�%�,@~U.
�Q�T���ZZ�2t[PS� %������� ���.�"���s����e78\�K��h
q�C�v{���~����������i��>�����v��dtU������5�/�N�z��E���.&� 6mބ���b��,}���Ge���hinAnvr�
�k������!+#k�Q ��J�@"��'���X��%+WcZ�,���C~|����@_'�I�+kp�=_�02U�F�'���h����q,�?�տg^r�z�x_~�p�de�p�d)��Zo��t�� ��{O!09
�g�^�����)"���}��Cx�g08:��!UZ:�/<��a��P>.�<��w(8�s�m�i���/��̃�V2a�|�<�TSH�9�Hb�0��]o�����ݛW�Ǣ�7%���/0d$�7�;��ҊHl����w��s���$�'���e��+r���R��>���;غy���ؘD��ދ_���P��7ɐ��΋(*��a5�#�����w��"�>!��7��%����^��S�PU��<��s��
��==Id�<�[���3����C�ً���k�����p� �өG�Fo�;�����u�%�r�W�BQz��$�����=�n���玟��ߍL��,�[�8��� ���"�J(j)W��
�Oxm������tUg��V
���0��g�G/�8�����,f�-��H3�+����������p25L�s�Y�0�2p������pv�s'��y;��]֛ǔ���S�h!!<xP+I(��J0��f.��{�[�J����cشi.���]��ɰ���9�I�?w����\b|���.F��A"/ȋ�/�ޡa��0
��k�!7݆�g��),9�;9A�G�������l}�s���>"�A�T��	I��`�u^�y�A�"Z-��'�P�0¦Z�\Zw�2N�>#�{f��EmUnҗp�6R��Hpҝ�����ƽn=��k	
k�:)��	M� �~
�DD��}��Z�q`��a|�[�D�+֭�r����~�mQι�琙�M�:���
�����ҥ�P�!�>�� +��U[*(e��!�dEz��a�L*����[o%�8F�y�����p�R�X~덛���o`7�i�*�����8��j ���|�1�QTex{:f�[B�IXl�`�����u�-,���0�B�j��u��Bo=�GP�N!���Է�gd�B��t�\22ҵ�P$bP+�*ϩM7����an�\Þ�Chmo��*�_�;�h��^Y�L4���=yN������D1�H +���޽iA����;��r"URI��0��]o�2"Zg0(���+�wێۉ����JR&,��+Wn��BL���[160��wZߒ�[�~���.\8>���p �T�ZBԹ�����q#f�ŝ[v�j�	F�(��ނچ.��\	T/�ʍ���K�D@K7��
�8lR?�6s<�����cĀ�s�b�L�#�D�������i��͚=��.�a�Q�3,4&��c���k�k(��C(��FU��C&Iv|����� t���0Yf:��^���2)�Q1}=��v�aO)`�1�;8��}�����E%��!�e��ta��B�ԠRS�d��V��"=-����i��ٙ�C>��䲗a�}�Ы��3�(/�Fww�UUU5���{p��7�J�2�IN#h�m����X�~V���08��@ϚDk�yļq̨�K/��.��y�H����Ο�8�v.�X�Y��Ĩ�TԠ�� 𣖂]�x�-h��v���&�ڞ�0h6���S�O*TedeI�BJ�+a��E]D!fU�1��z��s�Ϸ�X2����Bv�WL��A�[������5�!F
1�0uC=g��r%X�d҉R��N��-��b�Z����!����CQd��2WeA�`���`}�_R�Z��>�1.\:@���e��R
&+��������%�Ԏv/��||�{�o��!B��_���m��̨�����,M4��%��Ï�m��t��}�0x~��r,)b<����q�H�P��x�{���<�7$F�ҟ~�p`������<�$\ٕtm�_uE��m)[_VKjy�����$��Zߘ)����s�~��Kre�/�E(0��^y�d��`��)@K/����A��r�m"�A&�l���W04�֛71�'�p�X���A3y��ȐV-b�|A*���A~��	���`�ʵ1������
[q��i<���1�~���}4��GTbA>���˧��s�ǧ�2b� >x�5\a�Ia޳�������l3���e)�α^9GR���j\h����<����+��K$����3�ɧ���z��:v��i����[����iT3�b���ػ��N�	h�]��&�S����e�ج�K��ե�������á�N~��k��jT/-��!��U 0�v����LCԚ���s0x܌{|�#B�������WK���`/*�U�,f �詣�==�(�˓Ҋ�q����R��?z��Ê��I����	�%06�;�&�s^ڮ��ڮ� dMK1�G�����{)����f�����"D���K-4��)���+Dq1Zk �#D���ΞV������������n�ݙ�Zzƈ{�H\u�`xl\[oW�i��n�3�O�yA�MV��bx��d��4���-�	Y�p̣ҍc�H~Q�U�!j�m,��y=�P���R[����P}(/4��H`2aA�d�x����48H�NԔ��d[��v�Ot�wލ��3�L�r��eBh���`h9�q��t���sX�d��U�**����ḇV�y��Б�	�ՅȺ�4�)�1���QA���Җ�ge)W�� ����Q��T�w݆[��܆h��GqW
�m� ۧ����;w@4^�v�"?X�h����F�-�7��f2oQ(����a�
��ɏ��R5��"K����;�>��l6�U5���6F�h�C��D������Åŵ0��$��pv]w/6�����k��JG��Ay�"vt��C�S��Ӧ�[71�nN���7I��{�Y�"���t�2�H�m����"|��M[oi�����㮇gXL��b��hk�&L$�	b΂UX�d5�o�%UX�~;N;(Ž��q-�A�I���Y�5[&p��	i�X�l5s�v��F��J�7���;u����m1���&]*q�����Yz�A+��Ō�	��RAs�,B����t3y��PQ3��@��x�l\�g�UՄ��O����JVۮ�ҍ��7Q��B�R0]�a^1|���W��K�v1�����bu�f�p7҈�
Kʩ�(��=����sg��ee�
+�I�g��Nl�%�O�AvK�I�g�0��-#CY9֬�Ƽ��kj��:d�� Š*�X�=7���{�
4. ���SdER��7c	=A�����ើ>Y�/-.��oŪ���]���Ö�&i�5����o�F�ZPm<�N��0w>�n�Q�J�^�Z=ۚ�]PU>khV���U6����+�q��V�9MVP��'T�j�6I?�	j�mS�%�y�j[BX-R�BT�)�(�~wthh ��	>̋Eӗ���AC��`7�[/����I�@E�J�����L��Xڏ�ǚ��q;�0�����	
̑f������@*��Q\�����S����2��B!��QY�Tu�3����w�w�a�▛oƢE�$�(̟��8u�4nO����~�kp���JK�'񽧾C�֤�R�f���r���t�N����6.5�"y��������9��RP}�=��/�����a,�����S_�+�H������~�ޮ&��a{�O���dO��QtĬm�SZ���I�Q�O�W�^�D'1�������{q����#Nb��WB�=���_Bb���4t�:Cp�Ӷ"�X����w��D�c���SLƝ����Aq���fB�}���q��x����m�&�,���Gp���	U��[o1��j!L63v�~�˟	jR��?��e|��O1����/���O�8l;��Kg��_^�ß�M3�]ｇg��3����K/�G#���7^��g`U%�gϜ����;B�o�f��8��6r���8����+����~��d}���}T�9���������g��'���R'4���6�C�򃴩��d�ќ��z�׊���}0�#�$n�fGUYƇ{Q�U���f0�f:���ɏ���,Z		�@�q�h*��P]��es���መ�{�����Fme���"#8z�lݺ��h��f%<���T1��0�:�1��g Bv��{�`�[��e�ؽ�#�iX�$h1H#������sZ��H��T����*u��$ÏA�[.�3�:v^ma�+/6"4�v"�v�	����H�i��-�͆�l�����}i��KԶ?��B7���' jRJ�KK���/mR�5�G(�PK �\M!�ɠ4��Ox�1"���N�y�h� ��CE�����ǧ1^-rR�#i�1d��Ts��̣P����C^�bʊ��lwv�^���B��*�6������aue��Ȧ�Mr�&���`딆�)RTT��'��{�H��`��颸��砷{?�o��'+��%˗�V]��[�m���0:x���߆���P@V�z����q��aY�6� +W��Tb�5�Ås'�W[���%Kf5H��BM�-a�<J�@k7���Ƶ��k���L	�.��S��-i4�
�Xj��PW�`<lB�@3 /����v/R�҈�i5��p�Ӄ�?�iy�,^��[������<֋Qϐl�:������aJ�+��[zZN�"������Ӫ��������
�����J��+��o�e�z�]wݏ��Q� �r̆M����{b\h���c~�=��dш9��+	@��*j+z��у�)*ذ~Q�MF N�BI��/o�z[jK7�t6nܨ5q���K����I� TW��ƍ��x�,���	�_�����|$���5k�~�A�r؉D#>+�m��fP��X����l$�&=$��bJ�ʲ�M�����#~l�if�\I���L��[�?}Bq?�A�[]��&�!�IX����Y���u((ʧ�&�4�>2�G����.�_PO�]J�;��SK�|�=4�ˈ���f�X�22��OO=��)_ϛ;]��}��2��lX�AB�Z�Tm��#�'���X�f/�(h'5-a��>�Ie�u5Ӱ��;p�M�I�t
ў��������fϜ��o��6n�(�b`��j�(=j�e���曰v�����?��0P=�z���J6����Bi�3�MQ���� l-7]nz���#�d�Ͽ�k�-���%ziĴ鄹�X�=���+8r�(�tEŅX�d#j�)��4?4�9��+ǥ�0����m3�s��)Or�־���-��nD�=��l*3��=N{/��>"��BU��W`���R-����!>��}��=k}�P[)���<��_���CPp����>�?O���q�?�яp��aI�s���S��gY95Y���7��$��E٨���|��o�K8��gIrI�Ik/(��C��Ŕ���8,�]���֌�9)���v�͢����?]!ݴ����^ߤ�;8Џ��lL��������sH���CG�Qx�<�ch�I7��͏10<�lZ�ko>O��o$42�O��4��"/ہ7~�>�7^�s��L���ￌ=��q>��v�f�t\!��2���;�^~g.M��3�����֭]�=��rR,Z5��9x��L|��<߿� �:�u"��8v�/��������7^Á���n�rt��Y���g���.�7^G�AIA62R�h8�ګ�������M!3�Hou 0ڃ�����xP�N ���PښN���6<u��}?Jr3�(�豣�Htv�K��]_����^d��"L��꫻�~�������A�a�"^����X�|)�K�+�f��DmRj?~�	�68������%<��~���/z�F0���_�u��0-8.���A?=�lܴW�/K�����N�s8�F�R��1������L!T�ɖi����ޡu�3�vttɩG�V��JF���$^kGkK������I�S������$���n�˭DGv��n-�����5A'��ndk�u�HǾ��(���THYI	���/����q�w��Ҡ��ˢ�>�1\��c��/C���":�k�������p8.Jq0�}~8��#d���X��+�� ]�@�y"�M�8��"��՝1c"�@g�q3CC�JuIar���x�7�@�W��f͜�T���/[�G�alxT6�i0�-� _��h�{�'�arR��3Ż�Nݍ�����Cz��2`b_��=a�gf�b�\=� 	�1�d*�cv�,B�4���v��A���Ȩ���/��̍�Q"���]ʚB**�.����W�W�6SU]��v܁SG�a�	��w݆b�
U���Y�ūV������vd���l���(��%K�x�r�������/�|��e�v��3W���	��=�S_�y�Q;����~�V�8�����e�����¤w3gN�}�݋w�}O��,Z��;v��Z�_���߆7_C,qݺ����[��D5U,k\��?�0�!�Q���nټQ�#J+_��_|�o��5=͎��7c��m������Ř�{p��Q�ek�W�VF�k�l�m�P�à�Q���$���C�Ό�����
p��ں���|�{R$f��E��ˇ{�MT���B���}�����{����ZuY1�.�+*0K_z�oq��U�����BYi%y��p4�3���S�i� �H�,g�Ȕ%UN	Nr��>�$��wpr&L�3��8��wbӆMQv�5)�2��'�RTT�m$��׬�%۔�t��������0�N*�v�"C	T:;;��V]��w܎[n�Yv�:�V���sD��ѕոᆛ�/o��	�3=ˏ�d�jcgyE����7"y"��t��'p�S�#��j/c�Kg�bnuB�{�+�XWW���Z"�|x�0H~�ή���ۉ���i��X<��!,��~~�	Z����a��0�a(.	.��Ǐ��W_��&�|�"�M���C�;H�72z#݇�`¶z,j܌�yy-C�裏����&�uk�Ѫo��槒������%��mh`�֝!�ٱD?��ϱk�;����[�$�LKːNG�g?���1������o�����w��1&���}�9����x�3_#+274և?��'hm:+b��+�#_��u�?m_�v�Ţѩ�ͤ�B<��M&
��Ǉo���te���Y��(kɢ9���[a*3�k���{�[��⢑$����O�-]���_��KC.7�a�������_d�`��	?���&�j�����6�@Ϛ��v�D?ښ#���������	ܺu;����O�o����3':v��<�7���w��)�=�A�;|���'�|B�����c���kWV)��ٻ��y�OJG�{~HR�����f滎��<#�w*�����8{�$j�R`�ĺ�^®���;��lx���wp��1�ӓ�!���x��	���u�D�
B�Ԛ�Q�
`h�%q�������o������>211�A����DZ�x�����}�t}?�Ә��mȪΆ�
��axtyY�0��W�oF^��8{�$�c���e���N�S�0%y��u3fo�&9�L���X�wM0h����p�֝D2Q�ݳOZ��S��G��ўh0[p��(
�Oe�Ҿ�jm��<T�m/��`gB�d��D�F����_(��TW{GG3&<����{sL�Jmқ~ޮ��2��� F'b�LN"�JIs����MC��f�V\���������K��uI=����#�L���.�
g>Z�7J��7"ӑ	'9�ي��u����hЄ�	?r2�O��k3aU�G�n�]9�jO�ڽ��GX�d��0Mg>ʐ�!X�v�l����=@��@Ii�A(UrXA��m!�#�w���X�aY�tz�1zi��&!�y�l#S@k��]�ҫ�>�Iw3*����P�۷mFa��g��	d2'2IǬ�u��,����#SmV�$�\X?���%;�V���I2}�!LL�eU�q�B�uR��A�Gk�[�K)'����dH�wث���RLV�ġ�i�+"�^�r���P����`�)H����z&�3)܀E�(�n�P�%��֮Y��y�ar�Y{s��߄�X��kf/\�6�pR	�ť�."�Vd�����P���Pe�7��NՎ�p�8�������,�Ƨ�4z��1�Pii��V�NK*����#��q�4\�u�.jD,LC ��>���i����b}(ș�����L�+o�5�S��Ѹ"X�i6n�Cr���bV�<���`�����u�fl�v+�A�-K?q<�:tSP�D(��P��99����a��/��"jk�a۶�ƴ��L���1�l(����L��i���+a��)|0ڭ��`r
��j�斡�r!����-zņ�1��JÍ#���5vzNH�b�����D�Wŉb��G�����1���|aA��tza�f΂�YJo�!�$��"����Z�2��1S�XSyDE]�ƓH�ԡbŨ)Y���E�aY�S���#zO-n���_w��#�C�I;�PwV�ϫ*�p�NB�nP[>9VC�Az�ԑ����h��zr�Z�3�	�oo�.��b���	��3\AHظ\Y�_�B>y�/�a��|�BT̘���:*(��H���a��rQVۈڙ��RT�iFg�i� �֢J�W�@Y�\*�(]M-8��;p15̩Gu�Ԧ/c>pp�!���$�W��e/GfZ5Ҝ9t� z�1avQp��#��x�7�dR{]"�����pv�"^9(+�B�d�����F�0���5n�����Jx[���pD#�xi�؆�������_�.rs
eW�ۃ�쟱w�i^�5���&QYV��Qm�H�;��s\�S���r���&��vb[R!+W�*ߤ�����/΅���ݷw���ԕ[��b�dh����v^\9���6�5<��2İ`�vy��ԉ���h�@#Yo;�1�y�6Q�>�C�DZ@�3's����d�0m�N�+�\E����0F�Ֆ�[�����j�h�(��ڰ�`X�!H�]Y��&#�ng,?;�#�3V���ׂڒO�!Lx�6�C��BBjݞ�T��ey��.�5��=��4��q��	y�x����L�=�v�䉣4���q��I����'�xB;38���e2ŧk��!ّf�eeU�0���M����|�2Nu�>�#���c��s)� ��	����e��~e2��r�B�j=���¨N$%�7��BU�*�U���38~�8C[�ɐD�ɯ��M��	։��3�x1}^9�1
m2���~��E���N6sp����O�����W���GhS9�����fh�F��B=�1�tF"�؄Ω:A�l�	Ǚ#�**˩v��I?�9f��kƉ�,00�v����$���twu�a2A5>J[ջZ�\�c����U�I� [���Mq9dS��DB;��s���.`��t�M���I�U���B|�� 7�E(b�z��@j��ɷ͗.�� Yr�|�䈈����
��}Q"���4u�>�Ak��z�}(�d�&�R+��HL�R��أQ�����]�jװZ�Wv��*�Dz������EE�F½x*t'�
s��q"F���M�0>�l~_�1��W,��*�����8�	�;2��RAD��gΕ,UZQ�r�ޏ�OZ�ʺ*�/_�TJ��$W��HT�)'��R61h(�MIz-~�hBQH"&����`��	JUR3�sp�����?��C�H���¥+Q\\�c�����t1�.vP8��Q&�e�N�Ɖ�kk��=Љ+�Ȟ�
ͤa��u�;�P����12҉����n������n�?ŋ�����{�UjYNG	
�������h<#s��^!�]����r8��)��vWJ:Cvv=J˖p�Y�4���+W��e���hrJ�VH���Ӑ�5�cW��3��y�2l"�JČr���Kpӭwb����,�u��}��j{=�M?�ʨ������B�Z���Ȩb)�G��@��ǐ������o(S��F�E,qn�B�~����]i�U3KZ'#����v�f�j���d碴�^unK�*��\q#J��?$R)�

I�)G���ض�^Ri����V^c��������W��e��X��^���|ZY��y�P��9u��X�f��9�Z��Ɏ�����M~�*�x��V�͖����ɡ�3�\)fB� ��x;|���;�0;���@t���*��%ex�����e�KU ��mm�҄^Y^!�!":S	�Q��R���L]�ቲ���i����)�T&9����#|7��Ee�L䪐A��v���a;uI�r��[0g�B���)��x���9y���y���>KVS�!M���� ��*V�ЭEy�t�H?.^8��^zsf�0g��d-FV�*9�*�c�}�a�:@��ir3� �H���c"t��;@�_����p��
F�>��d�4g�盦�,�fιT�s�b C}���0�Qq�CE�}p��D�@���G���L�FT�}�3O0��]�r �/~��߿���b�%x�_FfV� ��U��j�����J=F�e]�!���!�n�}=�]8x�0�z�qy�̝� ���'�g���{���q�r?�.���~�=0��:��ݿ�.��σ��������7 k$���Ʒ�E��M4������{���?���@G;���3K}AZ|����P�����K����Ig�x@[g�U�QQ�c�Mh��KK����s��cA��̃E��k�٦c$q�-r"����;�&��<tt������'�r*��� z{�Ǌe��$	|�{Nۃ�<��-��_����?�5Ż����q`�.�JSF�;u �{Ƃ�}�;���"�������a���b�������Ʊ`�|&5s���F0�����;�p��a,Z���(�Z0cz)�m��J�p��Ҋ�+V�ҕ38��<LX�$�=y�$:;���Z�x}��L1!J6�6)�8q;�����2|s ���h��[Č���[J:��˻��db5�K�r����n|�{�Ѿx�/�H"M��jǿ��1�g�1<���'����?��Pag������vZ|o����Q9!H�[&	T�ư|�Ҥ�?܇��LzbXN�N!��G8���f#J=�4{�Q�h��`	�G{�T=L�i���z����)�����%��u�,C��3	�/��Q`Jkj_`\�
�F3�3%V��{����(x�C�r,f�`���|�m�+yGNN�4���S�����q����,��Ǒ�OE�F<���.~�c ��y((��P���
/)���x�Ř�ήV�_�r{q^1��Js`ɢ�x�M��F$�{&�a�B*+��+�U�����7�M�	��kܰ������\9y��8	���	a���OmĘ�q��I�F��G�-����P!�h֎2��m�������*k
�3�Z	��QE�YW#����kK���+� V�[n���W��c�a��}�3��D0�NW(��O=�_��_12:�����gPDh#qk�5�q�a�����i~~1n��a�	��.XK,?��_E4m �ӧ���1�%�fˆ�.��C�9�=}>z�!
���7?�i���_�K�\������bH80k�<|�s����ŬF��{>Cnb�������G,G�,\�k6l�s�q��_M#�!���,[��7�H2��`q��t��ǲj��a>n��N
߬\;�\-^i�q��h���7�����KFuM-����c��X��Ș���̨�5���Yr3r)��sg"&���9�y˭��>���ue�D5�EI�e���w��҅�

QTV�I��&,��;�n	�χ�e(J#7a0Y"p�j?��/a���L�F���{G�z����ؾ��߸I��r�8h��u�sn^���v�NlٸE��)鲲���*��Up����OO�&����L���"�ʕ�b��۱�q��<e��#̨��ܤBP���[oǺ[D���1��L�v0�~ҵVl��	�I�kL$�9ԖpZ�rR(��+Վ{��	������!o�
�Q?�%�D($sv��Ԇ��4z�Q_�*��´�*����|SK{��w�EC�ܙ3���>c.=J�\>w{�y���5���ؾ����=m��_? �p���Ý�oĬ�yLSv���_���_���(j˫����#���D!��0~��ë��F�J��������+��5O������7�x�V$����|�)9�C"e}��?�}�V^__ۀ���<R�IhU+�����r�䔊������S"5�	�O�4�O����?���N\�Er�nB?TT������i��o�t���FT���y�n��)A`b8�Ǟ�G��?�&�9���Ձ��v&~7��Ʒ��x9Y�?�>._�����h�0����Jl�����{pD'��I_��"��>��	�R/~{�<N��HXq�gϪs������x��	gjyiNZ�U<��_�{���le8}�8>x��J!�=u���K/�����A�H���|��뜧j�����<�����_zB6�~��n9�i�H#�:�b�ǯa�ݟ�Hq��] �J���A\�z��}�m�ܭ���ܘvX@,�(UzӚ�d�V�����C\W�U�jQJ�z��	T�ʭ�dW�o{�eWy��~7��o�(U.e�$$!!��$@�Ɉ`�����M�ƹ���~=3~=���=��׶1`r���"HH(�R���Vݜ���>�d��֬5�Z�o�9P��:�������N�>{�d����.@�� }<ee4VA���*Y�	�C	�"I�`jsz.vS�Zxb��4H.;�c<<2���r\��AIEa	/��BG
�G"2�G��Nu�\'����<�y���������01zmS��'�a��}=��c*����͗/+)�^Kp�:xr|��x14Ї��Je�F���t�=�51"�S�h����C�w��[z9b��nإ3�5f&���5�qp]��Fl��M�+��M�10�Nf��SW���r�͇h*���X��� u�7?O�¾�k)�I�:�F�mT���Y+�T4a�J����;���	Re�
�<	z!��$�n��(V��q�onzS]5bN�"�\8`낳̅���{R�N��i����Sz�c(-��D<���F8h�"\��Y��x����oa�r�O�*�)!��9����$z���A.n����2��͝�o��ߏ�"U=-�"Bv����>ltԆ$2�qf��}TEIŰN>Hk�����f��Tz�iY�����V�:P��f���L�����J
�;o�KO?�b��Y��ij����O�_z�63���e+��j�������;�|��Ӟ�ukn�'ϣ�3g��z�m/�߰����$��W�t�Ln�(v��D��Hi*�����4C�կ|�<�b� V���|<V����o~[_yNOͲk�b�[���9�M��p��_�K/����K��7߬V	 .X�<�=��:mP:���Wb9Q�Q�������<n��+(��~غ�o�"=I�I��clFK���I�?˃�宿�0m�#��J+��/)��-'�@U�W�� !� �
JPI��Υ}��kf͝C��Cu@~^1=�Z�t�DF�A��(M�~���E�X���*q�7SZ!������\�{e&��1.?�{%nY2f-��(�_aN�hc�X�v=�-^����[��lWO/���M-^��K��s��V���~�A�u�n͍Xz��Q�r Q�=��:ej����\{�j���e�3����m+!{I7��_|�&�
<������I5�Byeev��'&ep�Lv�j�����,�g�dC��H�h�,^�siij@�:�HI�"�	9�6�u䗵��{�Ĵ����53�KT���J�<ƅ����6���
޲r8�6�>y{v������b����Ь��0_���x��xbƱh�5�~ӭ�1��P�Z��pd�>���s��/X�[7�A�٪�������/�e���ɏ��S��k�3O�G�B�pj���w�jZa��uԯ�+���Ƙ�,�G?��
Q,�V����-Ξ����鞋�7~v�WmJ4>�g�|�~�.n�ͼ��_��;���`�,�66�re����y�~�O#���)'Ǔ8p�C:�!N�<�Eڵ;v�M[��w���W��u��p��\<}���_�����~;w����b�߉�����7�
fW������[��PbϞ9��g/�'�����O=�>���/Ө&q���5��?���G��>:����|_mӷ��߿ϼ����e�pN�9��%���?�e���x덭pȳ�9�x�8�����O��.��ݻ�ګ��96Ӧ8	w�_��_��?�	�%�}{?�����Z_B;��ON6l��ڋ=�v�����#��?�#~^5n�r�g���YR�+-	��>CY�?�!n�vL�����w�A�S�'�#Wp�\�㈍�a��jU L�x���-���O��~�cC�	��\��7������h�`&iQ�fA]�(��ũ�w�6�8:C��D~a�@t�8����>�OIІG�P�b��w����I�C�BeY��		��˗�*ǩΤ2�}��R�������K�(�r�Ϟ7f,r1�*�"t^���(����*<�"�i̻��T�Z����2�hZV�x�c�=�hl3W�ax�:\̤�;�%`��FVdr�П6D��\�hn��.H�$�K(������뵹�0g��{'�I	YE
!����4l!��^8w���t\�ЗG��
=N�����X2����i�qS�|q����X�=yJ��Mp�z����6JAMD/.OU���_юȖtFI�p��ِz�HH��\Ģ>̦���=�~�m�Lx�K�z|J�,^����`�X0|�7 H�-�9J�4C��$J�Np���7�s[&��o��dk��g�����LZ��+���'����zZ�;$��_dg�_G������*L�d�������
W!�wvj��8��G_�N��s֢�j���pݥ�m�/u#�`aٚ-p7�O�R\]�5�n����Cő�_�e��F'DUS��܄��{��WI5�m��/#/��/���þ��SR��b>��w�ܦ�f*�����i��F�y��:N#E4���{��W_ۆ|��r�_�!
��46Oŝw܁�w�G����˰�5p(HhZk+��~|r��ڐf:�+V������Μ=7l�����D���[��o�m�e�1EHĤ�#�ٱN��h�"���u�Sq�}_�1��3����X`���T���>�Qv���f��w��v�P5m����`)��S^��9{��ݔ@ۢ�(�m�JDqI	��B�M�%��%r�����ҭ���ڕ�[X�CR(��{/n�a-�Omm��?8��G����*��,\b�#��ϟ��4A�]��o\�%�,�*yi��������`%]Z��Lz	���_A���+���28�E:#$��6F5.�r�����y��#%�J�o2��֘�+=�,�2L��A0vC$`��J!�$����y��ǐ��3�+@���)���+�'1_7.{��p�Uc�;��3a)����N���O�@Ay�����u��;w�\�����i1�`��[PP=Mg��R	t�8>��4�uS�7��z�&�����s/h�`�M���}M!�ب`0�Ǟ|�ą�g�T_��|��<I���8�W
���踀�Nb���x��ā������?���WX|U�\��}�!j2�xtJ��8���u�A+����<ETS�j�|=&��L��eg�f����xiA��t�����6Y���3�R�����ر�e�޷��P�4�+2n+�v�zoE��Xt,ԅ^�U7�������}�W����@��%��tw���kyO4�?��(/��K��q��{ 7��CU��n����RgM�~����m��^�:Ձ��|��Ҍ����,&����UB(S�� ^y�.Jn�qa�����_�o��ńC�����=[K'�;�-6�X�A,�>>سG�2���	�em��ͷ�fgΜ�;;�0dh�<8s2'���Mw�ʓmͩ'�lۮL;4
�h���Y��,]s6�>Y-w億�@V�%��ݙ����45��cJ��T8��F���!�{u�)i]�f}��s-�FG�_�F��4LkC��M5wFKN\N�o<��X��i�9'Ν���9�L/l¹�'�x����(��ȥ3T�T}4�&��Ǐ~�Uko�����86y3���@�u�B�)��jcccX�f���*(��%��~:�>���R�
[��m޼Y>Bǯ�[�<�K�~��_��!�������b��==�}�Nkv)Y���&�t2��B��-q<S�)�*K�)����4"�8>�Ҧ���/?w1�H����4{�L�]AEA�����#��Vs��_�6�i)�KH��B��bz�|�G�"zi1�����sst8�,H._<��q�B]]=|QJ%�j���'�s��Q�����S�"h�V���3��¥�.����'Գ|	�N�R�]���/!�n��sڝ��c��y8��Ǩ���W%Fh+��)_�y��b'�f���w�ԊL� a�۵j������V1�����R�%�N!LNKp�^��>c��ܩs3hJ�������Q���V�kل�nݍ���3���.cx"����U�h	��U
���9�;3���9�W6]	���~I�z�$F�"�u�!e%St�{qY���-:d���{~��ip��Q8y��!T�M��E���S�k��.�>O2aCA�o�A;k/����{�.M������D_B  ��/�|3B���
l��%!����jnUB}��ru]�}���*��n%������l�̙&���o!�H᪫�ƍ_���T`��,=�6%�����O�MJ�ղ��V�iM��~jCr�r��ZZ��v"!��˛����(u��&cg�i���F~�f��@xJ�*�"�t�|Z%��iF�̻Q۴	y\�j�=~iA�c���P�8M�DgO�B�R*��˗�E[C;��G"�yN��͠���^w�V 
���@I��t�]�����I�5��֨��W�ꅋ0s��D��6'B��07"յ��x���y�{�GH����H(���؋e�V�}���/.,����� �vD�>��0�4��؄�:[]����a�źGÑAV�3Er��z*2�?���ö΋0w�L��4�]1M�A�'�KX{iQ!+��V"�kʂ��Pp;aq�����ϛ�p!G.��c�5q4:>H����T�L����S�qfާ/�����+oFIE�MHFC8zx�N�	s�[����5D}���v\��$j��Q����޲	-MMJ�J,�	|��>%�,+��}�5��Rt�;{�"�^����� J�h�_��"o}�8rh�z��|ǽ��ʴ:1M`�KO���������0{3��"��2�8��*�1��R�l�P�ELi
@"��ѹ�!��^y�``(��3�چ��7��GdՍ7�/���)6�&QSJ�H��dw�[vV+Ppx`���&t��ਲ਼�v�����Obb�C�����ǎ"��G`�)���e����I&4��q��>|�/�G)��G=��S�*�f�*���D ����m�����GU��z{��م U���ϔ������h�{�u(4|=���3O��Li�|r�>�ZZ[襇��}�����x=��!�}�-��|��r�'x������D�h��w���g�P��IgN� :��ƻ��gt��T�@F}��0����Qfreg'~fC�bq3q�Ip��1"� o~�3gcjyҡN�J"	���E��4�G�Vʑ����"bOL�t���W��rCcㄉ6��"��釟�ic��;5���F��jG|��Te���n>O�ȍX�`Lؿ?n�r�0:6��b�\���Ta!�Q�?��M�1�V�x���̹s��Sq��\�=��F��J���Ӣs+=�K�Բ�V���6�l���k���K�;�w1�3o��ph�W9���=���>��6�FS�� O�ҟGY��s�2.:.6��ʌ��a83v�k�P���f��	OB�0�c9h,���?㰖!+���c4&-D's�\X�@x&�Μ|D�#4da�|8U�3�6"���.g>�c�J� �ʡJ�:���,�+u��L�
���44����p�2����|�X�C�%���܌��z惆c�M_r�"z�.�U�j�U�K?�S�����ra����0Qe]��~��'t|^����ؠ���͝�҄Ӈ�K���T�i�S%ڋ%L:k^z��%A*���&�F=Z2�2g$Q��"�F���[\d�Aaݗ���1k�2T׷!m�A��;p�c ��>h5m��s����� 5���#ڜcra͗VÔ;U9�XNd��'i��T�׬��h�M�3���Zڌ;���#@#^1�w�~�x�|�ܰa3���*7C����w��ˌ2G1���Cx���1A��GX�F���:��ȫ���^����3g>nڰ�P6��?��G�,_B#�,]BT��B�@���&\�~3�F̝5��V��{`�i�����������Y-X�j�2	k:;�QYM2FZW���-��3S�?���D�����_��w���A/��3P�������~Ӄ�q���+-^B>L#�WE3������-��P��(���X�� w>0M��x����)֒�pdVW�Z���?^�1z�U^�Q�S������kW���9�j	:��o���ćD\S��Ԃ��kpO��|w�'���R;M�3��i�%!u�d:�7���e%hji�/���A�a��q�����(,.��9K��ڮ�/���2�$��>V#U�+V݀�W]Mw!N��Qo<�J�s��Sڠ�6��u^"�A���i�����͕�A�����`ks[�B� ����5|=�P�oG��ܠUp���8v�#|���s��f�&,X0�ŕJ�}�8���5�-��	{�k*���'����Hxen/֮��к��:��	;v/�}���9�|��5((�Uj׭�l��2�MU��o=�e�C��f{�	�����f��������)Su*� �yZ�@`�~H)}��~WF�U+���A?��Ǳo�.����l��n��TC9�R���p��A���������5�N���	#b�bM�j�CL��
ӓi�s:r�a�)svx�B'ATUU]ڽk�o��չŅy���{�pl�+��%�O����-���|����uuŔJ7���*�쨨n�f��ﾊ��3��������{��9y���8v��"AA����������� ��< ��'�c�6\u;q��x�;����W_��x����x3�K�����x�����+�T"�A:�O�o=B���3��no���h�bg'^|�9�����?|���"ʽ���� F0����qa���Ϝ=���wq���󔜿�ڛ�z�!��&�2�~$?b�r.J[�d�]��R��3���!�B�+JR�`0-a��<�>s�G?A��ҳ.@�4D5q���Òr�=�o��$z2iUF���J�:<ԥ�(20K>řC��ax����c>�z͹��[۩���:J~��wbX����edܭp�/�#1֏��8�*�t�����*�JI�F#QUE~
�W@@2��t�,S�����B�������/(��2����=DWiU7=�}:ݡ��@+⣑	��ABҗR�s�I�r(�&ʴ������$hJ���M��Bff1���h���d���G��͓�Om��a'�4�����:.��V"�c�S�NЃ��杚��KQ�6���a���<�:r�Dԣ�N4�����ik��v� �/��"�h�s��*#,���Q��9�_��9u�t�P{m�'�������u:PU^��קO���J�����DBR5�B{��M8s�KgJ	������"��M�8y�L�I��0=�a�Z�9�B���mhl�$�"�$"�F�TG�DmRGiy�n�i<��Y��@]bW&�=u %3�6x�R�"9�0�8J��d���蘚���g7D�;42\�c�*.)����k�cd�]]��a�����Юܤx�u(����ƕ��z6`+,bX�P��'��Ξ��{����$��QPT�e+nĎ׶b"���K�_���"-C�W`ٵ���{� ?8w����f��(=Ʋ�K�����	���^�j�n�O)�y�:��g��`��mX=�S[Jʋ�b��x���av�b7kӭ��7���"h����w���=b֜��r���m�h�ӊ�7p��܌Sho_�{��������k��du�4}��[���w�\|�OT�3-mr���H�<o�|��),��r�W�Q)�=�Z�vK
�܋-�>�B����������d�o���w��	U`���c� �H՟�j�����G`��t�hZ^ !��1k�"L�Z�Qy�ب$�h��k�Xs���؜.��j@/��a��|��Z].RF����Օuh�>�u��Ε�)m����E�'���TK��[�kP^n����*������f���'��� �TY�F3B���0���M�Kg����\[�5k�H�n��"��=c���}	,
y���g�A'��2Lx:�D��
a��D;3��~�
:���n\����yT�Pװe3��́�R26Ѕ=�^��B��e�Q^�H����|��i|�λ��XR^�u�o�BwJZb8r� v�z��S�����V(?��پ�<xD3�/�[}-�ϧ�KP�x��w�[ZX��[�-[@��iZ�i����Ocǎ�uzB+7sӦ/�(e��&���..��P�2**�1�}�T�����8q�0N�<�Q���Z��_���R8'����5�����������DҚJ����T*�v�S�kKJK���n��w�W�<��լ�h�y�JUm���^d�΂#��x�ᏹ�J� N}�E�N�]LI�)ڻ�yG.j}<<�7�x�n��0׋�?�/>�Xx�G��3x-�Ö�����c���aJ��4��{5i��w��ήNe�/,S�8�����t:l2W���i���KJ�l�$���嗞�w�)a�'��G��D��B��Dϥ��w������:���_��]<�����8{���"�|4�"����t�|��:���a��_Rf>m��9"P�m��B�Y2��d�d����"h�U|[_z9��p� /�H�W��=y��¹��GIN	�ʌ!�8���Vf;Ν�#�Ok�2KB��}�ݨ+jU)���z�a��Oc:��|
�8�Ǘ���͏��u!@�U�� �j�'Ǜ'�'L4�%tܺ49
�U'�o��@��x ���"�F��_I����RK+��
�+�U6V"^j
�V��I4�����=\���"�� �8>6�q3�����B��@��-�ڪёa�A�X�3P"�C��e��1�M��F�X$fSTٕ�	o��=���~�x4����:�A8��6�y�����1��),�Y�A7�����X�N�.�D܁kn�����
���a�ݙR�v���~C#�6^��@���><ooqë��b��Pҁ�>��,a��uz��OmFSC3:.^T�1a7Z�z5�{��?ZZ��-����;�EA�s��<=�
���`u壟�'�)���RY'�E*q��q����h��%^�R�"mA9Q��[��C���ryPRV����.y'��('�6�1)!�Ni���~���fΜe?|�c���h����]A�1����@?L�~QZ������m>���T4��+��~�����N,�-J��� }��}�R�u����[�h�$���ʼ��{�ڶ�2C�bo��&%�����W`��_�˯<�(�}�t�vǽFP�P���ݏ���?�g=�~�Zl��dL�����k|�������ƍ_���p6V���|O>��&�͙���7@Щ��R][���m��w괃��z̹�����Uj�&��W�c�����޾��a��(�J��.��ҿ(�rf�g2e���bY��䨽���������bH'/�ˀ�H\�/�p��z��#�Z-nu(��D���Zq՚��H!E�4�bP��L*���~/_4���݃�pHI[d�eu�<�͇�j$�6K�n���%1��s���I�Y�IY���;�'H���L�r��J�P��q�R���
��?�6�@cP�	,uR�P�DT���Y�/Y=):��LH��}��\��is5Q&S��T{~:�2�Bhs��jGc�L�F����"���P�Y}��w2��d�Z�83�/�3ڟ�x<n�'l,"|��0퀄��bI���j�#G�E%F#�H��h����l�٣��P$n��r3�hLXO�2KVS�2r��-+�J���3��[�� �n��K�N�y+U�H0N�K�
���#�\�d=�9KϪ�~���Ji��d /�ɳ��g�qKi]��	�1f��RZ%�C8ҙ�F�%%Bbw:u�����}���
ad�;Hk�1�Ŭi]���f�;�S�ϩ,�ذ�lyq�i|Ѯ��I{9R���ňb�g�H'���h&�����>�I��f����t�,G2.!{��.�FU8�L|�j�Z����d��%干�R���ް^��M���+���j,ͪ)����Jd,a�_���1V��6��hѱ��
D$۩�"<�c���R�r(j~CR���Y��[�7�T�H���j��s�Wnd�ۓ4h)I+JѤ}YV]u_��K\��YG��?s6���d0� �5g?Hk��FpM�Gz��H�D�ɂ2)��D�ȶK&!���X1��!hu,�����T�/������$73���iլ�H��SpX�W�����r�ZרF*�'�Ѧ��,����y:�E(3$�n6��*�t�$�U0�!Le�Dx~���?����3�a\�=�R<R)9R"fj)��YF�Q;L�yM�H�?�����2�S�ZG�6�%�*/��,�$ӳɐ�TF���xVɤ%#z�eC�&��h��B�F�)i�8a��LT��p�dO�xq�t5e�Y�4��� �HkL)�-�9�\]��疚�%k��Q
��b$a4��}LFC�n�P�%���2�;mnJ+��S[ė l2FQA)���!��	J@\�WZ,�m.��1�d	�e�}R�U�hlL��Y4a��ɞ͖���JT��f4��P��V��V�~�%�͓��eyB���@CM����0*ge&�,��nS
V�=!�6�(��V��&+�M%\N����m�c�){r���V=�Z2!M:@�)㽍�g���<��h��l���SFH^�'>M�Lk ��"���ͯ�˗-�H����ƥdI$�f1e��E	Z'G"�v��4�9	}:n07��z,���0���D6�������(�:��0g	�-��[�ƔL�~fU��o�Ȓ�g�g1�\����L]D.��#o��n��!�ae�
XR՝���	rK~��52�C�C���ڕ�W�UfL.�*YAB"x�OArH�PB
�~�n� �gx{��Љ�7nC�C��J�Xm"*�&՟�cF'!pL)}6w؞�FW��I�Sԉ���J�T��q��oS�#��()�=1\��g �� -q�LƘ ���;�j8[&e�6ibIة��«�1�Y���QR�f�`ƽՆ��OSv�	��k�Ôְ��%���%7g�^UE�L\l���M���d�yB�UB��%�/SH��@ea�H�G	��섷�ݐY�f���� ?}�'�jkk��{1�;���H���~K�=~k֮Ess#.w_V�������*נ���DB�TJ˚��Α���`1bf���J\�c[6C#��,�aQ| ����&i�������,�tTE�|��,n�U��*LQu*VIc���K-�ɪQ���VIb�<u���
�L��^�ΞM�%4BW�+��^��XZ�RY����r~���O��,S���dl�_D]�#f�+�6��[��}zC.X�C�)�e^A�����Qz̕-�-���Ve7)���o�[��������R���v.BW�]Q]Eg2�q@O��c+�����BJ�UՖ�1<b��i��U$&�H���
X�����0�6����\�.r<{"���A{R���r���0S`d
����ƷR�����ԯ���D�'
@��dLI�w�*xoA>b��z���[R�A:�DN�d��WR�57n�#GJ`'���W0��?�C�D�*eڶ��ɐ�OwPA{�>,�0R�eI���+�ܱ���ֹ�?<��Kt��D�G���@�C'N��w]����1b�8]�K�-�/����]h���>K-�G���e�/s��AKK+^zy+���:�,�P懵kVkX���cZW&��N�6p�|�ZD���,[~�Ny>{����S�j���C��$�z�i����6��y���;5v&�&x@Ǝ�/���jk�t�VoW'��JU���D8�@҄�XFa��ֹhjm�fG�6a`Qν�<�K���S�+��Ŝk�Q��>�!W p"n�CY�%�gi4���H��.-.����Ȱ�T���
}����Q�p�C�TU�D���;:/jΜ�ص{�Qyaq���ݶm���Ŧv��G���v\��j����D̆�;g�,�����
Y'�R��X���2���vC�SҚ��PL���^�����]v,Z�ˮY�g�}A7R�nޢ,�߮ �:�i������^���<��!t��,�t����
�?���2@�����0g�t���3�S-�P���A�X���1���s�ry��l}Y�tҢ-m��9���jA�%[
)�3)=2����y��|����(/�R~�KbZɠ�vӰ�yJZS_۠����cZ?��ܦ(IYp����S�z�Jx<n��cǏ��R�,�r��@�W�	��M��z�|��|ٵ��B����)k�������M:�UF}��6���x��T����Ʃ�sAw�������J�dȽ�^z��8H�"�Q����#���8���%����jq��)c̻����nô���Nj�}��q���$�+���Zf����ȇ�uG����\ a���)ʬ#�m�g�!�5�שm[���*�)4�g�Kq��v�j��m:�j�P?�	'O�5�qʘȐJa֌���J=T���,?���Os3�Z�)��K�0�vJN=\�j.�8��D32<��ׂ��J�𡃔�B�&ȼ�?Klұ�'yj�)Z3��9� ?7Z�U����0�ՠ��^ͯdL6)��}}�1���E�H���&q�<��� �>S�C`��|�?����v�bj���f�Gy<�Dy�8�:���>w��c
��*�����1]�S!L^�V���4��+4f��j�yq�W���K�mz�N�i�%�>>6��J�湉����Dw�yC�#��.^��E��8?W�gk�SKg��sq���_C�D���խ�\���U�E*�P�tڡ��n�P������؈��M�=� �OYI�xi���]�gQ�S$�l�QXI�	���������b��X$��{��8nps=&bi�����.��,��Գm{u�:�fLB�l6ۍ���?ߐW]E��*���k�@`����1�
���	������:ih�E"�uq���p�CD2��oQI�n@k[N�9�c���C��)��6f��gR�r?���'N�U
V���H�J^~��[�abC���ǅx��Oԡ�g��k�'���c_G�0m�Ltv��/ �����Ι7�Z<���>�&�	FF1w��.%��j�LJyLZ`!h/�s��{� 0:�MD����@|&���T(@}K��K�-<6	�6Я[WS]c�FS.����S���������>E�U��Ӆ�5Y�y6��csp7�D�&�HaIE�������nqX����MI�y3��ݘ� ����.9yW��/8`�R�R����k�e-Oű�G9=r\f�@؈S����b���H
��ix[��x���×z^#�gĖ�1s�L��q��a�R�!h�
��|��$�:62�a�Ɔ&r��4�K_`<�51�!?m�@]kơc�����0O��N;x2��5�D���;���r����*�~{��o��v��E�i��Y�j~���¹ �o�/�ǅ�N�?4�ڳs�sxx�Z����i��A@��;ﺽ���)h���{�k�C���F=<AG(A�_����f�c��aG|ia��������'�L$m�� ma���!�OTTTp#k0AH,(F6���@�d��Iw�Ph��Yhi��v� ����rt�sM�6�`�e�,��L��܈)y��Ր]�NiIծ�ղ;���ŒՁ� 1<]h�Y
=�@<�g6Oy9�*���z9��٣�'���ۑW�����&U�#z�on�\_{�A�<y�.��M�᾽�1�pxtd4�皡#�}��J5�q��HQ�Q������p�8%BB�.JR�V �O�P�Te�Kuȱc�5�"�'O���8q�O�d�)�,�c'�H��H/u�2v��'En$F�C���f�8y���oI�P�$��F�@M�q|�(�58}��r#��\9r���QGwr�pR�\8w���n:�|n���fx(�v9�f�:�"d���fȵ��8ymۺn������/9\��:���h2��on�\ӧO���ZHL��i`��6,�%S�d%�����uZ����#�o%'�0�K��eq%���k��RIY�ƙ�<!��]Ւ@N�<Fc�y�y�F�j� �Pd�OI^��O�D?���T�{D�ķ,f�ե���Ӛ����c��&�g���i��<�V��%�}A|�G?�M�gW!j|Ҏ����\3n���3�����XU77�-�V��_�l�p؇Ϟ?����IrIa)��\J�8R���d�cF���&љ%���NB~�t�ٜm.tخ�~]����C��R"��"�]6�E�Al���e�5bm6~^ǇkZ7�o���R�'�AX��y��J�����႒Bu~�{��Ǐ���g�,+Є\�"�!(�m��8�~���]=]�S:ׄ����X����G��1���_2�f�PL�āub�DX\�y$��T�$��F^B�^�����,甑�#�L)#�*FXT��y�b�w3z��Ň�d�o���P.�gI��l�>�I��J�fB���%�(Er �*J����s���͚5���4N&C�eϑ0�\_hC�������O�:y������Ο^����1��f��jOfbvq�bј�)��x,f�B��Qw8�R�	�I3�i[ p��d��&c�F�VɆ����R�&z�����f��ĸ3)���D��pZ�����6\I{�G��$M3f�%�d��CC��ϟ;�"�.F*٪��t ݽdɲߨ�O_�"˦s�/�����yb���'eWrr�Іl߱���.� ~��8���q��҉WO�b�h?��4��B�d	�'��|�>�h��S.}�v��W6ac�ܗ�Ņ���	3����g������i���	[,�S��ۤ�B��h$b�j��{�" ��j�rS6K^41Q]�0�og�e%�p�\ΎC�����_~������/r��MAaa!MSd�'����ĉ3:��m��3�$�k�p��t��5�W.%�R�#�vAD~�H��D�DmIY2k��I�)������:}F'4,�EL��'��o�O%C��ҭ��c�R��$eˁҸ2{]�''�85Q�\�1�i�O?�z����/�����K�l��clb_�Z�`֮�n������S����{n�w���6d�����uen9/	������4�B�(���a:��&� =���
�1#�����q-X0�>�X���4�Z~9�|���ِ�/\�)�U�ڋp8�g4�����' ��7����u��!�9�?'�q���!�/�Xs:������kC�']�]C}���}�����?3���y6    IEND�B`�PK
     ��Z�p�Z� Z� /   images/0c8b7e0a-6698-412e-96f2-fdf086dc4925.png�PNG

   IHDR  @  �   ��t   	pHYs  �  ��+  ��IDATx��I�l�u&�"b��<�=�y-If��6�P���@�T?A��/��#y`���75@���M�-lZ%@���o{��f��ڈ�y�#�B���ʽ�˛'3w;�/��ĊYd�ENT \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENV \d�ENVN
 �����y�����w�!fz�߼���� ����������?�����o1��|�)�>~���;�zݹ�������Y�t�%�����R���o���~������o�}�ϯ�~��"����w���~�m�����.�ܦ�����!��7�S�^뗗+��v�?���:�WY���?r ��{����|���W��{����Y�����)�i�1�o���.�_�/��|���p1f���b�)�i���w��:��_%���뫷�'Sz5�CL�⣴������>���ܕ�6�G��\�s���t�ԅ�������|���x�������x�o��
�/���B�s��\���r�����?����A��ǿ���U�������S��|����������@���������?=:�:��帯*�/�&��{_��O��
��O����	~|�?��3������5��}��w���s�d��5 ���/�+������^����7W���>�Rw=���0N����B�]���s������!�)�I ����sх�Ot�ãƻ]�w��G��.���,�����R���k�?F x�����V&pA�������	�[/tx��ns��1�b�~BL�Н�͘�8������9�r�bw6�ݛ<���݋�l�os�
y2��ur���z��ǃs��o<���;���zߟ����	v�1�ex��NT+�ۿ�b^�K|�b�y��������C>� 7�>�{w����M1�n6�����n~��'�����o��;(3�����n8��S<��_�廿��ϯ��&��w~��+�� ��Ӽ9��n`<��Wp�
��/S�2�<��Gp��p~q����7o`��_��������D���_�����{4���$_# �l�X>��O����Z���?��?�_��_^lƴ޼z�W����˛�����1�k$f���il! ":}�'� �� 1 ����>���p؅]J)�)zD���X�;�ԭ<��GO1<� U�̀O�b==�%}G?;D5:Q�A�# F��xKD��T��\�N,_��|���"��l���Lt�ߝO\�T�|,�uN��!A��������︷4]&2��{8�d���F|��c,T�������p�������7�ʈ��v��c��R��Nʻ��q>p�R㈕��i��X~JX�xS�������>.��m��~����>�G+ o���u3NHØ�XW4��x#����](�_m�r�'8,S��L�����q�g���HπM��.�=>��q�v�Yw?�������O;�=%��S�v������C7�ٮ� N����<~8m��O~r�V11��}�{��'�_ �����A��_@x�?/��z��7��v?y篮���O���g��v�g�lv�����;9�?q���ti��w�W�.w�ݓW��'_��~���4��'�K�kT�V"
� �s�N��i� 0F)� �!�pWE4C��)Nހ����p�z]	tX�ؖ�B<.|�{������	g�zt$ �������x��D&�Tv>�/��$סgpt]�ށ]�@��o�gw�(z|0�m�Q8�<���=;���9f��A>Q��5�zޮ� �s�hn!:�� � ?�i��c�ޮ�:p#X=A�RV�ߵ��<GeWGmG󇧉�	@{o��Y�c�kjR9����/�u����L�tށ�����	�+5�w��!�q�S=︾h�$�h�Ł���'1�p[�C�V�{�<`���0��=©;`9�k����1�ݺ_��.����G��~����?��e�_ �v���_}����0�/B��P�z5n=�s]7y��ms�v�7`'X����L:��M�c1ލ�_���i8ۏ��������᣷��[/��߻��S�ę~�;��7Fǳ�0
>��j	�����H�:&�Ա�W� �X��D�"�C�LF�
�ܕm�
b�V�Ƀ�����J��N�f�`���V�D�:��,�Ƒ�r	}�y��\>T��7Y�^�G9_�aH�ʿt�r��ßo�����nt�G�(��.%�Sٙta�D+#O>��^�3��ef������MrjS�4��̐�
�ήG��� \in'<*d>R�@��Q���,1��ԃ�0g�\˔�=Hi��nH��zd���b�HƓ�<�q�H4�e�2`꽛���G�w{�z����U���|�����߼	�n��a��0�?������솿I�T�߷/��޴]�������?D���?�����퓻w��a��Ҹ���WH�W��a5B�j��]�|P[���j���"�c"�l؁:v+
g����v�{�A������C�t;�sT�6\+��	J�=�$ǝ�s<�2Ƞ�~��T�%�c!ތ;���t	ꭄ����z���L��)j��ں���X�r\Ǆ��I���mx2J��Ot�(Ϡ�RP���`M�y#D\�;5+�Ns)���+�	#�� al�g��F3fU��,X>G/�I�	Ҥ��y9�߼ '[
����sJ�ДY�`UR�_�Nq�=]�$"�I���ts�0T'pN�ы�&�S�5��2���/ve-ٜ�!L� g>�	�g�6M@v=�|H��;�}�U@ \�o6��W�~�����ź�xW��)��ϯ�O����'�_��ST�� ��5�'������7���_L����Wq�����n� H��ӟBwu	�|���y���n�mw���n|2���v7�#�m��.�js�&$c;G�㆘p&��tC꛾�nX���i����?}}s������.����爙=Be��M��"*!�WrWd�RhxQmV�&4C@�|v:��
�|D� evt2���8�S�����s��x�B=(�mg`'<����W�� �\������RD��@TZr�\>��-�� �P(TR/��Dy�k%�U��G�;���:�����M��O�G� ~Rf��5\��t���Z�Z_Mg1^h%��pR/��rc:�=Z��'�& O5������]H�E�D�U�0H�D�="nܸ�ð������<_^�������%~�0�z����`�1"�OV��!"���T�"ow�N�6i��i��p��/����CJ�js�~��	Y���_[F�h �E%
��{�oϟ���|�ś��ܽ���v��`�=<;L��a?^��z�S�#��Vb�q�	��B�vHa:ɪ�7c���p��v��O���;ߋ�����sdX�:_��H: ������\���tjWZ3r��Ç��B!��p/�H��r��8�Rv�HnWw���ͅX���Oy���N�2�]< �lTYi���Af �o��q�ƴ���2W}v)G�K3�g���ƎO�N*��^���6����`���7�[��9���)��k�ff����l�T؝AB�>�tґN�=Z^zޮ3��S�l�[�-�{�6kw@��{��.��!���k��/W��Pi�Ժa �{]SJ��]b9�Erˮ*�p�Z�n�>��A tdE���|�����r��;�������;��Ϫ��k��� �_}kw��z���ǯ��|�˗��~���7���~�E�v�+|mv���C:T���D%���"���_��Zw.tt�C�V��q���4�.�h��m
�l���*����%
8�).�����tR)N��j����2��M�p�q LuD��&}�3B�`96��F'�+(p;��|YG�h��gX��Z/\"f3��Zf
xX��@'&�=�FcV��R���H0���o��u�X�ԓ]6v(�%�۔˙\fe���ƭMR���?�+�)�C���˱2�f�X��|��'� �0T+�ԡݟP�4Q f��_{��C
�U�ݥ�9��_�x����F��8�2��trMr@a-u��^'��vXv�|��k�C���U�5w�u뛳�xs5^!����8�1��;�5�G���g�%\�߼z��˷�o�z}�O�x��w_�����n�b��]S�X=l�@�AߓL]�ˤ�Mc�:n3S��G�m2!�`c�c��#�s���yM���;&�b�6��sH�tU}<B&���µ��γW(Ke(�����~.�P\� �[
(�ﴀ�j쮲T�k��P�[j2�
Ol����f
��/�R
E�l Ȇ<p�¡j�BP�:?5S{{���9�l�J�
�N.�g�+YJ7��*�5����}vߪ��q��Z�K@�P�� sd`�ggV�l`=V�+L��42 b��u��Cw�����K���!�;��#E� C`�4�L>�M8 �ŘY�2X�K��;��l67gg�w׿Nc�j�v�6�����?�����������6�ٟ���ur�< ��U��|}����������w�ٗ�z���77�n�O�x���c�t��HۣI�q�J�yo6� ����z@L�-�\�V~�0���	9�$;Uy����{a2:��a�L%5�f�r(��ƚ����J�AW��*���V.u��AX�@�m���Fgθ\�nsZ�\[�0UG
�5<��s�7����D��J]��T�
 �sv��^�'�:�[p��o��z���U��S�	�g�;X�45m�j�J�MU���`���m�)�� `��|�6�J�ψ^Tz��tU��瑩����
�9K��<�㐦��	�t#T{����Pb�e�NA�A03�`��98�V���E��)�F��%B�8?�x�rp�U}�v�����1Y'��ȣ��������~�՛��}���w_�l?�ݎO��t6NyEZ/�;�Q<����:�bRߢ�/�*Z��h�B⎏ ���*���}���^���X�����r�1�ܜ�u�1�6�W��6�̙�h[����6����4���L�S�|�sfcԪjf���vV�#nC����j��8.�i�Ђp�ח�
�3��!�6O8��ֶJ���׿�ͼ�o���ej��.���N66a:7���˵�:ٙ6 `Z���zJ0:_�k��D�8w� $u&@���L���Fדu7Ő�a5�S�)"�iă#�r��� L�mD�a@�����7:!hN��j8��~�^�����Wi}=N��ڥ3,q$��+�?�я��5�=|4 t���&O�����n�� �ѻ���vH��=/C D��ě�q&�q��������N�r�BBB�^^���P�K}�l.��x���d@��t�6�u�k���s����w]�i1P?�Am��P4 ��3W��U;G��e�:��m`P��Y�;��}ɟ�T"$�D|#�á�A!��g�#�;�zv�g3�ۉ{��x��3�7C����0�홏� �1���+�[���y���s�J%�[C���n�Iq>9����05���U��{6EI����F9Wl�	���]��[�a��]��[��si8����N��dov����e�rUv��R����w7�����������'�ŋ�Oήc���]��y�����>ہy�Q�; ���3�?���c���o�����n���V@�Èj�#c��+N�ò�/�����0��d �xY$^�! h�ҟ�0'�.�}�\�/2(�!QpJK�j�an��=�,��Rn���2 �����Z���
�� �awe||v�|cV��0T�o>	(;��U�Wmz11���x�׮�cg�)���Sj�"����:�W�{u
`�ʪ�.

�ur�h��U���$���58v�^���yNsx��:����� 7vA�<z��2I���х���ø�0���pS@-^,h��P6S�^�6���ƴ;L�n/�8]"Q�DRr������k<��f�C��j���J�C>��w $��ַ~���mwyws���0}�=����p��E�A ����<;�aL�u'3�/�Ol�^��r數�_�]qb�`��ɠ��[�6�k�[��]3��V��JITm3$�'P0�r���>I�b�3�H�{Ҙ��IE�*,�eCv�<Z_�� V�4`��F�d�<���س���ֿ�- h�C�<Or�dL�IL��i�WS��_�v���뙺�O5�:��������Um����of	�q�LD��zlJ�N�R��H�@؋L�7	/�ymO�1��Թ�|�(�yf�e�2����m��C3�F�ڙi���z�0�<�1S���)����.�Y��.mSt��w��sG+����G�������p��9^���0�g�g�以�f�r����
I�%� ��_���u��L���&t.5U��/�IU��\��t��h�U�����8׎��^5�V�
j������տ���Y��\��(q*4���QЎ�R~a3�Q
�s	��`!/J�yI`Iu�X��וjr
~2��ʼ��׺p�&��m[Gۧex���h�Q�4mV�o~�.P'H9�h�j���7���n��Ե>3@u4ى��A�Z�`�K�;���:)E9�@-��#B@"�bc���]З������z�2q��1"Ǜ�X�~�7�C՘�ō��z�݌ν��q���я~4�ɟ�ɣ:D�3 f��5��M�¶C�1�sTW�䦐�և�Fbk#��,��F  $���2 "�cԆc+(JJ�+���WLڱ�	�qTm�*����Y2#m&mG}H�N�=s�ؐ-(fΉ_sI+�,5���d�#�j}4�qH.NT]^�e���$Cǫ�dxИ?1�S����2��j.)X��C�M���,���'�u�<����{�,����q��W+�d���R_"3cЅ�'�����$��ͼԀS�l�8ʦ���9�@[&l��"om�+�%4zJڿ��"���wp�/��ʢ����)��Nb5e�#�>:�~�2�����Z�6��ͺ������q�ߦ�?�ͻ���<��_ �Z��K�OV�.�n�j�6���O��Q�L�q�Sf Y�+�}'�^z���#/H8L�S���]��Tf�`_[d(*���+)S�3�1��ϝU�cG�����g���\�b-�+v> ��19�܀�1 ��:T�q'V�r� �#�=��D��d�"��� ��|_L�\�ˊ/1K�D�e��<�NM,O	i�c|p���\Y�m�M�W��6L����=ZUz�봽tB.^�#&�@?*tL?�>+5ҚvxȨ��ۡӑ@ �梩� �u�>s ���I�^l^��غjTHjv�\��#�P��6l.�WO���sԎ?���AH�u���n|'�(g�_�w�
� W�=�h�e��@v>`5�M ��L�3�������/�Ob�SV��DYW�}���c��v�ʺ�l����%� #H�t�IU =fZоB��5��:}2gNC�y���^�M�n�z�Ǵ�˚M Y�33�4Q\� �x �"/G�x>@V؜8�p y�Լ����MJc�Sa��x휧uf�PHl�-7`/�Q�v�gcgY���9���>��Z��ر��� �1(Zq�p�:=J��N�y��s[_���%�YW�Z���gz�q��1�j[,^p{�dKx��:"tdՙ�u��V�8�?L��y�]aw�6�/�)=�ѽ�Y`��V���(a0����0�!�nJ��������JA^��?�X�<_V
 @.�ӛ�k���3�\#�r��Q�p�.l�U6Q	C��e�U������&cW��
�)�]o�y@-�"ו��$�`=B�����߬�����~H��d9�8�+S�Ҥ L ����#|'b��/�7�TV-il�94n)�Y���N�Q����;��z`P+�}�6��\���\�1��X>���v��F�*,�U6�j[@�����v[���(���Y��6��
����Ǥep�r��/��n0q��5��$q
t�qBu8�8����������!�k��.=<��w ��6��wCNn������,D�	kp�+ר���w�<l��VLw� �k�V0�{UJ8�=b2�Tr��o[�Ha�ny��,�/������ـ�{�\��ٸ&���R@�V;A7c�r���}eK%>�a�P�g��rgl��Ff�	��� �����c.O`6"��J7�WLf�N�L��P�T�˖xͲ����[�y��h��R,@����� �w��8�bq��_&'�S��o��Pg]���ͻ��K�x�[nƖ�c��`�V��/���Ƭ�����-M�+P���h��SzZ�>��G����v>_����q��G����>�4�|����!N~�	�O�y!��6�b�G��-��D���cVs�M��
@=�
>�\4[�^T��N[Ն"�0u�?����|v�K�V�)?��c�2�����t0��y�L�n,V��f�)�J'���vF�������s��m��j�s�ڑ�ơ*��@��D�9�[V^��$��t�^�nmhuo����3�6���\3%Ȫu\(��Iʦy����N�:K�%
�`���Դ�ՁR�� wM0kl{���������G�tZ0�����w7����X5g�&�O�W�/������`�Bm��<���%�3Bf���dʎ�s�#9|�r��I�w�� �����nqf�`��MdI�����#�,pf��G�&6V�@Vpv�k���� �[��g�2X	V15�\����˷S�*Ievn�������=�AUˉ�P�@/�>�4V�u�����3�� j=e���\^��6���e�r�Xc%g0�u�tp�Y���� H�@C3e���c��$ӿx�����B�e�\;�Օ	�� [&�\��ff�|>�l�3��b�r=Y�'�\VsBj&Ѐn7{j��jư�Iݽ~�t4m{X����׺wkǬ`嵭Ծ'm����9�'f{!WS*�(��1������,�8	iJ��W`�c����_bK\fd��C����86@������O��z�S K�i�*vP6#��kݳ�D^�T[(u�� �T��!��<��g���F�~l�,�ql��ҮN��r	��29s:��������TB~X��U����u����6MB�\�����*`����76,a�Q�O�>#10e��7�L�	4�D���X���m��k��r:c�IˡIl"S��Q{^F��[�+�_�}��8Ŷ�l���j�	�g��m��ٓ�l:������6���d���멝;�3����(
��匞Y~��;Z��}+�3�S�ވy�
�`}^ ��3N�x��/��y��# H�]x63�ґ6$u�V�s���ѬEFuo�伵w�|�xց/?��| �k��"�{v��&[ͨep�|]��x���}��N;s לZ�?���L��S�X�(�o�n��xSb3-���K*cgk�Z.��+]]9sa�Y�i����a��+�y���g�# X쳹*�PT.��i�z��A3���z[��v-y~�eeB�����lQGqR�ҋ�`�u�̠�4��>aWy�TX����l�������׀jv��u�y��If��}&�	�N*�T�jLż��U��5�X��p�xl��m�rgS�N �z�v�Vl�tbF�,�I�J�Mm�u�2 
�V�67����t�2<��3���ԯ�8��������L�s��A�Tz�l�gBd�N:ab�~���a�K�A0w=opz/�fv�8 ����ƄŔ )�$T,d�I�<�{95�7�Q�{V��M
j���Z���?����~B�5�T^9˫c�]5Ir�%�U�g�2�C�e��[�*�n���u�E4��=�є�j<g<~�+���}u_-U���>�Q��<�aI�)�h�9�U	rebK�I�F�!��.c�����T*oy�c?��o`<A�l�8O�W����"K�*tZ�kG�ꏫ����O*�����t;S��~�����8l�8g��2��Ω����5W^�\k�q�X� _"�GVS؛����6t�^N�p`?	pJ	��$]f�e����.N&�5+ve�-R����y�z��6��ni�b�׉� "��2dln^��*���Z̲,���Kx�Ԑ��NXg�L�QN@}���s��T��Ʊ�`,�6��_7�7)X��s��k����r�f��R�Z?���@�b�,u�<iF�D���t���b{���c�4�v�\q���&˦��9y��쉧��C=О�Q�f���-�SƂ.e�Y*���9��M �1�t_)3u�y��o����V�'ߥ`�������V�:�/�q�VX�_����G���p�Y�%$0�Q�{���^�+Q��,=�4I�*+vc�Tߍ%���5�J�U���h��e���/�h:kǦ֭=����f�z�5=�����/:��8iL��i�}��[��9��T�RL��
�ځ��2��*���U��c�����>�`L��&3�܌)�@��t�Ic7��Iu�qU|��mv~>j ��M�6�dM+�s�P��9�f�_o2�0)�e=�k�+V$�\!I2XlpI=� g��
�}"DZFaA]e�U'i�e���T�g������z�%^M�ƕ�)(����ҟ�g����A�����I|]��$��њj��ib�܈]��O�.|�]Ol�n��>�6 ��b-3�C��^�S�k�DP�s�
�[��e��̚�u�� ^O������l"�@m��T��ԔM�VPϩ�8	mqj�����3�ve��aG�-���߶DSg��~���T�j���=P��\G��Bb&��D[�Urp���6���b7�d�s���!_������^ �M�t%6�Y6~���(5��q�!����ֆ&�̘_>����~a���S�y0��Z
e~`�M��f\'2P|���A ���� sl�T�2�$ko3�uc�`�L�g�V��Ӻ�̬>�tlw����r�k��e��e8�z���#4.̈́�ֵ�m �+�Kp�e�z��	�����Y�c3� �R�5����@q	X�6G��m_'�R�J�x�ì�Tg�k��Qe��+�=v(� Xy_Ak�x�����W���b�r� `�hz
�6����|��s_9���aw�Ɣ�3ux�ޝ�R�o���7��Y�冀�И>c6�Z��tL�ܹ��P�qv�f`(s4�5�p���l挮V���q�D.Fy�F�D�`-�g�J<―AŎbwV�$U0�@c��͵<������2wf�ԅЃex�U��l8z��V)JrZrR�U���:��K.i��mae��cn�U`0��$���W��S�����,�Xu�V�I�7J�&��{NT�P�1���ȕG�xn���r���T�}K�Q{�;���S.s��	���T�@Y��&��(���O��z���Z_��^/cC92Pԯ�W�; ��g�a��	�j6�M]V#����3� ��������B�ь�같��l�~Gs
�5��)�֙��j�\ם�C#+�e��*���9�u�� u��1v,hK9�܀�o�z�����@V���	p�5p�x��n�o;�+o����-�S�gk_m��fə��<��w~~�C�$6`̲FyT�QL�A��MM�����I�-QM�D���Pr��)���yT)�D�W�Gu�-u�?4����Y�m(1�-I�&�_�����/2���"�ē;�J3k'ҵ�2�7�X���@B�Ô�����r�9�{=�Ƞ������j�?N����l���֗7S%�ɪ��*p�K����Ֆ��zN��J���5f�>��$i�j\PC~��U�6�<�I�\�晽C��� i�Y$����<M*�z@!)�/����"��Y���Gu��֗k�w�uj��z$�� ��p sf*�g^��CP�2Xi��A�sOr�eE�r���W�/5�x67�����O���0����+Wm���Ә������o1i�
L[�Fu����rgdD���7���
l,�l����ok���P ��ɺ:@�ωO\� �f� -���9��1@���5�:SK:Q�n��i~��t�s��U&?e+���r���*����Zҡ̦�վD����U���H*01���R;�����w����4[���%]��{�&P�j�w)D5�������l ՌPePY����h�
#3��m������ܳ�Y-�bp 3�Q�@�#33&�3�m��IZ~�� h�gQ���'�[I+���(V�p�Y��o!Z�2y�e���YE�b�J��0�+C�zX%�3�����ƻ�i�A1�p{۸-�58�.v�<�<
 n��O9�d6����+c]N��pj��W6�5��)���7�X���rd�,@�?�f`/�8<o�T�z�Н�'\ٖ�٪���J�!6�#��)\_j���L�	�uh�f�d`f�����|��,���5m��JeT�M(�2�V�m����MK�A��m����`��V|��
�}o1�C��d��E�+�Pq8+�+�Ak�7/p5�F��l���&Cd?{������>�����L�NK���Y��;�ȣ
ܱ㭗��\���j���^(䷵I�q��o%[Ǆd������w�γ�h��$i�R�F��ł��A����?
)�6x;S�~ҨWm��l��	��l{S9�:���i�>�L�:b���)���3Q�d�&Z9J�yՇ-+�1�2��@%�[��V���{h�98�H��Rg��� �ȳ�	�:����5�N�'�)�n�8� �*{�ˎ'�<�������%OO���U�@P�2�k����PZ*0�:��1r �T��k
6�������dS��ؖ�Kߓ��������oYٞ}U*k����Y����:�C�� �$�(w�.�����s�ܟc�R��]}�L�V�:�Ek�)�1@��������w`��-27����rn@�@�F�� ڬ���9��ex�c��S��v��9�_��c�)w�~g� �Ɉ���Uפ�������<WR(�GW[����������>91)�-��������=���6�V�k�)���V	ez�54gp�PۯLn���l;ͪ�9���y���x�}��mB��7W� &�H�&!��������3����*�M���S�N�9��I������[S�%�+�U�]S���ߵ$�� �u�!(�KE ��+�$I��M��ɲ���$�b֥�\h|ʄ{�6��w���mH8�Fd��Y^"0���~�����;@�6�X��43��~we�5�J�"�l?��e�)��N+'N��%@�뤚'^5��ɵ~I��[X�����w�SO�%�
h�3O�0��0��I��l�'[q`{��V��M��.��\Ê���P{�v�K@*w�mg�D������)kc��:�A� ,w]K�e�KK� �٨�x�mc-p����N�٤��K�N�l:e��^*�*��-�.��
���Ρ��������6a����]Y̥(�/Ο L9�ƞ�vڴ���Yb/sY��W;M����p�{�z�u�-;J�Fk�s��5��F��ը�5Z��3y��� hpM��;g�֌u����b$��WQvĢ�Ȓ�A�HA�8P8SM���x�,ȕrWf�A6h��,��b�؂�) �udèv@#
�戉�0����(Q���Z{�{���n��ֳ�t�����&ZNA�ŚQ��֘8ԡeW4<�ق���ƶ�̀@i�g.�c)�NS�aD������g+i�]6����kU�u��(R����AC�f}n~��F �����J���kS�����-%e9�M\T��v�3)`։�y�\�B���zU�; �:�yב:����ײ��TYY���A��3¬l<��b*��f��(Bb��Q�6�qʲ�]� ʗ&�-1�i�U����E���=�&@�ݎ�ݯ7ЭW|�XX@a=��N"�����Ô-)��`q�"T#���$��,�2p�^Ifa�F,���S�����G\gt��Y�y��͗�%ѫ��'�l�#jL�%k�~Q۷��*i{Z��5MQ���X07���>& �J�8 }�����?�gSb�R��+���^�X�� ]�ǰX�1�A��9��*����a�M�����:IAnx�WB���9���<�;���/h	�&��m�m���K����x��`�4���a�,BbgH`	�mf�0$��3�׈k��jGc4u�����1+��\�'^��l�֖�R������j�:ylـ��g��C�>���y�t�j�Oʸx8�$�e�w�[�4X��<����~WTQ������r+��k]z~�K����;��,��UUԒ�+T70���@W�٘��4��Z�N�2�Wy��o-i�2�ȡ/��u����MH�xX>��x$T���zL��n�	P؛~7�.����}]�=t�j��v�W��՛��l�0�V�ԛk���le�z���c��l��LP�+� ��[�VOx�`���n�8�� Ũm�v �TW�`��Z���ÝA��S��
�eLQ�)��!�)����w���bO�zx���&D�~��kN:0�7�g��e��e�te�{� ���#�����#U,p�Դ�Ov@
i�d�J��������p7��J���d���5W����2ʙ�6ԁ��g�[A���t�(��$�!Y�0;\3���$�G�̎�d��ն
��ͥ���*�3�h�t��vG�����T�Su(��m2�	M��i�����	��#~�,iI&��ٱͫ�w�s�� ����%5iWK!�	����ŊpW����P��YMt6�f��S�4�?�F���d �R;��|�$�p#�� �����|3�s$�'Sιa�竬�֜o.�j�/��}��
�-3�p����n�kV��F�;lOM�_*��!�K!Y�^ջn@Uw�Pl��B|��^��#A���^'٪y�$/�0�k��;���=�,��.=�"g�d8�Yr'V5��{gl��_�F����BD�´�o�p6햛Х�����x�k+�d��7H���f�V���W�G��7fm^-�۵����Z�2�-��Q�િs�|N�5��V%N�s5��K�I�x<2�l�ck���RƝ�YueAv�uµ��r�ժ���8�&){˸�-�+�T�2��v��|e	�����X�ȄNTa^��5!��p�Epe�C(*�L*�
Oe�*sѼ�$���Ձ�fF/\c��g�����,���*��%�y���j�fW���N!ר�cR��n�VB�P��o�M����@R'��i�9>�n�i�M.*�UJ�+��+����V1�ă�&��͆�;�����f�Zw~��k@��Y�s{NQ�s���|�*t�Ml<�Ӊ1����n�G�����[E��+�g�FUs�9=��XE/h���l�����eXN�v��U���҉���0��9��ۙŖ&a���K.��d@��ĝ��9#�'��@�s��Ugb�Un�Xc/+=w�[�ly��Qs�Tﶟo.u7/�s�v�Ϯ �k ��0X};�4"�,3B����D/��AC�eB�	�*��u��$�6������-��!�z��w�9�����D�،�	�y���7[����R5�e͛z4I������V��7;:�7�?h��>���VD�W���q"��A��g������w	{��>U�;n>;��g��lP�أ�v:��������δN���Dפ���V耢�z��S&Hj�D������������i��F3���,R���� �&�	t�/Rrj�W7���`Օ�zFR]l;�e݌<++��ץ% lG���ǀ>�-j�T�DM�9|�N6j���$RaA|���u������Ʀr1�G�wƨ�}5��0/���m�(sj���;?U{���mp[�1�c���m�^�-�ݼ^g���#1@���r.Q��<[�$_��ѫFᔙϘ���������x)K�S޿��ggZL�`d��?7�=��f�Ԝ+7�V�Ѐ��և�?�ԶL�nv�.ر�A��w|�x3:6�α����$�	��A�����Y)}-���ҶӉ�e �A����¾�A��U�-~��2JL�����2�������Ɵ���!��T�Nv`c�P�:��=f��	ΰ]�s��^��E�mO�C,����C��leI�{���A6<�|��T��~-ːŜ:u�8�Q ���(˱�lU�����u�ib~��g��lι��͏j�R{�W�4`�h�����s���	��Y�t.�p6yLӣC�{��s	�Uuo�Բ�� ���
co$��aft�B����f��]� �Ѳ28aE�@�&X�u�+,(�q�^�������8�����C;Nd@*p�Y��+�R�}p�[ߛ�ٶf�����"�*� �5a�xeY�T���v��1�ƬLm��cu5G��By�d�۩o@���@[�#�|N@y:��?�-:ɸ�&�I�NRϒ��-9sI���,�k���RT�ov��&5	؊�g���kXL���+nNf�/Ε�4�j�C(�u0 ��g��zk+�S Qp6w��JOy���N���ړ��P��]5q�r�+�	���ѱٴ���T���'�3����b,��R|���b�u�����2�z�6����v����}^���M�<��ͶI�:xo	@U�b�b����O$�&2���O�Ie촠t5�����5O�p�ڷK8��\u�X($ƭV���%��~8�QT q�u���9�ǃj����N�԰#Wcy�GI��7�b�]1�ѽ={���Ak}�<��ܫ���S�@��4��>k��e}iWI��˪I�u�(��j��`�HK�^�@���h}jn@?7k��
SH��ӂ�\N�&kG�G�5�횘KznW��i(P��쭠�f=�s�=&7c -%m�0@����fr�D�z�lB� �{����	5HG���bFx�!���� ��d���f����5����\��v$i@�?J��ӕ��O6��Di!�nL:���)\_�銑�޼�7�n`��D �*��Ť�JV椏�Kj�ھ��J�AO��F�w%6:=c"���3:��x5�~H�FQ��E�4�i5��P��$T��`CW���	����#�
�s��@��:iW���1Y	b�AR���
�`�y	G Tv��c̓�T�\��ab�n+K��doK��+��X]�̕g Y�j:�f*oA��
�n�j�37�|��Y�.�7�禼�ǖ�������N�DǺ�t�WO�㤌>�g����8y� �]������@D��ƑW{���N�73߾7�:��~g�7�Q�Q:k���M�Е��H^I ��,����\�A�+��2�-�o���a�	r��-��XDZa@4 S���s�#��F�++���$`pAY����b����$��i8�S˪C٢��O
�𢆆9l���HAWĈ�@�+;JǏקͅ(��K`LES��?�NBw�w�4+`8nŕ�b���di��'})[��ڙ��O�LbA��JpS6��f X
7À+s�!`H;c���pv�~0�����j�0���o]�կ�ݜ%��*u^��sm��{�9�����CM��� ɓp�=V>`���V���P!��q$S�t�8B�[�{�1��ja�Z�D�x�ɋ� �9<�Z�0"��{5�K<fE��7��o|O��1\�^�[T���m�\�K7�A_	 ���T�ƒS��*��J�&��UUU�)���j�-6%�PT��ӱ������8�b�sN�*��K̷�`���&J�!@�k��QJ�>��2[�*�%x�H��=�O[�5o�O^���{���v�
ؙH�^���3�����+����
�����wO(�\*Y��J'sf{P�_���!`P.Q�b��Х/���*�[�l�F�mV2P�/k8W��vd3F���� �
�mN��G���.�H4|���xY�ů���5F���N�~���]��X]I�K67���HfbkǬۨ�ZzN.kL�Ƨ��=���#yv��~oҞ���/�]���kxv})�&����`���STGg��J0��r�]Xbp�1ee"��^q�	�" �]��^Qd���k�֏0Y~qhɨ�BRkm�g�,i�aKh���{�Ld��ڱn|B@mcgu,�c*AR˸Cם�1'([�p�ً%A7uJ�I�����)K�\92㝩�%���? EK����[H���\�����BN�r6�K�M��(�$]�ḫ�f��bm�A���
55���IG��η�k��Q)���S�Ù&|
���w~L��`��!F@�iB3�5V˭��ݻPO��!)������c�#hk�t�2��ڝ���ܐ8�P卨�N�[�� ��x�5z���7��������>���%<�:��3��8����H�G:Y8Ԇ$�dB��Bj(���� L����
]`�ą&f�*1� '��	䜀�p*JR��W'`��q�(���,�t�R2�q�5�X�W��L���o)�	Xe�ZձNT�B৕5���������c�Yxw�U0��ak��^�gr|sUf���z35��h�h$���q�؀��!0-%4�qb���K;�.l�Z@�W�<W�?��)�hyv<u����P��bI3H�}Ot̘W_&G��L��6G�b��UQ�G������2ٻcVM�k��� ��c��'*2�@7E9N5d���._�R~;��e��j�#�mYP37��"��SO伃�T��]ng����~������И��v7^R#/����߄��!1�ۻ��[��(�A*K�P�#�����M�K�!1wfv xY^�ɡ�Z��H��g|��_�3���u�`����x�=����H�AO��&@����+�F����M2@٥-�`�!�k��G�m�9qP��+��i�e��]��֞�k�����91X|��퍍�G��� ]ֵ��]�^r����e�V���3M\��4�T�n����U�;��rjڐp볮Dqh��`s_e�T���`��N�z��rٛ�j�>�ƣA�.��Fc�vO{v�b5;c�U]��r�ΩlF���VW>��W ���>s���}��@�))v.�df��Uk]���`�i$5x��XIֹ�\�m%jBR��:��͛k�ZȁIV�.Sx���Gܲ�K������a�ݻ�	 (yE�ί�q�s�\/�\�f��-�ݏ0p�&*VdP�;���K9�X�Յ�d����F���[ ��|��w:o�}@�,y@����Va���=��`���5(٠���h!0�w�sy8�����ƞ�,����l�� n�c�,^rf�~����6���p����i����x!�B�6I�%�#H�eǘ��͠�mЕ(X�;�gI� j�e�`�%j���l�o�l�����ZQ���c�^2I4���M���R�d����n�"��Α]G���{����0��`���Ǡ�h��w����b�A0��@9O"ʚh0�^�:�uL3�P��ǧ��?0MHLB���']��g�f��t�U�T������&z!Ij�KSI����`�HP:�D�����b��6��MF E�l�|cN��l���6��J��T
�|g�Ff_�V�;��~�+�<Eu���nx̛xw���	�Z�KOt����L��_�jK��83��0�:WR��C�zVOӄ��� r9	b�F���w�kTM�d�\lr�@��	�B|��s~���%N��#jJ�%�d���v\jS�$�R�38Z�@�
`� b�+n?�j����S�����J�#f�A�/B]����?����I��}�~Ug�\�\�%�P����|Ӿ��e2�Q@}�X��-6KW6C��X$�H���jF�I��(H7��,lv��6�$f�l��Ce����!Q��XI�yC�3�s�<����'���8�	��&���ˍ�1؈�3�Ļ�i�f��A����6�Q ��%i�.���ԡz1[T�٫J,LQ�Ԅg����4�:Vk���2��I�t��;8{�.���g}�O��`�l�;$����װ"s�������XDe Q��y��`ϻx�c��c`6��V�"h�Q�bT�0��V���Ã�%�u��?�r�1Ҏw�U��2 �K۵$& L5��'�$� �<\gٰ��A�Ȅu>ȑ���:f�!��%i[b�QW�8	���' �s��4���N���EN¦���N���S4�_�Bge�N3Ɨ �Ң�ƚ���N4ӄ��k��<��M�W�|��J){@[9�	C�W��`S���ݏm��N��:�>�������Ы�E�c��n��������ٲ�:�9�qtil5N�aI:H��������SY	P��Ԋ�K�&�{jPdi�cX���6& JF*W��&��s��ԉ�Tpܙ���EՌ!�xp���~����0�!]��V����s���w��y�, ����>,i�x�	�;J�Oe�k�c���%��>��:� h/NidC���_y؜�`�9ÿ{y�����!!��L���' ��D򷦱J
lQ�2��F�Q�-�L��uC����a���m�`�&8 0&u)$ ��k%GBT��g��\(m	e�O`;22�+�U� ��kZ3e�up���g�6bA��j� ����Y�E-ع�Lɪ�FeSj} ��kT�:]����:YW��[%x�3�V�8���&
ld̺]/gզ~8��\�����y�"���dghW�أ���g�8��9��-�2�e�I��C��	e�pHN�������6*/�̐�c쓨;�VUoG�	<+�[!�T��������`<�ʜKӱWR���hJ;�pP�c�x���3T��	h�]#���ͻ-���`{�D��T�γM�ly�joV^������f�>�+d��yS�!�#�oQMDPA5�cy)qê�4!�
k�F@FF�٬��l���s��q�W� &�5oh��z���1��	�XEb�+f���1'À 8�����->��v����Ƀ&��	��5(��)��:sY�BI<y����m�.K�$�[�Aȸ������d�K��9/��mk��ee��'���]V����� 2vn�@��4Yւ��-@�YX Xr.C��PG/��# d6X��d������I}c�W�և�K����ʎ](*0�RFd7f&�:�{�4�řss���O�����g�As���ђ���-*4�	��� ���lS�,�ڒ��R[a`�
5 ���\�݋'�')11R�I"�j�� �Q������9�np�?��Cx��'���A�V��/_�8�Ƞ&���-;X�8I�yQ	Dh�& ���		z��m^�Eg@A5�`<l�����:?�52�M�����|��@�<���  y�����		�rl[�h�qhCs��U88�f~ o���@����B �����Y3��i��;ޱױ�/Q���ȎFa3^�e'�h(z��Ֆ,��j�affP���v�k�5'��"s2�\�N'z���L#�e�`�NӀ8:��XI,�d��j��
����i�ē3���}N����l4cI�!��iGZV��=���}��ܖ[^���5|�l�j�b�f�*�ϕAe*G��B
k'�,
 Ϥ3d��6��!u�"Q^I �t��԰�3z�9W2�8�Y;<�)�t�q��$�b��w3U�غh6��{{��0�����Vkdck8��b/���	npЏQ��Vp$@��K`�A����a�^V��h�PTs[
�y#2@�;O�>��xq��~���3�"�;[�9�6pv.�oE{���Sa/p���;�PMjr�g׉���5N� �,��b�$�'��@*�92=c}~������v��v��{{{��;��a������"  {f�NUt��8a`ꘙ;����T!**�Il�l��ˡ�_0�k��6>g���ʻ�Y��0,�(�%g��x	�,9G�ϼ��Pl���( (m��G h���������fh&8+�1�ֱ�u���]��_��-�"��Y�sD�:'�����N�d���P��N�o�����j�G�AAa����X�"a4�2,�L�NN6���G��~�vr����K
]����osv	�P-�G����?��j˨�^��DqsQ���4��cEK��h	ڴC�{7������� �O�^��|����g�*�=Q� ����}��r��8�k�u��:���Y�$'F4�?��/5i˲��Sc�գ��#�,��9�w���@H!BER}G^F(Lp`f����|��7o��)�6�ݐX]={�}�fgY��z���@Q�X�#�z�����B�.�8�/�1jB�b����tǤ@X����\�ז�D�a^W��RFyY+4��u�(b��pv���7�z� Xf ��,��{��4U,����'V�S�̶��k"��)Ê�ݨͬH5 (3]n�׆�u��tL�i?�n�U�kRt	�1FP����-�Oc'Vs������iPv� H�U���.�&�[��9߂�Oh��ݼ��_��
ot�A�~��gO�x?�Uw�*��0�dK�$�]P�z�c,O�C�&d�Z��o���O�ყO��g����^��>��?y��;����j�^O����q�&+dG�]���N��yc������\� ��e���C8$3M�7�����X0"���Gf�o�����^]���
޾�p�-�҇Ab+N	�j���>Ͱ��%���v)�[k�����TQ�PuSH�n9����W��s��J�c,]�rv����K) �fs3	AC&��ے�9#�|e_�:n�$���aL�����JZW�aٽ]3!|�o9�	[��ݧK�`sF�?Ԗ23�7[Ba|Ҡ	�8�e�&�uN|z�'�\�f|5u��-��O�)ȫ�G��`���{v�İ� mr�P8�:Zz���4x�S�-mÁ���+V���^^��}��'��X<�N�3)r���� Î7?C�y݉�>��{ӰEp����>|z���Ǭ�~� ��_ל���d#�{i�YJ&��ܴ��6P�QrWZۙ��!�����B�
�	i�ͭlr�֩W,N �K'��0�c�p�O�Q�?�����~���|�Z���n���6������CF ��|\�j,�`�8T�k�tuV�����:��c80�x`p�f�1uY���`��3	��jU�mè��[XB������M�ifw���RRA	w�1B�)���I��N�J��vf�q���a ㏉ �i�Na�,r�Ն��e�6�s�.�T�c�5�f1��Ķ}%ﻫ�y&�S�QZ�ڃj�y���B�;v����D��99R��O��))�eG@����q�SE�N��G�M��CM(�����t�w�&v�@Hec���l�#�;��p����2��%|����}��>���3Tu��~X̵��F��acA�YU&�+�˲,�n�	`m��wp��^�����ɩ�©[��~8摂��ƖyXZ_�D"�����<���sx�`�
���7Ȯ�ܢ�L�>d/%f|#�B@D�$�*�p�s���q��2k�(l�
�0餿q�}�x?�uj(����t��E5s�M�^_�7���e�<�K�!�j�`�$;PS���|��
L��%(̘�y��YL�Y������u��9�I���V��0\9�9ؕ�7�DYDkSp~���,�)�]�( z�,rɠ3v*a4l���/j��U�"p���y������
��s&�|��oGI�xp���� �սI��c%��: �}#�:�;����mVB��%, ӕ�nI352�#gG����3<�)2�o#�������7>��W�p�����	��%���ŽQ�ǒ00�$^�l��&
c9����Z4�7� oV=���"�B<(K����.�O��ک8Z�����m�~/6���ߟ?���n�«O�^�_��_����o��i`{��G���z�\�^��T	kf7�Dr��@b
K�p[&8����dѮj�d���J���҄wʣ]�H%��:]���l�P@�Q1X8��]C�d�p���z�9dT�Bg�)
�A�%]��4�HQa-b�Y�	 Ȝ�P�br�ڲ�ϓK�
�
R�='A�u¨��FP��l�j�U�GRî��q�'e ��c��3����F��툦�Y�C~(����<�^m9,�V(���n�b�� �2Ѧ��A����8m����И;x��W<���-\\\ �ZI/�C�X��8"�Rf�p�ȂP�}�@����'��}����f��N��qfL�]�$�;4�j\���@�K��% �rn�u�eO.]���p�j��/�*������*�'�TX��?��M�Oo:oy�mw�3��s��W��W�_"�_�ޓ�~�z�L�f�@���c�~aCK/�mc=�2��|�x�N��b�>�$F�3�'��p)�' �~jW]a�'A�[�ɞ$��KV'�@�&�-pR���t��ꪞ�TX�x��}��Ցc��b�Ōa�$(%��=����2����K޿
Gʉ��<�5]����Q�`���RT���<�2�$���ߔ�~j(��������]�@֟��3������G�\J�:�ۢ/���U5J{R����DfB윲s?���4��;��dI�$�cU[�=��*�jjCMs�'����/�)�o��� �����0 �ЄYz���̈�p73U3��"j��8DFS�Y�������ȓ����wo�Mi����Ky�����`&�^�R�����{Y�Q����}�/�/����}��ky���LF�?6s�X��|s�ŶXr�%r��|w�D�} ȃ�\05����m���{�N޽{'�߿�S�Y�N���(w��rj�����i�di��d�݄��b	�=a�@$9�^�`�2�]c�A~qۮ��L����*h�Ok�g5קƘ�x��-S��E��i�4�V��y�=e�{ee��I�
�2n���^�[;��1���[&�D����Qm�F���U��S���n��x����Fd.)6/+�����!���:���_Vj��Vf�>������J�8�vџ����h��mJ6�
ό�oLo�Fa X]}"�~#���'Y�����Ƚ��h� �V)�f�$xfp�:ӫ�9�w$���!�t"|޲R�Y�|�5ߘ�ìgo�X-B�͋�54�4M�53��*nN6 9���k[�Z�������ͧu�����]cy��_���������W_ɗ�iN�.vm�i}Lb�a����&cV �bV�P�bp֠fN�A�ޝ�{����۷o� x1����fE��[FO^��{��˞����n10sXO�+2Ȧ&��.�/��``2�{�gi������߿5��Oo���%k�4ɶ �l�Lr�@EY<A�AЁ8�NP�doj�ٙ{��)Oܓ �3���V+�T�V ���k7l"�������Z>���p,[ J�|@U�`Q�,q�:��Y��>����( ��?�!��uN%m��,A�4x¬���u�MO?������.���r��\J=љwݜF^��uh
���f�E֐�WbZ�I���W0���5&قh������u���1L��$���rT�n2�'OoX��뤼��k�G_��*�c3s��IN���g��/���~%�Q���o���YZ�����oɒ��T͜9�Gz��+ث3Ѕ�B�E	:8��W<>7��Ⴡ��=i�Dk���N�cDzu�Y���{썣\�'�ߥ����X���3�0�����&�^�m�,қW�>x�n����_}������G�O����1n&��H?Qŝy:ڦ���*�m39[���c����w�f�C��Vn�z�Y�%	,���]�O�-��x-s��٣�}El�D��sWJdl����Fc��9�u�ׄ��qG�� �A�k���sd �4�sb6E���?C�,i�UKq3���#@��	�c�37yc3$z,=�����6�;�`8k7#�9��|�����(�~R�)��Nw�]{��������`m4W9	�m����cL�I�еNV�˩���{MyqkR����կ���|��E@���bL�^����mq�P��+�'7�+�t��� �S��#Q���Ã�ۨɫ���>��*[�����,��r����g5���\gv9��ہ��B�"�I� A��
���nd�$i�{��|/�	~w��t�\�6��A�e���i��M���1+��a��V��V,iw`@.`8�&�*.��@`�Y��Z��C�B}�2���L��@�R���.;�-&I�8r������B��<"�v��9غ{�w����ߧ��Ū��ka� �=ɜ�/�+ə�2(�j7	|M;��-,++[)ۃw3�������Q��[��I�����S�C�;
c2��"5���i 8wI�
~c�'u����W{��F����h���MD�7��v�TG�d�l������V��7o�����o����|�B�~�}})w7{�,��2\�0B�Qq'������U�W�]ծ�H�Rq=�3T��A;�;��C�ҽd��E����Ԫb�W��1����Zx��8 iJ���.��e���戹��Wb���ql_��q���-U��֡�}ݩo����W�(���;���7\O�^�B��j�xw�h��7�{tAR��tn��E�/�GT� �pjV��]c&`t���G�/ (����_���i_�2�`�X�����eu��kb���t�R"����A �]��:�	~ ��r(X^�)�"�_ ��tbYf�����H���HЏ����T9�}�3�ξfH"�u��zK[d
~�	Z}��\��7&��d�|&� -�kL�4�G�͑�
�9��OHKl���'HQ�hS��ѩD!��e��Z�����0˫�f4��_��[���o����J�n�;3q3�ðkތFBXI�|37�V�2��r�y���8շ����������l���&�,ﰳvx�u�=R^0>�vr��G%>Ln2�b�`��o�\L.(���+/Fӧ��W	���A+wv �igI�Ǜ��@o�ζ�⇷��N��Q��jU�"�̗�,͛�Ԓ��Vol`�V���"�&�0q�
���MW��"��1����a7g��d}f�릲�2/=��n=1{
�]id�s� �{��Ng��8P��C>���3��WUE�e�19$G~�(��br[ j��.}�
����ʴ&v������|�?���_�^���"V_��w5)?���[\a��d�� ح���O��F�'��a�o,mDY^R_dcJ����yg�4g�@3/A�͚��i5ev�����Ս|՘�_|�|��]�SP��k�؅�o��W��E2kY�6&[�t�r��;��O��k��C3y�����}����4�k�O\	ZY_�!�:����qr��T[r3�=J��6�R�sW_]8ꧩ2oD���Ug|�c��A �	��%j`C�~5}�'��������O?����?4�b:�u~���l���͋F�b���.�a�� �%�� d@-#�E��96U�D �.�l����n�j�p�_�m3���!��濔��g����]�N��ٝ���<9ޒ��3����$ӈ�! ��\ޖs�*����# �U�I�R�#�G8~}�4�2��k�c��o����z@ ���W�,����b;����ބ�$�q��U�zŮ�n��ꢗ�-���ei pIz=*�Q3��^���'9�������W���/_�����|!_��k�O�\�ϕ<��"��e�u��2�֕��ypZ��.�V�c�gM��� �}co�1@��%<Cz��&�� @��I�CE��l]�*@Y�d���������J��+�K��~9r"�f��������bi5�/�3���@�juN�����+9Ҥp���E��|~�/�,LÔ���%����q��hs�T�]f5N���.t-eO�)h��O� g�a��7���<�37������$bH-OH��q|w*�q0Q�BsS��C�qd��}������w�u���c�̸����c@��^�f��6q���%�KVl{!;�K����qGt
#g���6����]��X�&cu�K�{[������wǽ��_��ז���W�-����������
�ؿ��?h[Y0��>MC�.e���BƷ�`h�[��] <��{�^N�7�X�.���1n/��(�2�V�e)殊��������&{�4[�����8E��	�a�a.GO<<����x����7_��������Z���ŕ��eo�:��\N?f�2=WߦX����l��̧�3�A-8]�_�j⛈�Q�Jx�q�a*��D9]�t�z �G���b!+�F���Y>/uC��1���9���>XG�Z�mW�K��.�)2�N��E����c64����^�E�(����jg�77�o����V$2?a�*$'y迤����%�r[��;n�K*���I��y/���3�Ox>��j}�4Y����~2�R-P����+�ͷ_ɗ_���������Ʋi{��-��?����2��f�i4�ҋn�w���h�]�����%>���U��:���s��|�	I��%ߘ�<��ذWHԈ�r�Ձi�5�t	z���a%���%��k�m���k{��움F�/j�+c��G��.�R���(��,(2��magTk��fg}y~q݉x>8d�#M�k�'W6(�{����b�Uv���L�"�}����RkH������c��z��?���O��ݧf<i%Ⱥ
��m"�:wK�Oйs;K!!����C����K}��G�4�4�\��%䡱ݠ��aO��b�qR�@�~Vcn朐S����ڋ�|����� �C3����(���������7����o��o,��1?�FJY��b�4Ԭ^}SaD�	G��`ĥ�S�ʾ`���RlC� �@.�Di9Ü��{~p�Vߴh��_FN���B\,U�g����^gTĔ�9&>�����v���\�"ޮ�[��y�^"���i��d��z�:��ʥzt�~h׮ͪ���V漻1_�,�IV�k]�,ww@�F��T�ȭN���`�<��D�#Q���|�d�%j5*_�W1-Hmb�gMFҹ.���'Lo �+&�=����k~��@m��?�/�����_37��m�EBb��B������d��o	��ƈnUN�`,P�0��bu?�)��L�u�v7	R�fIپ�'j?Oڄ$)���W���ʲ�
*0�3C5-Y}yGevG�kkJ��~����_c2V��S����&�.��, Ҩ�O���(0YS*�|�FQ�C2���u6��b�X ldd�a�A�	:	�h��HOys=A�E�� �$aΜD�']c��ظ9�L�����X[&)���̃~�]o�HV�;h���]┑Z��j��;y�x1����d�<i0aV?�Rv��i����d�<��pTx����«W��&p�>�$�́� +�Dd{U�_�__:u��/CoC�:���h���z�\w�=���N�_ ����a��/�
�~��L/�!�|PWm�QKܯ�}}s�H�=�x�W�|:�L��qŢp =ۅ��3n/nF��Â6�]q�*���/��M���3��Ne��h�ɽ"V���u������N~��+��f�����_}���]v��v��@�Z����^BeӖz�2IH���I��jU����iѣ�z��Ճ�{����HNf�3��'(��ST�U�n �6v�2��yf�b29(1�,@�;����(�93��7*�%�W�? H.�����o����<��vZ������N>�ڸ��5��Y�b-��Q7y�u����Q!x0��A��\���N0��7��9�K��T{@*/�c��*n��s�q��(���5�bD��I�O5�������;����,�W��S��]�'K��_%j�s�����袅���<��'�Y:4�WS]�D�WT�L}3&\���F�`wi��L�6 �A�#R1���L$���_�0m�����7��j�BٟFz����Wo���m�7*=���9:X�=y2WO�m�[k�
6`o�`�SصL^���s�'7;�C�L6K;�� {g��L��	}��}���M��s�c��r��jx�`L�c�L0�v v�Q!�=>~��9��^�.Y��s7[ؓ�/':�y��;�D4�����/\Cɥ�a�7:؅c��u��66mA�y��`�4]r\�,�ٶ{���t�5�t!�`㞁!8�u����Ǯ~�H���R���O����e}���Z�G�}����a�"�4
�a����n`��7Т��4�K����읿"� ����d�&XFw͔z���m�S���Lz�L���&�?�i]�t<b���
���j���onf���������|���;�Em�2�ZΒ0��Y������`=x���.&ṓ�~�Q4o�lg�d��:���b�#�aN!�ߛ��K�xx΀U��)t���'r��n�3�K�d�"�{b�.�3�3�6},�-�,L�d�ԆQkym��l	�%q�E�9�과hU����I&Ġ5��k��: ��������8�����|��T�}$̌�w��gst��V��x9�޷����\Dx�9양�*#\m���5.t����`
v������_ /�/�Xr��e�9�,7�K����+�j�����惲�B��8�\Y�SN��%��Ӊ�U07� �)�"v��G첲YDl�MӶ���� AW���xC��>���d�|sk�_������!�-�U��E<��}V��agm�ig8F�(/$�/0�'��2;�͕4�O�	�N_b���WB�̰�f�":ؑ%��������h�q)� �p @��B?��3�w^:門nB�ǃ}�e�$��'�1��k������F�\���f��hlj��@g$R��� 7�"�����c�a.G�"/��A�iN�mq?���'W�����U�}ч޿s{��O
"�a������u0�s��:�n|��B�����G�`,u*�(� �.���Vz��h2��@�~��ꢓN�1��Ų��J`;T{�`�	��mB�"d.[�Lv�#�k���=3��`�)RTRjW�6ߚ���0dv����Tn�;yc���s�޼0�ӦGY(���ϫ09���k�+)2/ЗU�W�:�hۙA&r0V����� �<�a!S8@��V��_ �s1��l=z�"##5%{�@�G��x��c�F��a�S6sЂ���5��G��P�������l��敊��~yg�S���5m��h�H�s�~/&�[|��:��o�����F��7C����v+��g�vp�k���G�%���xEAbxF^"Ӽ"�OM��E-<�J�i֎y˴=�|���/���+%�?�������2�l�]���iR=��(�7p��W�$&dyԴj��
�Z�aE�;{^���SC���i����&]�fcB~����&���״/��l����VL����e�	��~�u��^ր�$���?��}�������˶�^����?DK㤢��-Ђ�d$%��cJ���s1SKxF�0���l���X�P�X`	 ����&�RX"Y��������6 �d��ܪ; ѽ ���&Ox����C���xxRjH�D���������GS���/_�����g����L���(g�{1�l5�q�:aT�
���h���I�3�yQ�2����-����|�;o<�MLYv3�s0G-T-h�n�a��A�)nl��J��2�a�G�,���s���?���'��>����������S{u�T����I6J�\�N�*<P���ժ;����	{(�M����+ƨ$�K��4�̓i�o�⩳�f͝����7;u��*ғ��H�P��}|9�m���5u��ҙ���뗷�g���=��SY ���G})[`�ZٟV�h��
��FS]��WU�K(��3o���V�_�J��f�Ä�.��*C��"��M^3�������� �Uaz�!�ۂ\���{C]4"�z	[*R���Ψ~�^���/on���k�(T0Tu�z�vT�H#i�[*L�pu�FU��`�j��u�Mܔ�3}T�?l��x/ ��;��frAvҙx��I��S��O��Rh!Lnb5�İ�* -#|��B���<�Ow|4 $�{�������e�o/�7�����$n5�W�'�����'1_����b�&bz4TaS�%�uh^���M�
�mN=��*0��4k�J���i�4�uZ��Q����Gg��i
�g ��eWk�Y�/�X���p��WY���*:�؆F|�y�~rY+cZ�r�9d�G�dĿGT������j�7y#�b�F<������P�qɌ:c2;� ��<3�: ��Ϛ�������$6s�H��H�V�E�ڌ@�םQ���p��ayM^��б�!�"J^�Ɏ�7�t���Ъ8�C���`�6g_ޟL�V��V:��k^�Y	���j������8v'�� n�X�����uG�{I6���,�iBpS$�e� ��0k���%�Fx�D ��R�"QJ/��|��������Úu����O˷?�����e�7�^�i�k�l�f4Z�QV�C��s��LA#�Jӛ	��Q��[�7o�:��݌���Ń�Qe��Z]�3�2���N
�M��3;��hb+CO3��֔�
A�Ŕ������<y)�Fy߼z!�^z���������R	����g�yU`��ї���j.r��'k��9�(F�/���'颥X��83�߼��Ǵ��1�zs��=)��늤[
��I�o�;�ef"���^�ן�cls� b�(��)u���Ӡ���/�6��������N~h�����bj>���掖����@���ɥpX�^CG�l0'ҘW�%L#��I����iIB_6�Ybh)V�)�y���u��a��ֵ�ϵMN���c��[L��O��'���*�\�����73O�����������ߖ�~���{�� ��M���?(�K���Y"�2b���Z<��S_�r"��Ldg@���4ʚ^�AVZ���}l2 ꦋ&�MM}H^�f����A��#S\��LS��]֜�^	�&� Xd���\|��9�_�L�e������!عV���-G�'L�H���+��8M�2e��ö�Ì��p����c�4a1G=0�q����T���Y��2��E:pPF��Q崭����}�3��2�ѽ	�0]ʧ����-�/�s�Lx��?��wN�p~4U������5SR?�]U>�AOƸ�5(qNa�c���Y _�W���Hj`f�ӿLU�v�n���� �&l[s�{���M��w��.k�]Ɓ�%|8���0#�}~�^�t��h򉏏��������C>�n���Ë������p�������������/�K�5��C�R�EJ@ _Kٖ��)�c-'"��S_}�uP_��e�ӟ����
M��a'S�^۱�7.�.�d+ �*0))��C5GM�������{�b�?ۈ��)��UR5�$�詬�/�Y�aW�%z�� &+��yGL�e�4���$
��y����iك"iA6L���`/)�n+*: � ���t��"��侀��5�_n|�������Q��.S� �}�;�����l���,��)�{�Vު9�pi��g�C5=��z���[�蝎k�u�4e#�:�{	w ��\�u�x�`�������������,�Z���!�P�a#&�>Z|ƽ�FC��IJ�rA���M-N�s���w���O����t�p�����o���?�������o�r��4<h�3�=���<DmQ���^=*V���f+o4r����&��}�������ie���1AM^���� ��wre��Y�	L���O��s�/P����Kz���m3�^�ʛ7�R�~���ؑЅb��p�ؕs��`��)|]�lA� +���`�j*37gNlق rM����ɋM*����{�z�[4��<�~��K���}����o\�5�s��k6��M�栢�w��������\�O柔y�H��pwX���*2$^3|��g0����*!��F�`�rN_���ǎ�
��8����n߇�[�z(X�H��k��H�!��)�ml#jfi:����,�'���?}������ֻ���o߿{�����L���2SҜ�N([h@�yL#�(���s3`Bg0��
����3�b��7������
sV(�٥MD��n�J�� �����~�I���䨽V�B&Y�Z>���o��=���ݭ���i���Re���G�>�j�Z3�O�6#�P�B�+X$(E�!�> an*��e����U8r���POH����Z7���٥�i��`q�w[FYɊ6G?����lK$X��G�},p��6Wqwc�o?<�	��ѧ6,_�� hLp6pH}��7� ��8�=�1����>aZA� H��9%���B6߶w`���쬑� �/�5�_��U@sXUd���a�!�H�0o����Fi�m˟uW�_��<�O��������������||�*JU�oc��Y�1�U��3�1X��K/W����$b���^�����	a��H�{������'���Q �f��3�1�l#��
��mS٘�t���t��ǃ|�>@�X���Q��ôJ��&��&x`��h5s��7���0�͌f�KDQ)�}�6��.�P�7�T����ڏk���S��� �=��;��x��)�ϕ����Nq]-�t�z�S+΄�5�j�z)_�y�p�?Y�E��gw��F8_L�̈́o󄹛�:�dj ���F.��zD{������Z0@��XNe��X�C�Y�����0�̓m�-%l?e;69뿬�e���ÞP!4u������
!�l�Ow| �����7�w���>�����F��ڭ�5p��4+U�Ǜj ��?�Ѫ��/�1|!�Y�	� �:,=�x���yqgb*�/��7"�)�
�� _����+1T9d��*�6�v�T^&7�UA�?��]�Y��J����k<$<�����gҒ��MQ$��uP�a �8���td���kBy�Od�%T�ӫ�{-� �Y��@+D��i�����)n��]�ݕ���~�9�7UF��N�l�Z�>J~uQ�Hȱ���*�u{{����-�PŻg�?}/��ŪC�r6׍6_r�?㹭�0ԓ�]�m���>HO��W���\�_�W�ɡ�8%�j�a�D�NJ�w@�@��H����.Z����	������ֲV���8���4 ��Kc���)�q"�۩-�|���R��|��E�0�J�K��l�
�vKt��<�������e���c�e�"��?,���rk���eyu��:�˸��@�%�V�MTk�3Q%�����s�& TYN�ڢ��4j�aw3��р�fo��e£&D���6B*^�x.��s�	�{�������G�F
�T�ξQf�4 j��Z� Ml��t�g=~��� ��]��<y����N#^q��V�{~�]W�(Ev��qP)}��� �F~|� ߽}�@�1H����U����6Ŋ�W��*����B 䙧��(s�M�X^	�}�(����iBb8X��wE,�A1$��6��l[��)��<�,PJ�։��'mC������A[T쫪�Xe�wm���d��d����[���툗49�:�݁U�ki��"�3�c�L�M4���FB�"��y�B�������J}�b5���7�[�4�kTz��~8��U!�"�j�2CuC���ĘIT�	��X�Jvݶzs{#o����O�d��\��*d0�S�>���]��mU+�N)X$߀�GԐ�ZkD�G����m�� Ҭ�{
�# �??9�H�Ӗ�m��9{�$�k�\��%���I�XX�Pԙ��jms/�{qs�/�9���wr�ǃ��4�(���|s��#�$]�7w0�\R L܄�� ����ʒ��JFh�_}���
��O�\?���O��.0����x�3�Y1�J��w�	{�}j*�ڜ�,�����Ī��$��������X߾.�rn0�?�i>[+�<%7�\`����8Ӥ�!����,!��C���y�,o&]�F����{�xX=�� �Ӡ����C�Y�N]|��<+�.[�5yc�}�ޥx�r~���v�W����Ec79jε-��e��U�����&�D ~u��td�����$~��N6!#-��<:x��.�D&8�b��<��=0q�c�aD����"�4|�)�ȟ]o�F[�)�\I����+��㠵�/n,�SS�T�{�hC��:�-bi�� j,dc�Sc*�2�
�hK�ŀeu���1%��
@*���������h|�zi��y ����D�yS ���}�T�Tn�"ȃ5��'m֥�uӌ�R�I�%��q����G�W_��c�[�:��~YX���~;�zH�KY�J�Rٝ~!UF��T��A�4���(�P�dm��ׄ�6��-��� �L�>���/��d
|7�I���v��Պ�CSa�N^�1?��{w�k�i_79t:jt43
��������>F򺯌��w9�����}9��~�}g#oS^ 3�-oA�ߢ��Fן�w9޸x����QE6s��붩0�XYg<D�'D��Q{�>��Rr�@3�_*���rj�o���V�� �+t]����	.a�V��{g�.B3�H�M�/=LAD��3��j��px7	��a�H�0�+jɱ�jR�Üj����T!L���t#H(�j�����=���ٱ��8��2@�OB�J��u'�L&�,�Y��1��A����t�9�4N)@���Be}��:�����t�Nh�LN��q%\иGϩ2GeC� <���~�f�S�)���~��"�H�}�ƫ>n�����6q�F��K��ڛM�����ޟ�煕��p�E0j�g��)�u $�c������m���Cs�^=F0�l��������}��)B��/z0eO�^�f܇�� ���{��1_�~!߿���*�И䢕!�G��[����:�����LZ]�O����/=_���^�>��\���9���=�k	2�+!ր� ����y|�R�5'���(�LϺ�K]����k�����t��c�
���փAK��ׁ�΍q1ӷgi!Hv���?�rH>�R"͢	�2; V��D��D\��U?du7u�����������N�UK�*��Nn����-�7/o��a���eAS�q׭1}M�T�࿍�ؗ��6Kd���Gv8,&q�t!����L���`��_�H�u�����9�U-�O�c�^���T�B�&t�'��:x>}����)�TA���r�O�?E7#m��b	�[��7�������r��ƫ "�y���E~+����
�gdxn�T�����#'·��:�C�������e#����mG-�d���)�gF�Xu6kB���<����^ͬ�������c�mdn���֮��(�=���������&K)jv]󸛇Ɯ�Q�k5�mGzI'p��>C.?j/695Mf1�U��f:k����X
�¶�8/6�M��t�����s����F}߼�ۗw2�<Ȣ�hM�Qw @� �K��e.�/X1�ˬU��#S�m�5���S7�]�̥���h�^o Lp�&���?d kkv>��v6Gߟ�wf?E�����ٲ�k���c�f�	D)*،]@�:���=��z�*��/oo�ׯ�Oo>�?|���x� g��Z���u�	�l�;��ڌ��t%�����Qs���\�f4yʗ��5��� %�1�S�!|�����3����cl���Z{kV�\�П)��73�����:b�m�KR���~�eW{�J���7t�G��� �Sܔ2&4�E��.�L�QD��#pH��EL�]2ڎ� 8'��iD9i�u~'_0^<Y�ܘ�A��/n������4��͆���셞�@�>���a\
v魙)�}LΤ0�<=��2�}L"�B{ahW��=�{A�-Ӣ�>�Ӱ�F��=�㏕!,������?%��q��d%��uixI�����s�{a]�S�T�S���ɘ�V���mc�o^��/~|o�	�<��Z_��l�VR黵�
Qr%6�����ƕY7�6Y����%��P?Ha��ǳ=�o5X6'ΰ��8lo" ��膲�o-pMq#|�C�JH|����-̟i-p;��.M_�Tm̓�.��?�˒.K�f��2�f���%�f b0���{JX�>�RBg�� ���B���F���;m��ny��n�� N*�B�m�]/Z&�~_/�wg+�S��|(2�o�Ý6m߇i�9�}�	Dd��	@�+Bpm�QVn}�G�RbƲ7�N��&������k�E{:����1���dh&�"a";�
o�<�����l��yu ,H>�g�j^��>>6�7���nE=l�7���h�����ct��yj�jCu��������.ؘWԡ�5�W�W�!:�M��}����WŰ��c�m�A@�R����]����<激�'
9�^�X$��4C_��͝	�;D���;�u*%�������W����,i}�O�:�lpx��5+1���u����%��M�D�H�*a/�����.uK�t4u�Ҩ�3�%�&FP�^�p\;��-JBSzm[rl��Q���_6�ˊr-���TG�`��-�!{2�#PT���W�y�����Y{���dm"5M�F2� ��Z��� ����x�?M��	��ֿ92w���V���͌���Z��̏ ��/~/��f!�e�>kfJ�ԇ�&�,��܇h�P(�̵�� ���F�2`�'(5O�Λ2ci�	7�*��{���9�q�z�H��ܝ���5��`d�3��ˠSh\A1��[���l�z볔�'/�8 �������"o�������{��R�� �e A�S��#�I��	15~��x����&0?�C�Q|Gӻ��).P����u]!eTab���*�a<�Y�nd*�8Dn_6vp�B����zd�N{G5�h
W�ZR`���T�Pe��C�D���<��ߋ�ASX0]�	��}[�d|��냙�K;?��"[JX��P�w�5�*�M*̶��<�\}����e݀W�cs�-�U����D}���'?����6
���N;��vɢ�$i�Y�B]���E��ޟ��.54 y�5��G���{Q���&X�+es�]����<}A�~�G��%�����L����-,����C&��L a��O�:�)�T��al��\P�?���wo���	0�7=-��!(���Y�5�E)�P����H7��7�N�]"��V�L�m�0yQ��Ia�[1킬��x4���f��1Y������xN�×��L�u�� ��S��C��&�c�&�{��W��n���z<��h��{�p�����Mu�������>�Y��o���4 ����:�� J:���1n ���@kq�	U S^;s�y�:�2�U�޷�Ƕ�d��Ȍ�p=D�Mܣ<m &����S듺ҧ���r��M�������㏅Q�*���Q��י�������U`���d7�ƴP�&bY��:�����?>j�=�	�`��f���Bxr��`��߲��7��◱�I�p�J�����"<t-4��m��R� 7n��Xf�I<U�n�;���Rnnn����5f�Y!���0���O�h~q�M�� َV��<�Z�&��DO�3�_���Xݐ"bwQ�Ͷ���# j�p:ǯR;�E*(�S�{.�p�������ƒS�lL_5� �~Y�~��"����*�c����P�1�vw'��5�>��ڽ\�,K͑��TI�0�G�lJ�}���7Y�y4i�{ΒB\!=��)0�k,�ę?`�@���tU����9�K�Lu�S��j3�Z^�sn��c?|��(v���Y���'�i�핫�(W�`����emv��Xi" A��n` ��15yNUBҬSq�5�&�I����j����쵑�no��Yu���pk��Y�>ի�9�#\?{;�Z��B�~���� ���ź�) X��BY�.*1����� S��	�=��̑9��~��Ǚ�oW�������-=o��-%@�����&���@ �������FO���=Wg�`�	,O74c��~�v�J�1aV���y�;�����la���e`p�Y
wG���8)��E�|f�0ixf�9����	@L�﹡�fM)vS�[�&�68M��	���ɇ(����5���ھ�1��>����UU:��x봹��z�Ny|WL�������iBU�Mn"i-侙D��M[7��X��������������� 3J�X���7O^cIy+�������,�=�W�}�v09��������_���(u�kf9�N�C�� %�Os�j�R:�b��lg���M��{�3����k��[��V����Wc�݈�g��/v�|���V��g��ӝ6���Ȉ;�m&pcz�w�zr�f����>�VZ&�V��'��a]�P��J ���3�^Y0L�K���I������M>fu�}�����(�����G4���u�Y��e�3���Գ-y���U�k6���x�5n���6���P��9E� hÉF�_V�bϯCg$���m�����x< ��l��5�����1@m���`L�E�� L�:�uSh�$&y���Wu�}��ې$�q}&�Z�Z.s4D�8{"6и������ �쁙������.^�C��g���L����+�Ǌ�o}+ͅ����{
��Z�6�ws������0��j���=�BFX�.�IAQ���K+�Tɤ��,N �*@��t�ţ�}c�﯏t��Í �t]/��O���e$!�Zr#X�膴�r������ �};�|!���'7����3L;��b(j�7W�%�H�>�#.(_�ݷ%�i�T&�k����^�dӉ蹃�%<��Nk����b��n
�"����y���k42y�8�F�U��@����-K�XFf$뇁�G����9e����k�Q񹛺|M�R_����x��n���~�6�,���=��^���*0|�(_SL�C��mR��F}����z�8�q�����s�Ho&�#Wwi����啣)�~
��b!\�SJ�B@��J�íe��IÒ�K�����Y�o�i���5Y�d*�4=�H��� �w����E�\��T���.�q�����	��{�~�E×�{����9����F�AZ_JO�+��{���_\LoN�C��(}����xR�X���Rc�M0y]z�b��؎��P�3Mk�m�cHE {U~k�����\����_Z�_L�r�ӌ��\@�'ϕ��G�L�C��e��z�+Y��Q���>�I��3u���P�2#����W�g�s�l	�E8��j.?�����7�����Xį�����kx۸+��{�/��"��=T	�n�it�9}�A���c�Ok���w�s^�S�������Ž��d,�g��.7(НÛWya,�S�"��9�:����K5�L��V�1�w�Pf�zt$o$C�������@�.jg�=7�H挓@H�k�lRg�Qy3�	s�z@����쫏b"�c��фv�Y������:+u_�v�msfM�>�%*q����9���_H��~Tl�q0y9��	F����T�Ԙ����z�y�祽����5���9��1^Z���49����)#�Tl����69,M���h~��P���!�n/k=e+���ӆ�/�-�5��L�{:~�k<���>?��K̗��#�F�.�Xg(
Xj�(���G{���<�C�M��3��.3&,�Ls�O������M��i���R�	�O�� ̏��?7��&�?3��>͹ۦ���{h���W��z�����ψ��Sj��cڑ=P�
0�5��ի�cy�����9�	c��Ά�& �f�_kZ>��asI�9�`�t�gT�|��������5��_�S���?����Hߴ�L��.ڔ4�g���7�!��'��#��j8y�;�>�g��3B\�7��3���]��lEp��lĞ���L��Ԧw��DpU_<��'^�O�|����&J`?�����9�_U0�- ��I(������>�=��
�_����E؁��LSyV�\�u��t�˟�a=e ;�Q\�}cҷu @fX�w�b�~S"	�EJ�D��U�q�_�2�V���U��!"�E��b4|M���k&�#���)��������Wbu��
��EË��+����+ֶ.���fUC6�>s9,=�6�ZV����,�vc��:c�=_�����]�����~b��h��nH+�&���3��A��$L_������a���櫽�,޼ۇ�J	s�hn�!d�Ϟ�M��ܸa<B��x2VW����=1��A��]�'J��\���~�̇���ٕ0,��>�k���<	�#�zۯ�;dkLH)h%?��ٛ�p��Y��[8�{J��k��<X���A�]b��C�ol#�~q�T�m�G�}�����|�n�Ļ$e�IuVX1�*�6ޛ���q�՛*�i�)�z����Ap����O���꾘N5�D�s�F{q�@d��L��]p6	J�n|��/�������`�ZRgqr,󡭡z5�Tc)�g�WV
�xk��(	�E*����q"y�D���`�X>`f:H7ݟfI�����x�p�U8�p��7)�0t�J���M ڽ�K6���@����4�:`;��bۋ:�ʯ��*q<_��m�c~�U��nD@����[j����s'Ժ��uf>�m!�\(��骈�tH��+7	I��s7�	~|A�M�8�ޡƪI�y�¹�>F���@P�HNR������t@�x�r�O}�"p]�\K�5��!~;���q=��zm�}���n&<K���b�|��װ��A��K�8��9 ��[�ҴZ�t��	]>��v�4Gl�Ӊት^잭�J�D��
��'s���x���_=�����>��L=zD�2��W����L8E���Y��U�U B������0�HЬ�e���O )ݿ7��� |@H`��K�_ �&��~���{k�d3�T��؀�s���zvBu����t����q?�).)���;��>�1с'ano7�*�GS8�T� ��<q���kj������� V�]���y�����B�ns�����x `t����|}c��۰~����s��@��P����ݓ,��rH���{yT[�.ʜ����������-�ٺeY�/��ѳ$!⨌q�������~j����ӷy��{�M��=C�ǈi�.k�9����������d�>vq'F���a� �Z+�U�p�k`B�6L�>RJ0�-�[�������������y���*{���r��x?M�&��J�!*�fnx�x D�ˆ�2��^u�iS4�%����w��K�NF�;f7(����Ϩtɳ��r��l��xn�S�㮇K����OF�ʾ�4�_��؟��(��$�Γ#H����kc?eOnܶ
�Z��0�H��d
o&2���l��G�&���i��$٘��HUjQ+{�:��ԯt��?����⸌{F�$mY�����qb�@>F"YYb��ً+d$�J�bm"�H�����1�7@p m�`�,���a|������nB�����c�cd}|�k��Z7�vy�� �~���W$�#z�$A;p^l��H��P�����"��?�����4&�Ǧ�]�ȏ9Ai�4�}iȉcï�(UF&=�%��S��p��IL�9����	�}��پ����������}���0?L��4/���ZwUM`���߬a'�v7����ן��`������3Xt8^�qCfe��{g˷>��lm4�	㍔ڂ�s��d=�z���W�s�\0��%�K�5??u�C�z��4Ь�R��ո�
��Ο�(�{���=r���\��i���	�����)����zK���)��6lNv�
ٮ�i������=N���1���V% �K��v�_6943��Մ'0-s�T@�ȋ̃��+5*z�0����v��?wn.��Ҝ���D@�-TK��b�x�0�j��#�<s$��b�K$��n��x��+F�%�Nym�l��E>��q �w�����ߥi-��rZ�m�*�>(��9x�&ƀMԍ�G�\Wl����_����03�AP�joJ�����$~v-L��g�����d����9Uv�M�ś+90�b�d��I$U��YN� Q�X�,&v��3|�1u+�/	���ɷ�Jݾԧ�h*G�8�	9���w�w��2%�B4|�5��9� |���0�/� ��XB�:E�����A� @����<�@u ����dd�.��Zt��_�G~/��M�̯�آW�s�Y�C����N���Y��G�R�~��z�*X�0O�WK���@��P�����~6��q����5 ǭu��\�bb��#3ܛ�ּ�S�,�g���O�����$]�2U���E=�y4	EQǹQ��,[ǟ�e���s�`ӳߣ�suh"hV�)g�AUgkx��.k� ��ۥ�|TZ/��I��"���]�o�����ʅ(*��ꍣ==l�{#dS����	��H�х�� pU��{�p��~>=]��
}��n��Ȱpk�~n?U2@��5�_���h\��T!�7�����m0{ze��X����RY;St_,��]"��b�*?��3P]= ���X���l�2�3uf0!�d����^�+2�"�Yi���b��aP��֧^����+"��$���ܾk&?<�UC��Ֆ��$���R����}{����~��״4�S���ts�nԡ��n�@�������T0�뀔�j Xݙ��0Q��A��DW3_s��gؿL��7;��Y�'m��*�
�!+�M�T��p��H6�>F��=�@� \u������N 㽩�� ������'j8�zd�k,%��r|��6�s|~$i��㥽/���g|���^��5m����`z���R�҃O%f�66R��xb2e�W���s������#�xZ�b
��L�������g�o���V ���/h9�;�:���g�F�����ϰ�O��N&����<�{�@ޖd~؍�@s̸�ǰ�Ʒ\��r����:>Z��ۿˏ%�.kn&ȮM������Fۀ���5ę�.����@��fu3T�-��4`���܇㉮A�k1�v@[0L���X׭b~��>G�`d�>Q�=$�ĥT$Қ�HO�J-L��a�"9I�oq"8��;����o7_��af���S=���t��?�'��S.2�\[��#���9��׸� أ��&w���w��6U��͏R�`~u`����*0��m�
��f5�蓜O��ۯ��WࢷwP��Wd5���t/�T䌺&��e��!�uih����(�s
��M�7�:L�Xs��j���Q�y�����;�'ø���:�ZR����5�Q����e]�U������4<�d��_7��Fx N]�m�T ��JƃI��9���S���Y��E�3�7�RS�9�r�eI&������z	[2Y�t�+�K�h隭�Λ!�-TIh
y���ƙ߄Ɋ�I�n�"�6c�w��[�ʌ� �����O��>���)D�r`'��q��`�Ε]�Ǯ�����[]  յ_��ї)܄<A�����xioq�r��K9޼��q�@�i�]���
�zVw�Xd[�,*��X��@O������� ��y�f��AO�qqބM=#�K�]R_B��n�K��uv�����>�x����T��l2zt3�
D�I�O}|�D�v��xj�Y�����Ԇj|b��F�LD������� 5?����$�L���M�H'��ь��`fG�=q��hqd.�f7k��N��~AJ������,��>�kd��Ɓ�2.\7W�8*,�aS;�*1vi2��M���B��'��4���cx/��N�~3����e�M%��#�3&H�[�^� �},�M���3�[Mߓ�@픷 f����m0��
S��L�Ϳ���D,a@�a[�b���+��A��u{M66��M�4	��3$�N�v�}�ӧ���:� TVQ�+�����������;0B�j0��?s��x�G��rn&p��k0$;Ӧ�ő��㈯���W4��W,2��C^uµIk�X�i������u�S?�����<�A�B��1��d�������5x�	S>1_TvY}qkr�m0ћ��;F�hn�����R��1T���H4����<�b=�!�����e�����|d������\��=�C��!�h��+�L��G C�w��B#ܰ���]�/Z�YTb��ţ��D@��Q�QPE���*�� @w����Z� `�D%}S.`��-�7j��	���Y�d���9����ǔ,K5�`q�y��x���������^�{mL{�JN�l�7�_�	=�_��� ��J��f���5�ォe�M%��`�q��h��ndę�& �+hM�?o��@h 8~�0A�0*"��a%�O�b��^���J�{�	m|���nt����b'VTth�&z ���R��~;ۉ�5di$"�G+=Ȥ���j��Q՟9�2�=�4DR�Mg�E�l�z>?������uc42�fm/��o��tY+=Vk��?/P�h�|��*O��&�o:�����L�㼳h��a�#f֮�6��f���B.nl��&��,`�FD:u��HpN�V=��е5?�}� ˺�y��F��9X@���\b�`V%L�͝L|&��H��,�7|�I��|�F[���h ��O9��FvJn�����.c*
���J��qsƁ�ݺ�K�X@�LTw�a�0�~~f�f�Vٛ�Y�zz���>YL�dWc~�fϮ0�KF�p��~�k���An4�x�Vb¨��:�b��84~�ʀ�3�Ծ�`P�y��*��q,� �63n7�l?25#�=%�ϒ�� �[�$r�Δ� ���я��������ۏh� �ڕ�{B�@������/#�̍s���3QM�4�����]��� /_����[kpe�mX�K�M���������8�c|\�J�R�!ǜ)��	s�&�6�?���	�g h��Ԣ�K9,�c��Z����m{��u8���n)W�a}>9jp���~�6�քL���i� �i��G����m��͐1T�W�Ķ���I����@�9lj5T�����-ɰ��2��#Q�=9��o�?��Wc�<��ϳ
�Մv������`s�kױ��Q���iے��NI�o��X�hfH�,؟��	�AY�rJ�@c `B������d>�l[y߬��׹i������������$�s����6r��gӥp�0(�s�RG6��{ �?kK̓�����J�~gp�ep�Q^޽h �M��v>��ri�}j����mr��4���!E�21ـ~H u�FxiAB�A�����r�-q�z-���v�bW����%�ƻQc�Ɵ�9?Zl� 8�M�k<���H�'=>��^�/V��e���-C����1���2,i�v+� 9�>��i|�@�
Y��'&�l���4�pUT��H��YЯmr�Y��6����Y�=�P9�\�o7��{�k�y�DOǤ�f_�Q��>���� �`�끈+ '��ǈjE��"�9U[8R��j�t�����2	w�g�`o��xe����8W���L>�Aq�*��z
�dl	�u�h�/C�^�ߓ����G�K7*�"m~�@�������^n�r�@07�uV2�؟n��w��xl`�A�����^s\�Z���ȫ E�t �{�q�������
��	V�n����v!�_7#���{� yk��v��M���#r���"�g]Fg˧9> >~Y����P/�z(��i��u���`�'�#��t��5�H�ջ�w�Vt�E�&���/@d4r�dx��%�`[�V�bcKc']T���AX�9��~�=��	�777&��X% J?e ԃ��n����xr�(���{k���d(_a��`)��D0���Nr�,:��,�>T��EF��U|��UD�=%h�Ly�u2�R���\�K�{U��c$H��{1��MF����M�U�o����j���7��vt���c�����$� j׸��X����]��V�9�g����Mb�L@���~�}�$��tm�4Mg�M����(rA�#l�!Q��58�%_�焧����L�\��U��"��m�{�˒<5�����K������|V� $���1�R_ǜ��w@�ax7��jP�ͥ��  v�"��T�!>MH^�(,�ţU��SE >43��=fW]U��Z՗tssg�whg�Hu?�~�Ҝ
&!�3��<E�8�d�q@�
T� �Y�/'����Ou�-l��������P9���Q�ˮ�!�~&��
R�=�*"*�c�}��ulx��kc�j-z(02!zl����7+=�eu���Z߫��K�n
|v9�_��̹8����^��y8k*T�;�К���-��2_��ߤ>���ۗ�B_p�^�py�q�:��oZTCEhH����-xu����%�p��k��EDc�"kp�,�i��~'���Է��=)�"��o�d�Q�Ɛ��i�|`���5P�q�o��ޒ��s�3��\�^sSLG�����z�Ǆ|5@(P͍ݭ�x�H��� �/ma,���Bp���"׀����v�T�3�I��^��G%%��L��K�W/ �4
��2y�b����$R:jh�E_+,|�͚�)%�5�s����x]�A��5i0����n�cc��㍱d�s�x����s����T�T�L�L)V���Cxfh����M�VAU��$�$���+ ��u���Nǫ�{����Lߓ�{� ��{e^Y���F�tl��	��f5X�f��y�a��Q�������ԯ%XX��V<�s0���u��ٖd�;��*_� �������ں����A���A.�Bª��u�ۆ�>��}��%�/�,s�}��� ?y�,��R@%M��xd��_�n7@w<��,�G4�a$�N��< z�k�n8�V5b.&��pQ <������'9������OE5�7E(��Z�^��Z��1��C)dzl��A�{@�)�@�v�e��:7�t�,��$�.��æC�K~_��Y_�����]O�O�TͨGVF� �A��U��uuS�מs7�ս��0!���'��E'���6O��_9#�k���d9v�kxѲo5��.��ml߿���~x+?�{���"��R��/d�}��� �T�բiyVF|��~p6����A�MMxo�] �����x���]b�4�:��>�y�ܭv�tI��;�9>\h�-T���2M�٩�:j��].�k&� �m{|/���.D��p#à���;��a�T=n^��*7��d-��,�C�p��G!P[0�GPG:�73R�Ӊj��.�<��(���V̻�E޷�}c�wmn޴�+��TK[Q�E�
4s� �qR{JA,6�p�
��5øqd�hb�L��[�\"Y���5ìvs�K������7�?_�&�)?5g-��{8,1�{���ᾥ`�c���ɔ��%.h`�=��p��Pr!|3�ٙ�u�ԝ�xq�ߏ�?���g���\���������Vj9i B��X�t��8.M�^��*��*�/�畳���DN$U0�'80k�(U(���x���CJ�X���u��)���� ��1��͹%��Om�6�J������ߊ������K���'B�BmY$&m�.��dv6��N e�5Ӧ}���\��&�2�%�뛨�ՑC� >�`H�\�ü�I�mKðZ'����-���)�73X���"�-4��M) b�_����PÖ��N� ���c4;�NX�݂�;��f�C=fB�@/�Q�� hA��K���\��*�^t�>��	M0� ������n�O}~�e=T�83�co��E��9�y{#�kʁ���V��dck9*k@�Z�C�[�66����o6��i X�uP�d�Y�(�ߛ�¡��n�eq�db���i0�SQ]uCh��D=�n\X�>���|$}K҆�WE	gB��e1I��m�dzB�h�� �$��cc��c�y��SIbil�j1���㣧��lC>��_PEƶ~1YG� Su�]R�	ǖ�����@+���d� 8[`��BF�~��, �?����!�r}��Z�E��������45fM� Yti��q�R�ĪU<R��8�@�І�;<bz�v,'�)k���qU �����,�S����dPb�]����r�tdbo4[�P�U�ws< *�ӆQ4�ח2R9|���3��;�a~p�`#
�aX�K�(8�yBB���E���5٣�/�\�><Vu��uc< ���l��U�m6 T�d�	 �)�V�2\N�N����ִ �?XY�sw�dͩQ!Sw܈�[=֩��=,6�v��� ?���@X�r$�h3�u��UQ� -/��ڳ��|�x�Vl��4^k1���ޥK ���2ŗuH+��b��,���p��-����=7�j���I�"�D͞S<�= ���\���v3�����󪴢ĮaJa��Qڐ(zn�G�D������� "  �͕��7~�J%�2��Sj$�J��xޣ詗�)�3 l�g hp[g���`��lO���ϧ���*џ��1|MuQ�DAµ�<�\ӯj�<��oߙ	�R�<-�������f����=�˞��ep�G��֐�J�(���5 ��dݐ��ʨ A	��<^+6�I#���m$��`�Tف��h*�:�E�%����-�뇈@�ִ����������^���5S�6�?��s�����0��O�N��F�J�������M��&_��Β.D�X�V�M� �}�$)`zl�i���p�Z*�F�6ɔ�+[P3X�b���_�V5�*"��(�]7��9��c�捜�g�����UȈ�i���t���������V Y�	&d ?���-b�j a((�i<l<t��E~�~�1�*<^W�(z8'��"uX�8��B���?G0)��W���	.^d����	|���?�w��4#`ok;��|3���e��Q�_h�d�v/W�$� �Ec*���o^�j�n��B�+�.0�--�k ؀�m$�v����'��AL��(�̬4NB���y��B�c�j�cJ�b-y��<P5�o��-�����s֪��r��d�Ɛ�E<,�}N�͟�z�˪CV~�fF1����?�0��R0�IbfQ�l��BA��:�9L�.�/U�=\ڂy�n�F[_��L_��l�F�-��pc�g��������Y�0���nLg��Iҽf6#r��Զ��d=�C�.�W�d:Dg7�Ez=���:��ߙ��-؝��J)�z�)چ�����S�AS�9�h3��MB2��� Mb^�ޗs����������o�[`�}Ӏf/'I��,P�����|�N��Ǉl|�A�i�~)�q�Y�ͱɳ�4UK�W��d�|?���_p�>���a��K��#ii����Z��\��~�������eN�A���xB���<���������I ��1�!��bb�o��o�64}�M��O5Ln��P�P���>�Q]�� �|h��[��7 �+��o/=����i����NJ���YS��g��VK��.��_W����Y�F�۰@g���/�X��_ӿ7�I߻z�W z�&���+]�!V����o � ��u�g3�8[H�
^�VZ�u�?�{/?����7e�G��X1�Fը�|h浪,�����p�V���c�)bv�P�1�B)N����}}L2��H�r*@�@w�to�O������`��Yk��*����un{C����G�~#��?5�WyG�v+�j�#�ؘr�&ːm��^�z+�^�.>g��00;�$��q�э��$��n����+�GM����U[�ZdM��{8�����N��Z{:YB��_�TJ>鵞��i�s�ϱ���� ��w��0���I�R�	�Q��`�D��Z��>$hO0�w.R�\��7(?C].��@$�@-���T�ϱ�E]q�K0��7�w��'�'���<Rs��t�w�W�{��v�K����*��XB�d�0磦"@���ԃe��I����Q-�`��C�<� ��8���A`��Oh��<b~���q����󶾭�,'��L��<l�1���3�����v�FvUF��7��N��c����ōl���`:�%��$��,�`7�H��`��#�vC~J`��?S#��2��2�r�X Ē�gyq3ɫe�����5�"BY�^���,�W��g m������1�E����Ɏ,ٖ��13����f��X�q"�x	�Y�iZ_PR��A?���|���H
*��'>�5�y���������9f��݌ȸ̲L�፵�Yg�}eK��Z�:�]mZ)��𰼈H�p�`��'t��6}��n�ɉP�ůk�OTa]\��k��@ì-�.����(I.�o���nv{-��
�ey��,<����4GJ1%E(��\On";mRi$2�����1��^ɇe3~c��_��T��}`�χTK5����.,��r��S�-0�w���S@ݬ�8H������$lfQ08c�`�$�
��`�.\_�i�b��a'�Ivs�	R����Z����P���|��⳻��ma��;���|(,p+ H�VXҤ!JU�Q1�<ʃ�:$W6�DK�i���:�/lA�Ɵ�9�e���w�%������n��O;��)���>���(�@ "�+P+'A]�� R��FEh�		cc=��܎7��pu}�W���Tg�h`(����T��������ڜ�QB�l'�=j�Eö�Q�0��p�[)O�+1�F�����ʠFt�X0�<o1z������M�'��߹���k��S5��6�b�<V'�::�؎f�փ�͝�9�3����On��W��b�]=��� +����&��VB'-IL�UPbG�Y"B�}�o�z�y�w
���r%%g�9�:w� ��Z�B�,��S�Z�&�uc��Ͼ���U}�˫!�"f9���n0f��7���+�)S��Q�4i�o���֩��+����w�ߜ+���wU���.?_��Z��t���ko4U���.�����>b� z�Lr�����.}x�K����M� ��jB7�<	�H�����L��'m�b����hx,z�8	L&Q�L�Ӝ8n�'������hF^�\f��N������%� v�T�7:�X��±?`��b��!�D)��e_n-�	�~���",���8���>ɐG�b |w&
tI��n=�2{�����5��_?7 �u)֌O�ЙX%W�k������5|�z5�߼�m�c=��^L����k��n|	�iz?4"��C&���f�hTK+U�n�H#�E�' X����������f'Q��^ � j����+�i��[��fK�U��I)ć�ۍ��̄���j^���mR2�0���.1hi3?0-�]Hp�f��V�{�� �������<�&y�u�ny1 ���H~;�Y#8A�6F16�pѰ/��VLk�t��t'UpX�{h�!H^3�=b"Y����WO�erO�_v��4��]�T��F�)8�fBA��7�\�{���1�k4[�n�6@5X`��l�>MpQ���~ů�����ֳ@��{̶(��Oc�m?4�GyK���i�{rd#�>I�qu��6Pw�7�d��0������>1 ^��~S��-d�ԡ���	�dQ62���_k�$��ȳ @�ɟ�a^�4ƣ�|=mV��zk�VQh1�����-������)i���O�F���׵s3!άJx��G��[�V�eZ&ޤ̈́^ae8@����ԓ��;\�v�k�8��Wh������/L�+dM��/���|Y�bηwSn�L �D�X�JZ�%A��� ���%m��Bm?.��n�^��T�����F/��&�Ws'-����ޠ��ږ-W_n���#u��NZ0J���&�*��s�
�: ��t�06mVY�g���'��?f~~�77R.s
�Y�;�B�SumaF�;�$/��l�����k��l�Ey�pHmg�x��&t ��u�"��6G��^W>mى�Ś��N����V?��]�4D�+�^ '��Y�bƱ�UW�b$`�V���Kѡ�L��u�Nز}�W��E�x��U��s�K���eh��Sn�G`�DH�����A�]*�o�p���&:���94��F��$xֶQD�s^����V11W��(��]q<��7���$��V�x��o��E�(���J�2r�8��a%��v5vOޱ����\�a�v���4��N���B]_��q����-�/g!/RW�K\���~��� G� Νh�DelpR�Y�G���%D�Խ=mL6�b�"��?^��'���[�S%	��Iu�qGW!b݁aO����g��qhTi��a�q H#,��B���G�w�^V+-���e̥Y�*�ڠ�c�ãؒ�r�E�r���+hv�l�#�%����1˅R�~��s�h���n�����.:*�e������M�D�����f�#;�B����E$��A<*�w�$�x)�\ga�ĳ�6����E'Ԕ��g�b�űzA"��r�f�	�E�h/���e1M�5�/��7Y�T��������'�e��|����> d��L�᱑j���7��/`( ��H�n(}�	8��fMz:�����ќC4%K��C�������A��M��Z
 ݢ���j�� 1���[V��t���A?�Ů/܅{����O��v�W�^ ���|�ׂ�y{�Bi��dHZu,�0Z��(�Җdi�SR��p�� �����]�`P1�3'�N-Tkf
�$kk��*��93���|W�ކ @
`�)U&Ӆԝ��$wO��K0��Mc�s*A�0�%��m���-�UA��>)O\}��2�����MJ����� �/a@���?��=�����ǵ�ď� x���M;Pu�u ȡ�%=�,}���g������w���;��C/F�q�-�7���;H�	6�,�,9%Sy)���O�x̤�=gK��1���@����%=f�ڟ�\fL
)�� 6���k ���Lp�)-��|�l��@SIf�eI�0��t��5�pY�k	v��l�u@r�44Ð�X���Ƥ.��]^u�s�V��Yf@��"P(����_&
 ;��dW�M�Ǩ�YYV�����ܤA�5��?:)�yy;��O{�nᛳ3x+	@7?J���S�)�#��b1]ݲh���I�#5F�
!/B`�>[0X��)*�ͮ�s��:'��@S�c�b%qV����G���ooW
j���O�P��%ϱW�ΐ�'�q�cR�^I�4R��r �7���~�������Sa�Q�,�'K�LЅ	���c~�m������ˆG!�*�6�kO�ű����C���r��R��0�U��p�l:%r���vL]ܼb�&�	o��Hu��ͤ���d;v$&�����,�����~��1������ (�F�bYi�N�c=п��`L�҃�P`�/#��X�u�֏�	�7()T�*��n�{�C�Tgc)nOh�����Y+	����
T�d���V�����'�P��B(����_��=l
rV��c�7I���1�u	�e[}-���"�蓒w�\�x_����iR}[�BcSͤ��ۈ���R�V,�7���5�Ea`�W{.�/g&��Ƙ��j�;ϔ�6H�p=���K[?$�g3�:0�QT߾����{�]�����v�1kv��\�]8����5�#�a_��ٮ� s�6���	md����.bj)I��I�r�t����(~���,\S���H�6�N|���*ƼY�P����=�ͮ!ʖ��4�-5"J�B���b	�ŭ���@��b x���i����sd�22�%gI�M�̛_XF����y�9ƻ�}�������b��]d����[����-��Kk3T�>�m�5�L�D�I2q�x犻*��� �o`3XB�r�\U��k�1�Ƞ�:e�%���~a�[�*U ,ee7M�,���"��o����r�����y[����l$��� �xbw�lB��ŭ��-T�`����%�w��G㗺�h-gnsft�b�����K����}�>Fx�Z)�9 O��'>R���=W�+b��^�l�/ ���a{&���')��	@t٪��H�f�q�K�s��Q�!�MP%��oڞu�����T�ɋ�Ͼ�,�I�zs؉�ȋ��"y�'�5"=:t�F��l/V��/M�~���_�>��q&��Wù�Y�߷zv���[=�4�I)���/�cg�(��uO�hfO��$�����5=��(&Z�@O�J�=3FY}�2�l�|Î�Ȭ�� N��HX�L��Q������x��rHU�E���r�gp����O�3c�3��Wˆ6�%jjuI�=�>�n{�יa����hp��=��*#o ������V����[5m	R߶�Ldg1����QǌOF��K��V@\R���j�ٽY��F�O�{������������
�Xh�n�����-�b4��'g�愥P���"rB��oy�s�"K^�����a��f�%K8D[(;3�jm�m�+�bi�陹-�$8��n�x�?��_,�Ɔ�%��Ƹ�yh�@�fQ���t�uI���3<�S�ړȃt;^�:�XY�_�r�����鯱��$��$��z��X4+)�1@d�Ր2+ �� �y���>Su�Uk�R��5��R)9k�,���0D�f�Y�2�
,�}��5W|T]9ju.�B7�������� u�j�C��7��`��%S�1WO�)Ef7W�eܧ�#���^,վ�_4Zn�ae�iڔ��!\L(�n��h8���[CX�L�>8^T5�q�x��Z.��2;����Wʢ�^E�*)�{Yl8܍�ۿ��~����0��>�(��"n�Js&}9�C"<Dʞ��������4	>H*~��,w,�IT*5�{�3�>k��٨� LW���R�gƨ���'�&�B��[�k���q���Y�Ú�C���t�X�q��ƻ��l����L� T+p�?����k�gp�V�����"���Hī+C�KMS`�:�(���m�9�l.Ȗ!��K&&oM�6����,�~��zN��/)�c�$+͚�In!tST�2�����SL|+������̳l�����2�&ji��m'��5�2[�,G-(�;���In�u�I�b3x�`rP wYA	�/�y�u"��5�������6��iڀ8]����_1fJ�y��I>�ʗ!�fTM`�.Q���?�D�c:UEL�]nvc?e~�{�����ϻ�8������ʖ��!�V�R�GY�rԑ&�my_��p�g��xS^(��f�5�	��7� /E����-���%�����#�&';E����5|�i3���]�X�
�0�T���y��C'w��1�>���ʘ�z�3�1����v��t�����?��_�XPoà�u�����P��)ɦ�@FWV�Pw!a4aLq}又���p������؝�Lo�y�[�G23�N��#�|��N2��Z�a�r�:�_��_���H�>%S���}���x�Sr%{'�5����<�$�9�c�`n~/諹�K�e��F�ͳ-�����<:	�af� �_(D&y�[@��"?1�@� �ˆU�6샚�l2U��4�����4����0�c7���Pl��]a~��P��ӵ�2ݱ����"����Gw<�&r��`�E�\�A��z��� e1ǳ���x�q��l�ҏ�{'��El]c�ɜ%���0�T[��|7�4 ��%
Ѡ2��84�s!Y��u�'j���5  �wIo���!I&��� ��('��G6�Λ�������U�=��o����P ���b��*�Ic�xFf���º<���ȖE��.|���y��R��������S]٥��<�l5M��0�L���2���%��7E�D�̏�/"0��>We�t�*��؆e�����^^�T� �R�_��ٝߏ�9I{%�
̙���ۗ4�vF�Y�D�y"5��&;S7@cTv4�>ӉW8���
��&V�oEv��%���#̖&s<֨HT������s�6����{�-�n�0��������|�z���م��t�E�ЦǤw)h��h*l�����פ��������s)�Aj��˓T��k��I�nȊzq�P'1�&I��N�`����N�U�jl���:��(ǡ붛W��6�¢�u�D��=}���a(��� �����휷���0Η�M]��4�B�'�F�b�U�b�Pv7�F�T��B?Ë́r�}[��7 �,;/�C��.�8���Y�-����r��e@,��P����۰�
 ��'  �50�nk�2G�]�0n���,��p-p_&ݻ7����("����������C�~�v|��SifIV7!mj׷�x�,p�gs���z�l!i���@�(I�o�I ��I7+�7>n����VWr����l���$
��i�J.U�:���(�X���`��������>),c�|��EǗ�rK�^�N
�R�llk8(����(���-�<&���r�ATg������A{������ǳ?;�>"Oqo �Dj��̠7�}Bq},�8W��APF6Ǔ2Byak�:O����3�
#F�/�շ2����_��4�󻴽�������ҷ;)��]7;��U�IT*�Eu+B	#�I���H׬K9��E��=�����>af�]\b��־ٜT�L�=���� �AS
�L�ipwgu,�ÒL�s����h�5r����9�B��8��]��3�I>�
p���oa��A�u�	�b#3�t�rƹ�H�,�9����Ԑ��Δ�֭�}�cfg	>l���y��:ԢD��8� �����eb���jզ�b�BD�/P]����"0�d%�i~UX��������-|������K���^�1�f����&~^�7���46Z
e�e\��Ѭ�h~G����5�U��CYP�./a��l.8��ζ[8��8�3�.����y2��f�o%J�Y��R25Mdթh�MON�VD����n+��+��e5�G�L#�W��2�j� U�ky9
�G��}`{���շ7����^��������u�B�ﻔ���qم��ZL��\��z�R�@V"��%��AxQt���,#��C��l���T���V�ob/}wǽ��������(���
����w@��VŶ��7�J��P��w��f�2UԪ��g;I�:��#�F' �D�:�dP�1e�j�z��;bm�E�ĉ9�jᎥ���s6�˫��(�`Ry<�(�[�� �F�r��s��_0 54X l�DRa�r��}�BU�W�+��n'W�>1���7E���Y�W�`�������6M�J�l��Q�\c�L���;v{�⎚�b���P1I����<cYPwea��n������8�.����7����R����P$�	�f�8��V$�z�;�Ŕ����j�h��u���l�:G⯏b#bUF
]���Ԩu���C�.�.y�D��� �	N�ʑ��׷�>�����6>���l��8����l1*�r����0 z�uV�K1g.4�d.��,��{ƫ��Y����N�ja��z�`��y"��YY_Y}�Ca|���l���'\l��4詿��z�6���OjH�e2[�yс�ngT�es%N��T�&Z�:����î�gk/5(��W`O�.�(�+����;KI�^$����з�o���Zm�k)l8��ZP��R��I�7�6�B���ֹ��8��}b�Zi�,�ڨ�詈��B����|_�����vR��Q#;�s�G���:/�ƌ�������6�E�%�-�xtIX��8b�D[\��P��t��n o
����:E�����\��7�[	�G'�/T'o���#9o4���]���t=^2����$��҅�y4OuZju��������=ۋ1��E���_����}����v����l�geD���s�GU&�C��e��uM+
��](#R.-�2�0�n�If �`e_��%����+�ֱ�C������M��  d�IʊG&�Gq s� s	m����Y��2>�~����Zt��;�I�1��{g�"ޙ���O�FJm>�M� ��Rn�Dt�vj��l����&������bbT�q6�Cc�ྛ�cZ��8�*͘�g�O����h�&A~3�X�lQ@�jnJ���
�Ѯ�c�c��x�7���wG�,�q�������0h�F|�r"��Fo�EH\���J��$vt{�u4�?��ɚIƧ��������p~���q��Z�Ր��P��kt�r[��m�~i3,��������V tKs888�O��\�n���x�_���������È7����n�q�ܕ��
v�edv�>S�tf�ĉ&{����RK�Bc0�j�\OP@�N��7��;y�r�ÓX��f�ǃ%/`�Τ/ȡb��M�X"2DDB<:a�D�wo h��b�z�0_��If�S��̓~d1Q�G���/"��/`7^��sv�A8��ˀ9M��T���Q��Ro�&08k�j�
��=�r/��.:bJ��Ey9����#���d/I�U'�����L ��=/*�:T�9p����e9?���ۏW��K��"���"�r8Za}E�����JiJR
Y]����) �Q9�F�w(cz�>��5���ue�� �����,i\��~��п9��|g���8�P:^\Y�v�8Np8��'�g����$a��^�?j �u�F�l�VJ�Cx���V>��З�ڜ$���`1��_�����_ \��:]~���� ��Ӑ���>���;���C�;��$n'��M͊$�gR� Q]�`�Hg&tL�Cr��aTDʎ�8(d��_M�����y e'u�avǀׂ���`Xg�P��=$��wJC9-Y�M<f �I�:A�F�neyw6��mo!Z$�!11i1��jE	[�S5��J3�n@HyV3��(�'���X 9�s��d�� �&���.�8o���2\�s�!�k�,�O��߾�Վ����ڍ���V��,�~�:���'�
8�_ �<�˜��S�[|0G�J�v�v@-�.�qw��wB?ʢ�z��nS,�@�(cY>���Y�^�P�y��n�������b���s��5��H$�uX��ȩ����#_�,%��Gr�x��D"s�"W�Q��Of�s�^��_f�AiV���P�E�������+���J{}����:��o��ay��7��9��M�S��/BSŋ�6�OW0$
IweE�č� -��R�tְ"�(Հ�X}�$��AO�mK��Cy�cK����\�c���L_�?�
��7�:�W�t�qE�Do�^GGU�b(��hN�e@cŻ����Z�0m��w�Ƴ��ΌӐ�k�D�^,�	U*������S�3�p��	�B��/a�p���X�@(!̓�4�&G��4@a5�<Q!Ts��-�	<�h��I��P��V�L�pUD�O7����J*����jW�ܔ6܋ث�'f���#��M�%I0�c��-�"�ŗ�c}2/�.�4pἁD���q/㚌q�� @��wy��77@�?������$��\�S2��ԅ�P����h{��^�Fb��+)�W�f���<��G�</Xj���6<3N�$�qx(���At�s��8�<�ב���F��LĲ&d���}XU,?y�1c�h�1������Q&#���$&6Y� ��F�I`��L*.D%��-�)A�K��Z��jf�e��eqQ�^�Ӝ����(�����O�$Ovma`�{����i�W�|С���ʌ�V� 1�qy7����`�4���n�z�Z���I�M�4��֣����E%��*� �h�P=c����]�A���O!���T�.�9�tݫ�wl�O�&x�d�p��)����+�	�&�N�s���R;�mQ�������������午�l��͒Д��v��r�����QE��.	44Xm���|p�L�nP]�83/�E̝e�5�	���-�Y@ʾ��s� /f}�i�Ho��]�h�,W�.
� {`�Y�]��$I����h�[%�����i+��Y�a��S=x`�ÿ�4�1��`s���������"�{�4b֌�2'��u.΃]=%a'���V
�8j��&��UW������4�C�U���,Z�;�	���5Y+��#A6���-j��+�;(��-�Ę[���o*q3X�PcI��*�5��"�����ndp��T�W+��d��<���q����_aP��sw��=�C��W�RR-���q�d���X	ѶgY�g��d2�[�L�l5=B�d�q$�a^�/��J�� m�IB�l9Nv{���*�ʵ8���=D/��ӄ��������Eo�}�f� w�������qU^�~\�*KV���'����j��u�`�O(.�ui�2o�l������mK�ʫ��veA�-@%����x��ŹqI���8��j��αt���"��A�O*�uQ3��A�R���j���V�M�:�F�Ax��|�e��˽��r ���T�dcS���c�{�e��,b�ԡK���L+3� y<�ko?�?�`�a�w�Sa߳�����e%4�u�ox���Y�a�"���Ǔ�d��h*.2�.���D�yT��n#`z���*�}0� �&�#��	������`�Q#�L��М���~�/�f�������wё�R���w �v\�e��1(C��b{��Wb���aT_f��E�cQib�� ��([ڵпM���LEOZ���0<��D?��_�P:�aˌ���$K�s�w1Z�5�?�E>HQ)�eqJ���P���������fsaN��,x���Z�Y"�3�5o
�1�}��|�Rr�|wy��D�7{.L����c53�<d,��IBs2v�*�RK�f?OP�R��6rc��Ӧ��'q4I�>�Ef����c��5Kr���bu̡�q��8�B\�̸&�9Gש�Y��s������}�jhR3r�C��� Nڇ�-��K��_kz�mz�^��;f(�^S}u=E����n�T�
������N=H�EeM(�l6�G3�_O�2#�R�i�� ���y��h�n�琶��I�xkt��������L!
�U�/��B�;��e�P���� �ˉ����w��i��:f~,���J��x�=�#��Ru��ikii��Y���$���D��$���A�YX��
3:�ݶ�7ۤ���7  �IDAT�_E4�Q��Y�/�'ejj�fv[��Ę"��EYi?��?<dW��G���%�<�����AИ����o���e_�n;��A��MT����盝��D�WD߫�ݮ Ȯ,�q����!��$�oi%ĭ����3���n&֙Jzͥ���%����\]�6#�I#���y�SL��,M��U'�`��^�M��6<e��*"�G�(!��ʺO! �q��)��)�P>KVK
2�c����$��M�$b	7���&K�����W�Ö_e��u�I7*�H^���k�^ ߗ�X���H��o��ɒUW�D��G�HW��rY��єE��L�쬇U�v��nf0=���_��Ȧ��%����&�1�uN���H1[L�*�e�v���+dD�ɘ���,n��u��՚�߶f��5ǨRP}� A���D�P2�q\V��V,�su�����oK���my���N���h=��Dחv�28m�a#}�02Ĉ�/K;� (��<m�V��� � ň�:WnsqW���5E��a�ua�9[��.�>��A �s�	��kql�D/�1���y�s��+�g:>@-A���0�Z޲0}����Yt)�NV�
9��Xyg���F�{1'�I=�,r�Ȓ�Hg���2��]C"a�,㍔�"Z�|�'��t�ee�
c�){��%ډ+�� h���W�J��n�ɪą�ף�г0�Ͷ�3�Al~SS���z��?��?����8hˡ���;��I�HJ�(��gfPV�\�\��� <��<g�m%�L�(=�q��Y�s/��̡N}�L�c�㩝�u�Eʤ�Q�&������:	���<����i���tRip��!{�`̨��OK.bs��G��XBI��=[]VF@�	q� � ��Ua�E${w�û�ޞo��;P��_֤qXeHIVu�N,�_�/Si��j��=���޴��ZU����L=�����KʘgKKϺR���L
~�\@����*�ǯ˲H^ު�ˢ0�����-�Y�FYh�Y��_6��������7�t���Pu����k�	�,��v u�2�)�A�Zc	!�l���e|,�O��A�V��ֳs}��d����`���HX#j&>,�7�I[�<�GY��ryG�9��ԺϤ}�l���\ڪ�AZ�~�;
J�s�Q(�
��+tU1����?�է2�'���i	hϲ��`Q�:,į_�����3g�(���53�ҙ^�H_�Đ8�|:S��ڛ�]T��:lv�CM约�;��Y�`M���=!E���+���,�	&cc���9ԑ6���y��"�X1���Y�U?;�&�q�t�n�ff�"cY�o�=\@S�ߛ�ov�f�8���yz#.()�8q�AF��'Qtr����d��z���� �����������7���:��7 2�c��䡗e�
���~�cvx I$1�hk����	<ע���!��|m�f���o#6�l�<$i�a�4�<�)��ǍA�5��fP�ڙ��+�uߞyF�����nO�+'e^0��Ga}\�F�;��Ŝ鈘����v7R�N}��=��Ma���A٧3��'ikN	����0ԕ^��!FP�J�%)�|	˴�4�3��(>\�l��f6�f�1��2 ���ҹ?/��M�$�M���K��A�ЧI�ƒ���I_��Q�ep!��0�9�l
���� ����l!�J�)rv�4��4Qʓ+�
5h&���=�M-r�
PU�������t'���*��&�4�M�?�<���w;SzS�����e� X"���Y�|\�v#"M�2��w֎:ar��fBXȓ�R�ϖ�j��}6�<�i��{y��Fa~�e�^ԙ��0
��nP�]�8^UE��_u:׿���A�3��M�2���4{�@�GG&(pK���:U��`Ʌ��穴��D�g��E��%Ǖ�����Ζ0i)����y�f�7�.�4��-҅�ez.�� ��D����gRs�z&�8�g�ʈ� �n�L�L�P����'�*���)�u�	���,pX^�4��{�X��BŒjq9"��BA$��R&��ƛ-�oyQ���zA��+S� �V�(u�YïΊ��et&�I��N��g9���`iN9�,?���J�U���sx��ڌ�\4��m-���n
1< T�\*O<;r���oM VR���퓺İ�L��E4f����?�r���g��8#	�r����:�"�s�`'���͵��к����QӬq�#�8�����8��J��Y]@�b�wϢ����Ge�1B&ey2 To	Y�³���D5ocD�D�P���������Z�>7���7�.X��FA�
�΃��+TO����l��u�-*��9vw�_�{��T���8T3��8����%f��ߴ+�wÄb'�?r�,�<X:����!�)k�li7"J�t�O3�nPKqD�0	y�����B���ko/
����/p�g��|)�_�8	�T7en�N�K"b�Nv�R��1��O2/�$&r�-���u���ժ0����x�j�Bq�v+f�+ f��T�d����db�Y�Lw'IO����n��H�Pcw�"j֕\�3}�[�mx��V��T�~�z_�+/wsBv�C���"r�'obи)��-�p�O"�2 �osV �#�*�7b��l����`ȌP@1)3tF�-
�}-�ͳ��;0�q��q��Y\�fq�Q�}gu289������g�H�@�Q���z<�����$���H��4�����,�y���[B��;o�Z���l= �#:/������g���P$2�E4�<��R��s�\��( �3�h���������;�c_?1����oP6�:l�A�ru��-["��-�h"��R5�I�1!ʜ�d�����We�|.�7i�����t��j#~f<�g��1rH\�Ս�e'�ugo��;+�TV���H������5n��Ё��X�g�$���l��M`b�8�
ZfKP��;�G/���'�"��L�{�����|Ȗ�U�8\H�:��R��G�v8YL�'��+�:NU@��l�b�`,�w��S��	���s� �@c�
�E�T8^�H�#f�Κ�5X�� H��G�0U�|����0��?r$�FA��N�����읲Yȭ��B�܉/D:�α��-�������V�o.�@]/�&h*|Q�tZ/[�v=M2ݱ�6�X�-���
��oV�s�+���J#'W-�o�*�wy	cy/��gS���eT Tz6,�.�G��d��j�R��N"��2l~���wz��7\7㕷����}�I]�EDO=�� �E�gyd��$���uj�G]}Xl`x�?+�b(�X�Y>#�;+��%TQ�G���,P�Rt�D>������	�$�l8�?�2�Gkؾ��#�rO�������N0	���i�&NXmXߴS��'�Y3x�x����\IZA�~̚�+��^�,.1���ǌ@�$���@�������j���Q�����7�<�n�6=�H
	RGs�^�<=�e��-y�����S~!���c��hᾞa��S��v^��T{��I�d���PG1�x��l�-���z�����X���F��ቱ�-���E_Rq��s<fS���
f���h�V_�C�?�Ǖ�qf6�d+ze+F,d�*Mef�&�9~�$O-XȨSp�+Ȉ�� ��
�(]�)$R_�Myeq��T��j#B-�d��Ğe���؎g��oa�++Ҥ���O{�$���d>U�X�HE<�p����pb��2�:�,vjS��L�0&c���)����L1qZ�������	P��;��.��)�9[$�M�QX�E��3˄ɞ��tbJU<q�ɦB0�R�6�z�^6�S�A�y-�^�Ýj�#�b�-M�2�Q�|�1i�Nݥ$q�1!PK.X"0�E:(�2�cc5,�;��W�1�\i
��lץ��qR�~t ����)�3Z�V�\'U@��L�oR2
iv!6� ��ֲ?��U��{8k��yw+�7^_��ע��0S9g���$��'u@4�v�*�Z-��@�}�q%]��9������^ ��\��x�����������)�J�9^�!� �X`���~u�T�t�]X��v�M�"Ys��8���{]�\9z�~N��C�4=q�1x�B/�� #�G���B�� 0���TQ�mU���l����A+Xa���<�b�uX��~}�a�J�c�X�D~��%y�? �,:B3�ũ&gw��&q.]�+p@M�C�"�'uP�V1�Z���ؙ�h�;�B��,�[r �qbƦٽ?R�;��2��2Zٰ���ڍ|s ]�j7��>�-��d�An�w�C��r4Ե�k�vFr�*��R��%��ؐ(�@�7��
 NW���
��*LsЈ�m�/�~[߃�V���>�6[lm�����⯺wa��G�(ˆ@:a���K,�L�l��ž2i{s�� �rD���g��.
 ��4�*�Z�0A@�Z��D��u���0����R&5�M�Fl&�%t�./~��Y>!M?u����1VU� �4K�4����YZ=͸��n&�Q=��*�(p����Q�h�	J����𤘚س��;�l��r	�8���R��]7D7!��Ҫ��}%]��ynTp�n�X��9M�mi-�m@P���t:M#Q���V��vNӣK?���>S�@�Au!�
j�Gn)�{�{�[��k��+�
:��Ϗ� ����������
�5��hq/���Θ��ۜo��:�t~��o�����$!UW!��w�
�2;u̮h�o�,��fk�j����kx��G�|[���� j@���;<�L1�ݭ	PI�KY�l�\���)�;k��a4+��]�����,Kv����V�z@��$�1�jwv��|K�8��,����Q�6�a8�h�8`3�0���*���!�^3,ÈP}���L��5ZT����,<�m�vm��Ia�D�4$p~�r�D�6��HS��B_����.�oO)pУ�8��,:�=������S�ck_���.nzm�'���:6���rW�؅�>�����
�7��H)�]�"��c�w, x`�/�yA-��rN�m>����4�ɥ���L��2<_�C�`�O}T|$����a��G� ����O�{�����%c�2�j�S��z��ġ�9DT��x��	]w%q��p���V-�mb��Wvc�.;1��M�̓�Y%1��Fs�tFb~�P��h�u����4[�+a3�C��͍uj�z�-�������O�W�p�S�}2�����2�Ɖ�'�_��!g�&��g���|[�׀Cڲ>�/��T tP�zf@��m�VÃ�aS�3�C�ϫ���*�{����\��(��~���iSh��YB�A��"���Y�6u�(������|��bl�������!��	��+g	$��x_>��lEI�,
 J�;g�ѣ� RWL�f�E�e��>p��{�>l!�Ka�d�z���0����]��vV��0Oi���_��
DW
r'���:�=���qO(�Y�${˳"W<�%l67�k1��t�P��0B�)� ֠:.�{����0�8��Ьx@�ܪ������=��F�_(�A��~�!�Rw��}��Qƪ�ȃ�R��5��K���ԑa�V�_�}�z�[)�}$���A) ��D�J�{�שˑ�\���C�Š*h�r�fj�}u+��-Ү,>��ks��.4���@��J�R�O���3% ��8�<n��񹰿���q+IY9�J�8}2�/��4�X�p�UԔa�("c���۱@��so�.M�W�T�Xy_�?��u��Y^�����.��~7�i�'�@L�}>�u�2��I��{�ge��V��)t�t���T:X�sN�zQ���d���ډY�.N֠U�$��-�����}ȔV�Q�M�w�,�O��2����ţ%t�~ i�׊x ~Gр0�����k�*^u���^�i˨Z�S�]��?q\����Zpl~0	�ZZ��(������}���\�Q@�<>�X�m�8�?��������И��=7V��_l?�{\t���R8��~5#gq�\~l�( 8�D��l(Tw�^�X|�c"����e����6�Cg��T�s	��Y��m#����&�`���ܣ甮y��WO��� ���������+�3��4���G��E���q��p�0��x�,�p%.��.��Z_U�7�6�;q��AB�'�*h�J|����# j�p���zn��y�k�U���,��9���z�	�� �>-.�,���yNMk���o�>>�K�@��� �j;Ò/���v�~y&�C��㭂�.AeS��� aP:q���������;��:�w���Xu��������1�<ƥP��i�U���p+5I��������vn�⻑���#�y晚�A�mcQ�������Q�_ �'�8S����竟6�?�s8\���hތ4n�iJ�d:3��n��8��|M��z�d��̑���tFٱ�����2�}Ё��$�|�R���vr֍bz�{�o�q�X)ƃt�_4ǯ�]_-�i�No����+�<����-����������V�nA���;-/�����"bt��U�E3_^e�h���ϧ�����N��S6��mT�:J�Z}5�Y+���?j��|W�ۋ�G}��u�����R��s&��!* ����6���Z�=��H\�����RF�J����)���v�� ��
D����Ay��|h�·�k��D��Oe
t9��Hzt�FD0�O��
]����N��]{s�S�GOy2:z�>z�t�&BI�W ���N���nt�}x�N���1;��8<�f�MK���ef��F��In�����5�U�
*��Q7!1��f����D`+sK_��>_���QBS����;����ӳ7�o/
��9�;�|<�9o�8����{M��6f�h�G�Y�4D�Y��sDܡ������J&�5~����{��
��`}W%�V����Ή�C��;wr�����e=�.G�����xr�c����O��`=��������[,G����en��M)D*%�{��,Ղ�SYIl�C���J�o!�]��̅�y���(���fX����-�s��t�X].�dA�pF?��g{1 �ۿ�����n��`K��Mi�3T�������ֳV!��B�ėBx�A��w���7��;�(��Q*��R�zc
hh��;�B�|�s{���-�{
���|�=i��5V���9`���{��w^��%���o�0��q�z��%lz���JQM}ouB �J�a��Ո��9 �y�AB�d�JZ~I���ŭi��� H�姑�Z���'�"2-;}xu� 'A���A{��g�����i��4ƛ�� �V/B�;��a�ϥ (p���H�R<�6g�b�
h���Y��-����8%��:h�7$�D/3NyF?��O;�⺮�X~�(+���Z�f�>op�C���v���F�2�{��'��_��r�w�C�@�������s3���&[�|-����ѐN-M�&��4C��aֳ�=S2B�:)[|��'0�򈺝S�4 �`{�~���?�9��/��KӼ���7�q���X�J��nl!d���"�L̩�3���svB�%�+gm���˱��Ef&��JRK����F�b�U�qi��o����ۭ��щߞ��[�o�/߾d�-��>Y���w�1@k���~�]щOt�uO���&���\�̯CV�ְ/K���Rw2@2�[�I���������&�NݒV�g�����v�/��H#�e�Q����µKu�R��� ��۳����D࿁��o�j�����|*���0�C�%&��G����<�B:���q�6t�������Lӻ�Q�ˌW�@�h1��rYɶg0���0N=�R��g_���?��T��S&��S��;"��~t����P�{P�/�;4Ƈ�&��;�脡%v]���f�ܶBV#���/��Oh�]��W�'G��oп�t��| ��L�@Y�,�e�����i��ҠZց,		h�V$]55��ح����(/�I:�^J@f?Q��v�O��o��7��}A��asss�v<�o@�m=�+mn�U�ʪ��m��,~P]�Wr�q��s.�	�qꟙ�,�i�=f6�K\^���[H 9��[�#��w�Jm�"�$��ŭ�#��k��c�|;�O�Ή��%>���5�|จ�y�'�~-��Զ�t!���G�Ἴfϑ�0���6�'n0���i��`~duS2j�
�4���1i$M5%Q[~]3�p�����N8��	�>�D����? �v;���w7�����pVX`G�[iR��\X4Y$��\�����DR�r�مR�i+�x%�<ux6E�,�&)�׽y���tZ��F���Y�Y��V�/ֱ}�w|�2������1�~����+�'�~}-Ʀ��6�[%�ɘ����OMm�H���x�!o�[�u�!�z��8��Q�){v�h$m��(v���?g�z�H��6�����f�c���p�����z���mow��4�$V"��W(�Ȳ"s��<Y�6)�guh�q��l%&;6|��}�E��Jہ�rBOЄ#��\ r]U.Z�.`�@'��M� ���7��&���.(�O���1N��������c���~]�=��zgaqzUTw��CѪ޵�Ĥ:(Q�ǝzLPB��� ��������}$+���AJE���C� A�	�ro�ufs*�Գ�K�C����E �g��~����3�ݸ-"���~ ��j��@����������Z��V>�g�PB�7�^�J�;f��e�$�a�O�H� �F;؋��wz�c�o(�ӕVhQ#��1}��9 <E�C~~��@�����5�gB�-4}�x�{.���6k� w�|�-�>��ݴ�o�Ggx����c�%9�E`��i�D�D*���z��uܱo�W�/��zR����o��`*�G�a���a��%�����$p_ym� ���:˖�6�"s�:����2柨�SA~�v�=n�y*���S/�酚�*K�c��Sj�����DM��̎���Pv���=���oS'E��T樃�kXz%Y�IӴ�Z�މ>r���=JOx�U����\�d�| a�ԧG%>��ͳ��	'Z��k���7��Tp�����&���bE⡳I�������M+U�������@������݉�-MjB��D%N�Y�����Q���YLgh����f��i����/��>���0m
��L�<��܍\�t��B� �ԟ�kg����3��f% ^	L�`��-�G�
n4�B.t�s�I�$���^�Gƛ��S�?�v�
�C��:��L�߃�6�ЩÞ�=�|Nm����kGॶ�����	��07���RA���TT,��P�	 {=��(�g�RBݘ0�[���r��	�>q}��m	������Y�&��������(�S��j0Ѵ�0+}���/	r��x�)��s�蛴0z��,k�<b�M{Q�:�T�4�^둏�au���eRo��B<]T�B��l�ۑ�yz�R�ӣ�=�B
����o�1���=6rᚁ>�_)M�z������u�h{	<�08��(��p��1�:�nk�.GEM����P�z��*�]bX��ⲥ�R��hK#�`Ҙ&����Z10iي�棅��� ����L�y������?��wx��L�v.GDB��$鰡Y�x��"�j�htQ��@\|EW���#�<QPG�!��LE	O&�aA�_��_%��_������e�Q'n�x�����TP��[�{�\�Ǘz2{���G���r����S=�?m��M�=�=��q��EjowZ��R>��al��qlp,+�k�/,%����0J�ղ;Y�����q����ɝ}	E/�,ti�mɹ	��2Pzf�~��/� ��4��"��@�^�Β++r�\>1N\a��ڒ
�9U�ClO����ˋV�/�ͨ,=E���L���
�{�\X?��ΒS���z/K�wü&���L��nA��d{!��S��~�͸�x�s;P�v~�h~)K�{S�i�R�~�����jtHKi2 rŰ4 �_��6%�:�V��#<��s67gEbc��f�,5vr��>���o�v�|Cg���R���ׯ�/����s���)����础_�g*�i�z�IZ�Y���[B����b�������]o����BEۇ���>vvb�&X���.}]�գ �9���O~��rg�|[��B�����p�E���B������;֟^�5Il�,.0Y�^6 苬��0��4m���eJ�:Z-'G؛�[���M�Ð�t�0�����?�^LHS��1�E����Pb�2ª;L֙�W��V��i;W��F�d������.���U��{`g�!P����?����N��u2G�]�y�����^�B�Vw�� ��|�Rwt�IhXlm��nY{�/�%I��N��9/uO����|Q�r~-u�vu��pp��!p��c-`O�4�����r�������~ӱ~�0���Y�-P�ZR��x2Te�2@\��
�!@� B�]���b.�T[��Wյ��.��Þb ��k�ީk�Y���ߛK.��*ǟ�x��>�4�mN\��h��3O�8�#��yY��)~��h�Dm��V�QA��f��c ��$1�9�� ?;���;F%�"^�V�~髭zV�g�É�/���E ��p9��8��<J�w@KH� �N��K]��}[�! 0�AD7c����Q;n�V�η���\`���������ǻ��&.ݷ�
W�K��@^�xH�О����nx�3�w��4N�Ӭ_[V���U_��p�k*x��	�<�f6]�F÷��`��E'd{���I���k�"ҍ�\�-KJ}�pGn�c&�Yˀ�6�O�
�ۮ9�7-��,FO���$�- ت����R���n�R��T&��b�ub5m_���Dz�`}풿�'0���i9>�n|v��&���c�������s]��g�k/��@��ҤN�&����h�d˲q}�f^��[��4O0��p6�*T[&1�2Af����z?���t˹ H��eTu�G'!��uQ$�Mk�:��ϒ�_y|ً�m��"+-B���]�-��A���N�� ��\����[qfu�p)Y��a���zqr�gy�m-������1��Y��}Dϧ����1-�EG����J$�5��<?����O���]������%���y���b��E�{v��>�����z<�SnꤐQr�%9pa2�t��'�G�XWgeO�/&����WGRn�z5�WXr���j�
�k�{u�$�ue9�OU&z������c<�[�����%.� ��o���x�z��\���-��/����A#*���p��*�>4���c=��'�,涥�)_��YG�\�X��1g����z,"�&�\C�G�s@��.]:+�����2🕶ۏ	;N�=)�?��,D�q���l@���2SXd��nz@�PL����fR�$�����v��ӊ
ܩ�[�ܪg^��S����7���h⮸��9e��~8�����`M�W.Oѭ����v�:"v??a�w~������m�}6�c��)���z��	���:!�_�׵HR��A)����'�QK1�x�+?�Y��g1~L�8Na�~���7��,�����e�wm/��Uy���%��wi�R7���������Rrۀr���܀Q���aBk�#��[;\�n^4�S���o-9-�ce���ޏAw=��ʉ��{�v�2&��}����w�X�y���R�G��`������L��뻑�ǔ'@�lR Lz3���<�?�*���"���q��9e����� ����t����4�M�����9����"���z��* v�Q���O&���� L.�~��i�N���\��2���Yۂ!�~[����
�~��o�Oo�w�� �<�)�;�u/U�2Ͼ0\�R~{Ǣm�Km����t±�u�
j�|�"ZZ@ˋ��k��u�շg@s�����Oי#�9x@��2Ve��`pzCn�耍I5��){���2ґي�u�j7\���Ofό��/5���n)���~OG����E�/ޞ��}bةm)��+���W}�T�GM*hgpAB>� -��U�RILUR~WV�;�ϵ|m��9I���e��<E�ko���(��'�����ߞ����{��/qU̙����P��s�-���~��5��:e+�}��kr���~�s
<"�s�`펩����8u0f�uu���t�w��c]�S�9\���f]x}m�x�%��B+4,�e�vI�������EnsK�fP
c!�|�~��	�|��*�z�@��-��M5L��׈̞F���[��k6��ߞ ��������ns;��_�
�[Ǫ�K�*J����Y
n��0�	#rW��o���1�nu�t������l��/?O�+���+��Dm(`�+�=j���r#����	�{��Z����9�6y���+��|Y5G�j�!��k���Ͼ���m�LX  �X����C��/�Si}q�0���*�D��QB�1֑Gm���3����O���e��97�ݰ��4�RX �9;V�
����[��!ƫ������*�!֕�t.f�@M�0�f�k��)����5��)�3�����/��U͹��юyIQ�!`�?d������N_�'lw� > ~-n�}�J$'�tJspti�U�Qa��(����$5��'�Ik$V���suz�x^P�3E�?c2=���+�S�n�;rȊ}��{}L���D� �%����ߧ��~�6�8�Ӝ5���z�#�;����ݛ�ZkĎ��w��I�g��`Ȁ��~�cB& �P���|��z�S÷��p<��kKt5�,�z���l�M��z����ӯD[���t����N@kܕ���:q��x�������Xh��-�	��&B��a�82\ԥ#�%�>r/s$z���M��<YW/�&�z�!N0b3���63�f^gS������g���s�60�.ĵ?����b�4K�{]�w���g�ΰ4 ���h�	xt�
u�w�d�$v��=v�X�M~�F0���'X��E��*�Byɘ\�?%j4n'i'U{�澜!��|��q�3;�N��~����mxt�ŧzIg���	V�/!�$'�"5kd�S�]tto~۸'����Os��ģ�j�s#�O3}B��qԁg���4�圸`�0�HZ+�hm?+�uX��lRFgŎ�����,�(q�F�T&~,�Me���#N�:��*��-�v\��+`��������������g)A�N}.�����9��Dg�fݒ���͖��\�c���������.۪$"5��"!x�#���EU�:#�G|ݿ�ֲ��Yơ��}ok,n��E�k��X�W�b��w;�#��||��	��~Nb)����'��ۓ��)�sq�1��񱭶Z�N޵qIWo4{��������p����$K�EV��p�s��&�w�����]8������� 3��U[e�s�i���_W�߉�I4���ײ=���U^oJC���r^�h�b���8 
\rm�<��<^��Ӑ�(�~��h��t����)�?�@C�Ҏ� �3��- 
�8bD���M% �'85!�Ɨ�^��w�C��t���֠u�=�A���ҳ�}��!ط-���>f�w�ֽ�N>Q��nm��F5�z��V���#s!O���9��I��1�� �R��Cc���!�D��$�!,��,zA��P
�Wߞ �����)��\"�8��d����Zo��[��H�F[3����K�q���~�Z}��`4WY��t��J�<"5A�����.j��o��^��N��r��؜��X��7�q���x�\�l?�����}Ow����~�g�Z�w�>h�|K�;�?<�����k��� �ݖ�r�p�r���ډ�lL�@3����$b���HIS���]�pl#��e�Ha/
��o�~�yr{v |����B�6C�v��c.o�t����@a+\Ji��4ʋ��o vb)$�њ�7FI��,_����L��	Z�"�L��%9{8ڧ>�y��wU%�j�դ>�c���%rޅ���%�.������7kѣ�����k�]���rw�*�Hs?p��I��{o徍T��Ű�9w[@��#ӼG��NR�'i]��*I	#����Z����OM�}�}����2�^��o�� ��B�~] l�X��ʸ.�X����v-�A��Ⱦ���\�߼//@����+z�S#��,�A����_��O�:Zp���5�p��nY��S�FǈT�z�Zf<FX��Դ�qR}��	���àq��\��a
w�],�Rk�z�v�T��}^�f��T�O8���'ޟS=:�k�r�Z?2�?
/:��,����y�pS6&K:�)��Na_�=��bk�4*�傆� Ѧ�"���n/�f��?��:
���ZA�A
V�8�Th �,0�"<�n�0z@�	�:���Wӭ`�S��_=�\�Ā�^�U���W���Y5��P�������Z�}��3���ȗ'�˝�h��?�H+���CYp~������6��ދ�E7�>9�-�'CR �1�!�"�f�����2��G�jr
�]��&yn&�y�^���`��?˩��U���B"�Jpx7�4pE�)-@D	N���%pŬ�>���a�Ҿ����z�F��Y�/5�˅0?q-���|������V��V�GX}X+�+@��/WC�k\>�n��s����k�C/\I��N�~��O�V|u��],��ݞ�P��k��g%��5sZ��,�
����s�Xo���..�z����x ��d%en�'r瓸���K���i�_��w�ܚ���^�������g����G��T�_YB&	�������E�,/�]�:g���X��O���o�N�'s�TGh��(�\5��8*�8����G��j��.�N	l��䆛�I�)����~∻��V���>���G8���}�?�9j��y��_��μ���ú'-���ұ袪��P����fe&N��B�ߤR�n0l �C9W/���װ�	C�ܳ�j�T̮��Br%`ڔ;�|���^�v�3��ιH�ٖ��? N��}�1�&{I�gf�3����7"��uZgG�!+��JJR����U�xG�����t�&>��0{$��}�w`oD@s���)��"��y�^j{n�T7?�s �b��?�w�q���d��.+`������~����I|�@��������쯀��VHM�r���Þ��q���� Y��zjP]�Ȉ�T'���o/���Y�~�v�Ș뺊:�0V,C.�2�LZ�@}�F�i?@�ed�r�1�&��. �7�Z^��3�܈�qe��4䮑���Њ��0@���j����"�K/��Ƚ��W�+/�}�<��������C>���{�չ]@X���c*����K_AM��JR�\�63�3�#��Nb{Eꂹ������ܛ�)����rD�EO��I�w�k�^ ��(��K'"S{���b�Y���t! c�"r��3�]��C�~VJ��刉��4�w�8l��&�V0Z� ߱�������H����&��bY�	�p� =�Dk�@����x�N����dz!�i�)×�
����H�����Ԍ$?�AP��ru20H
7)��E�ͻ�2���W����5�x�zk9B\�I:҈�~qW/����*�X���ο���/#�/�o*k�*�B�R�*��0��H�h˾«�H6�8�}��t�pκB���{�˹�ێ�PIb�yv՗pvDU#y���?;~퀕�቟m'<bC����j䢄���ހ/O����
���n���#��s��zMx��F�v#�`+���9+k �����R���2�g�3t��������)b�3bH��Rt���6I��.�!���; ��\./K=�ױ� ��\	.gYt(l��J"0Z�S��d*P��e�+ �/`Y�
 2d�X,-8f^�fW�&�,��u&Y�\O��^��j�	�ӿq�Wkl>-���GUf�D��B ���*5���x�֐�u���Q��?����n/k�WqSd1���&�o�]w�5 (�o܋5� ��dN	��A�O�H$3�>fIH2��]���Xn��T_�rR_D���� ��m_���9��AL�u�LGP+U����ɒ�6r~�d��j�c9���'s=��A�!-R�i�itX%h�V��q�Yu���@�ſ��P����uUo�8�W�:�_��d�b�d�����W׏_�	��v���(����I��G��(�&�bH.ǀ~�.`f��)�R86U�>x<�4e� 3@�K�N�$͹�I24�2W2j�/�y��3@>�]�<s5���bPC6�xa�Y��P �i�&B`�wVc'������@-��ؾ���+fko88�=w�z�:��c�$p%�k2��Ei
T�zp���-7|������ݳ�"d۝���G\��u�mu�Y[��T�\��ge�J'.Mw|8z�Ցq�f"A%��Ow�9@գ��JG�����<�:y�ee~~"�Q-��� @�X~]�����I��?�������/������vsʙ_����;ձ�6�5�b2gM@�>iR��dJY>F�c�d���V�{bŭ����5�P�E�xaI�=�Ìz�:�B�i|�s V����ڤNã�5���ET�~X���-����[}n�wi�ԾS^�w���-p�WV���<-�z���cC&n'�G���d;��ؕ���pT�ޤ���$�T"C�2mf1� ЂD���f���9(�Kr��g�\�da�����g�?+�_�	���Yt|��I��(���ٚ�"����r4=���\>nab%nY�R�L.%'�!���Dfa���)�ؠ��� �j�� �?x����=Ɩ�t"� /�_��`ӆ�}sS��u�����w�,���VD��9��̬�,���@H�AA�Mlx�z���3�H#{���x�3�8�؀��D�Du��i�D�^Y��q{G��3"�>�ެ*f�%��}�#vĊo}kŊg����K�~�Н��Y$��ж��X�TØl?���<lA�R�+�:3�h1��E��,���EtjF�l��� &�8{_"�#_��g�d�g/VT��I־�E�x>�6x�����D��8����I������ݗ?�j�G��X�p�I�������!����)i��Krm e���05� ��t�?]J�_2H#�ԐD��2�X��S��e�����.��7�XkGt�S�Q!g��
x�*L���	��l����R�\_� �ա��Ϸ����%�h�ҋ��TB��񥆝�.i����Lo��p��ab��U�ʢ`�8�r?��W���b�r�$M,<�)O{$�wL ~'&�q2	���5
�5UV�Ky��:	=���B"���q�J�Ġ2��g���� R��3'9t菭�aT���ݶґi����4<�6����$�
�3٧�����x�b�j�u9�N:9��3�-���e�rX�`IU�E�,�n����R~���2�E'R����2 l.��5�r��K1�����}�<��{L�ϸ-�!>�V��I)��-AZ��}<j�ª'�-�r�c۞V���X�?��{�ߋ��%Z����2��W-$+�

�:�qT��@��`�L��}'ٖ��%�+�ZG ��p`Q���Ev( �9��-(L>{��0�|�����ػ�&�� �m��3�n�D4�K �L�-H�m�8A��u*$�C-+�͜�'�������a���PV�@,�*w��l\8r�Տ����M���K���S���E�"_Uh��v�@�b#�r=�nΞa[���u�_S�E�}�þ�a������u������������e��a��E�V��=w��\�\���ey�5їSs�\ۯ��7~m�,��O:����G~?dh1E�/�i�13,�)%f��_-���TNŢ4��xe%Y���$E���B�4���`8*�����L�3�/3�,sb�@�%��O<�*X�i˔h����,���j���0S�T2�08�A���-�݁����n�
�k�]�yi^L�ALF��uWq���	��zɊa�o�������/��jN�p��dQ��9���=wƽE��9'� ���%y��v���z�iW���>���E~��Y��<~�~Y!�dU'_b(,�� � �WO_�� ЌյqrN�Ŗh]�8xɑgj�sJ��L')��|��χ{� ���o���$?�؏xꯐu	����Wj<�]��� *���
�D�f$? �����\���2��뙂�qP|jN�%kki��ȏ�9��U�+�3���{Zv�43(�l��2�
�'����5��2���׻��
���7��`L�5�����Å�,�WO0PZ�}�������\��b#����$��т��ɖ?�\��byK`h�m����e�$f���f?b~��v2 ����FE����B��˷g(�s��Ys��;��P�:<�buM��'gc
4E"?�/{{� x=|�h*�wY����4"L��.q�����U�-R��[ʆ`�A�4>�����t��`7l t�D�82W�\f���W�O5��ڜ�Q35��N�J�Ӓ�C���β����y�����߼�"m��u鹿o	�g7��n>��d�N\�q*��ݎ=���/H�9P�g�*�3�\?u�Y(��ٕ�ښ���݆�T =�����S�����Ǫ,C���� [�'$�CO�>���%���I�L�M���2�,qY�d?i��Fe�3� �weA$��D֯�>�����JL��b y�̙`�"Ss;�}��!�0E	*��MKARu���A~���,p�>�M����S�ԕ�uF�byN� [W#3coZ�@�ĕ�����*�,�M�Ӯmq��i��d~*��l:Sn�]��l��K�V��O�9�
'�3�/�����/�f����o�ϱ�B�=;��k\�el<0Z_+�=�lPrRKaU�,ۖ�\ZP9��5��򢎭��0F�r�I�����$
7�  y�	r3q1�g,�������5�������'���v:٣	��Ey����t �y�q˕Xc�ϗ������	�e��c����D��y���4LL���8f���(�36����'����h��di_XZ6�-��W�ɪ��R^�*�����O�_�U��N���t�l+s�w�i�`�� ��o�äր���/�3[�V{߇���}��o��=t�z[!�J���5��2>17��K��	�L��o��R�i�N�N~�?6|J��K|˚e�F���������_"��� ���  �1KWG�u^���{G�4Ts�,����6�dY�������C9�밽�U���w��\����Ȟ����؋h���j��Ɛ� ��tL�L�(��f.�Œa� ����=D�eո�$fЫx9vB(�7���AX隐�E�Wg�sMi�;c s�[bbȨ�zEk.7�ڭ��
��2��5���o�ݳo!��yu�|�QY�y��Ϸ���3?ԭ���{OY�~�V�(���qrŹ���ΦNd=i��xį� c�0������L�����y}v�y�[�B��r'�G�?@N�GA��ڌ���T��	�flւ
���u������暉�Dx�_�	_��j��N�j6��7�Q�=>x`��x�9��C]�tqf��Gg�&6�9B��:����>@
�?�����2Y0����B�K�v�q��� �5|�s�*A�Ōʅ����s���H�ځ��9�h�u�Z��4V�+8x~�ܣ�~}�v_�t�2��������nkG��V��`ɚ�?p�[�ny��)p���:)�,˷��6�U@�>I��Bm��TV"�=�2U�`2���y�o�zR�󤋉�y�T:���/�y�̚���0�EoT�3��)�Y��ɾ~^��V*�.cň�������ї�|5� sǹP���lx�s��:Ħ�A&R�^�p��<���S��AY�$:�%0��x�)C�m0QN~���Z�"��WF���W�E�)�˚Aær3@��Fim�~䝳�|�5Я�u�IZ)�>Ŷng��B�r%����Pe�ͪSo�b+�_Qw~�������b5!/K�)`Xp�̽����sW�}�W��,��k>����f�@I�\.�� �v������I��?NyE�Gf�M}#��3����p��ST�/U|������A���Bp���?Z2�^� ���fG�?��}�㔀  ����|��E�މ?OL^�NT1�i��
���Ls
 :�V�=�;D���sbS3ym(����+[^4��u"#�J�������^��:�%��b�i�T�nY�uq<��"�Kg/K��g��{���5{�^� q_$��1�/piS�6��O���σ�r���.*�d�0���ӝ3e�%3�px���R�V��Q-}���g�g����f
~����t/	Oi���m)t�Rޚ�ċŦ��ϕ4��ȵ�dC>����cD@%�$wC��g�������el�l.0�"�dcA* �A��ؚN�o���������/�ǚ��v�9���3@�o��{�l3�zY�c������a��n�(L?�ڽt�����Y��%Ӗ�r) +�	�/A�\�yX@�����Z�m�,a�e��
s������V��L��m��������A~����cW�M�^�ɺ�ڭ
�l��V��ZøK[��`h=�Yua>���ڭt�l	�afl�X��S4�3ɨ#-v4Q������C0����g2�d�$���Wٷ�Vv��p:8��+����B����"d��.f��� 7����?�/{{� �u��NY4�c���ߋI+Ύ\�8/���˼�G$�
#�~�T��A�u?��{d��׏��[��^��^K�9b������(U/vQ�ZPY�
��+�y�x�YVy�������� �s^;O'�
��J7�R�,���
z�nm�fݕ���ǻ�JM����NOjI�����2�ڨ��d 64V��9�N~YyU�Ŵ[��ܰږ��1ظzZ ��c���A>��Y�X���)R9�{�وĘ�*�,���a�l�i/�Q���I����l� }���t/��:Yi1t���[a���Rf�b���x��}��O�{Z^z4�}ԑ�l������ �'�S���(�� oB�G�@��"S{��'��Q���mq��G�X�P�PC rr�!�C�-�{�!t|dV�!��/C�SY�D���� P;"�����+�钗���)�#Ѵ������:Y3@w8�&�j�Z�Y�B^�k2,�*h��
���;}����3 ��S֬�=�`-+��p �e�έ�\����) V�,2`C5̥-���m��k�TR|�ƴ�~S7��'��Ra��J��A�H$c�NEC��3�yB �hȤ���X0d)Y�w�H����}~r���>� t68uYUW��A-� ����%�(ƑO|� �U ���dt7��p��9ARc
]�t�I��"�A� E���e.��5	���c~A��+��|o���v�~z9ƿ�H�Of�h����i���'�i1/T{�`JJ+,g'#״�3A��Q�9L�$e�w�^@��S���𢍋���^u�����P��!aH�!�C[������, ��;K/��kn�X�,/�E����u��-�l�v����V@��o]u&�0pI%]H0p*aSL."D���#��^�Ѫre��@�gLUh�z�s�i`�f^Pq��D#�sq=��I�-�Q&��|Neɐȉ�B3:��gz��E&*`;�ؙ�j^��ga�~�y�֗<'$�Z"����^���i�SW����͢U��S
��e�^O���;�K���+�E<�j�O�D=�롤B�Ĭ����cZ���� H�W�g�G` 6�+���,tN�S��Uz�ɴ��sX�2�Չˮ�2��{;�um��	��*��jV>�-��=wu�>��(j>��Dп��a�<\�[|��4I���,#�M��觖$���R|SK�����#���T��#"�� ^����Ɋ����,~ev�����H�O�����Dnt����@������ſ�A���>$�R��b�?�����Ҡ�?��-:�!��� ����eo�,&��s!S�xȬY`DWq%���K2���t��A���D����R@�f��(�sE��I51��y���z?�:�D���������Κx������?gW�Ŭ���I�U�y��>j��vvH��= X��%8,]���Wٕ]�d{m
���N(�����/�[ ���:԰[�qS}|k��u|��W������I%��
h�y4�S�$�1?���6�-Ϗ?=�%��p�
8aR)j	\�r�����ڟ�c�j`�����<yEQm�i����K"ia�=2D���q���he�@����I@O�mB&����fJ� �$J�v��.���ZDļt |����?�A�#.���T�E�� �ޚ lFF�l���T��n?H[V-#�c� ����jE5��d��Ҁ*I���F:�o����:,}�+�ʀG��f�¹B@]��q��z=vP�}�_k@s ����P���� y���wb��ʌt\ `���c����rn��Uy<�ٛ��>w�;NN�7Y��vM�-C.?�:jKg�T����T�r���@�0 �m`�ݢ�9K/ �]J%��������P�����e]�J�F ��f���EJ����<�y�^��[��2i@��z�[��'��A�R� ��gr1&+ ����Ŧ, �d�'�9�}�Bj
1䋋�{L������?2P�$A��uf@a�!(���m�8��)��iKy�,(X%��Ǝ[pe���U_[�Ya*����4t<�4�B��\����2���@_B$8��E��t, �m�8��h�:�AC8e�������Je=��0�9��D�0�����*����������Y�u�Fk��}�]�^�L-3h����0��nsS�gAS�����~Ўo��B8A����:�8\�G�6#���<�\�J���̣�6@�s�Y+���2��
w�W�5 �y>������+��B~D,Ǿ���ߌ�/M)�u:�ث�]G�)��W ��dm2�)�0.;�I�%����_���K�_Y����n (�ń*��~ќ`^��}<Q���Y��\���9�K�?���{;��,Z�Ğ�f[�Q&階��z�"D������27	e�p�2݇}�<�R�!�	k���~����`��E�V��X�9 l�껱���~���v_C����7hfX�לl����՗3�����x ��Z/mq�fo˖ۤ�9���t30U֪��S �WL6stU���0*bK�;��ڔ�:�	����2U����HJ̍#1h��38y$@�G�`В����ʁ�6���-�`�2��f0�ĸ��9���{6}mTW]LM��ճ����ţ��.z�N]�{���
2@�@
1Bքl� ��I@ŉ�aqpd���$��F�'�{��F�4������<@��KX���6 t��A1��	e��Ri`��	&�T��^�-x�R��:��~���s�v[�֖@�:i��}�Z?a>�E�Ϣn��I�N���3����r�k���iAn��+ ���������Ȱ,�r���Qj
�����7.�b*�1�r��^��OT��6!�?�w
Y9�p<N����i�,���W=����_eYK[����-�Ug��f�1�q�^�Wi!9j��'Xn��C5a�Ǩ/`�N��+� F����ĝ�,�'��z:�+���w��nR�h�@� s�o��P���.O�G��h�i5c\h�r�9��jfU}����0�e2��צa��� �fKn:�2g��f�''z�a]3s���;c`Ւ&�uUr�:�O}gP��ٗm�ې��靆��Be���� `e��۽ �����YfPn��
�O�D���-�hӹűR��/�Y9Y\^R �U�%J��|�p+ek��u-��i�����H� �7�T�]�*�*�������WP��)��d*=�`��t��?��Fu�<�������$@�٥Ս�Ic8BPޑg��d�3t&V�`�W�1�i����W4���]��.�ÜZ��N�c��K%�\
Dk�4OPe�������Q��RG|aI5
��U��0uA%W�Y�)l���X�/�t}K�d�6t�8���*����3v_�ɲ�����ygM�fs�T�?뻝����� �P�ϻ=|��y�r��M��Y��K�h6E�;��/���1�)�0R��鑅uۍ����K�����D2�CD�� 5J��y-�g��-�il���F#ȣ�4�uH�'�/P��k¿$���(����8�e�|'XMLR8���(��3��� �c�beO�`����Y7������W�ۮ�] ���d|�b�h�G�{+��:�:�15)�$�F�e+���glL�2��>C^i���L�BKIn������=�w梮� Y^�r���%�c͟	�f<��b�7]>�oؚmf�A�<rE�OZ�J{q>9�������s������뻛����̊�B�iM�W��K����_u�@e��[����D�΃fX�$���Sa�\����ͪ��2\S���E������hk;&�m!a��Bb6W�W�j</�1KD�`�Us�Y( ��4F��,!NBuCp�)�9?�W�{��̷���qR��d
'���&�RaQ5����&�9XE�U�	^�E�>6̪hhW��2��h��$
 �SZE��f��]pA��ܝD�{ո�]ڔ �{@%Q'�Px�j����.�v��Vހ�z+D��7/o���:n��[�ـ��%k�r�C�_ׁ���u��Q}�U��}�i�@�F�Kr[�_m����_��=͚H(b��U�5�/��<���Y�����r���X��2Z&lo`����R]FY؟�ê�Df���AP��0�! ɾ�$]R�p�eM��2N2�L�+,x�X�Rσ��^R����Wo���pL]wH�BaT���o���#D�����QO�:QM���z05b��f�%4pn	��Ư9$n3r�}\��Ae�`�gB��Y�)�ћ�Jj����d13
SiXk�&�>��ZZdOi��A�0@�W�t��ݔ���*
���l��{��z�`5\Y[ރ�k�܂���Sp*s{U)��ɾ��8��\�(�dR�rZ;���� �^^�,6!@��F%ǐ�`ʵ�����5w,D����S�wS]I����(=ź�u^W�d(�ſ1��!��wooo�z~��鰺CG�eE
az��l*���VѺz[��bK'/�`m�n��0�R�%*ϱ�N�F�R���: Ӽ�v$�β67#��J� ln�h\2�(`�A���\�o��5l�&�@�`$��}��ٿ�5�<s
���%D���7,�,�.�])�9����@T�6�x����R��OK�t���*2�C�֔*�U��@�Aq�������`�����Ɵ���(����)�\��k gq�m��;X���f�j���f�h3� �Dd��Âl�ޮ쁬��4A��c�>8CM���C�������nb���=������w�����?~LYh��f1�(&�s���t��hz��m���cI��m���٨o�`#d���$W�)�h��l���"�v��_� ��ڵ�"��e������]s�]�g�ε
��
��z�*e����{��k�_��L!��Z�{<��4��%p�*��}N0W\SW�%;�TXV���E_��Ɨ�~8i����3��%\P�U(s�g6�3P�v��͕�֓k���8e�ْ��e��*�Z�vnZ��\��g^�&1���#��J��'��򲻈��� ]�{�)R�����^Y2����G�$-gIEmH?�4qV�Ҧ���qx�m�����W��%�8�-~����1��8��ɵmh�k��ݢϙ��5��t1oڂ��n�L�I�W�������v�\������5����J���x�r�:��|s[��f	t�S���=#>' ڠ^�\̽����+��k=���\_-��S��h ���g"\��Y+�<߅Z��0}��z�)�\ޮ\�8�A��S���0��FR��-��G5��>�Z]f�Q|/��6c���G$>�HԀ��Q~�9wi�7O���G_�l�W���8�����Ġ-���i��̲p��j�蚙��e�1-�Bڸ(-�_��6V;bjA��Kl���]����&0�I�aY�\���u?;���l?ܿ����{``yl]�R�U��b���ړk׬�ul�p'w�����r�ء"O��L���v�[r^���;�onT]��k�e�Ȝ��F.�Lc�~n�.AE@<C��͘�~e�fy��&���W���g= SEV�I�M,�*u�X�c�l�������CO˞!�s
��>�4o�טC�������O�t��?�3�2�W����>��d���K��G^�6TI���r�� ԑT޴��,CѝM�@�r?��D���Ձ�Ld�"΁M5?���g>͟���g/\:��n���k�ݿ�Ź�nY���z���P[>�� ��}Y�S�X��`ZM��k@�ާ6� .��xEP����0�E�כ-�{�VR�I��t���4��/����l�Tk��*rmUU , ʳ�$K:ϕ׈g�| .#3���hz
���)�7��;ѹS����^: �d&����}�\I2)K �����j[ɒ��ݐ��p�����A�P��2X`Z�Ѿz�ӎ�ly�%�sނՀ)�8v����)p>�e��cw��g�s��P_�|,F�m���eX��[�A��ڠUK�^����J(Ϝ��_�ck$�B^�n-�)U�pY�Ւ���T�s-C��
����J�3^�}��wA�ϔ�|���:%���.���=�ttp<z�t0�C�dǙ0 �͈���q���_��/�u�^	�y�����d�B�����b9�����t��l���� ��朥@���3�t��C>�;����w���}_�mo�o'�	]�g�e r~�x�{����}�[0��ꆽ���bg���[@��}XUc��j�#�&�n}��Ku)D+�y��{� ���-�������'��[>�lA��F�Z�kI�ǩӞ�6(!��|��x8�1�<¿���SA�b����l{� �3�����@�5̽,~�Z 4�^��=�J��+�R����?E��B���������r�Y�ǩڻ�+� ���ܡ|�Ë�9/`������=^�W+ݝ;�����`:+�lGW����kݗ�j�{)���&Jh��|_�t���[[6��c:��k�D�:>fR�{:�}��:�;l���Q�N��3�c�k���:��k],�x<�C�`�	��&=��S�a�s�R~��ۯ���=/�h���2��i�gY��(��-���Um
�j=���[w����6i�S���E��M���)���V����1��t[��ž���xY"�VT�KUNt�ЎϬ�s?�5��X �*��BU�Q�{�5>�r�VkVε��#ڹ��^�v��m��D2����c��aY�&�N����6M��/��
hC��w�:g�w�ܽ����F�mK�t��v�)f��-����N��%�1�_��ܿ����|�"T)�1|�dĄ��n���[n���eQ^p�[�W�g�fZ�~ʹt���)>�{��R��)������!Mpv��q�C�AS�'�=�\���ʀ}�����V^}V.ͪĮ��B�-h/'�T�*\Y�N��U;)�u��8�<����3��i �C3x�S�[�~���#`x{5>@�P��jJSA�å�.j�ު��Q�p+V� �����F�^܏��CVމ�/�_�J�=</<������������/�fЪ �ʇ�`9]e�Rx@���~��Q^�����(�����E��r�,�=y��UB�ʾ�1)ayQnJr/m/�i�eULɎN+"�sL^R�<g��H
}HO���e����
 �g@K�qjcҖ�Yg��Z�P"��ש?��\��%1s��X��0=�������%�� �)�m���g�����z����ϵ8'Z~��`��Y�|��JW_ߺ��g�Ϯ6�Bp�ƃ�$?��D}�w�h��Ԛ��J�I	\bnn�����we{�;��~Z��y�&�YRw���O~����5=��t�0F����������(�W���d�QWH�t�\�
�㭙
%��=1��O��S,��|��ES?��'W���3E:����=�b嬲���U���s^�u],���ړm�B{U���U�J�8�
h,.[2�s����Q+$8�'W4��s����'}��1��|����w��^f�2�����6&l�-�t坬�����nZ�39� ]�������LLp�݉bB<�|������{H��o_r��4�X�֥���e#��poʦ��Ḯj$9p 
��`�"*aIϲ�6U�[��s��˙r��ZT��?4�!�\���g��uy�̫�0��3��k$�Ix�b>��Mm�n˞
�T�� �}����P���M�~�7�r����]MF����u+�9=�����N�ڷ��o��.�f��bu��K�G-K��b�,�I')�h*-LG9e2	E�-��^8{�-^�^���p��|`o�.�G�ŢY`�6�b����ZԞ;�g����#��'��*_�����f�mm2Vp�bj�(���L����bQ_���jg]S����t����B�3J��x�p}�����oնYO���x�1eֳtZ�X��0���V��sc,ˬ��h�!���e�x�H9MyN�����CH��7^&���`<'C`g��Q����l�841|g`��x1h�:?�>�1�(�6������0�{�|���j+�k[��n��w�~[3�vߝ��,,��y��j���1�w��e�.��3�|~;�PK7J���y��C�������p_=�n�L�� ^��YoZ�è�:M�Za���bq,ޥ�i��6�S�DG��Y��z/�5Ɨ][��N��mu	�@�˙f���G��c����^]�nV��@��h������m�0�P�v��~�U�@s
�c}���T#��^����C�I.��=yif>��[<
�e�X��YE)4���Fg�{S5>-WL_��{?3;[���=����W���O[���Q��|fo��x |��u��/��=�T�Te�\��@�Kچ��sa��׊�/ΐ(�qRu�|��f$B>f«�������7_]��J��lA�r���aô����:������@�E���K�"s+/��Yΰ���|��ɷ*�?�E�?�lռ�_�{�i+�V�P,i�ck�� X����s�쟾�9���]?���>��Y�$޳��Emq���T�C�-��Y,�rY��Re�L-�Z���\t�Ҿ΀�=O䦀i��5wR�c}:sN@�2{]��eqC}7��?iN�C��������S @�(��α���"� ��\� ��b�q��9{"��o�1�K$=4T�e�4���t�H�����Y��#/�9�-�����·���Z�Zc�� �(�)���\s��.�i��q��'u��|�����2�E#kg���}�.�[޻���{��^��d����J`�w*���j�!-��VMq���|y��lFH�и��P|�4x�9��	;����.�C��!�p@��8�qvC���k���|��2��"Q�?�fH�&Bhg�p�ol�"g%�AE��PY�x�El�@*`���s,]d���&P�r�`q�Z�XE�3 Q���/7jL�~��a�s����T��_C��mn u.�WL:�/�s�tv�z�鸶HVG�Ѫ<m,�^����|����{��^\�T���X�<W)b)s�ʜ�DH�}��I�t+�ߦ�9�TR-Eir)dy�ԛ+2S������O2�5��+��>�.�z�y�K|��I�!}���_u�I�d���,����qt���c-RgD�5��l�T���/�s3��Y��"�ˍx˧�{�k l�P!���Wy{�p�5�
���d���<J�l�ri�cھ-��tP�^f{����ٚ��*�ZN[��,ȗ�I�� ���M���ae������G)U��l��Bu�%�%.���ŝW���@-ns�-߫��>��dt��r�ǹU��X�K@Rh����X]؋���Zάʒ���{��������ھ�i3�Ӷ�������ui0]����]�+���a{�`~��?���98�$f�TY 2���m�K��c�]���>��t��p�� �йh5�����)(2�9�[��]h��6�����ܰWWz���}� nIi�hvuI�Ž���*���N�r�]hN2��
 ����!) �	����z-��u?)�K��m��I5�ϫV8s��C�OJ����,���<�j��9����V�,�}En�=��mˏ��r��>��V����jc���e�����¿G����Ț/���K��u�	}�<���jq�@G[��>t�s�4 h_e�~�Qt�`�<l�!=�����0]^t���t�v������0��1}>��2��2/(E"�tF��p��X�ߡ]�2	�7Wz��d;��6�|Q ,�mM'b�U�7֨��FdIg0_��m]�Q:o�E��~�����rV(�ͣ�S�Z�$s���J7"ۤa���g����C@߀�C:�]W�}n�~^�Uг򵕧A�N� ����,��0Y� &�vc�� _�- �I�\��L�Xr.c��f�d�y�ҳ�wp���V����0�$�*�
�r]R���YM_�`�!��%�� �-d��Zش��:j�"SK^�Oߣ�k�h�{�oW�g"8=2�h�n�n�h���vtp=8wӇ����.�����a��/~��@ۼKL��O�I;�un#52ȵ�v?7=��]�l[м�7>z^Ȯ, �0�y)������h[n�9�&,��l
t
\f)cES7���]evf�������;�d������죩l��d쏰�&A���j;q}{�0�H|�Zt�E���R�PS�ꡆ?eF%��T~_��5�6h9���;!8���0�d�\����x�;W�S[U5H@-K1�s�ʒW����w�j%�
n�g/�G��"�NAU-�)'Y!��!&Da��[��_�����x�3?��Zt3lGԴd��;��s,�3�������n�3��G��{���L����h �'dצh�6�i��%����ց��\�����J�PvT��j�^���V��F%��Wi�+y�̗�.���
 iO(�ʁp�faV&eL�){�nQVcr������N�v|I�:-�%[����W?�/z[2[��Y���ǚ���4c^V�p�F����z��"ȥ�:آ�\��֤��W6V}j}�c U�^�p��o�;�&��]ֵ�5��*�B���hJ%�^�~�0`g ��:S�a'V$�Ŭ ��x2.�B_�!�����2���J�����ͤ���IɞH�h�~rG�ciC�G���E���Q9ߺ8�a��7���o�ED��j2��_���]���<
�K,x�#ǁ�%;+�ϒ��9�P��Uʴ
3����q �KO���f�E�ўP�6 ����T��\�n_ُ�4[���.WǢx3S�����l�}�2������9�+E^�>7�W`ǀ*)�qQ<t!`g�x}[o��,��S�d�Bi/
�JZ������iuS�G���{� W6���ꙍIZ\ywSL�j���E�J{��ie����Oה[��2y-D'�eж[9�Z��ˎgi�r��U�n)������=���� W��� ��^ۺB�~U\����̏�0!gU��@p?x�����0t!����#2���R�<g��1�~J���TM�l/��� ��}��.ڀVfT���(�+81pГڲFY�^.�K��A��1Vb�M�҇Z������mV��?S�m hfl[��#r-���Z�b��f�S^�i,(�2� ����I�q���ʳ\�&>�� ��A�uסg1��dr�ϳ\���i)H}������_ ��qj@�����ҵ}��, O\jG5m���k�V���6�ʲ}�PMy��S�¯m�& �E�$���g�
�vܫ�B0��D�[s���\�5�*������WB��]ӛ�o�o�$�R%�E-��(amx.��;��}H���6}��;�{:w��G1�}7�o>}=�m{%>�a�����ɰ+3Gk�b7���WF�}gP��*��i�&��0�
4f&����F���L�\��P�u�tUpFQYC��C-�F��$� >�_A�1�j���Ņ�5|�\����Fpm���50�LـIA�Z>s  �ԗY Y�h8��q���$�)����S���f�a���g�Y�\�*�~�\:�=��Wjۿ�&���
 K4������~�yG˘k�ȱ�����e��3�L��E�K,��W]�&4�g��z��*�;����sPȲ��(3ݚ~ �����:Gy�&+�~����kLjf�z����w����O������f�p�&�m�b3���^��70�;`��˳���Ut�� ��U � 4�X;�@#"f� ��t��ڍ�ж�7;��л
[9qՑ� ��F�u���}}s��b��Dm'���4@pZ?2)ݞ%���rR�+ ,~;	l%��]Ncʒ���4��_�	��7K��V��6Yn�g� c"��������#4Z�D�op�� hj6����4e3�) �(0T ��6���U�k�
�'zZ_7@�(�|��i�-� ���1�'��Ɨ�>[ٛ�pZF5�w��E���0*���/����͗���������n:�s�p�����~�`�������t� �Tޣ��n�Z�sW��iQj���Vh|`��8�%%�k���W�)@�4 ��L{X��e�+V��z�F������z�bI�rR�u���<WC ح�*��),�P� �TM�����3sq�?0�Rݝ��/�?�Nk�K���Gg�?�i�C�������R	J��I�cJ����j>���;A�	N�U;�O&)��do���(����ԽK�LHq{J'���Ű��W%׳f��<���K�{��z���>�a<��d퐀�ع���	 #����������7=��>�^~��nܦ�}�_}��6��1�X?��^�̍�����,:��L�F�U3*�＄��i�<X^~���x9�lEV��҆��V��oP�&�S�&e���!%vi�eg)a(M�qq5��@=:�_����f����91�/�A7?wH�a�b���+2S�#Lj��q�,�2h}ߦ������۴mm�f �N-:�4�)��΂����Z~�iΓO.�X!�t����ZV��������2l,/lfs��@�r'��i!N���i�R�emBW	a��V=����(pF��݌��Kq�e���7��Y C��EHSx�O��1�N�+���3j�֜T`���a�E�[U�'�)�B�B*�6���S�3X�(3[�Ą��iT>���_�Y<���A���n�P���%1�HN�����L.�K��7}#xK��9�S�(�`�1���X�i u�uj�)��Aq�+5.�u�'診&�^�e`KiqѢ �����,��F
oT�5w�ڨy�v0����DV*���mt�R�����+K�s)��p��Ȅ9���M� w��v�֨7�O�< 9<�-g��({g1�&��MrU��C5�=ºk6��*U߽�P�"u�$�]�0����5^��	ns��p{�~��f;�����W�������/Cv�R`�����P�ؒ�X���yyR�&>�)�c��r��Ia ,����:g��u`O�B�=�E������h��U{�k?�"�(��X�����$�ڗD��ʜf��!7M��5TF��  �ZuN�o���d���f!����e�q)�U���j􇂚uX�a���]�<�%��9���0�A$��Z Zsܮ])Xg�oAP/noU������Us�ɵ�I�Y���@�q�R_zog��N�)�Uq80��1��[=Ǥ�º/��	�_M�_'�������7��	���B�K�_c�]�>��q���������������9���| ��KӁtG���N���TI����ѓ��bS�^w���)�峟���ǽ{ rfE��S�3����4ɲ9Zͯ���b�v0s�_9���{X�S^���@�L	lp�D�[���r?Q���Δ9���xY�A:��̤7(��|���=m,�<�� \� �8 w�\o���%{	��s�Q�e�,$}��M�2������)�g�v��J�[XO5��5I|�;v�����L�����X���=9�$(3�J�@�B���&��Πq^e������ ��R�1l�Ĥ�z�/^u��l�uڨYFER�Om{gP�����z-7ʙdzBó����e��P�����uy�;�߾xc�����u?�^: ���9�>�c~~G�D��i�J��i ]�i�y��ӎ�Q9U�Fc5�Z����<��L0Ioa�C ��>�pV�̎[��΋O,�hg�U鸻μ�)�V��4&�C���؂E.��A�uV�aq��$&�T�t��Pޜr�@uk�(��,5i(��Q��>-c��L3t�Q����؏(!��r�I.$<��K�١���QY����km��*��Z1�.�;���� vo���t������3M\nv�2)�X8皀�j��T�T���ԗ�?]�*	_�
4����׺5�ɍߵQ�ef}�0K3��6!t�?�J��C�\el��fBe��b��9�@����Ւ�ܐ,u��W>K���Rƺ��I�h��u��5�{�����S\t��i{� H�`�ٞs~��z�ʘp�I҄5�3u̳�;�'2�,�N�7��j�5�V4� ��OFq��Q` ����B�#x�؈�$�m�ȋ8+��D��r�cd�&�W:�L�=ɕ�A;rP�S,�/
�e˂�2I�H6<i�(�$�5ys�RN�B�(&�	c�.3j�^�9�A��85����K���%%@PDJ�g��a���EU�ÞX܀UKM�S�|}\m~-1ΨZ3R�ءB�+������|�sV�f�*t�q�B�#���r�nk�Ƥ/�Y֎�1���s�h�)E�%�\�l�8/|C����0��1�^�L*�)�uPu��8 %�qO� f
͗f2P�v�Y�u-P2�n��°�14�\t����@���KǬ�f�?]w���v�7܎��!O�xH�����%�t �Ʒ���'ۈ����v���]؏!N��,����BNJ�p%ڜ�!}��� ����>�"v����t
��,�G|��y�拱���1�0܌&^f�4�pB!�����-���w�UfS2�e4��4��J��N�n���H� �(�W�̰5T��fYb��H�h���.��Ó���$�j�3�JBF-�#>v�D�<M�t��֧ٱ2�&�|��{��)��yY��~6��#�]<X��9��;<;T
n�J"�����L鳔9qu�2��%��tB�+j�+I�X�Ʀ�U���$.�_���J�4��1�f�
��CmV�?�_�dY��T��uԜ� �:y@�cz�d�!�G)�;D��
�a��0ҙF�g���+a�c]_��t�9i0��IZ��-��͜g���t���� /4I��#���P��j��J�����8  �����v�7}�߅9�D?���O �����>�>>�c;����8<{t9��t5�L4rD����J��L i�毅���A�d%�<Bg'�g٥�,�&��m��{9n���RUW����w����L�4���-�f�3��y���bz;쁞���
w�"=d���P�ө�@����Ǿ���K�ɻ��L��i9�@�gr
�	��M�G+J'qm�g���C�Ph�5:ҞL̝�DHCt2"��ԩ�"9?�#���f69O9�"R��[��ą#�s^z�������C-��|1zq���S�d���J1�0w>���L%	aC'�M����ס5���sD�����
3���Хy�]F�'%w^#����������L��)��Ni���b���6UD�v�ߜe{#a�	����ޟ�2PyȖ_,d6?�r'j4��uN�ߣ�YTNg��$��@!Jb�� #v���x%���B�~��B���Et�׶�óo��h`;}��`Qb�ޑ��L���������z��Erwh�v��8��8�������/���[�a�c�����'o=y���v��S����f�����t/3m�U�J�BYf�]$s6���f�IJ�w8B@�W~�.z�)57�Lm�m���������ko�ɂw���ٳgpC x8�4ϻ�4��0��O�#��	��*vh�S\aP�1 �,� k�&�</���C�V�|��O����7B�w=>�K�Z������ԡ�w(t���Q�3�]c��]�uK�(A'�Aػ|�jO<Ƈ$HR%P��%|�y#鈊���ާ&!��q��;X�<���<�"B�H񃚾	_�a�%S��G�DM3��~��c,�h���"�f��Q�a��Տ�i�>�ϩ�i���L�̔��<�����x<^��l�{|Y�H	�>>v}���Ϭ6,� +PBC$�H�}~K�AP�4�#������6�vR�d�����B�"�@�&NS�4q*23�/�Pg��QZV7�l�+=^��i�������h X�u�eu�_:Y�gH�5�J�Q 6
�3pW�hZ^���NX�yYI>�55������C-�M�[,�]���+�`�'��� _����1��:�����r���r���0�ww
�t�=d��9`3a]���ͣn�H�s`�(�z��J[�(���QZ�?r�y@a�w���hx&A��UD�w��;o���͑���=|z����#��vp8N�)��;���x��I�_�����4
ք&!iK�ݞ�!q�����"�IĘ�� �x��sH31:?��8��zB3��z!�0{�q�&z��}L�pr',����܄�l;<�!���c�BX^��a�� qH΢x���xЈ��N;0BY<��L��k;��?��fNHc 2󆽇Q��.�z�n�0�d{V����Ǽ�?>L���oI��C`#�!yM�o�8#�Ƿ��~3]^n���ED��G'w��ݮw���&��"���e"���^s�����1��'~��x,�3���$Z��( �2V(�gαC���ʉ(����~d�d�$���W�q����d�"*,eJ�x`�J���L:	�y@��mx�������%��$��t�=�'�Zwd���c�L�%�����2C3�W2�n� ,*B�0;в��������Y��v��?o������m/ ��}��u��q�t?l~u���G��v�o`?�����ɏS���9�RG�_ ����&D1���+��89��M��*��D;X�F���8�d�%��v��=����|�IG�v�[6�=際�� ���G�y������.�a`�"ۡ��~E;�݈r�2\����#���/��9����.<�2k�c�Ds<+ǹu�8�H'�a:��葈bgC����S�@���nO�I�'�b;	�Qr"��8�9��؅�C@���/��9Fb)q��G{�d�& C@�K������v���q�bS2��$�?.��%b|�8���l�{5��������O�����ۧ�X '��b�'����,I�1b���v;m�m�d�HEg�j�1����f�����Xwy�w�L#��@�M��?O)MP��Z�]ϳiP�"I� ��:�m��B[�L

��b���c#����et
�|�B���.c{3�F����i�*�e2�3p���n�w�'����O3[/�ꨏ�Ds��(@q����3g���W��.s3��,I�W
��P���T��=/w�I��x����#V�>��.��f3����|����������g�K��ʮ�n���M>}���W�ؐ��z{��
����c��ϰ�On���a��'��L�9�
��}fOJC���.��C��nb� ������H�({#��� ��Qr�&� ����$9�������Ǜw���ܸG�Ox�����1��n�<�Wj��ww��?��]~���rx�vx�n>�-h�S*q�;��D!{��C뢃C�q��w�e0!�L���́<E�ky�ۈ:���v5�np�rdy�_C�7��}� ��W�#f�_�1�Q�h����=?�#O�u@��CI~'A����M�� �����ݧl�:	� ��s2{7����6pyy	ۋK"X�p8v��v���g������	$�!���1#a��^i���M$c�b�hf?!	q�u�E���lP���x{w���ݔ�����d�� � �YO&�@��K��q�aHϐ �:����/�ߘx:Vj�����*�x�<i�sv��,q��ԉ�n���B|�v'c����!���M�Hn����@�Aq�9�{�nv�(��0�� {��8��)q�Y�8�L��
����F��NMf8�g4w)Akz�//6�G6����4�ĩ�Q����!�Ѡg؄���8����9���K�`���x�?_c�	�s��i�~�gw��[|o��ͻ����0_!r\�y������"���i�Ѭ�^��d���?�t$��Y�e��@�:/&0}P��f��A;��J�0o!�w��Ӻ%(qG���G�O`𰇃���xx�9|���;�n[��������� �}���ܣm���w��Gf����ݷ�Er��Yn`����_�~���~z�>�\u���<`���!lQwdT��-���gw$��g�&~@��<t��%Y01C�[�aCN�4�#�;�w��Pw��>#Ὕ�S�W���Ra>���[0<���t�N��[���%ƺ@\��!{��;M�@�"�˟F
i����b�1��ǏG�z|�&��x@����]���K|�O?�v���w���f��.�eaD�w{9g��S�D��[� |�^����ݡYpy�7�U�x�i��lT~�@d��qp@��а#x����>��z�����u(���(����4H�aiB�tD��|7�=6ѐ�ͱ�C&{r�bYdEڋ�HQ��v\�����0�,��36o�wX1��pw{����i�����q�B�R��t�Q��z�DA�	v��Lal/�? ��"+�9��uDB�)2Yq�E<�X�G�e����&��������H*B���O.��M}���p��(������\��8�ݷ_o�G�K@q{��'���ŧ?����V�7Hc:���]|�&���7�k4�ތ1?��#4%.P�j@�!���t�)O��:XLa1��أ&ޢ
��	���G���&�)�i���$����dd<����;ȑ�0dz��~��~�/���~�9���t����q�w!mf���:\co��0�G�d蟰��b�h��0�����;82ձg���ko]����.�1�����6�����<ï�y���!m��2�5��&2d=b��G��"*�������,�Ð���n�?�>���cG�wWn��+������"|�����0��7�*f��@\D��o2�m�<&�~�?��f��"��e�ǹχG!_�o��nB�>т~g�v���	��~�@�)��?F��!�LD�ю%���ɾ�o�҆W�P�En�x."�EU�������k�e��7ô��Uu���ot}7���f�e-g�|Y���'���6��~���<�`�`x�ٗ>��:p<��sD�=*:7 �B���	�zd7��W�!?Bz��&�@'7�����x��!���G4\����g]�я~��{��g{U��obs>�>l�?FtA�t6���5�����0�5���.OOB���m�9�FEN&�j"Q�a�D^c�Zr$4y/д�[J���p9tφ��KG<�@���-I�D�LjI���x�8A	j�o�H?����;��|��~2;��+���;x�W�>u��߲��' ӗ<y���-<f�ʟ�[�p���|#����N��{��L �W��?�~��_�9���%7���s�����9���h��(9�	����{�,=	3� >z����.��~���|��~�~𣳹�^��`>��o������Ʒ�@���k�� �}����#��;��Q�	��������ã����������
��0n�Q�~<2�ݼ��Ȁ�0��O>v��"���}�`�ɍ�_=�������Ƨh^w�F�	W=�H�a��6�]  ��ӷ�f���]^���H.�Y9��8B� Fn/��a��y�����0�����Ц�s>d�v�"�'nL�p�Sz?�{u�c�`�#M�1oPV.7CF����Mv&�Th�x�u�Yp�t�vq���>������� m�,̳��$]��:l�x}��ǘ��Ÿ�C�i����͉�c��/�����y�)� L.f�:�ȑO!G9O�g�"�%"WW].C�#��� ��*�A��Nn4��;��E6H�/����VA-��f#��7��c]��Uoｄ{ ��aw�R�Q��@cR(4,ڑ5�Vg��^`�9�'O��3v���W��~�!��׿Q��7ry�O���U|-��=���~G���]|MЎ��O@|Y�ƍ��f�����G�8{�x���P�R��Ǽ'k�R�I�F":!�?bo׻#���aB�i���8�q��t�ܴ��w7]<<ax:���&>�?t�fz��"�����g�ff0~M?�	����c�G�~r���g������)��8"}vO{�.��A��#^)v4$�;��8{dD�d:�4�����W����Q!E�d`'� �/Es��M����#G�x�`�*k3t�)�yNB.���b�	~�}���£L��T�3OI�T]If=2�0{萙�X�C����`8����|m�X�뼑R��_���/��(>�����}��d]�}v��h+�%���F�DZ}�f��RSd�w%Q=�s<�A����h0��q��g���]@c
yD���{��`U��$z<�>����1�	��k:�ތ!}�u���O>�������v��^���m�����������'�����1������[Wwۻ����p��yN�a��6�(ā���:�;?��v7��>}�������w�dy�9��(Q7�G
_��C�kN�=O/�	�=�/������r�e�����q�|����'��Q�&��k컧Pbߎ�	��Tǳ
�hJ���m������"x���F��B{�Gs�m�����|��GV���Z�~#sww=��a@�ޥc��n�i~���{�;T��臑b7a4��㠦���s>��x��~������|�?�ճ>Ow�Ozo����g�����G�G��ǐC��;{���p�=B��W[����Æ�)��4��րfPj�8l�F���ҭΔ���p���E���/8��)��tg��@/��^��&��؇�u���������X~��pC
i<XB�h�����J<�s	��@,�ef�(� '�u���>����GaS?/L�$�����'��FV,=2��N����<  �y:�<�{?��?���y�2S]�4J8��/Ҝ`�b������v���D�=C���O�]�u����G��ڇ����#t���������t��wwW�|��=����^w|�͏�M��� �k������Qӽ�]�Ξ��͓?��xof_ǶJB�]@`ǩ�����v�Y�c㝿���^�����_�_���y�^�-��4q�,f}zX�i"R6T��x�(�ؓ�L��|�����/�"E1�5ƣ�8��Q�S<�j}�\�*�ýێ�b���}��~�v;�_��?�|�vT@C�Y.�4�ѥ�fYQ@奉C�'n�:���?"�<^p�O.G�|�ۻ�wx�<���� p��?�S���d�~�vo~/?ſn�&��}:�����I��ß:�Cdto=)�O��PO��|8��z���&��wZ��H1}�k�p�e����)l#��\��=��>�8���FMh�-M�q�`5���\*��xe���v{x�&R졃�f�Qc���-\=��$��.���g>��ct7�|#���BD����0ś�1~�;�_�Ŀ��hץ)���'���C
�݄.]v�|1���sq�`������/�v���<�]M���{�ڏ���e�2�<��=�y�����s���|֣�53�52Fa�� X�0fm#���b��A�űA�/����mc�Ɔv�e�c��b,VB�!$k$4I3�я��͓'O���{��Π)��s]��}'Lv�7O�<�?~O�#/(��{/·�ٚ6�23�m���33�lf(?�>2�rw�'F�=t3�YZ�٫�W�Ā��M�,w���S<�>���2�M�EP�!r)o���F7����C'�CB'n�Υ��{�����9ѣ" ө��q
;'��n���Ya_,L����ky������̫��j���*���H�jo��,�a�3L�azL�{����ww��3GN��w����O<ћ/�=@&��L]vR����}ޖ�C���/����+�RY�e)mΥ�|]��'��3�E7eY�%��33_I��̸fc��mؚ%�H�S���J��e,�]gs��*g���4��#����|<�;�3����m�)#��t�SS��g�94o_���U�祝~o`��F;�s�%��q���)8u�bVd����n:���G8�.��;K����*ݿd��rr�����������ߴ���'���	So�Q}4��_�[�.��%\���>�d�FC/�9�k�fR
/��� ���=���1��t�6_���"񥘸\ST���N�Ǐ������4��s?���%���_tR/���H���/ӣ�x�������^���r[�/����<������=�||���hZ��v'���o.���������,^�����/ډ?��/�G������?N/@ o+�R4(|~/9�}]"ʒ��WC�5('�Yt9g)���s`�c_BW��&OA~C�:S� �����D<���`S0�fT�,W��@jV���gP���@�h}�?_S�ԭ�b��W���ۨC�9mh�{�=������ƿ}%>�����v�nm��O��~�������;��ʕ�+�L��{p��E���||� �ϷU�&�a����f�ŕ�\���g�ٌ�CC 7!45�HC|���M�����p��n��"Hd�N������:��P�>t.�}���Ǚ"#����0�b�[��tD�׾���?T���I���U� r�k��#��U�
�
7���3��&�Ng�ګ��V�}�N[�;��Y�[H�I�.����੫BZ�v8���񋭻���U�����UŖ!�!��'�M���j�䞇�
��gV��N���6*���>��+MC����2��x�wL/͑��>Y�4]�_��D�$��'I}I����{O>�d���|f��(�����R�R��Tg����Ǘ	[a�gB�j�U����P�;��m��7S۲�~�{RPY���7F�H<���h���2t�>Q3&���LlaW�lЌ�Be�/���/������l�}d^V_�U��󲸏��J��<�����-�U%%��z�K���؀@�����2	�]�[���aL-~�$��SPz$�0��2=;��c� ���X���fs�H�Sߢѻ'����}��#�\��<���|0���N�sc���b'i�
��SW�Ъw��NGD{n'S�E�xQ�/Z�.n�0BE�`U���9]1��e�DlB�MT����OU�l��P�����[��m�mp'�	�͎[P�q��]�N����������|6�Q[�M/���e�8���ɖ��A��܈Z4�!X_}[��	x(��A>y��i��[�Ő*�/���M�H��%���K��j��h�k�A��r���_ts҉0��Q��l��@��i�)X��-�ٗjy�E"��7�B�y+��X�-��=N�
�Y��J��|l���e���i�u;�Z������V ۈ r����/�E����CB����Z� j�Xօ�`ʐ���Np�ؗ��-�`R�bUP[cwS�"�����w�ώ���l����E���x���#$�0��"�����0�����5�{_]�zRg��Ò,K���U��lF�<ȷ����z̿�-�����~�C����QNw�<�K��w��S������W�jz+������!�d|��'�n9�r����q��<d'�Z$�̕+Wҏ��#7�w�L��J[��kI��Dt�q�}���-y~��z[8����n�/[2m�{��S�?�n��(�2؀��
�� %"�>�~�,��Ū��У
V�M��pr����b|���[P>�F�aU��ln�b[��!έ;�"I3ӈG�8{Z��95�@�����H� S3__�2��ݬ�Ih'm�s�S�J���D��@o�h� o��`�O�w,s�`���E��$��>#�!<�.A W���ȍ�G���m�z<��{�T��ݠ�ϬaW�[9X'����v5�%����ZdL� r>����|�����2F��mk�o�{�O�l����xz)�:��!>�>M�_���$����	�[��f�N87Ι���Y��ۈ=�W���f�#��w?ơ8�d��:��UȲ�^�bM>x�9b�K�w�h<��H}����p������?~��_3��������GM"������s9)�5uby�s�n\܍+�3�6b23�Hȱ��a>��6׆F-����C7�e��Au��Q�m'~���� *ǼR񏓓I��X�>�h�[d�"�C_ʲjd�H���ȁG�f?�;������EAm1K�CX�N���Y|Tvɲu7�t"냬rz���2X�1K����8d�����ފ�rQ)���*.�X���N#�c�Ez'���ȋ3�U�މ���ş���W��u�o8�JI�����i����O{�1�b�H���>|��<η�յ��,�xSen�E 9LZR����e�h�!�(~����N��,�V�S?�e�����ZA��N ���� ��&�B�N�^@��,�����/e��Gy��5�V��*�kщ;��_��zu\�;�{���B��&�EMmX@�P5	c>/�g�0�d��5�2J�A/P��EO�x�s�e;\�s�Fpw�@���0f>�{g�ԡ#a#����ɱ��ԝ���Y�^:k�
�*���;nvR�VؐO��:�@���od����G�;��tx��@B�V>�e�˫^^o6�!�)��F"�����r	&_V1Js��������۲����;��yHT�5Q��h����룑Mz'�tc�F#�m��uˠ�ɒ�������0>!��[1��*��(yk�׀u!�J�'�[�fSU�.V�dCo�ܕ����[/EY�ҙ�����V�d��%�=��e1rPJ� �ψ�7;���+/�ż�Ekah/�;t[�ws��]�ub�:�����]�sP�_*v�Ib��f��v5�&�
?%�+�FI29���#�>��pYU������4y���a�/����C��a��@��[�9�m������ ����,�o�{ttt݉�n2�R5�H�qu�Ti��7d�3�_7`M$�<Ib|����]�"h�l��	?�?���_��򹓓��,r�oV�xq�m���fAe��P���ݕͰn�;|衇&W�\��'?�I�n���/���З-��1-N���~Z�
�NҴD>ꆐ�'�7���4���bRi�X�^��t��`��xi��G>����ЁlS|z�e��\��uOh��l�����j`�)|Y���:2�I��pX���Q�,>KW=��<��UuH �ҷ!<��I�^�����TF���Y-�җV,ߝ��E�g.x�L���lfK����½i�`�>�*mG��l]��gtET����R-P@� T�O|}���G�o��.��*Į�2o����s��ނ��Y8RmSNx��{��+pKm��[h���~���3�|v�e�oC��>ױ���.��ئ�H��ė�{|�G$���%T�4���8^��oCV��L�m:È���0)g56���X��j�N�K�����T�Zb�p0.�l!fH�뤷H~?n�Ox����()Y,�I�ǭ/:�m@I7T��΋�<�iVy��gC�L�R�7��H�9�w�(Mjc�^�ε���N����T8��-��H�gd��OOzH�3!~^)�~�<�XA����a�*�%2�=�"�-o��
�dy]oQ�3J�,ƚ<����A�=,�n�E注}��c�D0��2��Q�_��p��,��.���w�n��1�`Y��I�J�g�@ �������4�[-'�Ҵ���k����P0�(nXr����)�|���8���]�mb�-rF���#�[����-n�}P��nw�q� Wƈ�or�&	��A�+���6,nWg9	.�2e�s�O�)�34�g
_��]���c,�Y�I�� H��:D`��
 �Z:�k��P���p�&GnP�{�"f3�� A�v�/��K�Uz�Z��7�V�Kp�=���x��~�g8:>��<v�|j!�ȳ�/
��IA.	�Z<��
 QS�F��'��*{/��"Xқ"v��֌P�M�햊�	�����1�g���f���g�yfǍ��v/�������Nf>���0Rp3mm�$��G���;�<`�L�ߏ!:� �����`���?��k��ֻ�΋�h�W:	��M��$��6�h���ޔ̋��,���xm��H�ꬅ�ni:�F��|�P�����ƍ������҉;�RR9|?�|ѸR�T�$4� mz'�;;;�x�����/����_�1P�4,t�%I|S�t8,��[]�߬�'�j҅toob��
}̪j�*�]nx/%	Yv�oޕ�^ �$�"�a/���@��O\�C�ϵM�p4���*�� �˭���{h_?�7W��'f�:��M� � '���Ge�(��h��ȴ}��]Ptd:/ͼ,�T��p���^�Hmj`�VN�i�K+X
Mz'�E1�Ӽ��n���~I>�A�Oq������%�L����P?���ea��a�{�j����MM�zж���Xg��)0�X���T�1!�=k$H���+�H�Ќݗ\�zga�C�7R��%�]5���E*���Vן�-�^�}����ͼ��=W�������py����~ps)/�޿�B��� ��N �=B��e�;?e*-�U}B�D��:
���aYS�c�ǹ���p6b�qS/�0�a�^8z��x
���	�_7��Hˢ01� 1��/V%���:Wl�l��$���H����~..p62L�p��.E>�6q�-W��툎�u�}�p:�"�E?��v������J�t�ƶ�G��[U�'��皗L�e�r�`GI�^R�o�ce��#i�i(5���׾��Y��/�� -z'�t���!��������T�k�
�������D�_��H�)0}���`��w�\�I�nǧ�\�K_e��� �����t�՛7o�hgg�؀�@�����[�.&���W�CS��tg8p~������3C�NA$��o��g)� e0/���_�C�?%�2�~��I$�u*�Ds���.]����}�sptw�C���N�X��D��"t����t$#��X��S	����Y���\�r%������K/�t���G��r��%�u�j���YZn#W�!��˘����s��s	��D�x����<��t�C4u~#��PY��Yi���(v�+Fs�_���&�����+���˗/�ɗ����k�<88����ѧ�x_��v�������ϒ�aR���:��y3D�T��bw4�#��;��I��}/�5
z�����nz)���<%R&|�/Y�8җO��<*��dyͽ�'�o����{�x�28��W���������Ϻ�^��WU�q�|:ɾ*����S!�5�9��@
Ĩ�\�b$��"�<��#G���N �"��L��_�$p��������fgg׋d�.����K�.���>5`%�͔��Ǎ�G����O7�����+�xG�ɼ/���9�����R�Lr��X:��;H�h�� 3q_l:���V��z�<�.���]oJ�h�������7�����WՁ�]���8���P��d����k<�K������1�,��*R��v7�dI8 I�ߤu�s�L������Z��,ǽmA&u[Z��Q%Ղ��û�Ge��>�p0"mc�rz(�c��R�g��!C�L�)�T{��s���Mټ9����0��a��w��$'�ny)��§aΓ�ze����&Ty>�!ߚt���� �prˮ��Q�ŐO0�E����5�G�У+�}>ҁ[DlR�m@��q�?�� z_w���3SRxL�C�e�P '����SG��-+�f�3�"([��p��4bE<M�����~-!�F�'��qs4I���7��NmR�	�`.����� �
��p�}bl��
`}3���Ր&	�~M��i� 8t}��5|~��寴�i�k��9t�/���䞿vtt�D��s��}�]�����l���|�?7��X���N����nC�`����H� 7�bP�*�C�� �P������6�r,(��*x��rI�.N6b׶ �����?-������S�j����n����T�٪�L�.��}�C��˭��[�h) B�H󜿣�� \N�p
�6rW�L
�G#��բq"�9��!iY���\�KO�u��4��7W�x��/]s��R�k趾�����p}�����%�_I����*E>��R��������	����C���)A�|���IhD��P�=��9�*�LF�@h�nR��r>�E����t>���-�$�%��e!��o�Q�mcz'���X�������vs����7`^ߔ��`Z�R��}ҮE��L}���ͺ��ۭ�6��f�4獮���\�tú�/���F���,�wH�H֝X{�|�R�9�N�PJ�ӓ�@&��4N�酄��J�7z�?p6���O2���q���+ֶ�e����!����ђ�罔�� 5E�i���h�YЪ8���$T�����FО�j��%!�#Xx���T�j��_(K��,gפ����*;T+d6q �awPk������@ ��?T���<�~:hT'�S9,-�`3�!���jM�>!�X�%� ,���R�ڷꃠ��W6��1�@Պ�+�M��O��\��'E��{�oʚ$i�P��!�؂ǜ�`Z�g�`];N:�����z��c�U��tH�_@����Dr���z�DE�Xڢt���G���,�g�u�p=!��Y���&$�7���='K�n��%����M��_�1��ׇM]�t$�!�i��a�Bp��)sdqc���	�O�s�}~�,�	$\I7mK�D��sR{���<9h[��'h�a�F5g����� �c %�k0�p�D�?���u�Kz����۝e�N �+U�)C�Ȋ'�.����|POnJ.Ч����>�t`�±�Y���i���i������{�3�y���r*,����<;�D�y�<xx�v�K� �M���{b���k&!1��o����7G����c6��Q����|P���]T)^F1����E!�6�:�;7ץ�=�R�/��꾏��o��J�3�ׯ_���?'�z(��	S_4���W�$��B��� ��y�䠍�Rd6��v����������&�Dk����<>i��$�:gqK%�5	��y�ź����q>x;d�x��Z�Bo��Y����I<�TH5�E�'�ؽzy2���믿���˗�ܕ+�[,ʱ�� ��^�ӧ�M ��φ���"^x�K��������,�da�&�;�p:�@"���2�1Z!1�~���}n�<�$U��������53`%��NS6iX}]�����F�#�b:!���|�(�*=B�5U�,D��7�3�tz(��;Z\�t��]�K�0_�e7G��>��.j���� ��ĤŒWI�H�N��"��ՠm.��Y�=i�B}���x�1u9�P�n��:�
�r�D0�^Cij���,�w��ޛo��Ԑ5� _|�p]a�;��/�����,�p��֟T���b]K.v�a�W����3��M� �s	����t�z��������w�!���4�'��~�Lyk7Hjv��OVو��O�9��}�����r��P�\�|k�¿+�{��3-{_N˄Ah�ِ�M���y>���է˲�H��2����'��A�g#m�+��;3�lN=�)����W?7�\&\�x6��.?Q�C3��ڛ��w�"gqxh�vv�'ݐ���O�����Bv���Tm1�n*�gL;����ol���Ű�u>K���9~ǀ�� RLg�T��kZ��?%Z���/Ngg���MxO����{���ζ�>�m���Ҙ�0`	�oL�]�y��l���9�%�A��i%z(�1�I�ٲ�[�>��P�g
�7�4���WU�ٲz����=.>=�×���*�q^��.����*�ϴ)��Ui�k8�^
 ����o�2��a�npnr]����U����`�O&��+�e�u�_[��[�NgQR�K��NR9�?V�!(<F���[��!g�[��P�I�L��ߛV�3�^s���4�>�������1�+����@)���b���ߟ������^º�·K�f��Φw�;������A��.Ӟ�tk�����ϻ� Q|M����C�f����ΘtS�hL��Ƹ?ZJ����C�p�����֢�
�N �j�ͧ-�V?Zu�v�����3��[Y6��B��NZ�GE�J�t�$����,�g{�F�{��^N�B_��`�J_Y
��=��?�Rq&d����
�`g�����m���qH����,�Hv�;)ޏݿ�NF����׋���o��$reV�a>�-@q�P(=&iR[�d�|a0g�k�W�
��-k��یE�Ϫ��y �+@��eY��l���ދ��wω��+�b�y��]�Z��R�\�\�F�t�-rX٭��æU� jK����0�F�9�r~ץ��#��5�/�����|~6;���~��S!�_��R�/���A�~T�vV����@�z(��C�g�[lW� �&�4�"|�%V�,�c&۬JZd6?���a�PQ�P����Ȑ���M�my�`���� RC$�	���q3������S�"�ɂ�I��$$&���1n�����볊�������dv�M�B�+)�K�V��_E8I�a�c�Vu�z���ш����O����Ή�2�E$�J��n]�	�J\t�c7M�C��p��]_珳?h�K�^ +[��a��)D*y+����
�@�|�����*��X)9M��qk1E�e��5�A�����9�Ot��l��+/�3}{�ȱ-?t2)v�t=@0��R��O$q�)�m��P �"�Ԣk: ���d�p��p�:~�"׶���7�Җ���<���g���	;9ylr2�����[xR�/��^���4��t�Cd�$Uϓ�?BW��Ϡk`�zD�ӏZ͂��j������r��cY�>���}}���*�+~A.������W������j�P�m�F�֨�,�uY�띖��\�ՙN�i���4��N�F4oi�B�@�o{��%�o[.�DZh��*�@Ϣ�ȴo�����4nB���-/�=�Ϗ?(�E��l��
l�s#���4���� R�A�yj���V���E�����k ��$p:�3*��Y��'�R���tI�H�7�W��HTul������e���XS+p38�h1�ˌU���s*''�pBW�R-�q���Uй��៵п� R9,`���9��O[���E�\�����J�A����[��\�>���	":��,���~۟�mn����:�����CI�t�M���r�&`��U��e��s��������կ"
!ݴ�1;q�W��V�(}\���ѡ{<�H�pt�1��^�ڷ���\�����卢@E���
,��u���e��X�Ū0��"HFK��JHO9��\�;��¨a��~�=~���%g�����T �%��
��>@�ZN�C��MH�t�Х�ڮ����np�Oьn�8��&<�7̓���<<km����y�� j.�A�Pr��&lW|n���<����e�`���ご�ɢ�]#��	x&�Ɓ��g��.�A�C�VY��y���p&�@!nǖ�p���Z1�&,���$�kbx��
P����z>^\�+ϏaU֢(~o���!��'(5�2���������i��ևtMB`{�-���C����d�%5;��1��RA�\�2�������� JW8��%�˳7_o���|4O�U`�۴JB3��!pY���;��3��'T�JJ_�(��}Ic��}z'�Lw�{M;��Yl��O�f!��X�0檂v|�=S������n�:�u�}� �RY�N��}]���L�+�-�d��
\�v�QW�Y�X䩧��~�7~c|ttt�����r�*������i��>���x��� �w��lǡ-�{p>b�F�Tǟ,�!�<������&Y�N�~en�2��j_���B�}�eN65��clA���mKD�N1i��i��'���b�O�2��d2��v��&i�;nR~��%y��n/~��#D�D���GH����`z)�\Ƞ�xk�C��sV��bH}���	�����UR��[�As:���_r�I�?�����]�n��P��� .V'n礞~0�j0�	)j�3�Jܒ
W`���ɪAKY6��U��q�*����$�$��.�'��I�DG���J�r΃�������
�7���j�^�B�����l���|�,��7�֡��>�e�ݲ�� b�����/]���RS�떊2a���/f����ŧK*�躖��+�B(����R �ӊ h'�߈'	��aW��o�����,�e�yjlY5M��$�Orɻ�V!GS�k��,�_�Hu��j���}�
�]�&�'�~�'���	���=�'zi���-�E��A�HV��#�
S�Tzi�gJ��2��Pa�W��ȹ��������e	�<��W����	���Љ_�%!�� ��[غ�/�����G���p���︅���&��,�7�r�Ê�V 5�e}��������'�j)Z�D.�f10ڍ�r
�v0vcg��!V���R�&I���<�1�@d�����NN�ϸ���o��+�F �6��7�A꤅ErS��yؔ���f�PB�\����S�A�+�H�t��q^�[N������`����w��]��Ā�� j�@)�)'j�`�"��-X������!0��� gS9�����$$�w0��y>K�����:ډ�M+'O`z'��	gqHb8�u����?�a�2X���v,����)�T-sob��f��*������UA����;�5�(�ȿ]Wߌ: �(A��H6C*��p��/D�i����iw���߀ j��� μ[fZ��P�����w���D�y�B��f��@� gn[�a�cV���t��E�m�׃�[�:þ�Sߖe{h+����ਜ਼�ؤ�4���i�,?��.�X�-.������P '޲�q��ᑮ['[�5C ���rn�(:�n>W�L�UC�#'jc� ��B���n����o3z'��X~��^�2�t"�H��
�:1LcA��\cс~)U��mU4\ڹ8�`N�k�ːz�`�ٌ
��M���.$�G��j9OH>��r�)Jb�uX�0��j�ŵ�5rAT��M��f���^ؼh]e��a\y��A\���F _|���ŋ�w���_�����l�.�d�>��&	M
�#iN��/�yX�6T#��"��Ӻ���F���4ͼ`9�m�}�|�L�>����������/�f��&���1��'M>9�q��QL7(BVg׍��[΋��I� K��$� ������Y�Mg��訞˄��&H���!D�-���F ݗ��&�'�㯻-�G�U�#¦W�v��X�ӷr��F�[�|\D�������r�����-���B�v2�����N��N�����U�X���l6s�{��&��ܯ�Z��N�F�Q-xb	�I�>i���>�JQ�f�}X��n�*q�	�]�-9���*�LB���út,fY�π�� Z��[1��$b���>)&�)������J�zA���C㞹��ހ�!�i�Ji�[�"]�-��Sy�2�@��(��$*�^��_9=����<�2nZy�%��`� M�ʦ�,~?
��Kr� Q��݄^	`�(�:D���D�*� _��Y�nN^��܅o���0�烁���Q}��@��=6�r�	#��,��6X�N�}@�%Sv�A���'�J����N� 6�M�h�k�y,�~��1j!o�~lF�PW��1f�㓦<���d|���d�����7ݟ��6Z��VuV��"�R�.���dx�e@���P��_*B�����Ȱ�[���n��WHpτ��{A���YH���������~�=^5HMX��,�AB��F�͆T>������/I��8@�{8���2�ew�;�����	������.k�P�"na-^+����[_��o��$�����%��Z$�j2�&��}���[�Se��IBI��%�В�6�WȢ'�_~�k�T��	�&̱��O/_���$AZ�FX��|Yle�\�I���NB����_[��$x���p����v�ġ�&�J ��6ݟB�N�2����qp����b1�r!�26I/��?���a�t"��q�Ǘ�-T~����մ}�07�w�s��ևܐ��H�S��,�>�SȍH�p��<}'q���GZ/ZŷE�nЉ�lt���ڮ�v�$��@.�,��%�
I[��o2�ܖ����\nN��՚�+$@]�_���ۢ�u(`U��C���0O�sWZ<���	��-ق�`BVMA@z`��R�]U;ny��]l���'����*�U�ǳ�K�Q���%ǐ߾)�@�ٔ�l��jKPWА����
�G�v����HY%��NdQo��	��Bq�ӂ��LN�6����b�����5΂�>��k�*B3ք�벹�ׅ;��IH�bx����&�F )����2b;D�j��+I�[�]�s�h�e��by��O,"��&����l���nJo��V^����'A�m?U�G����T�܈"n��f^p�h�A[5����B/�ˌ��>�#tH���&�R cFj�rb&��G��;������W��,H��\e�a�;�ΗֺqK�+=�ƺK|�R�R��bdA"fz%�L��^��K�r�U358���
��%b� ~�(�-�lh�N˺�3[����L�8�in�܄�	�l�7`;0�]0�W�!����j�[��/�����x)]'�^�[�'���5�F )�MV@�k���C?�RA�"Q�>��[8���B}�����:�_:.��۔���3A������~]D`΃my�� ч �
�E�-d�xs�^Ѯ���ʴ��� fz(�]��������7�.��O����g�Н��O�������Ev<rBt�xx�#zz���]%�uȀ�[�s�7#�d*�9�<��߅��������Q���xV]�o���	�@������p�7cr��j�Dbu�_��L��&�ɿ�,�!�v���ݾ@�.�@��/�;V̀sOߗ���aȲ�-�EY��:�U�AB�{�}���mF/�����;M�w��m��i�w<�����i�w��-yO�����^bnoF/P�C[Ft0�6R�pRG�b}S�+쵑�}��)�� ���K��w� ���#����(��ܯ��	�C˽Օ|��Z�N�]8�:��-1@=��?b���Rs7��9	�h�&�`6厗��l�>�E�=�-w}�=?h�^ұ�v�z"�*Jw��Ͼs�:�/<�!F��El�}+��E�"�����W�j�.ϛ)pXT�������=|�]���!7v$�S�>�v���D���s�:��y�O� ��$
���Һ�DS �"�9�w���/:����ӻܵC ��cA=9���Yn	����~EBHWhW�$XW��yN�5���p����ٌ���S]+$�p�[b�nuݿ���D���>��@�f�J�%鉶�PO� �u	��`}�T8��r*"���:m�s��+$�9��ln���_L�[�W�ZҦ�`�����,Cps�"8�E!Fh�yt�;/����ʮ�Aږ 8/������ +q5��
y�	`�༘�^��I��JU�v;X.��"fz#��o�P���� �ֽ6u{׽u���̀�����j�F�"����aK�r�����)�T6�`6�(��]���.?���Tnwa�E���7�2y���]��بJDPҳt�|N�j�y����UjGӶ�X$����>�@�]��
$■�K�B�2������7��񵄻H���*��>6����vI,�!VAP��V���uM��8�ۄ�`dy��%֡u+��͛7^~��xـ[F�%�w�W!�ר	�hw�e�i��=��$x1� ��^	`���~�,�z�,�����î�I����.�ꎵ��N��T.z
���*��ǔ��O[A�8X؛�U��-����Ձ�-�v�*.�-��H�����1��|G6�y�\Y���N���I��K&*���f3�,hk<����B(c_����@B�F���[ݮ��x�M;0`s��R��Q�k�d�:��\U�q��M`��N9$�ȼ0�)�F��X� I �`+��@Ɔk�0dy9��tm����l1=�����bƎ�S�.&����������ԧ�;;;TČF��\>�o�NM��z�N ��-���J:-SlF�������}��B�L&�Ws�����h���홃�s��w{�����ҥKfߋ�4L�⋻��I��+�WO��,~{9ml�P��Li�p���i�HPG8��/zK�đ�$!����ޔ�`���~�7߭b�ڎ>W��]��������?'d�w�u�.�{��q�)���i���i[`�����t�
��h�0��r� ��AR��!!]d�k���ҦoI֧H4}}i]WpYP�X(��������SWp��#
�]�T����ɉ�����}��Q�N�X���k��6�{O����吘��F�,4�ɷ'�.2�c�Xߒk�c.��l�/���?���!-��sV&���h��E&n�g�A~���v�B_D I�vww�k���"�M���g#г��p�Z�J��>t�yWH��a�"|
\��̔�+�H\ AH�~Q7�7��U&f�H�\Uo��%I�g-؈� s9 ��}(����E��ɪ�����#�B�����DY +�mHoP;�e�����C��V����G+b�>c�t�`YDH�ʐ�,Ĉ� ��ܔ� EƊ/��B�|h��Mz�B�n��;ˏw1����&��.���S`�s�?��<�F c�H*^�[9	��h�[0�D��u�5�;8��Qn��a뮪�O��e�ߦ[A��q���v�@�#����h`|�ZI��ڬ�C����xkX���<m���9��䕤�ɩ/!���07�7H4��Ŕ }É��z�E��ȗ</�k�߁B9��*�@�JG\7 "q�dő��.�l7A'�@��oF�P4���Zt]�\U/�éi���O��=��$�%�п�N�҆ ���n�v�z��'�Ƽd�z�B �5'Ն�i����1?�:��+䭣�_%�r����o�23п&Sj��{�����R$}V���x3�x��x�]�Ao<�)�[�=An!�X�fNw��[`��э�S1u�����a��r��&n���3B0��B�".�Xͪ$�����&M$L�ہ�<�B2����yp'�VTg|���%%��k�t�]<�w� ����7n��v�
�&���Y���m@"~�]����c9�4�C�<O��W��w��^~��d��X�7�@!�Fk�]
k1P4n�xN���&���g���`�J|	]���"(q�D��e#F�Y#����J e��Q���͢Q���e���>o@�
WU���M�ul�����"gU�gs� �����s��麀l��p�9k���yrғ?�(0�駟��n�x��d~�M�� ]�\t��(���Q,q��w� 
Z e��Uyu�NC���������_�߿�cn~�Yt���[j����n���O�MO@m���!��t��s"ޤ��}/����^y����N�\������<��$�Gݘ<��G��y��Ю(�J�}�W���4�l�(]>�Ӈ�-�����e� ����}]�Z�t�n��|��_�����Zƃ�*�-��nWs���I̫����e�s�c`c6�[������i[�v��v�pkY��=�s1g��g�%��`0H��ٙ�f��CC�.�!!_R	Z`�R��[��/��T�u� .�v-����b|��h��ղ���ݎ�Hl�Y�wt4���@���ơ��G� ��'`7�w� �)0G��Jϱ��a���X�i�Jo�b�ɼ|u�N%��8Y�un<�we>�a��@�DP��J�،��dBan?�1�7�"�;32�v�XPd[�;����߯]�R�1\�;^ �9�|��$&�/����y≰v��X�[��Y������T�j�w���Ne���$؟>#%��aGY�I�	w� l͕>Z�(�f>���b��4,rK?qc�u{X���m����[�_���a/��mGhy��8�gAH�,'� �#�%���ل^�BYI�f��O ז�.D�����$���$>'��+����j[�|SsM���7�%(���9DM�������|�Q
��V�y�y9w�U8^�^LC�Y��Ka	���	�]��(J_)C�(��L�t�Z����	a�i' a\d�q��(�ư!�t�牷�{/�������~����kr���шVʡoHEN�㱷�$�O��	95��LnL�nD7��
��<�_E
���ΘC�#���}��u7:��7n�m��0���Tt�C���n���������g����o��ezW�չ��I���/t ��M�%�˴��p�t�[����$��V�w؈��pf��^u��w˪���E������>�7თH��v�#�rX'��v3$�,W�w�g����|����� Ft�?���	�k��D�����,�n��>�����g��zŀ�H/^��L&�)f��t����1A �Ϩp$��a�F����j�m�ӧ�4���>99��_v?�{=w� ���I�������~p7�}NG$����VA;��d��|>���<�	��8
ޔ�~x����o~�kE5�?���k��;)B�+�ɔO�����?�C�ƖV���'�Tm%�8�pr��N��;^ �{x��w��,�ٻn;�����[��k����qL���,�UBa��\�1������r��"d��ֺD���Ӎ:����X��N0�g��� �+�Iǳƚe�� ����x�?z�g~�&��	څ$I��f�̡/�&��e�����JO�<����Mn�f��L��F�Nm���O�t&KhS�p,���Ā�
�"vRA�ȴ�"X�?۽��{��{�ݯ|�+l�/�	�O?��U5���/?r/�R
9׭%�+}eg�xA�����g_/˓��:Ȓ3��RF�"��8��FvV�|�0�6�t(�'��M��"�rp�g�;A:됦����?�k�t�}��'��gC�x����?���pr��ޚ��(�8�As�Dp2������x�~ݔo�y}n�-�N��Q�f(7�8�%������V��p��>|m0�����N�����U76/�q��x������s~U!T�7����։�߾�ꫳO}�S�ooHo��_�b�A�̀��rp\V��!"H�(~ﬧ��V��*�_U�<�����_�>5[�����N��ʍ_���������6���}�_�DВ�>{�k��k�#��� x�q7^a��-����.9�׽��O2�QJ8�s���e�N���E��k�m�j��_���3�<��7�cw�8���bE�%McJ�1t�b2 ~�Ň� Xw�ݜN�_OL��_�L:*���{+ω��S^J�������>�i򮻁�^����ݭ��!2a�կ~�'���p���{�F_�������s�Y��pn �`e}�Q��~.px�'��Z���  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  �  `k�  ���;/��+~Q    IEND�B`�PK
     ��Z���Ȋ`  �`  /   images/457643d0-fb24-4111-9541-c1c501ab524b.png�PNG

   IHDR   d   �   >�?   	pHYs  �  ��+  `<IDATx��y���Y���~�ګ����5��HHB-�D�0�0�1l@�1����N�I��8�$�	��Ř��@�F #�}��h���ޫ��������=��ݪ�OO�T���'ݩ�[�~��l�g}z����W	r���&;^%�Mv�J���x� 7��*An��U��dǫ�ɎW	r���&;^%�Mv�J���x� 7��*An��U��dǫ�ɎW	r���&;^%�Mv�J���x� 7��
	b��������@Q/���	��A�ᄼ��2SD�!�<
|M^i~?Ք�9�HS�G�LE�G�_R3�O]NǴ���0��O���CAQ��jE�ұ[ݽ���Z���gh�֊�x|���m��)����s��b���m�6�7NS����^ ����t��JG�!�3��h��IZXX��:�K�O����h��ߞRi�4Hyi[���П<1���������������{��;r�����~����{jȿ���گ|�׉��D+m�����|�ķ�JUT��4�d��o|�k@Jk�UIq��&߰���R��H˩=й/%�G���@�%s��"����3���1B�%�{yaLF*�&�{1����l�ӕO}���������T1������D�)��k_���C��+z[�'����{?��46MZ][�j�h-��w�O�������C?�K����ߛ���qɬU��U����ÿ�K�'q��e��*�$����:���<�DAP��e�z�V,N�xf�By�|��L%/pŤ���O�Ա
�0H�iM����.r�킀���PȔS��b��k��T���� V�#��{Y�"�����k�d���n���4 �{���%ͨ�џe��z�̟>K�^����A>��?����7��'�?�3?�|����(-�F��O�qZ����=���g���܅K����{��Q�]�r�UY��,<�W:�"�����Ԟў�k��4K���ڰ�*=�=��2����3��ƒ1I���Ӽؼ~,!XE~�,|�+���XVQu�+�����]=~��3(bQSXr�O�U�b���|� *��N�%sG�#��L���v�����/τ͵����B�Lo����a�������7���)�?�;��?~����{_A~��{gHo<�V��ɧ�~��'������Gy��m^fO��U�Z���;��F���g��k����۬�X��cX�g����:V	��Љ�c�yP-��L-�/�����cQ�ȼ~��D-i=a
����ӈyq�D)��@����T)h��^*�|���"�p���/]�f`�[�.�3��?MW���4d-Sd>W�6i��f|���\�ٷ�1��~�Vٶ��>E��O�����6{�s���>��'�}��`r(S��ӈ��G^��<��2�'��	�o}!s?/����BXo,2/
iV��%�?��h��F����� X����"߄����� $�� �j�.�Sn��r���5Y2�_�в�5#�����0L	[��S�4>3B�s��N���#i��W��X+�U�� 5����S��r�O��_��o�Y�4�C����/I�����>N[�S�=uq����*��
?6C�˯�W��09[ǬTrJ(p��/�	Q��gde��AA	6`yK$,D���Ƈn�D^p._C^�%�i��
��ȰX��e�!W�,|GT܃1ghPϩ2KvG?�#��w�YDh>>��L��}���l��V���3���j
s�����<{�ݧ�����{ñ���>�}�Ol9��/��?�O��H근��L4(�;�D1#Fe�����l����C$��nQ*��Z����dA@L�$�)����A_F���������I*�J0���1''}uH̱)���`�*1U�1�wO����	b��w�8^�꽔�?o�S��D%����xU�i�{���K�tͯl�a}a������]�-6���Na�.//D�73,.6�t�{kڿɛf
}kU��bs��+�.���J��C+#,+��.�,���uF{�!���s�YU�aȃ����!Rǐ���b���f��jIY1�N��Li�g��DŁ#��Fg��IFUQ	�|f��[�q?��e��'&��o
ǯ� #H5i`2/
�:��e
����r�����90��%<E[�h���Ej`_��fH>�H�L�R%�C�4���XEAa�O�� 5a�eԳ��vx�
6�LP�a�Sx�=�E|�bL��1\?+=�6Ū/0b��R�I[�a�ɳ�)d���bvrq�i6dU��Ϩ����bU�h)���_��z�^���3p�&;Dگ�U��=���91	/p�D)�M��>K5c��0p���2�l�I9/p��^X���<�K�:p2�"��JP�*CS3�SZ}#��q!�+3��>���3j�eYN����N��fK��k{[q����w!04����!Z�8>W��EP$�O�+`��,��#���>��R�����ū�/0dnb��?)D��/ZT�noZM�Ae�4���%��R*�g���m_>OL^>?��Q#l %��Z	��F~�Wa�= QQ�hha�f|.�Ua�h�z}J�}�|2O��J$	�Fݸ/;K�lX}���ӂ�B
���f�����h���}�/����sW���@_f�$A*����Eq ��%ɏ"*����^]�m����\,����8����w��0L9ꋪc���ۥh6�1n"���<V�TS/��ʾ�ɪN]�%�=�|��J���Ջ)4��CV��q�\�����k�}:H5$'�J�A+k�R��0��ݥ�	�g�
��A�>�+�����;A�����Z�KG�R��m�)�:�;b�#n�� ���a���<�(����7x�R*�[,5}�[�"E�a�!aKx!|o
TE
|�v֟�b��d��$���Flk�)k}�)���Jn�s`	B��D�CY�j�Ui�)Am����^N�U�6)���R�})�?|=z�4A&�p����O*�I/c�Jx:uw-�a�P8��xk�5*Dc��%a}��xQJ	���0�孎�XDeE�Ϥ��"�O ��g!(T�V@{��|>\�����w���=�f��9�t����g��xQ$LT�Ѝ��%M]��1�t]j)13�
W�*���Y�Ʉ?�$�Z�� X�����
�e���"n�l��d���+�$�R�C�F~�O���r0S��I����p(�O��?�Elt��0 ��֕3��'���ya�&Uy��U�WгbC�hF@�	X��L�9��s�4�Е�~=�)�ЗS]B#E;m�� э�H�X�J��n�+�(�� �WF���֓QT\h=��I�@v�b�����Fg��M�m��x`VO9�.�r-�R~/j�י'ņ��	/R)?C������T�sl_�fm
�'>��Q`~��E6f�ˏ�\���Q�<�x�ӕ%�𾲨�	�yw6ҳ�]Ա�3���o������ ~��S���+#HjE����*qܬDx|3�2� ΐ�ؘ������G�m��m����H���|��6x�(7������͈�X_.��}
'jv��_�2b.O�K�-kh	��P nY� 1�I�7&L`V�A�Z��P$K�@�{%�	K�M�O�VMUN*,�w��E�,j9����-��K�/'�����,�8p�Ĉ�X3A9|�\�ʓ[��3'�4p�X�xA&k��l�E�x�{��:N_;w�J�3@\�4�x�Q�Ca6Â���g�☳�5+K`��}���[���
�;l�+Fed#�\것Ƞ$����x�2b��rk����a�$�T+��1@�R�-���w��I�D���ς~]��������,�_	A��}����:�� 7�HD��Hƾ��1b�NQ�~h%��p/Vo�����/�g>>�׽�t��9znm�FC=�����c'���p��k8&������@Sl�
���7�C�
�y�=��>@��~Z���pv�L�D��e���!XyaIA1 �@��Z�T����K"�)Q�+�oA�&�ge�@�Q �{*��q9�/]�*����*��W@��/ry�ǎ�J���Z�]F��L�<�_�\ǉ<x��b�ٹS��C�<s���������>z={e���<ۂ0�	#u�f�bd�C⥥��,>�L�s,a	5[1��M��`r�����:���N�7�h�_�0�e5j��IM�z>@��	Ū�Cd�a��i����h&�a�@`�l�*�剉��>+;�pRd�����]�E^Ė����{�>꽎c�'@F�uh4���Z|l$�e��7�����/X�-���|c����4��k�i�^s���_X���P�啬^�/�:5�������ӧ���:�<�Dh��6&w��2ڪ����6;{��nѹ+��ū�����+k��֩�p��s�4a������H �#�=�(^��l�m������Ȅ���+�c�s��3	��}QYF��:�~e��u�xyv���I|�(��XN�F(m���<�j�1��!�H������Xu�O�CøM��*��&{�z����;xMn��N���Da��1��K��Z������[OR�;F'�+�ʢ̉��E�ͦuxZ3,M�Ctϩô=���n�/<�5yml]u��� i�/!!%�r0ԛsjqH��j��v�b;R:���?�$Ka�bC�KPJ��L�]D�����WH���U���0I��Xm�w1a�5�ȟi �m�B^��b�����ux��)��ߩx�l7���������d�_��3���mo����ƻ��|�b%Dc�l���p�J6�/_������;n��/�����4�hщ�;�[��kO�O|���GI�lQ���eF�+
,�ݸd1��q�I/r�,����I6H����0�^bs��PJL5MAב�WD�l�Sos�yڰ:֜!$��o���g�ќ�%��ǯ�F��9sZ��*Yb��GYK�4�z�|���ʳOQ��`�u���M�Lox�-�`�3�F�U$ҧ��AΪq���̙3����vc���D�ٸ9sS���h��л��t��	��'?G��')]��Y<����a��������Yґ��8,��J#0]�c��B40��Č���I��)�0��Ue�'�|���L����=��̡�hHj��.�����~�C`�����O�q~0&\�|�&���eң�M<z���w����0�����F׫�*F<�7�{�=��3�
gg����-�t��	�����J"�^%�Q�v3����<5�i�쯾B��4{�]�-�ٓ�6�WI"޶D���Ň����F�%a�Kys�j����]���C���:T���>�y���p*�Z��`�L��d�?`kvi�4�i�I8ނ�@M�D�^b_D#�~���w��T]\���y���w��n=1���&x@Â�P0��b�,%�р�W.2C�����/	��V��ƃ-���# -�46
m���Z�N2��O��旊>��_�r�"EsǨu��1�G�T���x6?"�{ ��5[��4�G�XJE��v��(�r�z�uD�2R;���6��W��|���N��K�x��"�̚�H)��d�����$Hg�	�*,�m�\��oI���[﹅>�7ӝ��(V#��A"����Ujs'�'51��:/J�	�ı�"Jʉ�B�xTYZNdo�d�~|���]��FH��+O�:�Äs���[N���k��>UŌw���u{vM42�")69%WաJ�OR��}��������B�]MX���9��[��A�͆�,bb�X�z�Kӌ*~H�G������zd�0��K�#�o��^���c���5O,��x�XȜA�bEB_1���zEQ��^���x��\�d���b �
Hd�����}0�x�W����o{3�^ݦ�_�1tg�MJR�P_*�B��r�Bɾ�H��W5g:1
�=+��5K�r�X�JR�����)!yѠ�_��O~��?���=a��K���/h1g,-J�u�� D��)��6 e�Nx�X�4�S��0�VlhiD�����~�^�)jEi�n�y �x���h�P9!x����	6���4�q��JAt)\8�8"QAJ�C�YJQgL&������o�Z�ħi�['oa���D�rFj�\�8� (�I̘,���RU�tZ�򔳟.�G�^h1��e5�p���G�1s������7�𩓏<z�Ғ�7痌f���q����0�|�y��:J��Y��2�V�mQS����ŋ4<�	5Մ��v�ld��(`����MIe<�>���6�����wH�ԡ2��r@=.��xaIYV�K	�,Ki��,��p�m��c��C��+�wD,վ8����`���W�
����Z�o�;�-��#��g�L\vԷy]��\�0�/����,'�iվ��~��q٦Ƃ�4�є���/y�	.�o��3��"W�0j�7�hd���SP�Sѽ�9Nw.�P�d�uE4�?��T��{(6��p��I��������v�^l,����,W�b
� �٘�P��?�@�x������^֣$j���$�XM൳�"�Ƌ^2���3������Ul�~��4�Dw�d��(~����%��=S�}JH�@�-��[�M���նW���Xo뺘�EQlsI���1�:1��	bA�<0b>>��1B�lR���k��1`���X�ȩ��p"P	�����X	�	Ħ�]�،�����ܿw2�.�L4-g�%�7"��5����|?_ڢ���v�)��;啍n���!)L��E"�7��S$
R��ph����ܭN�&�d�c�No���O��*q������
839t�U�y6�AĢ�3]�����bB9K��Bx�!����r�=e˹�ψ��]E�(��I֏A<���
/��
[WQI	)�����])Euyr)w���aUb��f����n�'/}�a6|G����8�"ͭJ��I~����Yֵ)�|<|&�`��Ƕ���Ke�L^F$�?B������kO�*P��
���\�;���w�^��C6��h��1?�%,GOcQ�G]Q�@ D%�#F�Za�Ο#lcmK��i}�*��#j��6.� 5�XnϦk��,�;��8b�j��&�4����~�ˏ��tȆ:_C�
v��Ɍ��������u.�,p��x�\�w���KR9�C������{�G�`{Hs���Xw��GrΫl�ܨ5M����D�J�*�<I�d#�鐟t�=K�'N�h�G}�l-��P.,%��(9m�7���)`!E捹<�|�d�`��>F�/JH�����{a"Q��>������4�D9�8O����*�{�e��EF	l�����T��iP�m��rIE��0H�U|퉺������ٺ��b�ǒ�����H2G �������l�Y�>]S�̝��hv�-.�₫�봺zY2yIȜ�	�@�J �%R�'��9��}�K8_���aS��,�rm�l>U!��F]SVE�[4�d����q/5�6-̱s��#ith���{�X_(��K��7-���<c3����E����S�U��k:NQ�s��?\ku[���,�u�vU���6u�UiT֏رK"?��_>�i2N���S�5��@?5E�5�P_����i��o���1b�>�9|��_�J��h4��2^�1��c�H`9�3)��D<�D[I�G��6?m�zU]$Q`�T�B;r^�-�����n��1�S�9d�Ш*�� �k?n\15s�+�1���_x.�`qn�=i���M��:fu��	�Xl��l Jx����ZBCE[��Q6�ny�L*��5�y��d2fu5d؛��H��ύ�>$�����P��jKO���fb=e�?ʅ�kKO{Z(��ү���O���xq�(5`���:`���PMI�&�a�l��{[:BU��<p�b���C�>��.�~h�����؂hU�CY��]���iY�8c�)�|Z�jmMm+PL��t۹e��s!�	��=�v�� a�:5�F�6	���D�I]�Yig\�%<u�BIi�
�I�Q6K�th\��"i�!H�x����/��74
m�Gi��].��z�B,<�U�by�IՉ1)�P^0�	ՀY��s%��"���}(i����E�v��D���V!|!�T7�ز�<+����'�I]Vʄ�h8` 1b	Ii���
��r-=��1bQ�rFH�.5�{Zl�$�}D���RjF]�d}�'�J�p��xlԽ��_%!�A6ӾT[���ϖH����t�z/�I��F��x �A^5�\�ۗ���t�����$<GX��"%ZVbԕk��<AGF;ciS�h����uդ����z��XJ� E�2F#VQ|o�&h,͸���I)>;���
Ec*F)����5�VL������g��DRp��됻C��E��곪d��t��BE��=�UYŪ��g�aF�E�7��'Tll�!lH)��N^�dوz�2�A'����5��x*�\���9|�SbN�������v
N���\3�-Jҁd�,!����ޗ~w��E�����lLU�Q\e�|����I�
>?_<3�(t�r~>8�!��f')>�5�h�l2�����|��	S�ZJ��EA]��N:H2�n3aV+���:l�����d����V�nщ�m�EIJi�-��m�\JM���&Dx�8i$Q��ű�k��E��Ʀio�,333D�ͩ�����X|����������nl��Ͱ+�D��ҋ�*[@A,����� �%RN�n-�ڢ-+ł�˞�#��:q�I`h4�{rb�i�k3@�LU*��m�A��盇��B �F�Mc�؋����<��.P���3Gh��?��u)$�Z�hУ�֖x���|���֊Q�����<�/,S�1O������ˁd.%;)0_%�����F�V6�"�'b�ЏH(Z ���K�RL�=�P"�+���d�Jm�����^S���|��(�f����6���;��%%�4[��~z�TQ����F֌�����5��P��YJ�
�f���&��z"�!KR#DW�+���[��%Y<f�nw����URt�ma7*�<�̕�PJJ�Nl�
}����Rk��E�HOP�8fi@�'���\�gݠ����1�����]c���d0eXN�3���i�zj�y�H}ѣ��µ�3���G�G���T�TR�)>,�Dx�%��oetncB��Y�5|��m2�BYr��r����L�6�N��&��X�ц'���ϳ��qi���٨���)]g�s�������<�BeԡaR�5)���	ht:����/��^�4)Fr���\��O"����\�"�1����OR��X�&�<�P��P26� 2��F�=���L�)�3C	�$x\c ���u��P��[�m �
YtH��!�a�)d�)�C�x�W��6a$ac�"�K��o	S���9vP[V=#�3�/�*ې"�a)Q�C�ʖ�B�DH�oh�/B�5*ȥ	�vހ4Aؐ��q'Fa%J�|����)�<�m�b���y������Lf �Ѷ���N�L?Ю��Kh����ֻX��ei��F̔�1+�P�x�4�XR�!��(������}���R.�km H�'���gm}��x��u��9ihu��03R3౳�,4�G뵑�}۲y���DQ��.�%~�H������܇�ב�⇷-��v�\D�ؖ-�*�o#�vȌ�#�x���z�ڷ�8���5:sn��;ڠnYu��Z�x�S(i?���m
�~�4}�#�@��I��B�1z'�&�<Зg� �@m=��q��9�4S{��Dh�z�!3Cu/�bcI�J���U�W�:^�t`U�i%��1N�\a�C�^�φ�f���DTB��
-Ӄ3�F�oGR(� ʿ���
�MY�V6�>bNZ|>K�Ǻ~kh������Mz��Jnvl��޳pZ[�$~�gk�r�9Re#N��!y��v��Ae���&Ļ$�cb���9s�>��G�
۴<R'Ye�$t�Ѥm���ƱK5(�"aP��7�1�ߐM~Yue�8C�t"e�t�}J�l�d%5O��犡��]��q��2�ߢ��C\�����\'Ҳ�1���T�-^�;tfeD����4��Ej�>E>FTL� ��L2ӌ����ѐ�����Q�CA��}^j��ݠ+�)=��Gٖ�]��8U4`յ�=���O�I����J�֕��'8Uw=U�CD,�g���1ܷv�eVEeN:�A�~FI�	i+�����$W"҂��6칎�PQ�3w���9�PN��J2q�E9��g�����W��ۏvi�P�YT7
�}[�Tv��J��Y"6�R�\:C�^F�l-�;���I�F|׶��<CO�M�[��̐%�gQToe��1��v:~�i^ؔ6'��x���t�`�K�8�fOr�uc�r�6#%#�<�M�>ao�6���N>��sW�5z�;��5)�G\'f�F�
�~�K�:&%;Y�6)�^gaIm�C��u���3h���)��ct��K4�ҡ:D��%eܼ;�,��ƶ~��ׄ]Y��CŶ� %tnkH����ѳ��K��DuKe�J��T����tq�u꭯ӡ;ҥ�>E����(;RJ�#j�J�+�9��
O�a���FQ��� ���VJ�%���w^���O]��6)��-Yr0�!bO�Q�8XpUJIPX�%���gГ��k�F���Ϟ��j�H�QְAi>���[3}�F����|���	�*%��*����r5�b4�ズ-�8�8coy��a� ����k:w�G�{�=rv��f1e�.ۼ6�3��7��4�)��i��s4i��;����%�)s8]�z�R0�v+*^l��o��8��HB�T�+��%�<�@�;u�	�E��-���;z�T̷V���a�Ч0n�p��!!(�LP�6;K�N*�rm�|��lf4��eZ��ړ�t�B�f������A$�C�\�<�m��a�Cj�5}��2��Ѧ�f�(��(���]��>u��c��&�A�r�0A,>Rc�	� \�R��BK
�����[��2�hkkJ!6�� ��"&H��e���p<����ٖ0aUI�Zf,خ�}��|�e^�	��U����V2C׍�.H��y�/p`�fUA"hMV�Y<$�����6Es��� ϓ�v����
�����*�M6�*#�+G�t�R���%|�@�5�Oѡ�E�!�-��c���5�3�7ڴ�7�6��Bo���
=uq��XeL3�B+iSj d�/Ԅ�n�Fң���4�|��^�l^�c�*%�\�2�TR ���Q�р��=
�9����VLIX��Bo���A�eUs�)�����2g+vnf��_\�޳O�MQ����3K9�Z��͑��J��g���5��$�Q�r,l������h�.O��Z��̆t��,-�'�0�ᇜ���5��'�����+l��b�2�+�!����v�V����C^H��lqN@n9F��y�s�4��6^�JE��3̳`th(c�l��/F1��a��Jë�/Pc~V�/ǐ�e#�Z��d:�s���㔮��x��*H3��+rZ<v��[hx�I�ʒڧ�d�;+�洄OBf準�J��H�\���##:ā��(���2��	����,�n'�n��_�����20��hD�aƯ�6Y�l�9�P��e{13�D%�xVM�19��y�Ō5�Na����"�24!'�>�*�v6��p@���4biR�A��1��MTEq(H��*H�#�0�c�0K�#���?4�CG�V�#��x�s�ܡ�wi�³4y����u�=4�(���Vt"�38a�F�D�b/R(d,@"�j�3ҿ�ei�4Kd�7���wm;���*�c�#Cc�P���ܙh�=��<�i4"6%��7�ݰ5�mB#_"P���u�QA���3[5XJZ�A�e!�=+����S�4i�H����є�܅�1M�v��Ȉ�(A֟[c���zh�0�	��]�1ی0��qx���s�77�?Κh���3@w�,'ao�W�Q�EeVt��湐��ƣ�[)�V��͕6�]T�g�X$��<�]�Y �z!>�6mEI��(��,�4(�5=��΀2���NSR�BC��4���Uv�j�q�u�i�j0�6�������MB�N4J� �j���Kt���[٨�V�����SaNwD�%�IU��ǇM&21d�[5(�eӴƦ8��Q%\n�a�-��(�d����J#����&��t����]��N1��6��~��H��m��4��t���g�fW�7��H�m�<����!k.��|C��Q.�/�d:�H3C��6i���?�,���m�7�yQv���I�2�EhP|�2������jS����n�Q�U+d�����):�Jw���R5�VJ���vav�����u�i�~�_��3����6��B)V�(�ؠc,��� �|�p0�T�^�c(2��\P��T^�L��2�()�O��oDG�;���`���/3��>Uu�-�w�@�"�k�����T��7�G���C`��ݧ#i]f�.N#���_��'��2e�ܗqh�ǟ�6���~��0'8j
cbP�.���_i�LPTU4�0�;����*���3��<�g�9Mfe����@_z1d8�iS�;(b\��l�0K�U�ɤb^��]�����l�Sީח��976�&���[b���G�����`�Z�x�c-�C��K�[���ߜc�&f��QI�|�ʈ����$�1���s��vo�苿@��z�\8nhݰ�m�+*f���Y<jg��uH���˝��z"[����ѿFsL9�&NM��vs��@}��!��UE��&�'ڝO��R�u��۟\�������{������˨-Cz���a/��fZ>kH�~��)دQ��V�{��?�fy����1R�+iW��0L��T���ɰ?���XOY`oj��u����k�j�3�i���5g�������|��Dk�\\�yG=�Fsݫ�2qGf�LPU�wM!9�	R_�y�C��)! H_�7d���oG`G��-���J�ʫ�	��AR���_3�.��b^i>؅r��K�<�;�PS�}�Ύm!Gw���еR��q�
_�oޥ2e"�l(`��I	�*�G�W`��1=����Hm����r&12����ScC�����eN�L���;�0��݂�|��۱,4�lN�x^t)j���%��{��Xm�_h5�����j�\7�n]�<�(��ڜ�V��~����=/�I �(�M���H��}k�G�f�i����D�x�_���d���<�6д�h��ћ>d;![���U�nScuc뒮y�]�z�4O{�q i�﮼s��)���M���%-�,��1��U��3;��f
�c���N((�!?_��N���b4lQ�i��s�U��=A�v���f����Җ������x��*?� zR����\�Q;�l\�㢝P�.rغ����%��Э�.�2na�5��*�S9M��_�n�u�˘]o���q��B� ��H��ջ+�MOF���E�y¤��O�f�����Nޕ�~8��v�x3Jad�d�L]s� Z����W�5Jf��u����Ju��INO��F���dcv»�P�sJH'yu/�n	x��Ծ�%�SA��m�Qu������E^!mT�QMI9�2�������A_;����0nz�!��y��P�,�t���|c��!ʩ�v��t��H���9�Ht��^�i$խ���V=�TT4���s��A���Q뉼���f����j�oj��@A0��c���.-v|���O�ȗ0P%�[#6�UH-Z��V���)�j�C�Q��P.�б�gJ�I����:�(�QٻLj1� ��\��nz�q�ب]OV?�ӻD�Oܐ�����\I��O��k�����k���u�GZf��K��y�g�A�gl�E5�/�AX�%�F��*�Iݶ�4��T�1/`��H7�Q(�����x2ɱ}\`�dQE�����:e	�ff(�?�����yS�/;��qza+ѵ�G8=�N�]�SW#>	M��	�]�n��^�(S����.ĵ�!go�ծ�I�� Ǆ�9��W	cH�O��;dC�T��-'�j7(�� ���	2)sOk�����2��E3D��h@��%��Id�&���d�b*���3��#fd>�T��VX�u��rQfR�,�K�(U�?�R��:��M�j<��l��v=�v"R̒\ߦ��
�3l�ʣZXD��`O��ɴJf�5�}[��M�>J��	�Cek[lm.5�`;2`��X��I���C�������lt�L��ޅgt�*TM�]z]M�S��X���k�w��7��6�YSdx� y&�9X)۾JhY�kT��ʈthru�@�����|6�l+M�7��HB�;^@?�����_�v���Q�:f[�11F4�z�����×���B*��R���&"2��ڀa��i�|g���>�/�4��[���1;��8�>%���(�Fڪj����1�+=^���yғu�Tӹ dG��M2U�ɜ��3��#�1�J����jΨ��d�0f�Tm^���1�,�~��{9���/�{��E*�Iz�ȍI�7Oq6�F�Ƌߵ���/C/���3̻��� ���r�.���U#Vu��r	5{��z�#Dl��K������s ��ޢRr��蘂�R�S�5�����	RI9�������+S�0:	P�ҕ2&���lK|֝:l�y���"��+&nh���BwUl�Ce5��6���@����yҠ^H��_�w~�T!:�>�:����^��F���S
p�21�*������sQ�m������sIgI)�
;��	��#��7�N0�a�<�,�f���D������A�CB� ���ɶM���m�����ȅd\`�1�T�IO��]5]�����Ӌ�ڟ������k���_��ت�z���BN^&Uv���F�+2:�ʁT*�}Wi���lj4ح�3��R���e�f��S	����"��>��M��r�{��9j��F����-Rlм΂HH���������^�Y�H�S9?�'=u\��Ԝ�����EU�j竻]y'�UDM��.��\2m�14݄EFbD��ez��6K�åSʶ6�#��J�2:s1�_6�Ad�J�&��kc	��l�j�Fi�o4@�"k�Pc��D����ڹ����.:�d.z!= ��)S��>l����VK�h�Z���TO{�E���,1lQ�WwH��T.�W������q𭏣��u���e�ԗW�)������<��=�#;�e���2��??*QM.{ay�y����1l���yL.�Z�F���h!>�w�L�MC�Q���+=fd��)a;QLiH5����q�����N}(�	3F?��Q|��h�rhF�rkO[��K�е6���:L�"B����H�r]_���$��-�Z:����"Cm���\)锒��ȧ�������@)x�Xhl��	�v�:��D骬� (��%���1����J�f�g�8i�oޓ�h������nKS�)e�]������FҚh����JW��ɠH��n�T���6�5��n�n���E�ӈ5�����l	��!�X��t`3�c-AD JDm��L�^�^�\h-��'!��H��g`�2�3)6�A(��� =���(0��`-YC�h�O��f�tftG9&*`^��Y��3G���M�����~�c���ݏ�}cӠ��PM�Fw���ߨ�3���uhlZ�PK�4"�>g��M�,�)���mH�p���� �φ�_<��ə󑞵�Ҭ/&EtáC�	�0"�2{����$��l4���&�6es�65�e�+A0�q� ��4�T!J��c7Aq���s�ʹwv}�@�-������y�s�\��v,2�����%��T
��0=�U{;$q�j�����Wo�G�+��W"q�EZ}vC*F�u�^R:[���!Wu�F b`��_E5�C3n0<>|dn���Fҗ�0.�ƀ�R0�7��;m!ڪ��hU�zS�Sk�k@�T"vC"�L�O� ��q#SΩ��7�F;�F�ȴ6�*������L<�l���ۨ�� (�%Q`;�����>e�f7�aQ�*�f����N��M.���2�L��~��M�`re�NBH�w����S����h�^0�����EN9}�F7픀���U(��!�?:e�+�l��YX�^��m�z ���`��2�����؎�M�%oT`�R�:�@3�4�7��������~e�B��1����B
nz�%��DN]����`��zӇ'gx�V�Z=��)��>�� ����.�XJɹ��<N�ㆦ=�P�	��V��������ˮ����yv�jL~@B�eyUÙN[)��~�5�v�aȘl�B�StM�雪+�i)3����C���GEա��v�S�c��ꀠWO�&��_Wg˹�]�WM�7%�����i�s4�`����!�GOv��ݽ�w�H�o���\l���J�	��|[�V\m�&i��� �h�:jTY��X����5�yI��XC	G!�#�]��m��כɫ) ;��aU�>��z; �L�Cs�]�z8���M��l���G[ۧ��;� ����mM�Jآ�����+qvҸZb��� v�V���&����֫�Hd�Ξ	���P���&��W�_;�@�6J�3��P��_U.�dE�v5�<��}�U�{p`�DZ�e��?���$��^�^my�����)��H����s��t}��s���'ASu�ݍ�E�l�\d%�^);OKck�eD	��JL�S����f`�\#�,��gۑ�x�����������m{'H��"��1ö���;w6�eؖ5+���0�e胖^=3UB�� ����T�!��a�k�,Ƈ2
�@���a�8W�8k��#��s�j�6N+��Π5e�m�������Prj��]���BkZ,;I�@d�APn:�1��](�q���80M��������~Դ�Kt���}HH�=��&������!%�Kޮ
w_>+�GN�cf�1�C�8���JY�U�%�Z�4`��l/��ԑT0Ą���g�k�e��.��\;��:^�`�~X"��lI���*�n��B3yZЄ�v��[�D	�S��vt�&��nR�k
)��FT�6V�bu��Q�>�l8K?�����c{$�7\��"���+%�*�(���lh�[��RTb%!�ȥE��Q��D���,�L��d�LU6�!Ņ h����mOZ��XE�#�9���lBI�,Ɠ�`V�!:�u�r�Ũ��'s~D�1E���*��E#��]����*�K�`�-[ۏ����ټ���M JSU��=�2����A:(i���޹w	I�T:\_�O��ldҠ��F��{^51QU�-�,���4�
�b������Y|����a�#�%�)hI� gㅒSy��c�jI�~v�O�m����]�[U*#��"N���]L����
�n��^̈1F��ee���K���Ѩ`Fəo�KY�j��"��B�d���1Z�w¹܇ZO��U��7�n��F��b�~�;ﮮ|�˼���r��5J���4�*'���?|���>5V^��H��sSi�Mt0>�t����[���{�]X]���(�d3�%y.��|/dp��Q�iU���ZƋ�̡q�M�UUŞ� �a�z��IN�K��9�����yY&E>�n/���čyj�:�V���(D�0������L:�f�I�EA%퉬��E�1�3���(Z����02���Bb�j�Œ�a��h0���r����`̵v[!�ID�ɪV�/�t�<������?B�8������D����N��|��^sr��e��sWo�����ϳ�I���EEq|�q�0��7�D+�{���)[t�������GW���c𶮽<g��!]��Rۓ,(}�lmlG�W��Aw����X��N�JZi�ӝD~#�	�K
��66���g����>����Ӊ[n�{�/��~�ѝ�Yh'�$�����m!���Ac/(��a�GF�� �T�,6���?�k� ��>�뫽�����$Q���CjА�x�?��4�(e�,P^Kqb�Z^Lhx�����q�|���~������A���O,�"���P��fo�����h� /��2+�b�M���툶z���9�!%��	F�o}�A��?{2�E��d{S*hs<�aڣ��۽����~�_��xm�念t�{N���c��_����‿[�}��W�;��zF��s�a�����ŀF�����x��?�:6hk�Sk\��,~���:���>Ct�mb?�m�J���b�,|�k����K����o]�����>N�|������^ɽ�F�;��x�9��g�U~�������Vxϭ�����7��.�� ��/nJ��ŭ�ɭ��W���c�n���n�t�$�~`��Ɗ�9�{��n|��`���i��U�����\���T�I�~������l��C_a�rf�@�Մf?ޥ_y�2�4{5������6�_��_����g��TPZ[O�ïjҧv4��!����o|}�/��e�~���!,+�a�f���ƃ�P�(I�O��β�17��=�ı�̈́L���?�X�a�&�0�tz����L#�����V��g��A�j�~T��G��G[G6ﻣM���G2�$Ap�����~�̿3�?_X����>�?��G4���׿D?��?���e�n����5V��Y`��8�����C����ghku���fh?lF������ ��~��U���C:�6�g��{�g�'��6��w��mj�	UR���V�N�w�M�>Ӻ2:}���Ƨ�Q��bP�3����J��,2ny��޳���G����?��	���n��?{�6�O���E[�PX�(f�h`�{��P�'i�v~�b�﻾����>�Q��2n��$iKYQ�|���oȥ.|�3�hϧw}�	>j�ω}G�[d�ґ��x�����+냏~�����K��#��h�P�x��̥mZ�H��{�����ڮ�������6>�c/?V)�B��ǡ��D�e�l��1����%;D��3`�D#��s_�����h4�[[[�(2U���1Q�-b���<�xt��;�W��� ���'�^������;�}���{{ƽ�$8)0��
��+m1��-����[��[��h7<�}S`�7��vzi6��m
��qq�B��{�;/ʜ���i1a�K9�uѵ/[�����~��;?D�w� >��k� �Bc���{�/�EŁ���G4��O��>^SF����-�'���5��vM��<���S#J�ۭ���l2�+�cD�<�r�=DI)��Tf,�q�����s������.����p�C��;��6�ǎk�L7d��H�tPG�v�}�K;aU��a6��~en&駓�G�˱g�XC�ূ �*{Т�+�v�w�~v�<��#z�^ۣ��x>�eH#y��%�	T��B��A���|&D���F��ǩ)�j�&��5� �=DnT�~�U�FgI��)I�n��U�#���<����g�,��@�3
�<�,5ʓ��a��%��N�(���f[���\���M��c���z��ߟ}�#���w���6dNlH�爲�����=�EQ;��m�l`�)3�1�a��O �[��@a`���i�=���i�����6g�>P�O��|��/--e�����"4��l:U��w�}�7:d�n$�Z�wX�,+�q�������ݼz�z���޹s����$�1�d,�E�Iz�b4�����=�(�*FW���CA�4uU��AM&�1s�� P�Ք�E�����|��}˷|ˁ\�=$�����L� �nw��b;��w���+{� hz��ڠ����`��þ��m�-	����1����CQ%�Cz֎�����!������G�7����أ���RZ\\�dc.X�����S��r� I�����_��_�`Y]�!z@`ԱXjZ<p����-.[k�9�(찰{�u�,����;�12ln�1zD�z{b7�9�c���j���0<�\a5�r[�b�:HN��������N���%�cd��z����v�в��! �P��L�篷Z:�c�*�tCF�:HM�aL&�98�7ؒ ��]o.�v�a�]TJ�S��U��X$ ���sZ���<;�a�����ӧO�:�c�)ʜF�-�;�0ؼ���h�պ���͜�����������+\G:�*̡�Q�ې�Qf�͓'ON�6��w�0��'�?(�����.uE��/]�pa�Ρ�>d§1s���X�E��t�<V����? ���/~��<s�n9~������V�(O��Hl����>:�c_����0V����JHu��o��V:����9�@=:�ʪE��+?�\Ǐ��G���<���p8�~�����ǎI���\���^�#j��ލ:Ơ������Fm6���Ks`0�W��8\/&�0��Œ����*�Q�5I�oM����8s����(v5�3s�Zݽ{&H�ӦF�B��,~�דQDw�y���?X\^��z�Q1c_l� '_O�~د�l:&�]^h��_`}�jN��EL��
���9�c�,��˲�Na�>�6c�XOyC$n�S��8��P�gSy�
�{OYi���rMD'&�I�l5i<�~��^�=��!�o��m=d���(���'?i���{��k[;�I��_�!������"�gB'��][]�Bp��}?��	I��/���U������d<��g������x�}�7��.��}Ws�nV�n+U_t>���q���"�S�h��+i6���s��i~C"�@Y��1�4�ۍ��ə���o-��(A u2����X56�갾�v{�[Uv��w���`avvV��g��<t����z� �*ʧ��qmfJ�m>C���'N�K���-��\ݲ�#ѵL�ּ���vG�8���L�+�p�=�Q5������t�����%8��rNpn����؏����ſ����fS�e`%��%���������Yꋰ��F�x_:��|W���@Y���N�SbTE������?�s��t�ͯ�z�i�0��%��I%��l?��[L���!g�8C�ǖ��|io3�j6Z4??/\1��7��3A����!vE{1���}�p���Wˬ�#�<���ۓI�j�؁\��o��z�m!���m��ڤ;è�����V7 M��3A@ p��;lR�^XX`���p>� �;$�6��J��L�I�[�����~����^�bf<�.��;��n�ǾbY��P�Ϻ��f�fgf�?o�1���|��R�*Y�����?77'`�^`���4rэ8�a�KQO�����%��u�A���Y�gky��h�����5���U(qB�KK��|�*�̻Y�z�(J�HG]<���?u��(v�QBB�6�V}A|��)�Gv���$�V�%�j�Z��l���`�[�쫶��gY�I�*<�@�E8P�c�U�"��6~���M�?�85ۉ�z�����fMFcTk���ű�����pI�ڞ�T�=nD��a.O��ZUY��^�K�p�`)��'eL���Q���9;7"	�c�WLa:�s��c�s�z6��ڏ�TY�?/��}��|�%�g�Ot��1�F�\��A�.3�? n���}���pu��W�m��Ho�[E�e����P�QMoL��h4Ja�vO�;�c_��VS.Y3�7�k����0pl�������%��R��^�/�j[����[\\��uz��3t#�=��ٳt��Ev��+HM��w����r���e�ܼ|���b��b}�g[��5Y�|�E�_��=���C�Sy#�=dss�1�����
�.�]��~����E����P�q����2�)��A��
8���ٰ{_��C�?����׽�nı��Ch9�F��m�N�+++��!�b��^_�6�5�8�y!������/�@�d)�l��QL��.��F#��QǞb��CNq;��X�FՎ�ߢ��>�}�������:0����Q6(�C!>k��H�����}9�(����d�a�1R�_�6d��8�[6�����,oP�s@5Y���d��my,Tp���j{�Boı�*�L��%j����?�������>-,,ҍ:�$���A�����A�B`{�~�/6�ԩSr�'��1�N8�Ep�_�u(�C�6�>����a@&�z�1r0�3���)��Sq��B�TQ)�]�$�۽1!��س������R��aC/�Sn��I\���q��)N�Kl��b���i�&�]n�n�"멢�/��;t#�	�,����V�`�w��:0�n'R�⡋���VĴ�t��Ug��A�Z^��laM�:�X|�S��l>��%��o�jZ���9w&�d�LF[K�� 8"�P�hU%A"�s�ʮ�r�_�ʅ��n��� ��"? C3!�`��;�������}�sN����S�x�f ��9����#�Ǆ�JH�ۚ���J`�98���y�O��k�Y@�5w�(;���e���$7l,�Z��V�_J�c�8�^�O�Y�`޶�m��t�W�;���Y����#���֣��2=u�`-U�;��cn���U"/`gg����ӏ�T�tI@N�mc�p�@��9�X��YeVn�R��1���3Ǖ�~�^���b �t��8V��(W1�j��½�+xL�`'���ֆY�p
UR���VV��!�5�;LCâ�Я~F���Z�<���~���~Id pVa̽��
z�1;�Jl�ȱ�
.(�d{\5������(����ڤ��Om��;�M�u%n��fJ�"��C��R�:[s���X̐o���pgܱ� >�#I8�6@�C� �
���##�f�jq�g0�Q!J�A�y����g/"��h48��A�j�Ȗ�-"$/�T�(���X��N���x<w���yIh�����Y[���0^`�\�4/���U��Q��Q��b�9�(e{�YJt��U!J�>�D'RUe�LjQ�#~��!�������#�YA.o|�jG�=�H���%�#f���>��M���4K(L�.�a�/�8M�S���7���QX.�V7�|����U�"V6{u�  {��s���"P���	̩8B���=��j��A ?C�^�c��L��r��B��%Y�u�g�z��5�A�������R�Z�!K*ggg�u��8#�B�k��\I�d��:$xmmM,--�u�~�%�"f��X�L	/�U4�.�n�7u��w.yc7S�Yl�J6��R���WW���_��&�W�������q���H��/�3�.t�*1f��|H����U}V�����i�vo��D����RP$��J���)� 0�co6/�^��{��1�Mc�X%�1�=d$�^��@_u31�s8Z�3~^-�0VE�ΜIP�4ȓ�c��f	lt�l�FS����3A��4\sC5�>�!�����B�xp�Q�M\��'82A���Iqql/_�	 ��O2==�`3j�3��_._n�E�s��}v��l��?��}����V�kqސ����hPfb`��Fc�B)��=���%<y|g��D\�������Dȇ���r�a�����Fx��u+7�"�믽�H돴��	�Ć�x�V'�5�Y���� 6Ta�bcGY����}�n+���h�!t��ûwo�ܼ��8&un�1T�;������0r:�ާY�$b"�JV���mc9�L���Оq��*�w����L}�����t�c��⢰�B�lnv��ŭ[?��wt���`$�a$������x~���R�-~�u?�U���&k��$I3)���`��̊��h�ka�	���ǚx��I�Qi�D!B���ſ��~���(/[>�¢^O�)c���}Z�hSا=���yJ�e$؄�fx띅gr�q=�q�!��O�c��8O�c��8O�c��8O�c��8O�c��8O�c��8O�c��8O�c��8O�c��8O�c��8O�c��8O�c��8O�c��8O�c��8O�c��8O�c�	��!�    IEND�B`�PK 
     ��Z�l����  ��                   cirkitFile.jsonPK 
     ��Z                        ��  jsons/PK 
     ��Z|�%3  %3               �  jsons/user_defined.jsonPK 
     ��Z                        ` images/PK 
     ��Z�U ��  ��  /             � images/ae1d0bb1-db79-4eca-b526-eb1d648f9ad0.pngPK 
     ��ZJ��F�  �  /             � images/1348d1eb-e6ae-43d4-937f-d455f2ad4bcd.pngPK 
     ��Z���S� � /             �� images/0795b188-35ce-4b4d-8dd5-08667f88bf32.pngPK 
     ��Z����=  �=  /             U�" images/28e7f2ff-99bf-41f5-8f78-c92be5544a69.pngPK 
     ��Z��:�  �  /             Z�" images/8d902f4e-ab09-4493-932a-1f1db25b6d7d.pngPK 
     ��Z����(  (  /             :# images/4c416a15-58ad-47dc-949c-f0bec13a5bfd.pngPK 
     ��Z�/��� �� /             �"# images/b5c34fc0-5882-471e-a80e-5adb517f5654.pngPK 
     ��Z��_2�I  �I  /             ��( images/5f4f8fc5-f884-4b46-b794-7d87214b037b.pngPK 
     ��Z A���J �J /             �2) images/36e83e0e-fd9a-4553-9782-762f273f5010.pngPK 
     ��Z�c^��  �  /             ~* images/edd00682-873b-4230-8bb4-282089490c70.pngPK 
     ��Z?S�2� 2� /             �* images/da48ab5c-24bb-4ba8-ab59-39208c7b2ba2.pngPK 
     ��Z$�8��  �  /             �i. images/b96c8ad8-7845-422d-b49f-326b2968fdb8.pngPK 
     ��Z=�W2�@ �@ /             ��. images/14f4e0bc-85be-4a63-979f-9a3c78ebf9d5.pngPK 
     ��ZH��X/  X/  /             ��5 images/78e6be4d-468b-4075-9957-5b4cf1a5366b.pngPK 
     ��Z���y �  � /             8�5 images/483af35d-09f4-402a-a8a9-75c28eb4643f.pngPK 
     ��Z�9M/�  /�  /             ��7 images/0a03a94b-1490-4d51-a356-eaee23e4f5f0.pngPK 
     ��Z�p�Z� Z� /             !F8 images/0c8b7e0a-6698-412e-96f2-fdf086dc4925.pngPK 
     ��Z���Ȋ`  �`  /             �;: images/457643d0-fb24-4111-9541-c1c501ab524b.pngPK      u  ��:   